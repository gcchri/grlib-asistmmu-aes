`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T+jH+4FR1I5GK9s91kzV1shIHZT48KmVT7Hph2pYvu2a6tVFCDY09WFFeOIP0520
scgXoN4Eclhf8b0dWr6OT7AdClcQGGOnHRAkpxDy3pqzZ3QzL2VRsSyq6i5Nvs9+
tZk3OcZLxrsmhxiW3TEHYPa7HsiHi0YAza4FlTzOOEdxrzYFflvl/Puv410kLE87
zRL7l1i+j2Whlpl1gb4FbbpyPkiRcgTbUOM80fkeIKio86J5xR3NPVBnxie1A1HO
S9JVIn37OY1QUcOUEl1w+ennIC0ZL7qaIWUk1MZxw0Im6V8YjUEnw4NgjhpfHM5D
m5b5ZlAG1U/qg15S0jScWwreW1Jd+WVaaI0I8H4ObcBON43ImaYMCaUX2EpCUd7b
VNQOrq1o876Fqk3BY4RbP0R+tGbLJr/UJB8sVckOaXCWvu9nP3Z8BjNqZ8w/UaLa
zrQ/Gmm1aA+JSF5LLdD9mL+yimlSZL3h8eiTDEt66EbupvRzbq0zFK+9DMZqlM9z
nN7F9vdvzi/9SScnlJfxi6hIDOq5h+J4Fm0lPsYNePQRXBvQFhlFOrRoOm5A2igI
6MXRVem40n3vxl6aw1A4CNfUl/MX1YvsA2O+hhYAhRwRr8Wf+b1YkzgKyChjqLex
B11USUxomnRhKO8qdeG8P8to/BBUAktGe5noHYxGhYbzvlYwEddF8YlsavN6cja3
Kin/nVR6MCIY3hCfcuYt9fiLMFmT2BcWB68H+0trfEYtMh6/tQodllwhUsDVeS2V
yyPEl6pLxpSqGHkrBLF3JV2j5W0etSNUwr+wH+vYRZMI0gKlqbP7RW0jK4uUEVyL
pAJLGggfbGNThkYlOdXi4olVgwWGnHHgrL73YIYK2TIMUpZWnxaKoKyhGNYSL+8O
HK+IqVvqCFJMxKB8CA+2IDoFO3oBsGtTNxv2x2nftCT6LeRVToIoKr+mW/B1MPSx
FiAraW4fK8T2rfB9qkHXOqemH03OWkkfdOOESDcKqnPHrg90FN8mQYVJXZjODGfB
8qJkZJBaKHexj/PV+vghjIqLqLn03opmxQ1IPb7k36ie2fcvtiZengvJgyLd2gx/
9Rw1zz68WaXaacCj0/emaVV2aODJT1AhHR68V3H7XVLxqgtI+EZbE5rgH31lWQ0c
N+K7fdvg9DUlKSACFczWLl41KIRLVYge0GKHX7S6Dhi/3vtmQYmtuVHtoMBuxa/d
QRgWH8HiCnzAnQrPTE2z/M0PSjlXPsF4zd+l4zLcWEHgYTfkGGmvf2pbJGg3lUkT
uRrbTjFCTfrH0duiLqvlgnRs1kZKhewGsv93BHDrYWjEHWWDsrVjmz6bbqMNB5fS
82+JZYCGV13xOFDL5tsZuV1FdaF6Qxl1zQht5LBFK200KUBdJ5SUB4p0AwPgCpGt
DJ+VeWoOJHtAgch17k1hWjGpgtVekHbta9AkcSupH3e3oN93y9zHiFiZMev/xoge
gS2EpYaY8s/zkdslQ0Z79mybEWY/PHG1f18g1Zk3HZ9+l3zcfxYBeSmJRVxNZ+/U
Mx35jNxERO2mVKSHBxnfC0GSibgoToSZodInLDTt7d+y/skVvOa2N7O+5OkezLQl
m8xP0lCCTY+QWbIV9w+pUNvwVvuGc1JO6rK+FZr31/LXinvo2U8Tb3/VabmMqBtz
3QarFUH1jXqtdZ+wbE4AfQZhH3AP/3ok9SbkjG4VgL5fSLhsG10dBoTOeTEjUCIm
RBxBRDevykHCfve/IeydeDTWgdCMfCoPnQgbD9GC9pVWwC/8DRrPtv2fYZ5/9cHD
0sPIR98xfJumQ3I3kMbdyNUwGQCc6+p9jpbGCUSdtjM3dv7BTJyeV60taZwmsNZZ
VC5Cwhq+axb0cZQ2QY0x+idrDmaSE2qsWBupOsWUwQHcPdKVma6eVcM8jSdzWefd
lHQAQRIZcbqD3+/D7DtALsieCGMYZfJhOCIlmc+u4/Ylgn6O6/fkCFq5ETJBwzLM
Xc6UiqJpWNgw/NRuT2HDPCMFpUlE+2dVMd9AvvcH/n5oHmO0go+mGQeju7aB6PuM
VJiDMCou//lfzjHNNBWM3l8BJi+VKp+HqZYzBzl/2ixckJfsPu4D/wUQ6rokrwZ7
ebasSF3nhjv80plWHU+zoIjhlvLIJ4xhvD+OcFXPNR1wfDgyqlpfHs69RfPu+zxq
Qh4rI8EcCX3xCETf5/a91fkqpNNEIRequm+049G7gN8q1ZFJzsGpepHfiNP1ZpRG
0sZMJpehHgGDOYDpEXxNSvBKAF1A7ulgQ2hyhhprTGk0G1r3sojIOxOotXRrbcw4
Lfo2tjihNQOURICPZ96JdUq5N31XRdlA+tKmIesBWQRvrfBxd2Nm2c2OVow4PG3z
Cb5xIn3k1E0djQ6QzwL82m0O4AUqdbNQXI64ddoFps7LddBTLHQLPSZouktUVZlW
uO1U1m+5YNYP71ok6/9lTgStKafF2m860+iNBCzqgo4KdnTuxIQ/krP6fmHE3NIE
0pU1v4zZe3gqIQPV58u2sTfMLjd8Uzp2uFQYoiG8+epjPxOm6toaS/qvAUrQgiw0
6nzQnMDGJDNqoXpGmi/jrrHy/bB6FEHJo+N0UnlVku1IGxL2nDFOtd7+GzTy6niR
WNnaYbKVAclZURNJCQfbda+TA9ki+Vq05h1DMWIZSkOHBVStmmCt++KSFzz5PX5f
JGnh4Rdj4bl5ew/TSlWVBq0SwKDDvvN8BBy1avGFjfE5fhRIZ35uweZv2C4c670/
TVgSB/nPChgwQmjLrJ3qGwsPY/6iD79p5fb6CRQVgFr950VSZODdeuFJ0dWco811
VKpcq+akP7pgdgdsFyRpSdNp6jDVgJCFEC9F3B/TCqz/sb8dM4YQ+box6mp7ZJ9Z
YHC7tU20x0PAGQf+t/zaHec/ggar/0mfu46khcBj7eDZb0PmfyXNyzcHWJt9j50f
1bCNc7/wX9l8qMMJUEavmP3MxfAMHPBQT6UtPdsA5LIty68j3r5LwPXZAFh4i5Y2
5TAmTeBrS6nSncEj82X8WbRnlVLxwX2spizIrie+aTeEW2VBEN5xjXytRECEBhlX
7bka+G3L705+wsgsDon2Cbr3moax4e6ELwXXQ97EfkMrRQGAAv4M1r5l+bw7TY8h
YLHZ0TqU3Ii8mqMBH/MN8MJLrHR7HhTAKZHnX6DUFh0p/oP7fjw7SNEPP/cQ9mAd
djm8I5mFkzVcNEEhL/q2SmEzB+YQZAmvvrHccOw0xahKo+PUfa4T+mVu2YaSviN6
/Se4J0kf6qV8v0zvFgm2UhNYN7VE/dHFDhgOmvvkuLHkXVs/4Tk9dlIF9ShDcKOw
ACNDdFFn6XmqGEwLaA/wzqdNHjRmJ/OEBxyICm0OY/80y5d/ADVeUFhDdpYZHNms
YZH5jZ+8ZR2oy2ACELZworgKDWcogcO733zfvpCqA7JVF9ppnzprJ2pBVOthgCjc
KtWSAXg7vq9GGVnGtR4A2Esl8VIP0YenH/WSTMr88s8w9rZJVXNcg6RAUjrCEJLU
h8BuvtCijVJGzEj5VxPIjQYoM9A8UeBuQRVR3/4Ep+zUPtS18BGAxiKTKbRyAQ4w
dRdHcyDqbJOcRkt2/qxkk7B0L8XXHc0Z/+98ks1CEAJcHK9AF+2V55aJGoydGHy5
Tf+JFcT3/aPNAuGoiITfW1D0Z5JxsDPBmgXD6BwBOmULsvN20fIz3CC6d6f/KLR9
xaJHV5OrhqgDsKsHIMKhtMptZu1LBbMyU+qeQ91B3q+WCaTAcTKGbgot6XWwQP8e
C01E9Ooc1FSMD8I/p8DONviQfn5QGJHDu8R7/d1pwLf9ck9wEOtehWD/CrWmeH1O
msQotg7rbKhFylDT7nsSy82Iepa74qRjS6Z3QgmkKBYBAntRZFOIehCIzor/PAMg
oEFeJoTvyyVdeRYTx0MaDCMzXrF9E1SZOEDuWrW1suH1r8kNAZnzCfknDvVKdFPU
6pCUnVKHQ3TKxbgjCbMVobsYGJWC1wTtplERmRZu+z9BJCLnXQHs2nA+1wrlImVK
yGSL26g3lqG9V4n7Mc+YeapT0d9qUA1PmKH7qFU3sI6+dnZ6i09v4tEGjyDz9vjJ
0XyJAHmY1ves4n6W/Tk8NHNSFl8GIrHe+VBoo0uAwoQVl6tv6G8AYmozNR+niEbz
lqU6vEqCyZDTZjiAODD4/F7+rzVeAiKq49SgHXRZU+iTGNZcu7DRmsx4dEu1hcqT
Td5VoSoOWDYRHMqBq+h+DP/+PF2uoC2l3sg5IL+rTpqskovTSly8XYJa3r77DAze
itMAH9XU6Pf+YuTyAV+51N02TF0510dXzXzGhNqA5xfpvYiRTb4gYamr8o5rWwv3
9EvU36hPk5aQqab8vAVuChiUzzdx8eXsU4NOVgiGgHsumkTw9yZ6Ne2tBWvK7g/y
HuB5jC+/no/na/l9UbvED7CIVmASSmuYIgVFcilxaPkoFAee1LSpfOfq/pfKzKLQ
0YTEZjNJuMevtu1vbGN2UZ3uiZU23ISyF6s3XIz0DOMXWbjeHtFFV/txhrifW7CA
+Lu4OGS0bets5oszjK3+/TPYtIZ86JCOtac4IbhIDnQ+IyIPEINjaaOlZoSPBWRM
EZMCUpVjqyG4aLtqatAJ39saqh3TyRiiwfp00Hmw0qby/k/cTZvhQVDRCjaZyJbi
NQlxLKic3xm6vrx5ALLseL3J8wGzJ/P89csgN3yYjgYhIwRaSccDlsxNilBO9ev7
JJQifTjoIrAk+EKmMIcPSKPwzKyT9hmFvUGY6pf8wVbx5zjxFwVSFb0UisCw1Yzg
IqKTdZ3fhguv2u6Ddu3gq8jZyPnpJerofA2jt0BIDbEi7lCWc4C0lPz50/mBYr9R
mn/KZ6Yf9XTVWv0Ju0sEV2v4id98HB6GrOmbE+O6PNnlj1xzSNgyO+ToNUoBvMOY
pEhZ9PoQX1mM+oJzH4ACVUmYMDUT5Wx/jF9ccgKayyqgpPUdNClWzDXVubp7biPr
vK9wzRdKuVcXIQ00PCa0GjgSH1ewhFhHRdOxNV2diFprsq4hg+nOAx2oXJnrd/qw
dFOpRhXpc/AQiynr7Mq7zVX7wIjVAyyzBwDLSt7sxEU7Wpb6D9mPqbNznD75l0vq
Ya9qIAO+GJZQ7q49N5V1XjNkVO8SPpVky/R7lP7/NuLDl5HMnfqdi+33ZPtD+hXn
XuPtnrvzXB9cd7tBn7e8K5OnUbwXjpT6bEYOe7I9HIP3AbrBMZ4BnySTxkEGtZxW
lPJRD0padkahhGEW45yZBt47LnKXuRPge7v1WiaEQMKE0B/oCRhfeesnkyZ5XW3H
K6fzOAKHN1zevFPP4AhrffR3+v92TlMmFoJDBZFc64eXCOXMED7OdEpxzk9DsN89
TvvCSmuXH7LP8hl6vZBuTiCWjiACBmpTefsPaIms8mQ24TEL0DZAWYZHBhXa0x2l
1u1qkzpBmkMFsA5iyo1xqJsDpNDk7meGbHBQ8crgGtf2YI0jWVGwz8+/ZKWov/RP
l3RrENA+IWOqFhIUW48l9L6lWc8qPp19GLssATdrRW6VpFj9ZdnY7XOjshuMwATz
a+G+ac4oxs0iB+Iqs1cl1pQEkKW4v8EjUYWuUXfRquYFta/l4kOkL7a2KIYdUjxi
NY1DLOW/XlQmc9DcP+ozEsH4bZAC9yyD/py6T1Oer1AuQjlMGHKDwvllJxtOz0SC
CS2uNWLK7Kq9FbBRCBtAT2Qq0isqQ+rUECxTnM9j9xWc2w6epjFL8oPaDlCvDY+u
EVzOy3YefrgZMDIw+fRULCcJCthymMjoUM8V5yYBercniIKa12XQfw/KNNRtlOrd
JbyPCFyt2eLalz+Rg1u4fOXwhB5L7YZBu+XqC6GkbABR/cY2tT/zDQEpKnBogacZ
K1CtGflS+r9+FfuGTZrSPTuxFyBpCL71hfur176G0OjUb+kzmzBQm2Fre+1Pi/Rq
vLXEBphBT8Km4sXpjOrI1BV/AOkdlc09lYW9+tqs1HjFaPaUXZIHpoHRfHPL0uH8
WMHduc0GQKoDu+Eb/m94mZWGUKQB3jlxe9DU4NhFmp33osaX1+RiTjd87HXIjc2V
s7C6ql8v3ejervMKudNShl61gp2gZHEWaO2pup11S1OfRDSm2F7/fXM2QrSB8+Vk
VunqLy3muv7zTJKEmH1Wkj9APCFvYPTNsR+8hqZAllpdIiX++dctYoacA+Fy8EYg
S4/dykIWD/C07xnSaQHRucfEjx46WY05ZYIbjOkN7mbBwO/8F2kXkw3yOkGQOx5y
ayHyYjMcDyeRZLxStPzsNray+0rGZzq27f/VUlAgetG4IzhhWq+oFtB07nsWmtxp
7KnFpuiItBJvJFcg3U/az/JSV1hdXb9PWhtB9OsRb8A59I82pxnU7R4c90Hp9K6w
uJ1MHJjtZBMwfIfuB4m92m6riTQINxV3npPWv1AYg1DeC+Ijzgy++FcjcVygrG9G
mulsBZeJP0f5ZZqH2i7e9hoQ2hfkgZwUu1MztuYry5Z3jVhPbIbcEoUjs/Rm4w1A
bCV1MwQC3RvFHEu5cVynGeMh0U/59JM/yG/9/aGh89+D40blEvgIJIvakeAWo2qY
eSasnstKxWxfZ2cVJymtrwwWkUYCthP7o3JODlylSqgW0S72z5tzinIse/0/N7J7
aUSRY62LYcOu8nRO7KKMuoeqKqSCvouVUZ7MqFc7aeelM8Y7PBupF2CpmKVc1E27
lsZf9qpLSxc6zD+BB/kr2YndtiH2+FP18YZAyKbRy3WQx5bpDUyfmfLs9LcZ1rIC
LYjqoKY38C4XhA97PeRPmgakOhOP+j75CAHwPpprLCYtZssAr2uRsHhrGeHa/sbS
eUHZqdvv5NSAviRG3p9Y5jID445SQXAAnmNsrL1p2/sUe42sqDGLJruQqKGvfGt5
2eUe0TKZV4FqYK8pyWZYA6g2z9qDmMX8pu6d/U767s2tskt6SV0SfZ0YfNyb5DSt
e2XJcvfFXXmJZiiGZHKm2QjI5beVvBxEak86a5eqH9yheq02ljbLeTdxeGB9Y8J/
/tVXHG1AFj12PD/S3AW7W/rxeq3jc9PjIFdvHQbuaWEEovY1vXZq2w5AZdJFQCkU
kbqpErB4Gmp6/XNKfsQIrLHwnFXqQvEKURw2jn1YtPdEgUt7b/f6VLPFJbcfT1pC
igAE76zmEMx1HcPjRTkcxlbJz/pbIYCXH4GpOmeGergn3O4zE3FrU0mI6IbHcR1b
gDP1EcqJXMpXSRPWRoEbbB+EzoF/l0j43OJoL1S+dil4OP3n/xbONt+A7SZIsvG7
hUIHm8lHfhB8tM+Fej7p3f9tjzzi3JXaFiVQ5HsNON3bKcghSf773OzRXtmeLJP7
JVlhJtlJx/z9Sf99a1Ft8YsFTPSJDK9H/GG0Y4BA9ovtmQ+dVJmUhA+YQO08Dxiw
tYr7xuVu60CFYNbOC7SkvTL+w8al0THbE5jYlkXuvP5O/+0JctymiSVC2FK84wpm
qVu8W9Rx/tNTuqr/F3c7sJS4ajMDkeEYCPGaQRn7L0JZJ6LyEk5x3Lq8BSp8Lv3g
wBID01roQPcjNSlSu7fft6f4LXPEOinQNVSkQe5ZSR0/YZnvldhBDmkP0A/yqwWO
CHENRjrD2G6/Rq/GnN++QJkRAPnaRok1iPpGRPe3HHr+WFyvW1J0TtrSY8Fzr+lM
S5a/m79Iukye9VGiVbXTurJFityl2g+0daVer2jjOi+MBcfjKYp8NUMFI4XoD4U5
L2HyDl/rQ0hPWQ6AojQ1lDqhmc/q3OQtPW3Cwb1/9Y3fJRC6+z4fwOjYeP9j/0vh
9WCm7xplUzQraEtdPDOmYXCIk0u1+NivGuAge1HL6btVRkNt/7xfwAsV3koHzHlk
/FgeBPh+TO3RRNTVX1gbwA0m5oJK7D3O7XA0fKAKFaTE+HkSVfu1u8gu555ofohJ
n/Gre/T5yBm97I67trmMFDIGF7L3oBYsa6b0tsyddFwjI3VA6m0JWv4dSWGZuIte
HOpLmGdL/10h8az70abQ9Ap5k6LXWztK8Gkrju8gLmoN/CiFeb4QMiqVRoe3Tzth
4LUmETRgwxzwiflBjjZ0dyyteYhLmSjx+jPHrA8VU6Gdb395peg6gcScnd62MDDI
3QPPgRHiyTYtmgMarHsPgzRVs8E2/peLhsND5zN5SY9Ty2FiumNu8/VQ8QKw99oA
fpqreHo4KL9LvtWz+81ohD00t+V+Sr/Sq9CGVXK72MLnySykZy95zApkMaPVQdY7
sogQ0Rx73Xnzle825qX6FABr4NAjPw3v3ZnFfSOaNlLd29ZBMLMYS/5IDX7db3Bd
BxN0mK4WHdEg3XGbq7xxvvkjM4EODt/Rwxy92Mczw9z44PK8jSD+WW9NvM3O87Rz
FRSQItZ2oORBedsliuPUbBjbvy4UTtBEDy1wNy+hh1RdXPKXHEj/fzBo4taZj6hy
CkY6IaL7fqWp6GcExc1gDdWiAi6RhNBpuu5WxVSm+cLq3/hnZp3WVrUUtqczQkPX
ZnansyyvB40l9W01HJJBp1mklwtfUujEZ9IPkzREdXP4fl8FJO48dXw19zW+Wqrz
1ipf6u5xMw+mQTo1DdSY//A6XroSybvaMjISkOTt+zDqtRcNbxZ4Eks7BS95RoSd
2/waqvWG9x+RhbIPECny9WLJzu/aPVXHv7ZBtVOo2ssTgoxthUyNsah4zQuaxqyK
hBk4VI0SWcPUFPWkIrBuuXrubSOTPWPuWBF0pYF2icAkvpHNFkUQvc9OSm6sMJSQ
GCSRC6Jos7hbpCZHiBGKGB7PYbi9K8+ZSh4rsIFwmPDqsytIVaz15NtFcGkbcFiH
ghSmLt0HJhD0ZGwZ9C4WXFl9GnZd6AXCIoExjeTEvXeZ7nhqisdkOnaw3cQQ4k4H
ywnhzCrei8xv+Zja46usDgB4Cy+NRRh3TUqaGbJjmfpwSy52NFbzPw5P67g5Adbf
O+B03+Vo6RHk+3O9wQR01JW7goerlfx57kb4E4W+wGtyOvcg5YtXgj7tIShGQJ6O
AVeUvfRcXxaeisyErg7LnJG2SuSwGOtAcwmMcErTloSUXIWwfCni049j8zqNfsQp
5SOLES1BBQ+xvcRd6hbX24mbdC+R8q78VxqQ8Qau8kpEa/D5R4cYLlcJrmj1CyyR
V66cCp4ghPRFdvSGZNpUGssbOrvDvw+HapuAScIuWgnqe231PTo9xQHB3ziyfFnj
zea2of6R/fNcdtyeqRu8v2i70dVCEQLEPoeOCvAhC22geZNGq+zqNQ+Zh3SFoMP2
/INc3aBd/s/0fDyVTtb1GOf3ppa7zITDOxmnc6xN/yiRFQhKVU/kYCmq9CNntSHB
LhOkzzdad/aoaRKWuLO3uMyn8ndcUGxL5JgGKmePq86szUpF/MHXQ63NHr7lK2zr
3uwkVq9VvfyScXivK6ZBky8SM5ncrnU7/4ZKu0bIofZbkzhEJB7DRm99s2Oo/6Dr
YHeI0sqZwpnoRBnh9m18wf6vKYN2+ALhffogdQ9m1qf7oK+UgynZk/Kq2876T22Q
faBaWNnANXdsq7k9FI5TrlTRWXe+Ob4657BU+WQEtVZAXixBd5vM5sNIk+rIBE+F
wT1Ot77RV45ooYE9DF5uq74GE5yBpuszS8ued8e166z2cryhruY1twd/xjbESiRj
IX8zcmcEcLhRkuF6BFDkqsaCUlqb2eYeih7lq9WFId86pBOpYJvxByHXyQA0DrXN
yzYqu2aI7T/hQwEmna08i0FW/6EB8FzQ1JK0XkbT6iChTlYqd3NOGN0Tk4cJgPjq
+sK+xI7q5O74uPpyDHRxvcwzNoRhJpObh+KgJmBtAkU7FYh4E4y0J2OEzA7Oq972
SAlp2qU4toBpsu4asaeyBLWf1VvcHO3iJuCIjLb+afK96jvMWDhXZmpeNw7EekFk
DGGqqWXf+IJRShLdxmoyyu289FYgWwBkoyukE3KKizTl5vxnScCv8M5mPZmv728G
uNFVYQwzudzGkFcThnTocksOS3c/pC6k2xhKNBtBDf9abGf9eCfVzsEBsnzOVb6i
3GmTS8TQjPUit4j3pFzWoq38LyIU77Ah9syDR4EADSDCpvDgQpBCekWv3kgIziYy
QPYpbZ2NRGVQTRdZEc+Mu0rLHU1CGRLZozW6qs4IWm1BVavON8E76hshSeL96f8E
ni7gOZQwP3YhxECdJwRuuGwnhYgAT4vmVinuqXFwosziCWWcv5zL76hNZXd50Xjf
0x2jvWPTjoKkM/FWHXixyuzWf0i9NyTI6IY7l37DEw0ZIkoBV/WkCZluSihq0Csn
VW7jcw+6UyzXPIh6AqBSXG4OwQkxMaqqkm5P5PVUkmx5nctm1h2yrAx4o8FVVnMG
kqSRDLmOyRzQDwgnVcvr4PwPiqKdDNR1hZfpGmhVl1NrvlLdjcxvKJ0OhcFV0KLn
4LTLR1kXLtOT6oiIS+JZw7p2WaRuvvWBXNR2DHAIG6yXSHnQ3gUYoEBRmFVYBMGv
lk9Hy+P8MH5+EyFjjTyUn4XdSGDnaX+cUiCWxtNvEOMZ82Kb1HQqYyq4+BlZBKQG
0F236tQuuo/IPbbECyNpLRlyrbboGuAZhBo2Vf9quY3PIW0nek2qLmaGJOtM1e5W
oMa7/SydAH4aB4dpcLXhdNakGi6MtS07hk6kMDXw/iszPc0azE4fu2zNscTe7tht
K+f4AcvUHe6oaJLu3T5JzeINWSXIot3OhO6piXZvsIWsn9L6OFZtqipkIbL7/eif
ktpsLH+ejkb8r9tNRo7+tagilXceXutHazCg7DSQ6NifWxE0DEifsem6QQ39jqwY
RROfe2ta/CPdj+U881tKTPRFLxSMNHClvzej5dxIpkd6wKVKRaP2/yBjZSk5qHCG
agq+hKZCqS2eUX5eLT9ypNbYOSuXkzXpcDy9TeVhY07CLsuXWVzW7z5Vird36PIf
KM0UOrIa+2zKK+czWZe+1z1Q94qOnfKRdjfHgF1S4guUMCNvPMoDHpBOg/P16/oP
CxC7vkDdD6q6qd+0DRkfT5lMs9G7PjfQvFHpK2s+/dJPgSj9aF0XJxBBBvM2nZCv
UkO8BrOOwAtaEqS3hHKDyhlYscp69jF+L50EDHTabLkJqaEcG0ovW7MRnNAXbMc9
EkjvcpbiKF1fvAcTWXGQNgiHBDwcIM3ZBjBPcvQkGGlzHMhlDp/m9hmaAR47KJmi
nZkjHZqkwQGbdXoaMj+VSj+7h3qSqBinNsdphr97CfC918TnbbpkQIvFaVYSU4K+
TytE2TJ4FpYR9ejr+kxybicEjlR3+WIQIj9N4zQNS1iQuJAzmEsXmL2Y+K+lXOKs
4vIxEQXOXJVDkHxHYzxDW1rzqphwHXvYwV1/RbwaTUrDoPx94+R+bRPmrb4QkYpb
N4hFmFi+T59F0heZaJ/aoimJAzi8uvlM+V2Hb6eV0aHB9Qf50hV1GOFC5utTkp71
cM3bVwvEYycevq6MLqd4Ktv8pGMcgjEjnXHpCuoOud/LrPH73u8gCJsAgf9yPHwK
R8mveQZohdNY6nXCjG+8OcRHU+LPL1IYU8gdyInNGrHsne0lxQsu+UFYGtvMWnNX
SdbpGsGCvJLquJrdbB3JeM1GwmSJi7Du6XeWL5Cc8xD5oNKX7fYGnjDX3IRfJnNc
qVBLee/naHDwv7c3crXUsy/EwqfPBAOE7i4FzwxeQ+ANNxl6yo3Nh3kdl5593rs6
iD4xZBNGB2nFyqnjTXDT7fFDKgA6Oj8PLo1h7TdERLcPWoYKP8WE+DFIoWlZrlw3
mgfYiX+6GlpanXM0noMQVnk4rSIiI9WJJUV/gQY7y4l3/ui185VnlT8Dxl4jPWlu
ShROr+FZurOIdLGeA2k7s84azzkBlsJtGmXgqFifjZbpzLxxd8x2vyp0vp2fp/QG
nH/Id9DjS0zMqSmtQLAkF4wSCRE33Ae+bZlbPrwtG7CFOFv4IjMtMB2EsbHPSim/
NlDAoNNISRR9Uk+pSZ0q0KoZjFCc9UeuQCxyUtxXrJJTb4VTnMaMAezGT/QN50ae
0HKiko0l43O2SMMHaroYpb0sOxcfT7d2haG8d2TpChIIyyJ9WiYtbY8iZCMOj0ii
rhkoVYM6Tt4GpKrwOtDuFnFsOj6z7FQw0cRB9XWbB9ByVSOdeOBgSyqMevFwQdKp
GqFa+TWS0/RvgTG++XWr9MEWBp6n85O1i3zG7Lg79i7srZKVp/PVnLAfUicVFhcv
9JJP66bD53kTbRGiNBLfW/4GiaYSnCCux7JbN8tOMcXGoEvgWiYJujPV/jmOGkfA
FW9p7uqu9qroYSUdatPuUoj2cQDCIx1dR0dyh0Ni5ftTjlQgHuRtUQIE+cVZUxOG
R2IuqrKLgXypo7O3x5RT+pEPKp7pNrpvNDpPpVAeWusSPDTHUXsft4RAqSfRVuqb
0HkshEimh7wOmOfEmnIqCV7ep/ZEtkyiiJDpSg77c97rOGERZLiV2t+9uXeg9xXb
qXC7xWfXoAJdt2fNDNn21PRUT0wRYYVC2Dwq5MzLe6cQHz+k/fJqEgPM27mzrwRC
/BJmiLfWc3ub7Kg9hazsR1uLOVZlAubJGXGzRuz2ez+uJmJ2gnpv+RTwxgin3Evz
qbuyh+KqSSqY3q5yM33xWV0bZ91A+Fa0ekD+EpQv+s7YLgT+t9CWGB4XfWD/hiI4
rif3PxHhiiCj+DpViWwiXGfhMEOpAPKMZhYJnB5Smk3aAMtI69yTSrOuOEADI/yH
DF1B0bFV59oO71+JSDIi5cpRJDU/xz67ok8rfwDf2QSUY2l21oV71tFI7/ythnGe
96nY1G2XSSMbyXHp++fKHc8T04KkP1Xsv9X0Sg91rA52kPCp69S395ain1iu19cw
ZbPxI8NHr6DbT8lTxjFNX13fiRYmwuMHSAeSIA8tvi6Dl6XO/G2fXypUZWkn2jA3
qBahuoRUeFV/5+yYpX4xKFGKlVKPAri2SxemcoM1nNqIKguZjyFqLgn82l8FpSZx
0Aw+hjn3utJCDh0dvaMcdoCHlkYpPOD8r+4lGPCyGREjBfU6A4K9B5PKR9PuO+VM
Tz7rPc5hPdXOZBuEaoX+QRGnPfcmcV6XnaAS/grtFeJILjCrF5M9P1WGr90XEbJY
Vco6Qf9sOqR9WDVDV8D39vkUrZG0iBL+Gq2JGsQKzCOrmnzt937IfrvhM5C13/t0
5qngtZHAoBynp3iK6172Cc7H13E2V+JLmn9/20huQCsMuG/1jjA59le5OkO12mSF
yBY7bHiZrToRRaF1pBW1oSO2kNvzYcUCBThWakPf6P7GC9u1SMfDTt3VMtwvUcVX
57DLhUpK+Ewey9bvzBafJZF5YGgvTXI3qYTMkFOd9n8QRW7C9BmgVfDecvm+2YOb
wPje0iu+xJsesMXyCFvrsX9TZ+Z2VhUQ1PeLHXBp0AsDmPdpnkIZHB4BgCP7Xq3Y
jwg5T17UgqNlzh5Qu6ZtlCrqQ++rjIHrXS6wOcDvCJ+ObzhCFa7P0zdup4BG2s3m
Wq+BUTmxpgy86tY6q59UFHcM5kliFejAMJlk6h2jwy/Y6Z63zmIR+MG5rP13XiGr
cLcCLxncTWK3egZG7B758w+N2QYTayAy5zZigi8U0WWed+2g3GsjdWMcLxbmM9lL
xzPtFS0PW5tDYu8LaWVMMz/g/xIxK2IBnd63tOsN1OkHe0r2Dkq1vvoRmAWkE3iN
4ZB1KIRXM+TF3wy39ChxPFyhOT6PfXyL/UIWMkl1kpKG26wIGDoAp3dSUAg1QKmZ
JgfqGSn747jXeiDgyCEC+Yoqdo0SWI+2Y6R3kWfn91qSXDtPdJ7R9Y5Yk0Rfi2Fk
ANZXa8U6LtmGKyH3rB2Byf1ol+BpIbWLEAVzETCvofKHysMg9boK96rdAXpYWQKM
aNNJ7YQn5Lu/jAaqa3WQmwQKZzjaettrulE2hntuF6yHfiEgTFvXoVhmS7QjrZmF
TdpVARfxVU74iosSSdZltc3rsAXCU59iKWU+E3lkH03SYGUsBV55S1n0w9/8TbKJ
uhm7wZu1jOnM00aA66kUEWB73zngMqy3jcoADOaMvz4JwmZYPhuPXFcZ101dJueh
AXSCREZJ2oUxy/uS7Z5L/eSjBKIgMJNBaUbT3obRtm6ZKQbLnJSECABjwaZwaPfS
P5T/iCbIsLJ3AFx9UR37PAW+pqioj6X8osV3J8vponyiJl10zicivjY6shMSufZA
43i7k1OrLbBGWODauZPkoWo/hK1mbNvCdye6R/EQ0xvBrKvDnLK/BEaWpf0Af44P
ev7lss3YM37APhTqieXYhrUv+/dwjOCJQy8vZnkY/zpklPsbktsg2yVF9QMYf7tp
P1nUJu/6q7qk35Xaf5ZsxtoESHy0b/EJZ+tIE8njWP9JUh9J4gmgzzxXsbUU7T5Y
b721EDmbILUuq3yhw4B3cxOHc7dj23nFA0CsH1AKQXzqYGb+JW576jvyLUV363Lz
gLwmAAn3tjp+OaT+FIxUI/cnGhHeBf2j0/Le+mFTIFGPVMFGwAvpMEY/pT6FKsFJ
xabMx87XKnz2OiULA665lEvVfi/S4OzmP0V4x8wc7GmfbD3ZPaTO6tzpKyLbCOeX
QCVh4QW1HqX6y4dcRzi0c7eM5BKIKyEooQcfB3NEc7AVnFLk+j0BLJaoYZc8UKOs
MtaMkrCqBOs2Y+RM+JM2i0ggxp4s/G9y1mlzlfgXEpSrSkGq17UpuVOAOBjm7ED4
vo/3eFta7FJWOQrH8PBPKhEjLJwp+zwwbqupynM3S2hBrQotsZcLNfaAZslxUKjQ
nekpgBzbZaicSC1fOs/apZ9rOxKAvzMycoAK6ihhAJbTVSuvnOMWuxRCm9psZvS2
jntkPSw/wTMgMP3yAhYAQM9CUh7BfDNswim3pboJF6pVK7VxF6erTDNenJedK0DO
ye+u0QnfEjIF4zATWdEjFPv8MHG/bGzfcNmq1ItFrNISZDGJljMyoLguVZuagZMA
ZX4YatZJR4VWnaM+F6HMNatf3Th3mx/YwsdC9b2WuKwYRqo6C8gN1F6da5JN/aoA
KFT/HiUYJqiNWm+NmSCDV8heH0tjFsd4I3mPd6dI4wYHOGpBcXsiKD68hPpwdkz6
kd7seIBq/Ng1sITIeSEZzbDqlK6LPNPtmWJDZT5x27GxktDZaa+iG2LZPK328EQQ
suknd/Sch1mXxUMQOMA7rOLGRBqy6v0jIgh8wT8dFyzZpNL93GnP4ddFVO0s5W6U
/ZgRbOniLmrGEHppH/k38tOyVOhfgQyYlm8g8y/wiluk8PdJwb/yp8J9PhWf+Gh5
poQGvr54PXEJLS/bukz7sOEIW9dG6bBojmaDU170LFInsK9vbdZJPEdJcnj2ra94
jSEi1AvK0Xlz8lqyjn0QuSZKlDV3ZrIq/WkTr0cuWpX7sR6XrqCu/qQnoQBLK0zd
Zon6mtC1GfCwr8tRFdTY3zrHaEyX0Xn16TjxDQCjYnQkjST1w5nXcmLZMjUYuM4K
fDp6GTPeuLumZQFz0CyURMX4+8nHQiQqMdGfg+mlWVOcs5ovB+mmbeulbH2622MM
nLUZTxib1o3a33oH8T/DfAYj6dhcpUGrwEB0OSEkyEdbF7qjPb0sHFXqEfYzuyF3
lMRWMiuhTsn2+Z3q55Z/nGO7YCSgsuRXeGVXG3ZDw2K+UnOT7vvmZTgpMBRr8IwL
lQNb/DzydZeOzDUyeERYBeNHVEUHLbfIeH2CzIA3FBVS6+Mr/2Od7exOmS9dZjOP
Hz42FbEYcldWMzT1iOeAML5JQa9V+T1ZfeBtWgdt+f6kctEsGNVBU8AjLARDCMgA
NeA8VWUbcyrF+hIAuE+SscHuwUIobclP8LTvyvUGzmVd3vll7cOqfKwXKy2vDSZ7
0ZnntRBaU75M2LeNM3aNBeMZTDNiYDfuqr/8f/Mi3+OGp86Xs3gNxpRnkavqaOnO
sTFrlDk8oCvS02lZbYfWpXiALD34YP/jPhCKaBIhkQ9iMlXLzHAEw5JwnKYlXHEB
/xR+dR3TQ6WtM6ShW1cuuK5ssQhaJ+FR006rABXNQCTTXRnLDpZoR6ttBZ3eudnY
T491QhAqycJtoW3tepJ2IJw7fmHzXGRvatW4GFrl5nWMNc4P29sNbgIeD/aYF6TK
nw9t0UtAQIHz73HmczpxqQH3wfJM0ANTXp0Wu+teY9Upemv6zdmJS7PWh7fhTXTE
3MflvDtpwH59MdK83sM8I7a58r9QLaeg7QSB95kgF/kqbRFTimJfGSKbQAx3sYzj
sfpc8q8X5eRtSBSkbE2ijU2zE4E/u/6HU0ZbUISPBl4hoyJN4U+vsoLIjbIYAwQ1
xuQTr4JJ4RXJsBrr1sVH3mOYz8NxN2l6D71mw8UfGFm8bov4iCEHZlv2V35DprG2
TMkoiEn6/pCMJ2QzsVK3UJTT1nASqqWmkqx1tiVEcQtg03NScL2h9UxyDd+o9/wv
5zCRHPUT0rDNuqRkq4JKOhFFPIcpfRObDGIBFBU8eOVsj2hHjj4fqnlRtv2NF6qB
5PCQFV1zf03toUYs+XbFTSHJsW7U0ex7bzCIdVQJYXNgfbjhC2UvURVCFuE0Fwia
0HRHoPwhKBhEtIUENaAlJvOV9LkjBl3XkI3YKM5NsOTIYMUmOIP66FiKiqWATDD+
7ukyGJ06UGyVCcbYuBa+jwSPlwvd6MNw27kLGG17jBUkQ0GxcENi/5xwt7qHLMyQ
s2RWQ6Xgs+KSnO+DKEBiJ1hOVRZ9dnzIP3eDjr8vTlkEGsmI+o0KwtndCvzYByus
MokwuzXhRbpAgzKys2ByYqDjqo508KOdprMw1QnzA9i8CMFUpqYKNREhlRWS23d7
zvvDZCpC6rjCw1qg22w/tqTeD914AKOKKDZnxQJMpIend4ttjilAzGNTu/UduH5Y
Hg7HRFTcf5JYz1piOw3ByQwpH+aqo5qdGrqs9NtjSvXtF9GdY/CIPbGp5XsKpNSB
vfSjhmmC1NrLjJ+wUC85quSvwC9btMr90fDz3/AK6WKDtmkeLUlgMW9k4kOouXYV
aR58xuMIuZZw9S//z3w/6pEfCx34AcjSq9/bGIzL4UN9gIUF6wbIOd3kHNvEK7Yf
lZvBXDVQohqftsqWkJ7ZHechKg/iuIjgB3IdjZ3pUU21uM5cV3ToilBap0/CiagU
W6Qmv2phhTRIXNa75yIQCz+zBkp+QGqorMjO2f4dmvJSlpK/ZvPK12+tgYGGBbo4
CChBbbngREiiWRDw//4g7GH1hlMVHrbPPWc5sDqTWqDUnI/+OIwgsLV8L8gYD3Bd
rXeNEPY9KiRN17aTjPPnaYq4XFZruywjCo945iuyO+iz7emeEUeY3+C17sUNvJMv
CVYVbJGT7X2EGbeoeTNb4f6HJQIM02OX5GRpcwR0HlT5tJnsX4soV9QqA5VXa/B+
lJ6WlPnaAu0FNJaY0OJF90IVW2r0QmJ4MOwL+80BMD/5ArIhTrGHyZSbwHE4JPfQ
D8ebVKdmI9T/guXtjCLhoTJO9w2hyAiJXa9Q/rCnOFRADlL30DT8BvbceaCTvUHr
H3jXTgv/o+IOWmk76DtlnszOsAwBX+hVOzpgnxanO0qUTmd9iKSrGPZJMSy3h8gI
BKcFUdZHz5KaHITGKaUcIUi5pAqGLRDw0F306XEV0m2TRkBxxyJyJBntHASV2nyn
Vk16mBXdK4RxB7f9tBt4AlVQaXdFYTFcKU/+OXXtvHCcZ65Xe28Y+WiNHlHV1ZYA
ICq1KQJL0sPhsM1EB4i4sow92HTtfxwvT5BYJu3oXrsGuwfhT/Kq6fO5q6UWoGan
G4PN4KDH4Q+S1nmUVrhscRxIy+XO1dCLD0m+Po8ytuv3xuITworGvxV5tUeyfL3v
3s9N9sVvCFh5EW8zUa08Vs4IjMSxxFHQowzrjCVKZy2CDNFATkISoyY4/4jhLapI
FYXuHDzrtJhII8dFFUHC69imU8GYD+Nl0XsXqXxTsQS0cPr4owpKtyFXjAa7TzPk
0HWxVL/yQU9L3KcXzAQ7NheabeI36ckrCapHEZPeBIt0GXgaQVCyjhh3Lh0/oEjx
wpqnZ1MeVj8hmLoy3KhwY+FjhtlfHmZqQuTx0CK+i3+9Il07V7X3R4NeUddSl0lZ
L34P7ULMGNqDW/EspngKvjUHYlriTvAD0QDU3+RSzRf8tHw0dJmGTKtjugT0ojxA
ZDxgfEvvAJa4y96y1k5JoKBIfAhUCQ7Rx7HQ3LVS959MIBUds43lBWmfDsrGq6lZ
o5N+U9Ezcl6xpGO83iPmTs5irdPFhOYRZq6cTntLHEr/ygMUIqy6ldr92aJ0+Uee
rqMFnOZ9OnZkpFVFPo/ageFqQQj0YLCddIHlZoRuca60uydtyZIIdMberZvQzxV/
WhLlkM0tF4A1EStiIp9IVwbz0daW36FTpPewmqDiWqzY86KgdVn6wcutcILISpU/
a+xXrmhh0Msu2DYhjgi1UVVJe9esZIzNpUKptiuoLHfxJA9mYD1VYTjdp4nvHYxP
TMJO8efSHiN2oitre0UuY+g5A7tfOXWOjOVUMSqg36ReGvoFpqsMfFzH4ApCMA71
8l16DqVowd84jjuYKjCxSxkgYXXTIVbIxku0JNfpCqb4+2xxTCe/8m4mmyGFSH6V
h+b+BAqvEqzozfm9Mys8O7fkZNsZQ0yvyjcrEbo4XYGDKGhkhHSEI2UU2A/6GfA2
kmGqfBg7yRNSbBgYC9B9iG0X+m64DJ/qc8ZlsgwDGx1aO4kntyU8apDz3eWhiMik
jS5ysLm4Xsa0S5085/+4OhTeHBG/OQuSj+Y2M6JD/m/rUeIDpTAPs0OMH5bHTzfQ
mqFMyH1sRUqF5nBvOf2du2rzxXfd1mgX/YZVlCBR3YDUeicULXLs7UecrL1cm28D
AIiMw26BpscvYvKqnGDAMxhajd0VZubQ/Vqk9JQVjjbla1O0j80p3i5PDxvrg3nb
8/Xad7wA11JgG/3MeJh0pxKgBCfFAvYmNosqFw3YftfFAgnTk4FKE9QvchqTlBGs
LU2ywPEZd+26QJaVzDP7PvZnVX3J9I+8C3nmXzKDByJIe6zNGE5bk9gpS/I3Xv8H
gByWmbHU0Lp7050fGDNOBjfvFf32S9C0DgeUaXUDvaRoaaG5YqnkZPq8cZeoj1BL
uczkI1ylEhlUOZHE6HpK8dL1x3/J/xyFlRqCcZ9S1p/oZgytgspLaO/SlQCKCO+s
bRntOtdc9o0AT+qhTgeGbX6PtWnmzjcaVoSkFAG+kfIeISVF2qIhxXq5MwahOlji
N7c/TS2NX/+FoeYl2PZvgPXoqDxoGHr3shjLK2zXgbX+F6q6DV24BhNVsiXkrQa1
66DL8Yvhu7jxONM/BsHFuaEtNVEjkBvsJ3rp3knEeZCZ9EpM1l/IwWNd3ITN2qrC
aR6Ykhkrsxssb+qjtxF3hc9EH+PsBSKOnmOtyrghRR7M/QCtt74hX1hvaS5V4ids
hpbqRo43KUckDV8MTizCxVkup3wfNiJNNuiRxfQb7nJhdkXYaAuSnkOAQjujKTOP
bfp2V+pjHkrJDyFt1Ss2VvBM4u4ZMso8pRnkrSoQMGUFYWsJ4Zih2zawxqRekNQ2
lPtQo/ytDt0mGEvzitkBQGiW6QeVr7AfTxMeYjIycThMwLdLoEEycXdJEab89xB4
CkiwYlSs6azWxX+EsJLu26O8PBY1x27ISC7nIxwYFRgCctGHJXM+m0oUwW4uMV55
chFnPByZbVFL6zLTjQJCm6dFiEyQhfT1HnspJMCTspyul2auVoK7NrdW3qK2z7Az
zY/qssDogxscR09+mdqMBMgcc5o3etmQjhjmRfjNupVW/Xpw6PK4dmXLPaPP/MRO
DhM/VgG6xJvpr179yzAbbDFDHXTaRsq6EKPsLMsv2q/BHnVxF+6qt5kJ0OmAgK7f
IDNfpOJPutONz6T0exYAVs1hEQJ62aws3tRjkKxZhonJU/LKfv1x2aAo71RhANEr
XyoMzp17732w5f9TwR2rZld91ZHG4y0tphGAJbQZaaXQ7xjbxqqNtA5C5LQ1X9Hl
XTpuNf7SAEY04PIsPwJgTk2w4WlDk2+kjJhUStH7koGd+gcgFfPuQ5+lc9wqPkLp
vFVLzIKKYDHe8xHX6spsQVQqdHBsnzEDw7jBkwt7l5K+Ue/LFFhQwOKtR0bKA/er
o+W5YmWwJa+q2fThJfanK7ECUlprzB2cLzAYaWJ1+8y50vBFVdiHw3hgGX2wFXhZ
uE+qY+znK888bmzMpIO3zOt7/t8nA/01x51rIiXif7eyeevzdHeBLPjZxGZ1E8s6
/gqESeZKVKB0yIONwVO4cqeT8jFsajqim2vIO7Bxu66XQaPILBQG3+O+kdVLd6lW
u5lBBv5n6AzP+fgpDZlf8vBm7L5kML0guXFZsHgUvcW05B5M1+yI1+KIpbNGV4rr
pp+I/CKqs3VCj3oQ5kD5/jnT9+vTD6jg3mvlczNFnqp7tPu8HIV0dpVqyZXGz05D
lpRX4UByFZpd0MvK3dsUolMFPScvZPYz6ngblrxeme9IT28SZL2A3HTCMizAv6Kq
0mKbcFydOEjaucGCEXGwO33QV/txzBsQx9p+ueF0ucHGXhj+hkif+1smjjVK2e+N
BMiSfuSKZLvwzttnjzSBtuiPJxIjq5/M5fq1/4t9hhSqr3r0i0zPvG+kDUFCo3FB
DH80+K+M5InEUFwO1bs0DnWHnZmg8TsNonO6tAN/YC83HqQallk67Vh0C7wajDfy
TWtXrB0af0x9WCVvaNeVs9zecudM3+fnx+n47qP4AqX5wMKZKtpnvLhTdFIahqKF
Ask0O2Af/09G+SpTOR3i2Zcq50WT7JFR3I2sWf/DCmBHEmU0fkCZU6T9XZCH4BEW
BE1OK3Th+FIHq+ns4+UMYNcM35jt1PVdzEyWfk4X5HD4KWxTvt1XNqX2SMOCQA4h
hrOgyKWZjXLQIy85G0xdSYZoewhziTe2xzowwm8d2pyf8kRogZOfjamXFG17CzMi
UYEZOqXKSZwC4J9ZI2P1WdhS6iq9OvtSYmtN+4JfJRrPUnqCiIwriQZDOgcIPyV9
cRUH8HJfQ4xqm4jlyBmz0khrCqzmuCukElJeWPZILVEVubRzpFoqHFBiU23YHVLv
+BcRpsRN0u3zl+6O4Uk0/xUGF2uzvAds0Cv8oC+GflcVZWtK56HAc5MbOdNxlC12
RZYKjDH9tWjRPFY2qBfqMr7dugBW3aet8xUDvQ+iPbccLkuvhVv17MMqAF8NbXhs
6sUk37joUIoY3QuvycHy/oWrteLGwMXAWA4vTc1eCCrNS9ufztxuvaSH3U7HyPUw
LqTVwpnHi4UjCVAUB/GdIYZiC4bR2H9CVYfmjjYK6fP8iUptOAIBWde1WyPsVegB
zdi0Y/CpyA1ATQRswHUIxxUXF9s1qew1bFrVrwUlt/GyG3bhYM7/yxpGoBn/ogBM
Tf/ka/9LJ6GiSFepHThUKe7VQdcdNRlHaYjeOHoTslUXPJKizSHo7BURGFPH7A+h
fZyDosg3odAOOSTkmfYBVbV/LpeJCNmRf7SkQCEYcA/jmo8DWGsTbgrFuAi7PzI7
YOgS1JhJy8u9RK1ZAlVxftIAZcmb1vRfegzf42/1yQjuQaLPab6F8Tx05ZxH6ZQC
lakMLkar/aJ1I0rOWwh4u2SAKxIJ+EYQDBuZAqJfKqxyBHIhp1sdUZd2mv0i0IaF
ea3qZ6QabPWKC/X7KNp7eP+voL4aPLOR4ykP39CWHsndJIGzgFKWn1BcvJHiYJCx
m7Rl2T5NEB4/quT8q9hMQF/RtQkdsTYQYjfnsmNScD+b0txmiqMNCT3GJwyvtQli
xOizbLNkWMh2QSBo4eqvZCvVHUlVNnv8GU77ybTV3Cfghg/XzqkpwUZjJafg0kCH
zlrd5zeDnzioCty0BsLzpEj24VVE2bZA4gcnAFzP23rXhzzKG0hlRKJfvSH5Vb/D
tlDc/AkX7p5Zau0Y7g+3y/6jJfXdrUy6iJakKKiGxSMZXrqEOB41LM63um6qGJw4
eR48cGzByyB3/AOkbYyV395YUDzRJlHCYclNdsvNjTBSB8zQ1Y0HPSGJbbXVMq/u
YersK+ejpHYCrjpR2NqKfwHZf+vA++gEcVApTLj0cwTnEsCm0/mcyJuAphJZ1PAK
cP71okktRLgun5vas089owekd6QRWSGoEek/zQ1mzpnwQiPEfe1mHNe08SdhebiI
CCMwmua8HPedB8ezLkatt1oQ0Lx30MJwp5Aaed8DNBoJEL/YElI0hR/rnYDiijGc
bmyit+eE/1xNPkdvBo/s1WudXBz6GN9lZy6ovMg1JPxEYCEmDaMl7mQbUnXNjUOf
Hf9/s4iSgzoCMYyoFR+FznubOVc1UMbCxKYkew4/ZomYvZlJlnOwjIpdp0ttZ57U
uNngVTswGX/HLkYbKv8RTPqr3Q4qRuLqt6dMYsPWmNepk+pPG/f6L7DLY8doRHNK
IeFuZB6nllp3exd9I1BkdqDzBsejbKFQFLr7zOQRwLJCNxnaB5cXsTLWtSJ/YOkU
nNWynsAbPBMOV3awJ8bE9L8eo6igG7CKKgRdXn74nV1cceIu9Z43KY6ZAkl3lfgy
vBQZpZdn+mzdSMkhwUV+EVemWO2U22piCuhGYoP6yUqXWmOnW20uNf1Pygt0Fkh1
XHTqawySmTYrz1Pmn4Ot8mpdiDrNSVwBCdC6djYxVk+WTPxqWVIMVjMoLTns+5b2
BhR5LExvtGuImSdlZxH9Ywcwb6H6gvWzRDtxTPxWi5bSyQZKRlAoeavil8t/JiXq
pJIBD0/Sc2FxVBGggY9c5XjghK7JNaeh55b/3oG0PUDcVBXqzsE7s/VIcHOQx+cL
HE4IXyzBexVfDEYEMbony/td8GWE6uJ6yVjJv8EO6+AkYiCiMs7QZ8+L0LWqMM3d
uqWDsN8+SmkGlOOgJ8WP/aDo5ornTbL3YPjlEXf6PAvKjMbd2JfG2T0hfyGGf55B
Nz/ERSYt3KKz7Se487jXwc1UQGWNFAII/cd0HOdxXiJ/zsuSHRBwRSmuvC+wg2oF
jdFOmIpAcF19anCWCOfOSm3CvXK/BKJmcfdBZAbJIjmnsIkE3PpsrZXMAR0vgkFf
O59g6OT7DlWiKiZyQsApor55mIeJhhvu85TBV1GOvznj6zsn2FlNlQGB/XSRbYxy
NohRB+S0xcCPcwfjeSQ41HxC209oqTaMrHFqhO4xygFFbAeraw2S23O2L8JHOe4N
rKQnm62x2ysZjCoOHN4OBr3Kz6mS9a6rmiY47YKCcLt+0r/A8Wzne/rbnivb7IRD
yOWhRpi8ELwE/F67x4MFkfQ3RiRVnq9SFWKZ/eQ79AA9G5Cbnc+2BSwjaGWMp/Me
ylb0RSmNK2z9BQangVGxgPzwc1m2RDZQwcgUMQNEazGyeBwGnssx8eVEdxHzF3p3
xUG7H9HrY/RQm/Uie+G4jJO689Z8pkmowDAZ+7J3+J46S4RTWVj3cjGgpMPdZpuz
Pf308I9K8AFLTGS8BTwP6VIsPkTc+N6gO+O1kx9OaPSGzijmYD33p82x2bH6DhL3
nRpWtn7Lp9PxvmD7+klRwaiCkWSOqEulnYXFhvQNtwjfp7bB1xOhPzjDOjnx6ErJ
pfCinuPecloPHgqdJngXi3SSY8oJ1Vk9wnobay74rnQXkGGeI8c/e5TnnaBrVE2z
6fAm1Qr7/nOtNC0Nr+ym95eCbruNDuX5NTjCVwmpVAIUnqykr7cEDzvNj2zhJhiM
E6fGGYA0O/SWIjo7ZTmFp2XYUzSe/my06xFSYjQHOx94oCMTFKV4kxFcS+YWSQ0s
kUfPWEc7fSU9KuvED+pRI60nPn6MjntSRrkIQgk/0/AwvK8VZ4fSxS3wY4NZdfAn
LXz9RUxFmixTXnKsFDeSXhWwdDv7ARTLSsP0xAURARlc/Ndt8CVs3mB9mifTcikF
3F2+G7CtlUjHEUfL/WeyDPYlZgWv/e08m+P1nV7JxXisQgZJhCjwx9laPXR6EkB2
BDp6RS5/eMiXoVKqFqd+YS+9L+oY/AtsBtiXAyeqocUDQUeMnAYgCmP19hWQBkAz
REkDWeX93bQBfBlQBW4XDNBCj2VkpR0xUbmY1t1uBFtJeL9VQeSmClvFZ6Ji7bIE
OycOmfxo0L8YoaJOFUkWpKs3lvz5XJzocyCRcf+Opz/I0eEnLvmYkCaHlR6xm2hR
7NKYU1BGzyF3kMgJrwRkEUbwgpXmHCRt3NNr00YE+SV+FHMHyO9McY1A+IYjXTYQ
KDm9XI+nJ6h2SxhfFs8+7QvlQ47HA05N4GwNDT9Utge5umxfz0336WDuk8PatHuY
B5wiMM43zdTVmZnhKzv1zZt+Hv/Z/rwOUvkoUIbRAq2Ba06tyCicKK6wtlLCyO7v
3Zs6Fa7po/CH/km91Q1cqjMFSm1du1rYZIEIfa2tkNsC2s4gVTyMjVkMq58k/dRo
zBzO1341H+lr1MCw5YNXHtzkn1svJo/nthgkpPCvBX/wjmp+3pjiThH4Oz3s5qn1
fTGsOe0VT+9xcZm1Tj9+Ff1sVW3q9C18q9B8PaQ6O+Z4UYubuE8OE7zMUO9YSpGn
qgo3HRgbpGgUYT5VugkvsbavXIX3aczys5BhEg5l+KDePGYSlDwGtO5elRgXaSRC
D3hHr42YY6OEblqqOBiAyj4EGXAbIdZSWCCDg+c9jtYvJmikk/DuN8u3scAmYpaI
PhbmifDOzbUhX/FVELy5Md+/THdMn9RFjgcXNZRvBv7Sto5VgLoBqNdGD0ciUcjX
CUx/wsxC5JAScJrB+AYYyoCftTPiAuaNV7DZuXMxlILuRCLAM3/4nfGLnYBZgT1D
es+ibTiC0iyCv2oRUYKeLhsooRmZNAhcAnqVFH5ul2gXI2RVAXVCLh56aaIeA29y
aHun5VbQYDCpiGGhjHID398whBEL318NAmgLW18yQEwah7bKU2nh1Eo5P/5GTtqM
lxasdZoIff4P3BIhHtV+DbnOsJCxCz8dpd1BLWpvAGqrk8hD11X37VQTSvqbBazJ
ElH2mIUbdtIzIjewg5iZRIeRAMEWbkRMJZ9T+CYdSyHcvAlIKWr0QRzBp2DVtpgc
kw/6ZYu5FRTEXUAqUpKMTYk/Q11LvxWa3aZw4lW/dNIJrz76r7XnP84JHTq5K1ud
kJoCxHxyQUjfU7J/H2rcBuPRFfbN792B07FtjzZwQe+vt+pyecBftyE3QqNwfpYm
WvxsUYVfTdqUl3l5MGtiM/AV2R8IK13KF99UOLuGZ9uRiqwjxTU0v2WBQbooOdG7
O9P8VLs6IOeTWS2ZZWgR9mdMVdIR4lcxLeCDVk5mN6xrPZOZyNLwQoNXB2WesJ/O
JDZf9hc9V+JYSYYTYYUdIoaY1MZU9k+Ia4VsD03tuD0Y834gg4rMgKY4axYutJ73
8QjWbYjkisGaawUK84Dmklav+JW/kmd5PzGK2EeCJNgGExJkUT6Bz6TQl7Mtf6B6
EVI+NldKLLSTC0quuYpwx50KSpMi4scpSveybccZbmzQAtPZUO0kXjTdIHvrsGW9
xZskW+N10XaLUNYVEUYGabEF7NXolx9z6eJudwnvuY6xCuXb4dPVwHkmsvJCf65u
/Z9WFNOg8CNN17mhEKzNdnrNKMUIw89UKuwLI/MbfPvcZxVCBC35NlwoES39RpPw
e/wcjvl2TExMhgLw6zo21Nar1v+tizMHkJdQLugw19Wx7nUh4tOdciEPpjRfOMmR
lRrg8Ae39URBvk940npN2v8QtbJASXQ9dBDBIXEpG9UIH6/Esmhwl6bJV82sUeVx
AU5lUz3eq//M3NSbF4kpSyapHeFMTkaQ5WGzt2ObT4qGBvCHpIcfX+ZEWQ+HWRX7
mVyL+rbVhC36VlZ17jLuAWgQSnexBjVpiICMCmlJP4kvWs7jnoJvpNRsKL11A7SC
a/48tXjBrHyVIq3PzBaUff0TWKXM+3Kzcqjyoa68KHV9AbyCnMR2Fm+foZalCpPc
E9/NYqXiIIcZjMpq3BEF78ICLd9CaOCe3q1fHYU4U0UuWxVmX8PZ8MvvqN1DHNmL
50rSRz8s+jd9gp50uxkWvCRZpLtIeOFR9njGJGk+rRqquIEex6Yl1w1d3LDFFScb
6PYDtWLUymXef7kEk3f0sLWVmYY1Rmj/GuziPdjDeagtdKXEU+hYrnqnQ9JDRIgS
HNl094yQ4TBrKHGUVJ4rxuBKGXIbaYGWDhRTBzaaF7HURYtyliY2tNYPBigQdky2
e4KyvJnoOtipq50wioPTOleoM46XnLWIrXG+NeozxsVY/nMhI/DkIlTys3daOXgx
Lq1isoXIc4FSH4k9pLOBlJbsAK7hLzFRjyVPDIEe5dLTLFHu6Q7VywuzjwkLtLXt
NPzNEVLj0ThIFA2OqJfWkIjUVgBT6bw+0NDqE9BhtwbOCn7U3GdJWN6zQvmuNLK4
rf9AsRfvuSsxc84jkbRAsqGkCdaEqvX3RlGzhsD1+A4gU9Saaty78KgHRandI/ov
qn9AErM1vSBkFPQuoZArJTlBOldmxz81D4pgoqWNfkOW8VMXBxYQQezfEKGdNAMo
Rxz1Qqj/4lQPu1OT7ZZo+MJyy2445TllILnDIs1JyAoDZrmqAESxjX/f+Khb9aQy
y3p+6ivHwSu2ewFbkt5FHJFmlEPTD/2coQFU1h6u5p/A6hANJq+XjRjmGY0AWYXw
e2VDEd0YUbzIVQu2pabM5UluGOWo6OpkLnDni+Cm4DF8A9KxIlNWDQ+QK8nVuFQB
8cnDLQc2e712h+/3FtQyzfh2M7jDp/aEGuSwlJG8ggNU7lpzVZuYLZThzmHgJXF6
FWCH3F6Bds9fJxyfOU8Bp+BfL2hX98r4mOmgsVxnmQKWCCEWO7TE8XT085YvdToU
sKmcNf3JKRxdIGqF5ZYxJ2m/OQ7KCfHS47y4w/Mszj9RmVSpluw9jCAus6TObEf+
IQ95xG8GJ3X8YIHw9MwDPOLPE0XgxiFzZfiucboPKYUnVo+ykxnlCSRALRAoxcnK
N5x6aZga01wFt856moSy6to9C8kn+KYDZJE5Fcz/QOcN9qCQMKqb4uuGRMzfnVpH
n3YGuFn0gDXqGprTMa7IdfAmB/C9/X2Jv4fiIIfeEjVdemDCMjJ/Mlmd8sgcROaz
xvhx/ZQqBFGivHc8fu4x2h7rQGuDiOQc+lNjrpCbcklIyHdDv/4H5jxi3tYt/255
eiF2tzV7oEHt0UMfmbU1Opfixw6iKHQC65dGBn5nTIAhui/v9lUY+358oBzo06Tm
S2bXC1opGLzz+cKmt5EjxbSpCJzWCqbVkFKM/3TnaWZP2AxGjVyVYTsUGo37lV+k
s+t5YpJ8a6POCENjRk8QIaZ90x9GWFWMTSi/nLUUNRAwdS2FAGrQAvAcqA05ZyfM
hC0QcqrSNblZMINVBKWCTQJ3nrohzTTI4F8wOEoYW9Cu4HjTwD51bOOoZJegWYkx
tZ/AS9UxkAXib3/zH8yEEQIgIBmFRqW5nwPqY/Z5iH9e5PLpAGq0A7wj1OmGL5je
NJhAwF00rjLN7q6qmfMd0pQwE7i/Tk5+6wNpLsOdQ4VCmFiptIDZZpZH/j4CFn1f
TlO7CEdy5SDqeG4WOKMvnsESZ3rSQObuCBQwUs7KSdnBDnGACotbkfgYo7pSnWtA
Ak2G4zIvL6zoDmnfa+mp8RyVwyV3cqRU1tKjzW0mzCccET/fTEXRjFwOVNGH6xQv
5l6LtzbjmX2jqm56oCr4FfqGBF5XRJhOvwh0+c8qAqNJZ3bQ3K6qjECsLbPsYMoI
w/AEgFKqpPm+1Ja8x78bSpnEl8TftfgO27AgMw9uloWKwio/T/Wa3fGkdTP/+QGO
J23wC60xEgxGYRb6v63KEq3wetf0Z47M6wPHA3Mv21PGF1xuq6l6PGzOA5sMGO8l
mRt6nLILsgqBUV/eDfW4NBSe+4rBvX/02Pregt9GL6S29PoIFr+6opcwAYLd2D+c
msKqRq6jcpiCfQjUNeBBzTwASChL0k+hIkT55kcq6JhUP5KKe6a6YuU39cJb16Yb
bZRBXruwrDkZ5Q1bC5GJcvI7kSKhILvjyt+8eNQBCIOhW5ACVj0lvR3+3KhCiNxh
p6tra5w5lS/dognvu2TYEgrUaNtlz0ByK96/RK46bL05pe9SsbKppVI034I//2QA
zlcCsXU7LqIZnmK3nkZfAKYUMQJ64ADb6Oad6HK/DU1Gp8zOSHg1mAEI1q9QVCDT
40tOgVEjUs41qCjzR8Pk5NVEcgR0OgEUSQ1H9ePtssDNHBrjrAsQfgfLQHsNOIc2
Pz07d6+gzurmCjdnbOuRlev2serdF0KV0zw0s2aZMP9igoZ+nk0BPzdVwGNaRkat
1Br0Efsl1nDg4QUyJR+Kd23/AMG/JcMif1m66W42N0+wGVcEBGnxRUuuODTvjxb2
6Z5K9AqataweAZE63YNOhlJAYWCf0ZTBPLyALxVVvWGfhGJUk8U5a++vkbwDGNYu
tF6Jw+nPgFxpwvBnZufxOsLf0kKrrzFCJ5bEwqv5RXtpitzP4VW2aNLfhYKtrqTH
GUJEf+pcQn/RyKGrA0Ln25s2XgfWZeyVSdoYsrdXAe09PrgCPNZboYA40GlBDi/L
WYogDbx231/SWwptl53sXvEiP0TS73o7dhv1v06Nk6efpyj2TsQMRBHMAo2tRa6o
hPk5gUYZWf6vhzDHvUWG0RlhOgqO/97fp1k2BDeOtx1EzLPcHM2xcx94ffizzHuA
g2LxQpnY4lGA9Mb6XsfHg4gcmJbevqDVds7n6EpuOluy6AWGL4FJPpeaRm4fvsws
1WmJP+I1ZMt3knF0eti1gpYTvbJUcVGi7UrMQ94hFoaDTURkilFJIX0uURPTj96+
3Xyw0FOEByMIVa4BQJwTR2V2GYM1D1o+7akoi2PUQHxNbVwyp5hakdubG/yLpEpw
Gy+FIyXUP/9GAc8IoPRAI0uHUbXLZs68RsJKIMpP/8OGmBaYDEfCam4S2OlVmlp1
iAjSrGQbDcNoV0CM2BNbv+27e8L87cAJSNPXiNTpe9KV1pw59dWL6QCbZ0r7HukG
/g3GiT+liPp+j4rtchUHG6MEUMUtUVBJv00H00roUxdDezHyqqQGZ8yqlO8D2Npj
V+Tu5tdNFn1y9JEwlYsJOGUy+Nb5GxjMpCYX+ZgoOLjDPuR3dbL/Le4Jk878rz1K
Rj0zkLZx2ClbC/E3chHA9DQHpYX8yEQ24hsSs4U/aJM0AOoFfCFmz0h8fQ8sThfu
anmnodBi9l59JGSzvKX1I+RAAbqwI2Wtw3yfekdySoLui3+kD8Sb+YZxo+f2j/JN
5kfSgTJcVbWvaFQlA400jIS1IDBT68upsd7aLyqHsp8JIBz8xsgO/RJ76cQt61Oo
TBPkIA8ohk1JzT321Mz595K1/qCYvTh/4D9Q0BeYOc8YK+zpWt9vWerupLD2LqIl
0TN/nSPmB+jvVXGGDMAqiC/0ZSGKCw8LhrdZBoA3tfUPiCJwOruupDeDdNPNbz/A
fyzZItCGWnnyAsL3GpXTWZCaujxLFa9ZK0e1p+DmDVbA8FJIIGqzX4ofaXi1CY3r
Yyc75gpS2aQ0aQ17wpfcLzFwfsaUVWdXEa3giW3EC3ZNF/KDZyGn1NiwOxH9HO+b
/9v4618oUyj53S0qRQNhoI8HM6Rz+CCAR9PQpJBeX5fKq4asSCgicOLqeYl4iDU1
+RYD1YVjRp/LBlRc7a6OqDz1k3jekTH1z/A9Evf9wYggP8wsukpV0SLMIan7+ikq
Ma62qgUi46018KgxKEmI4jabrsAdk/lF3jNuIX5oI/SYOWZA4JMOqQrsdbG4uO6u
cyJSRnwV2Zo02qcOl7eSyC2PXBoV2EfoszkWYViLrFF937y5eL84d+3+nIejlDB9
KvhHtRc0NYJ0gAmG5ZJNxL5RiQTgoo38Areb0LA6ZGYvP4HayTNM+ItxZD80s879
4d2UrpMCqVFSePAhKj6jMi6rBmHvnbr/yO7FIVfigcoMe9nrmkLlXc96sQflS2hY
BFVG3Bg7LJGWK8BSPg5gn5Ilu+BZUtzUFXxe/XgYC95vpilxPZVf2Ss0+UaX1xya
D8bZ+4qWB7ymcB9GsodkF7IyxSg7K+CeZbW/X4apMzf4nEe+zWjkTtUnSbw6WCl5
kSOEqjzyjY+5sDVWvNkomIS8hMP8SC23DM2pnCETkga1OUda+MQS6Z1w1Aj9FIWh
WzaRu+ihboq1Ho7rpTEXshaEMy8ka8666KWcIxhxsQV9o5fFFr+8F2WGCBxy3Nox
lLJV/jiCJyPkMFt0q4u/xO9x1zGZA0OXkY37MxPs6V55RDW+Im2Gt3NfEbUtG0az
AkflTlZSkeL3eaaLeEd6b3yVQOBjKAzCMNku3IMaIJVcSc0gg2u4+8MVTs35aqhG
zdGS8Uqp4PsGaTZaA1qzxzRMpK5ymVz33KtXHak9yKBgKNUko6zw4Q6J0NndmDUD
qkLh4ulVUsdp2grmBkoNhwGs46hh1ojqFNQyrvM19SlIhv7rMnEewybMAsNplBcT
jmW9KcOcZnMRYiOuPT/2E7HmR5skqZNrXKNfCNoAZtYgOuJ1+NwsrzAG4WvIvCUV
m3tYiHXUl48l1smYFlHwGOccPBo4GJLOUOZtJ2xYDlJMKb5M/lQg/YEOahQf4guF
1BFVdLVghOe9RsWk2IZjbjBGnXa7NFV0yZLffDvgHgNFvZ7TeINw/05sWjhChbEP
WVg+rRGdrNKedEdXhWNa9kK6cRVSXZWLU/BdyLcktPPmDYmUjPLM11L7aA355nVE
cknQHjTNhgJk/OZjnWgbRiCyLY9DcvIQJ9I1Vi7nQqQNH+qqI1isfrO2lkiwPnSV
sFF/imdH/QJoIOQ+K2lr1zSJk1GMb9VDUxQEKFjSiDZ4YCDaZdaKqSyWKDGMVyTK
xtpB+E27rf0RWfeKFJzbxRhOfCFTDtmGz7z1LmqDed8hnqsSLUvM5BubtM6SMxQo
L0MYqSrSvvgT4rtg6lIYdTBkL+FJ2r/f+JXCMQGq7Yi1Nc1fME2rYzlMLd0Qapoa
qwkD3uDJFKVSsWNP/1FK1iS+bZCq+HvF6tdMFQJMQTJhkXYsyLVn27/6Vz0eYDtL
g0qxGczv0bXBBuVLKf1NbXOLXH4rxYqZV/qyjqw+ClC6jIV63tzdg1KbH0YjWP74
j7DYs1jsCFBcKc99+fCY9P84ocEMm9dsw9TcMn3KCUYm4wu3mj0/7HAZxhAgd3BH
6v7tSE7fH+RVHzAj+AQV9TogXmfksQdNtcHSpuySR0BWbChaVVuDHGm1irRcnqk9
JPDa3/nAVJZDFbf2s9ARgghoaUfr1Y1/vUcBPCwqvVm9HIstK0Vs0aZmwcodBhxr
TzDDdidO98i53PkLT+wD/ShPBeFZHhljYBn+7lrDALPXxT26NV3EefF0g1n8rWfW
EnGgXdtVzGmLJJv8Csvu36heLGTjxu9KKiEyakT1cfcUahdCIfi0SrDc2I+YXJ5h
s3rFgZJx55xoSSKmQfvvrr0ny1cjM+k3KSaAxYSu8uzIFPbmZlcJ1qrH8GCPzSRr
xK3LxmbBPj84sCX48u2Qpq87C1NW0hDik0hNIyiaJNX+RCeI0q7GidsdKUdumkcA
/pt3ClpYG1qzT+J5SeKV7AeYa6c9+aNdEuoLRVopMCHv9g7wljIR+iiRGvZPpD35
wC55/dWtydxBntLRKYyjlpT46eqazYUlQ1sDGT9KX1T14gZJzNR/zPPmP3ayy2Zg
uG5tgrMTV1YSx+QTT7rol8urZN6PqyHzuAtb3m/A58KUe3H7BO9707voYjTFfgwJ
DMvUfSXFIdOXs715/NRXfxzi6gtCsiclsslTJowoswFyExxoqoJbINHyambhvl/E
XNgWuvIfa/PjS6FHJke6IxKpVYZnl4A7C1QiR1K35dubELasiRdQQG+gtq+V8DOI
zYR+eCU+DpnmjSk3ZIfu6TPneI11TnT9Q2t53FsX8mG8k4e6TiYAtZOLX4BXW5cQ
BFXjzRuw1ohC8zJ5sqRfPcvTo4AjKqa1qFLOSfsPf4cX2ObCAEXHgm0PREKdMkHF
srhgbcq0dHzjsafOO0kpxsVXV2Wb9b/0dGV5bgfxHRK4TimVZfCLdbEM3hrM8Vpd
s32vFVBv0UF4XjVVuMAnzBPtFhd/aSfEh7M2y/dTO127L45uQHnfHMz8NJ13kBAL
2ynBrvue1d8VEJol6BbPUFFZUAaa6OgdUNet1xNlQ2Reme9V/Ys+5XG7aLojonJ7
z7AhkFVKSWL2QUGBuK1FN1YU8i0zPndfghqLChOxw4rK0gjA3jK/qtafyVBYKw8f
NINiybLAgFgimCtBBTwkQan+5P6cDhsoVSWiSft7ZMe/ChY8+DgG/msAYf0JSU72
OHybVv+cGPj9uHnnrhzM/XygYa5IBrRvzbnwjsahj4oTY9EPGbT7FzHtYF/SzRHr
km6utT2+YtYWPMeJaLIi6t2P63tiBYkLxdhw/yVhtAtIjomELYjy+7y4dawj2TuO
vIR7pujRciFivgosmK/KCQVtAasePuQAOpFCWKRpqR1MmMMO2beATJo7Ddpf7qTD
E2dMmXclNZIm4c4hdNFQ/MUhlf3N9g7IUswsAv05soxjQxbNNtq0Wx0vSJE/KL4A
UuK+JvUerUIPhX1PjRdwG2G2z7C93PYdhTM4PL4mWLpPT4f7xggEJmZjeTYkkNOh
fl4Sj+jzrVA+E3HlOdbGZyxMhXRtYs8SV/y9JhQo6N8vN3nQQh6/0/z5CTFbEki/
PeIx1pc9AqbMIxCBS5myGXItqXXhW7Ctsn2tg0OfNtp8uB9qKzYfFQQ2HrOWRYy5
VX5yhBFS7NwewSm9BIkccrngvqPg+AZ2f/9O7Psr86YbykWkGLATmkI9DJ3VMhgV
puPHhZ5CJD96z6HP4d6KhZqPuTrPtr72bMzKu3LiQ0kKDHCuYKfRx2y8WYDUv3NM
UXFEoxjdresLbipHIMF1mHSZ9i6ABFMQrOnW6L0ItffZjbeaygjyimu/2/dQMU2M
fSJWQj8yRtLgx2v8E2AywTx6de7nkYe0/nhaNRSvj/SK0N9ZTTBU032iLA/UTafa
aQ1qxiA1IdzkwWQMmSo+RbJ0fBrPGIZ1D5RNfO+Cin0yAst3NiY1Gn36QQ72+Mkx
AcqjSTW8vZBU3m5tqcJwWE8NAsGKlSOoIVwzSWPy98O+vx7LdPkk+A+xLPyT1JNQ
9EHhisAXDrVkAwNPRzptPLy6BahYXo0eznxlJrfHIVTrOTDCYVBu6n7I3NcfKmW2
chTgWDC/iBASIx0kr7FSvI5DN9w90dqgl1XHfmJBPzbWyb6Df8RN/8U4WDQDGF39
vUsA3GC4QhjrWR3TUIt0rVmCZOJ9JSbiUUfujZVuDmAeaUMuaaRvwKbHgP5QpXE6
OBk+JSrWLHrZFCbroVqjatT5at8MNrtqmcJTRm/2cGWmAvYvaUT05XdbATq4ifyX
TA6intpkUYs3y9Hkc8xf2ynpNe+AMbFYOq7yeZ/7NqfEtuyygP2SiWcw6JhDPnXQ
djEuBdRG9yHtjNZtvGJaE/oyW6E0jPzW+Bs+sNrUoARbA+3MhU6MkiejCwvWXtRR
IKkLX+2XxIenvKzW2+ERemnxetuVXJjw1VlpV/hH40ZuwvvA9503CWUuE73I2vZP
PNMoWw4/UArqGpjGT0y8McYa0XQL1XckTx1dRIujw1sMI3Z8NB0R6yE4YlgAiS3K
PL1M+SD8+EgX04jI17+DUyzDlVRRHE6znO0JA1rnjPnBLAVZHGvPBKxu+kuaKk3K
a0pfi1/TL3qHL7MCmcjPHyHqdOga1rPWw3ArMP2aGwAZy9tzqGZ5fgDR1wQ+tGUv
QR1ov7IzwZO6ydi5/p44liGXaI2GUH5Q0zKW7DV3Ieol4klNE2DQZS+NK096AhuX
eqwZp3Fl3FVaxib0IkyHCwMeeQT4cGpzV5KcImBd/K0rVlgp2ppCljKZkJheEyW7
7UcnCVr9uPZFwt8KCCVLX+J037MC8j2zOWVxvS7/tDYiOVDCVU1mvHBEHB2vn4xx
nhIZMMQyUXtJl9SLb81hq0TqA0fyf9iqzEZxMIA0gw/ZxcUl1tZVWdI89RDrpT8P
xkUmkchQ493BoCofyAzRcrl+ftK7cXTXF/S2dBEnax3MeGFBOFjBgs8nAPP/Izhr
qszAIqTZaJjeHlFIfYlwOp3CUahfUIj/9MlfPPtOF0dn9aYuZvMWF+9bmEayF394
kAIvwJsZxgN/EwGoZbS+eLUZM4+9KKP8/TOk7rjLGoU9Zax7nhIyjSn7TOgv2JrR
642CsM/MCICc3i7R7KJEV8bJnIWIDXTGL+/177IGqPYgp2vf7vIRrPVgiYp09IwI
wiQ9bNA/i2HHslyA6brVm4ow+8awYHPPSO1TEYBefvUUNrbAfC1bqP+VawCuI0ix
TStzjuxUR2JsKbt9b3V0DKT+iRPIAWT7h0eB0LMGcY27pLr9IxFcAF9VpOBbYath
BokdAEMdLKfJSj5/qDiUFkjsqHasO+NJ3UfeNjfUOseS27h2vl8ZOxRysTylIsJQ
Tgv9tdaFoUv5SXXFoE9Wj6eeYJlFjF+lvYjowuWsbZiqIqpSvmnajji5FqBxByQ3
mMTBdwplyajhPAzxrRV8lXqDsWipHfBUOjtezvao928Jsfx1gX0gC7IaIlNpRspD
m/kjjk2WQ6SjagVR2xh6XXh/fVxHZ9P7M7fe8jJoXcK5uw0i2JJzHBh/WC3hHNyj
pT7vxoYGH6QNLZ0VSSEfPXfaSmSeykVNWzFe5bOQgP3ZJFo4tahJJu8FA+p18FWZ
AerRQdGxFq0QZTT73wzDtHQJMBLxi0HPwYBy9XYUPRssmLtTthXwMzEyTmdsStmd
plyrTVNAXASU+iXmoFN/qDLmwLiNEa1NVm4G2lObLdcxlu8ioVqo3sHaZeIsty7Q
gKwhplAQ1b4P/NpsxrtOtZ1kohM9WvdS0ewrbD3N7pWzoXV+F1wsXVE3oCIVApVg
8VnlMIjMlmbEtDb9Pr3pJ7UlpT2rPh+YidiU0OjchLB2Np7NIIU7gs4/GbvFefJv
YPk2rO/w5MUOujeYP7ExTqoDfUgKRtrQGwWn2qbrpfR40VQyMAvDeg0nyui/1qEk
I7BOLXruzpRW6Jx/MjdYK1uD7AjzTcGhhsxVUWfGS8eOG4h1pve2BXoToA40g63o
R4z1r87sPed8i8bbSiO3/AQdOu4KXdybmltXbDAUo0r4u8umIesu6rPKjjNbGbyk
V7zAdlHLELir2MBiw9YlGa6lAmYoKTFk5pc/XKun+VZceqantXqBVdl+JUcMlwDW
dc52sF339fC6G+Du0MApQJ6wwyu0zImVnP1eCR7NUgGfOOnobIdnQz98JwmJ4eqQ
GMJ36qRud86wEC5JHvPoIGue1o9IgBcEtnBHDiXXuEcCHpoGUrEWn0FWtCAKDV0/
/rMdmGca0Q60b94mgyQkO4DKxdAvy0r8UcH90wyiOG0n4kabjj5zF+dNpplIJhii
UwnCmxdOsVbGbnqPoFyVMrG4DSR3Or2CIAhlHqqx2QyeK2kPM2dNQh+HRfiYfKAE
z9O4BT9IvqhURkLQPziuxiK3pxvjd62+dRJWGOPJupaLDH2u9OPKfK9u72zeQPVx
9pJ+JwTJcxAt9CCWzqPZyphyTRr5n0J09FxxpnApJ5d9tFVO2wrR0x1dcPE5GGDp
tbXsJD+MXycsYDjuiy+GiN61By2a4YKQTRpA2V4b1Ird9G5TU1U9lEdaw3SrCNVF
1LQtz3dzsr7Xx9hQNM4ZGOGBXiUm1taZkfVpdo77g1GcXygjUvWnnYSWdHVlfmVh
Jw8h5q3tsEDJa0pDjGxclRsQ17IYz98+88NRtSqed6pmbOPvyfNAbOITLFJQtTIf
O6dqRbWcnbN3+TvTqNiRjQi6lYIiW8ITunnpf3UbPkc+MRi+saRi3Mo6FB21oOnZ
fp8HDMMECo3jWEW5NhW+WWJTsfru7UwxWKmDHUmrLGODi31puxEGbjcdPKJO8eiW
h0IIptl0CRSRDoQKGAeMn566Bocn+zKFm71WrAeK5Y1KfDyEZyunOiBtV6ilAWgU
unSA8nWMMdNu1fWgynIe3wyJNrNJdNWsdG+3cXk3KemajQENYiXWOw8PZzvXBUKS
Tq5xXvjJlAFpiVFC6OW6NX7HRxSCeaGFg5MTToQZ7fXA5pNhW9JrRZSdLZMEFelc
LWgdtr76quQ+fNhAM33S+/1UGrm5xJhCS2S7kBlHh6WXlejqfakOrn7RBF2ZbmLp
Xm9RTg1s5YEh/zx/CbbVyYYaHLNPx4BmsagZH0nAOzXzgATS7B2NB+l7U6hdyHta
JUrwzZDaPuIrOdMZDw7Lqd2wqrTUg1UY7/PkTenS2GQID4JBYZfBM6uIFqLo8eia
xHIkKhvw4TjKaTQBegp9q+YnEvkPF1EvjEuWuEe06dua7fy8aK1lJIEKRoS9F2qg
n+S/mI6H/CpSubkCoMA2UMjklfh+rHWG2KtRnbOP4hEwmyNoV3LjcPIkQGZhrEBy
PQYS8Zvr0/EeE091q7qjQf+ka0yjiF8vkgksQZla9MHv++ouMA43Jm6kPwMhpDri
fwjCWKoCaAtnDdcRCgsPCQCCDCI+jTfiVmcTBKpQxjxcieMSpBthmr4TgDkogPKT
k6GvVr8NoGaE1UDZlKT+Z35NGof8SJX3W11CoVuqkjRDh6i2PSn53OL8KAWOEGG8
ATILj/md2s4jAcFekxmOnnc/KBX2g/5tveA+U6euzw9H9dI9IfsKdJX3NtKfG8Xx
0pTfX5ITXrgGB+fI/8/KiYgw8VfQbnEqYH0GCeISK/4nzUcgLUU9VfCMmy++AdB4
aP4dFbPyoULglYsKiecJswYSWdX/V03Unutw20reHijlVA1HeKSrTQSFldfDbJ/L
LOr9rEzv3r+mf1a2InQYuqxfPaGynhLJ06eRoCrrqWfmTEICm1nLcFlJwCWD1OOT
3b27BJ9TYgBgBy/NWTYdRuZlWOnsZ8acvXEx9Yc4SDexEfPMCV+oIMipLoUPWObX
77shLd8TH+6oY9B6K+ioZ+RVtmh7ll53+KRjmvNxOM7/98aByG2bzLfa8vkR739e
m/oczfVTmPb8XgUXyeAH14WCGNcsuS+yzovfijJ71QzZ442SnQWJ6j2Se/oE5zUD
BjHxIPmxEauoMs1lqVGPMbl2JC5QD4CRhfvLIJY8cxR1DBu5AjYX5QvsnBLs+vDo
Z+kRwzsAAGUoMkgLZelP91ykciIIK0aE5jqFWTX6ytxZRfMRY/OJVSeuFeKNvoN+
DZ9JsjujUydSymdEwXLZnV/VoKyVTFbwDQgMzylLH0XNUS6YQJVewbDsZ2ZyaTSe
VuOGFjGtONqQb3jL2wO0lOAkPAb8R+furdfw7ccpfvrtc/8Wey+D37lIKQAug6xz
tst/lO/WWglxo26LXS9noFBky6cjUSe0wfGst5RXDcvhh370vzjnwXQATOJWNBUw
HESZhnFXxQRdHKikX4uwNs2EK/UmpoteMM/RtUykuwTJTUWtOb04SUFZ7n/2N7HW
GVgpoOS1xOhTwGZfpzZ7DYol9jl3jwK5f00+u14t2MlKQK8Ig1oppGL9lMMohRhL
rn0gYUD7+VNSswdsbhUjhZNpBc5YTLrmvBRxZe8N7YaMDFX0LwLHVNh9TMtkXNC+
vaPTdHtF983kx71Iaxr/pWwmqhyk6n4iALHw/7R5mNjtCMxl/aaPM/4EksIHMrxa
JuIfL70fnJxkW3PgTJrgeNHP7g2mEPEwy5g7WysCfn0TGint6+Qe3lZvx1cnw5K2
+gvsJoKTPv2VrPIK4EFKLfdXzCzf+3/Bq7dTb7IziM3kIhXRYGOQEINXcmeM5rQI
luEKi88/xKxhFeas755m/2JbSMaOtZBV38H4ucFeKX0LxrcVYUTLjqOESWv+zn69
9SSx+O+/FBBvgS5esii5p088DX3pfyy89vP1Vi23CLPm+UxhSN9uIBTqcW/opX9j
I/YkQ8TRU8K4+65/kjkBLa07dpztQOHQTzNRIMQ1QA5kc05EToj4mhF1ZiD//g3m
I/UFvn/iAdbnUdHd/0XpwdY11zXD6Fo+hkUuwJ3jO0vJC6wfANDHmMI60oykspDT
RapRQq93eIDNgeSz4y7yQb+X+5fz2znsZae1ZW7tF1oSLHtxPlolrQN25FO20uTr
+IlW5dm236tDDdSh10XZ9/i9jiQrygi65YqyTHYMskTXN6/iSMO8ZzzFq8UfB8u3
GJFVUDZFn+1AB6tkhhiM5jR/WChncpzq/FaK+D2OC+dImHTXuXrqannH9WZyoSTk
g+Xga2I4Q3RJWkvQ7ifP/I0Y0r31/AuPr+AY4SJuL4Fz4XfUWP9EchT3j4XlKRGI
WAzdSWd0rHkHFATYeSP1RTxKyG3oLGZBCS53k6Lsqxy/fPxoVj38hCjkMW1Ymi/x
6q8LGyeEbUXTSbevzTDEha0JwPhyhImK6bpLOP8mIZQswju9/t7GuJp1+XZRo6LU
/wzLgThJO9R6Lra3zObgJ9Rpd2UpxOM4/jWylt8FrBckZ9BEk4m5DEv+DQzwnyKe
U03ZEiFdvOIFb+uvu6DoFapmL8GRcdOstDH+RaS/wnloSryeoPtmPl7NhxcKSeAZ
fVvVMlk5+d9dpskyqNzBIp5jRckoHVv1Oci/FKOt55SKh4G7f5FdSdORvM0LDq2n
0vTbuczicplsZbVEMOJyJbANjHGZTpxXGXGADhV7HU5VEuU6OfHRVgZNz8e7d5y5
ebPd9eOTJ2GNlWedLtp6kUJbpY1jv4QYXyh2Jjpo/cMxWmlPTYm91jUYEjH/LBlD
XFkglZNi05kWzLhVc3wRtpL2nCo/HGzqfylDu8QQogAPKFbjtMEcu0KPG7EDADrw
wf18UAu7+CTIRy+vnSvkjvC2J3gT4gGJ9+8kv8jQVT4/xkkZzFv/ZIFUQhxL21Ti
wsvI50uCUvzu63kg78YDq/+NWbaQYj3yoruIicYok8aBOqofWD1Ix18OMFHqhLs7
cYxJsBdnphQPT6FkmSScSCABGha1gChVI4PZDs7wRWILE6QDNgaAQFfrqe73SHih
SmTbPplYzDLFuIKQHMeZMcHBWX1Kxz84jB9wQc0J0PstHctWcN530khTiMDo02YI
mydttTjdqc/I/FaoqEcoEwe66wtAfBinBulzVzL3zfHP/iGBV9OWjShIftqm6Z59
1Ned0YwyubNnK/s9sM1AOc/BUUk9xtQ5Gq5eAhJv5hPw4coMzeiaImiMyFxb7lV/
W41WppH+gNRzk3f1jAW7nGsy8TEFqcwsxqW3X3WUWR2xMKKrPntBawKMAuYnvrqQ
EweIIG9M3RvTM1ItqNgw4Dk29EG0tfeSNUVcj48CU643i3tpXGKyz7gyWHTiVCGm
RnmTXyHDj76PsFaW0frWehkNv+32OBhhvcH2p1CLG2N5o11Hux9Kt3/H75YAmXSi
H2GKDgJVjh8ohjV82CcLmlYG37h9KGnU9uefQz7oqXRFwEU0MV5FxvzUlFTKpz9N
Fk2r4de6nlRrlqkSDKt9iI+BeaWZ6wl9lyoYrE3ukpS1WNt78W2pNbohB0bbn+SE
crgPekxDjZnIQUsVY77kW0pcBbTN2IglIG8ecBDIbV2DaD8hvgTXdUeZAlp57a5Q
v8JFAqP5coPtJBtmx4WbeQKEEpC0b5BellOdsyHoMnSpyZ6P3NRZPWGud9pdHioD
IGQdgu00mxz8P/1vgvQICADYLaSLsO7Evl80CoL6qcmIlOXQLcHh5I9OZBC4wJ1q
VcbqJrx+D8LZIJK7cOT9xFhyjeqpc26/NxyGlgYKeMc27HM/Yh8nTIVktb9UABua
TQoOHVUEqU1PkbC2ZUxUfeJwulCMG4qFQyeM6/F1hqwmsmHkkMrcWtX6LnNEWnJa
2NMxOcYMKMNpmDDTZFAMU/2p+4jG5mG9ROQAk4iV1VVttaIx0NQP/8EcH9VfrpRQ
PkyR2tYFIp0d63nZjEcoKHsJEN7Zu+dR+69K1lLjWv1HfbWG2OimowZHRf9rtzsq
GvZAXVvn9CIOcw68s80QhckDuh95wSRTIBMN+/Hl3q/a8SctSCV6+qJlNOUe8wx5
zfFl1QK8ilrHZgAf4ii7yMztcKOhoGtTrAdrld/xgUdztq4oEQbah1i1/xZ66u5m
ZGxH4uJff0moRWi3v2PUSCrGvjAgFdgKeG82DfeRcreoo+PECwaHpQ6xeE53XdBX
Wb6eDZYbXdiqOMqq/hebiIlrot4Ih7FR9eYhJxhWN2YHhL9F1VdctJa7SJa2ekHe
jZ4RwHBlYaMhWLY5amPNkjwv1IKzGKbmNXqsZPs04xP5wgo9IOqO4QaW1LTj2fkQ
A9cJSnlEbc9wiiaAb6XNJbCSof6MIHjpoB7bblDz2Ji6uxx5abE3GhbKrxWrHxDK
aQD2P1Lia/nKeRHq/ag/nVmg13zanuxJQMR2TKoIK2WfSMyVAfaVdy+KIzTecG78
dv5iR4Oja1dzlrETFNdUUCDm+TPDwRez5/w3VoPMrn6XOmc9mlArHnrmXICaFqwf
D8VvExQF+D95xLeOM0Bosx5+pVBqqivpYwFnOG7AoFqixjOcoki/50dVeQ6TWwBC
rw75tfuR/J65G5hVKPSQXMsTOeQAr4sJHnY9SANNgEepNIkrexnG9m65Po/TytTE
eLYCLXPyxQ4yg+2dh4jEmdUvEFjMc6O92b6+EzdRnF7Rsl3UEyIiivLLG+my9xvO
t7LDGZG+6sgNe9GN1slt+vhPhdOo8m5iPyNak+uXbIzXN5z4eIvSKhvQs5Ixa55w
00QUD7Tf8OqPqwIpiMbh6sA5idICFN3odBAi4jMJm6JSksZpk8cGahUzjzfYrOm/
3GBjSs/7WlZ2+G6DI+XghBTE8gXG6VMgZleEzYiZOS6CvxyV8subyqgpkuiXUq2K
qzF8+GyNS/7Gl0FyJVJ/k6tK+3Fm7LD2cNYWJb5vF++LN//nKETD17GRpkYrDks6
S8hgjSsKz3L6pLBfLrtpf/naBRWoqHasRFPi3icAfutoGcakuIw98m+4F+vIf2/3
7LV81zxe2XPg3a26wPCTPx64EvLB12Co+/rIOJhZI6v3Y2FSPgAiNDEIKneMqWHT
P22BS9TeBSGI+CZbH/GV3SpBf2GYlFl381b2y2hW67oWSzfHWOzrOAuj7BZuvK3I
WtYftZknbtkmTut3hu0vjdvTiTdI1gZt663eDnWbVccoMVs/ZeyLNQGK3uxg5q5K
qcSRn+Bkemky8SHjzLk3CFX5Y5j+dfHahM3ECm/6iNdOap42c20Foy+25gJTh93g
Av7t8wYA4V6zPimAjjFyWZmnG7N/VqVY/0InnFKv0aZtCDGArsctAKv44BD0fGNg
jjahR+5wt2AqLabsA+U0JvnYMuPpy0w9goDZ+fKElEsQeZ57pt9w4y+DnkuBnrEf
mXzFkEdfnVNwRxacHibpvbEiW4moA7V8BvJiiuE/BnyvG3VOPP+ZrvmNWW2/juQd
Vq49kIncGiuR60Mf9D9RnppkuAdSZT/FU9+aN0FxYkX2HrVAsTGGdyEAQJ9MFJHs
lI14N7wv3lsnXsMthfao2waF/rrdyyn+BwL5eHYxjSNHIYBQUIz+ulcalDFZcvww
+HLuD4UTs6cnu00wfPgHJ2OgoQqquXBUASdHOa3lW6Vjz6brBYL2Okq06om8xDiq
osLv0xpjI/PddaHdJvs3T0fnEaPXtFgeCShJLaC5vgkrueY49KFFX69Hf/Upm8PY
AS9S5xDwLK2jUprsTD0qlMD+PohXtNAWmwSitbiE4wfKkxww7kkSI1XQLrgL/fDJ
SDs9bYiivtVq3prg5jjptzEbVjTImP/i4XCqJnZZn0f6BsfaukgGieMlHlwl3RUE
fZ7YDTLZT7yyeWCYcasGBEYPjSJhVg07onWNlRX1sxiB3cioIAiJKbMUfLG19NWy
sI75p1v2lWfDH4bKOzeDtLGYzm6k4Uq0bz0L/0NDFDGcAPe2q9NFEuRDxXIv3euX
fxf1Kw4IAiTnXR0ohaNfB5ekP8sOXr+S6dqTu1edpet/z6hiGOpJdRMVTf9fbABR
Z/ZutP5I2ucxjg+y42JpQDqaK8O9qFSm68BZq1n7MkjGPY9QI5tnH17g21B3RCCb
GGJLiSFfl2ag/OeUwwSXZmPym5eNDA/fbeDb5dYDhMcraHQc8YBl470755azr3dq
/WEEzcpKNflwr5bFhYZE49VznGveDMLCKEzH/NkyNg0zxz8B1C2TeayLlGJEd1pR
4eVD3r3qfT7hDBFhMl/4S7mC9hGduYBGzAPxngi9L0jlBMIWwjMCGf7+3kQhI0dO
IjGfd0GeuY03uUVdE5jAZcJLHdVbC/U4twlurcdVJutkzJhxC1+9xd9vCfDs39Ns
Gmpe51NEx+/OE7RtQdmIrd/QBNO0w9KUlKW8Q+nRGMSX118NzRs/EXCGpXddLuXq
kVcBSsKbdgRks38nnjY3bBB40+U9yKW2CWdPGkBA5A4yXrh8o274dzzTK5+RS5z5
73zEKiszyq8dOTx3l9dn2Yr8TfhJtyHxaXo/Dsqp1IZblDSq25HJlsPwZDZJEqod
g/SxlbR2cyU5vSsWjjaZmPclYFzJD7ef4ywalIy7jgA1x+IU9JR1kMPE3HflhlU3
NJxywM7ddY8b2NFxL9tATaY/pcOYnuoO94eOvWsj5b3yFZz9W9jDgKI/MwSspKRD
iaDNDCz2PHJjPbu6LVK4ekorgxzq7wd9ejbcatZurIYj2Wky4Dyk4uRK/g/XmKEg
tWvtCfVwTuFbr34fvsgjaycI/ZXiYNjTKjUFTZw9xCH1YAg2Pj/o+IsvZPDq3g3b
tF5f/6gfAr3hBXdq2QkfixV5CGt/GfMwMc2WXM3ilaHC794i49XJyG2G3VV1qhA4
9nb6rO9a53HKj9LXRGxFYpZ0CvzQ8Vd/qK3GMj1WeWnE3TrT4Z2HACvVprDViHd1
XkgbkuVB7TkOdnRhc5+thEG3hFYCBr8iwEoLPD61+q2oLf6XZA6sADb+R7Knj84m
4o3XwClAJafRnJdGSZ3EzatQzh9dhxZJkt55IUe26U0UrwlbpmfllRaPwGkRAzvN
oIt1cRJ5sGXqY+v6Yq2+fWu2sq0z3v1gJtToeahuYJJcNaHCWfvAraQ+J0F2oiNJ
UgyODwKFbcMF/LOxJTipqxfsh2UykiYX8UhlcKVWCcjGVMUAD0midbZZA0THgO4D
haloEPOnJgucm0u/VsuyH5oIGgHnYsrMw7sR+1nmMoXSVmG5TeL34N598uXitXPA
xqurbKF+aRFXnrwPP/Phnzzn5MvcFiKsZmUrutCKiag+uuymhMFCB2U195TKnFj5
FvsP5LQr5/UWSGcNwPsHND6TsDUTn1ujAhojjwwx3Dxvpif9d/KUAjPopeMn9+By
yMEFrPqiwURnTbHhn0FQSGzw/Q/aDpV2h2srHVeYDxifBOu/EnCVzedKSEAoA5ck
UNEd8xs09uBhZdAxk4J4OPu66ieqJUdhLMXb7TZOAoKbkyoQcCMUn9SjesTKKGju
1nUG90ljTGUFTV5RqJUNB6hFByWpd7AkUmRs/D7HeejxUCru6dJXISogfb1SWs9j
6oZwDpyqQLeXY+PtPR6Px7a1ebLswbwataEdiTWi70BVJVgcnruwLVaoN7rYiFCf
euulnv1u8dbt3kwQTIGd0UmNnQCqxlN3NNcSIrnV/3NUcKNX9C9MPq5/eBf8mnzb
h0A24IR+Nm4EyL7qyuDOBbxZ1HM/Om7q0MBhx4NF9+piM8JEkl/kM2TNkD5aTFRk
JWlwJ9t8pUKj2AnyQKwH/jwZPfhJIXMvlLxZThoGAYPOueNWIfOUPabOHcjqVrl5
G6OroyUwYIneVXotI1SlMZhxD+UGTIalrtCD1dp4l5f3p6+cRDqLRiNEwOg4Wy8L
TjWDUK8u48+AEC+sBm2Rn41F+Pqgw/fX4yPyY6eAeqhMOffApKxX0px+IeXU42pk
BYgZ0NKGYA5EgF8pssQXVm7gPjOZ2fQqZId1pYbUiv5gTacCqIWeT5wFPY1o45d0
92QOKFa9vnKZGs1Xb4tlwfvmy8zYrCkju93+MEf5mIMAZmj7+MEMZmV7MxxJyMqt
lOAYU6qWfs66qWgOckoAtGfE5PjkBOWK2uZhcoMcmrIVST0yftvqfFcItOxYCPzx
5jsSvgWPA0ffeQUoAHmKcobx12q1mFeZmY4SL7mYSsggFJl228clQGH8mco1w6uE
mF/dVGgp9vX67y3a7l5+mdtGW0u0JOuCrhaCD2qzh8bfMx/dyrpcK1YXoqWdgJyt
4+l9NwaqbIq9Dsy/Vjes0oNsP7KLFws4StUPJQC2V0vi9qVcVrtTxLdvaPHHcWol
Mp550WDR6sPbh2NmSWMCf6FCenWfXkuMkA9m73+QsRhjDCC1j2mPhqgtwB1XKgJF
hwvR/8jyL+NLaMUTyHw6d+7Crrb/0fTc922NBPFjObQOvv5xoxvvMaPJdeoWTD07
HdskvF9uxpD0l7IRdOhAs7UH+Y9ZT+rX+YKllP5/7DwWt4HzKmNkBS39qIjXV9rg
9kuI5pJr2AG5zl7ag39eknJ30TRCLgWge298d+3yYWmQhhvWqQ70IB2458gFcZa4
djAa9bWldDBI8Fkaw9gGr3I3YbnDqXnhho2Qc3p+0hLRxQgzHKq6XwuWRyT6iarh
3a6ix0Rt3wwY9117T9pzgGet+O/5Q9jZmH8Be7sMEoJ2RtILgfafph233ygpLnIM
SY4Q3YPe4eDV+oytHB/7LZg76rYKoNK8pnmVoPjXOXrzmqWTnCSm9+El868lu5EM
cHHrsb6UoVfYipbMDE5VwQFqYuiCQsiwAOy1pGA8ico2ts1UgaoA1MGCV4cvVtNc
EUQ7uyitSaWHHEkLierQUwxVbcAtZuXUvduGTqWNlWga5j+8KE+9r7LiISHyaWZg
LRqIM51Et8iVrdAyKPbyw7Xi5O7RW+vxtN95OV9A2TZh1bnIETZ+89/PPytv/iEz
ajmIcmriJm/yd2UhbleVkPMwUZQ/h8BBBXq1quhvwVpt2JGrrhwRwhKYIouHjUn7
KIUqRVl9nFkp393Kb07NRKKnCysQXvxkX39Zs70fTSsIHo7yrj45bIMrsiqLPDdv
U+nEohhYef4Yt8cHGceVqVYLKNFPn7uGKVB3rgFDae2S/12ToMEuSO6bQ0knUefh
UqqTDFZfWRL3belGniQsp9RzSGdgL51wdHqRHW7qz7Kijtp+5KsIcTCTlYP/8iIm
kvogzuiPbeUlrgBcEWfJZa928w/5AP4nZaD/4YXVYRpeQpahz0JpCzGFN6OyoqR5
/sFIavTI+tnsugFLFm9DNnVspLuwdwStCxmvBcIns7OFu8OQ3YxOjjt1BlH0RTaX
yCuFKjNxLc8Gxj1Rt0Phn88mJHapga5NmXVmILtFjSsRYa9J4ggByaCdNyOFVRGx
Q/4ccDdZ0KF3u8AHSTY2mDK5i1FvVUDN0HcuarctLiO30CT71ABY7I4pYeTvK1B2
irNm/0qU+f160XqO3Lzo5lslPjyPvodTwlKmf81UidN+JFMbLci+09qGTTTawa/1
ywW03eDzXoU6jEVgsjGFPNe1/g0JrQsF7kF09HQppGjo1oZtknLtpFx3ZHvbwI1n
h9ISooy3u4RZSb80pRF9WOITCVxybd6RBPCE+pqDjse/RN3UAURArv7PtLZSDXox
1MJfnpJTj/16RcfIDN0KQyqdLw8kSMfzqbKn2Nyp1DzZREr5uRpTBZ/T74p8+qyJ
rfEAkJxNpNRKzBYl5HmV4kP9eTKv0FGiK3eRlH+m/FQf5mGaJ/DazT/zdEqfINjZ
ldZ3mBJlhPf/XQHgr2ZI/gS3w7VsFAiYB+qNLQAXqw30eB63LHM9bEpL0zG7J0XH
bp9I3eTDG4DwEWRd6BtY4LIkY8n0O4WUsXl9KpZWK4MSxFN3xXtkFQ1PiaDk58ZG
OgCiRIHuwxI2fIB9iiWsCIkSsos3MvK1zz8P+3x9CZKut3pFzLtcBNrFcpeGZwGj
GezFmDJBgxFVXO6ydhRKztm2AC6bfctgv7InjUp6XHo0emf3NhN1SUywsHbL89oI
TAGGo6ysYhK1tnLSr+czN7sckPBrJF+e6s2nliAIh59n2HbwSyAFs+ZRmUBxx3b6
1RuUFtGj+VvmqMI3BWvQf0cpcwJkXj62mHIA39KD9hIJqCW7d+f1zwSmp3ytpfrp
NeOncIJsWCahYf7kkJppkJ9s9FUFoAFWwGAO1VWTxFa8593AOS3lWJEvrFckK3Co
oOJ/7PcQhYZCUToc7Uk/woYD/pOWNbefBAKyjX9xld8dTLLVvrPzKqRK77FEojUE
MMOwzKE1A25liabwIR/0YN9vQ8Jwt/aUbTfdXRShxQS3sKSg/WZ7QrMS5T+YfjBS
5QYIc8CBduAKTImankk2By1RqWoMiRV6wE3myYAnDUUAWlzrklLvqhxD3NHnPYKa
+E2jVw5baIj5BuU0XNft3ZQdByABl4oH5BH3dQ1W+GxESF8EG5ZmL3fFbbIPJdc8
1+X4vxMd4FxLfyOmHiwKWeCOxaxUtzIgGbEgrSk9ChBOr/1ryVOLkyEKkd+8Tt+0
mMFesioOtd4oU9vhxPZzHD+x5Wl1aqEU1Y5oqO+L8Tbzmw2oWghFgapMBHJAUUIR
ZeUEGEIdYPvtYzSWaBRHsJk9l5spj+zknqQc9EjemMzo5rgQ8ZbmD+3K5XzF8nJS
7jLOUMScoH8H0EuiR6gcJgfOEJ2labZiz7+TW/degmaweBZJhUpgvSTYL3uyDAoQ
7xdbBpGF9a12e/d9e/w+L3H3cqUwvXE7yvhrOTDbr8RQwiApEokDlsZr/OUO1gCy
3aw2HTmQpTaJbeBeUjNr6vnAj8aXUviFVl2hnq40DZHEUqrKAyZRd6mZmxGfoJcH
rzfHrfuaeQ8pHseXGC9O1DfBh7afd3MUJpYVmQDYOqOHvDVDVM/C9gMLAmSNRNSH
nInkfLwnxOIEDF/gLoh1rRsvDWNxBdYKH8CsZJF1/q/nhNqpiNUCcTuwKW09QBbB
9tSNKjygU+er0Q1rkEEAat0yGi5orx4pq8cERpvDCwIXjUNHXEugUkIkOwk71/Ab
DOFHJJCWwBAo9clL7DD+3QeX7HNUUiaDNLNBrssAaETbcBe0Cox+vbjOtWbFZI/w
/5VarbPEZfIPlMl6j5PU/i1oWKRXY459RqoJ6qulkyDt+76tiqrlqReOO45nrVKo
k3mzvL2w2Qx11z3lyuUYysHv2T4Mu8ZffD8RRabhQz3+e1ysDK6m+cjxZnSfpPrS
IV34nd6wPM56V1vzTVLU7GrfbnPLO3MX3w3UPccVQggnLF24TbrrnHRzhKruUhF6
YsuNtczji1yRjAj+XiHXjL+5LE3k1DTX9PU9R8au0v36BVPIu/vHEEZf6XfJceth
AQ8ccMYchGibev50Q8xPKqZXec7K52obkqiX2M2LDReieDhyTJKvSTgZj9I2R39u
TiAXNXZHnYMnEvz2cHT2i9r9rxPTmHj3NvxIaIQPO+j6dXB0NJDzwSchpawZc3Jo
EfU2DvNmByV9ZPppwWcSjKFUMfNYJpq/JUKf8lV7OmtfwDvvwdOXdUBt7PMgiWMf
h4fueJGoV9ncJWmgUkwejDdXnhLUuKt0zRdSeh59LdgAqdZxjYiwD4Vt/Y5BBfmc
GgPOuFyfM509IUi70nD3m77wHNfQv8GAGe8Czzr4wCJ85M688k2ny42LRMxLbp/d
D5WdD84HK+BPg4755an9FJSMvYWa1I/tPmAV1LrDJM8iGu5GRPlAHH9M+ff2FdCt
whkWK0LmZ8KddKV3XJlZA+zETXYAX8Tcm76jsTukCD1rQFe0yGbNvGn4sA7EwvGg
SEjDY7gE5CPTy4h7q6IihEBp57PmxV/+UMj/nXRE2wsWXTmEl2GF21xMkJUHQmR6
Tl2cAIaiBhuMI9mX5g27i5gpAddSXZ65GI0uJrA54Bpn2JnbIxnRbdRaBAVtsLsn
Gq8g5lld4vcTpH+zj8jgI9UEpjeo9HU71NiVBgXvNX8IEJJzJtVCJeDeEo3y93d7
9qw/JBd6YzFF9OpAW8K6EPF/5mQHZ6YeplqrMp8z/0lIEjOGlIFLlHkY5rd6Ims5
vH45mE8ciXj0ixXzCFf9FahRo6eGxG2ZGUHpXiqbFle7awjQthnsPPycvXljYMiI
sRi0yrt6ZP23OpEVn5CYOhNSj8Jc3obOVB1Cz6YJUQtZdW03gm/L0LjGTtEF1yIG
TXDadiLdfjHgyBG9uY5MqlfQem2jvGHI1tY9OwyN8SB+JmMZDVZGfwlAjc69v21p
+zN4M68bar13haYWzUnN27zyd5K4bOdoZ1lvZ8wpVwvDQ/xZB50Fn7sOiBiS6Z8a
nDpB/BXplRM2JukPhbvGhvfVqTYvqdOdTcBbGCpMFWVcDYtfHsG7uBxFSAM+ohHs
bW5pyoEAaqRmMLskclvnsTDu2XnrDoMEChB5nOrtr7TtZavCqvE5pW4wVGlorV7c
i12pzdvwer0+8wS79MuWiNnjptzDT8lGMiaykaE0kjFpuPiZFXVJsjAPdAIJp7yq
spHCihNgC4gz2/JliMacrGwSLn1BMNarE4V3WZ5yDUKQPGAyWyHbf9jeGPmFa0uf
CSA/6D7l2NJ1u5b/6+11q6v3mIEb4g9WnmGOmoYHiqjTyHCNmMysakHXnesxtYGA
jjMLZhcxbFkxD4J9GXVSdohpGi+Peb/rb/qWHttrGaXjLYGLUcEldpJiR0dGfWdb
ehkzSdu2lh9WPFs9i3EPed29W73HXOv+jJuiNy1N9or6pf8ldI6HE82SfEkgaauJ
gn/+35p9y165wtU5OutSzXuxiB7iVydo/2opD7+zT3WJWfYBSb06Eac/hwO0RAvt
jx/YwR2PIurHCyJyVriiVtvpOaIAkdfYkShhILhRt+vxnFflTMYE4Btq33GmKqAt
8K49NjXTEd2A/dyhdnh1oT37rRX1boldoUNYucED5RZ1H4d3s4dPvo7OuZ8K2KtW
/VX2eSSVfUeIsWC2q+Nx6jOAO28uboKr2onsnN+Bdzc7Mn/S9JnGvHXbdI85NRe9
hBRJT18iKVWoxDVNGDEl28NDZ/xXLQYplBbajFlwjN++rAKsAs7doein185ajgEv
pUB6bGw328kVF2FVE9IcUA2HXCUrF95g7DARbaExvPEwuGvlOMmUajw8iGiQxKaM
g4ZqTxni9m0zvTRE8eKAGECyI+i07ibj6ZUiOXv9Nu3dQa0vFDU7Zu1+v1idOegK
m72WjKjWBkUBgsBUH7VDluOSHLGt8SfLoou6xMy2MsO5tyOKbQCnyy9I2mSJsu71
yH6/ZnKzkwac6Hp9naOPgebMsOJ96JDu0Tiq03twGpMhL46bdczBOxRKZa7FzkGP
Wo+0Y91GKNL3WoFzyxlH7PL+3vtZpKflAGI6ii94KMFrbiJsRC7/8rJNyHkGn7TQ
8aDOkd/1phPejnuLkgiKd1521P/WNsML9QGuQTtRrxcX51uZd+0DUX2LE9Oo41zC
r4t1wN/gZ89A/NVg2lcAbZokC3ZwGwJ/87XQLOLjA9ZPE1DnBuYExK/abXiIAy1y
UayAwkRLFw64TRxt2NyL/OMVP44pFocI38gmGUgP22DBQ0aH3SXLak8tPQdMyuGt
C0BghyuMXOTM6/ERbOxebm3bF/Zgd5nUGilTsPwtuX8aUMJ7AAyw4brzHmLcqrjj
2biD68EJ7AhLki3jVsH1BauaIihWFfAtASeyo4yRzTSHolLJ6n0Bt+gnEcAeXLNj
AskE69u6bZLv/k6rU2fkzLTpOzLfuWd+1edRPCORDUjOmtCOP32+SdBsvzGlUHpQ
TMHvOQkgIB8vvO6/MJaYf62my9UXzJaqGIZ5ebg4C20PYFabiuzafvGVtTZJQtkw
H2D2jM7y4StwDINjR8YxSg2VOzjrcZiA/d9Pq0DVPQPIbl/FVfqFjJ3cZcW4k9oP
brtpl52cPRsZ4iOjexIctQZX4BFMLvA6bF9RnxvkIBhGqZz76X923WfrUkeb8rQk
2gzFpnXmDKdKlSWO5R9XK72C0swWAF/j6LfUScO6jleeS1br2s5rJBl/6naX4IhX
X41tLOQyMxkXcLT7/JsHUSs4eYr3hm3ETQdAQlh2E5BIxomopr4rdYoyqbdS0H+o
vf3HU3ngZO2IzNw+eFYrZHUpEzbCdbmTsXr6qyCagkOcjTa4MTZ5bOyRo5j6tSix
Dmid897t0Ictqcii+OUJaoMfhhlzrIBEPORZAz0PRaAtUoFPpD0KLqOuap18v/Ih
Hto2V9SbSIl3SGtGIbCzt10Oku7vR4riDmTnRpc9r7YsXjPSW0XBG94og5RSJ9RC
BFc/DZS64U/strFpVHEKGQZw5oteh9OjBmFHvAvKBzZ8NADh9fTNrlldGfP8OoY9
gcM9Usja25AqGkgwrK65WVo4sWs48OTyOZlENcMKQHgojcDCoqwv6ZXcwH4RK5FJ
IDQy/nbAlE4PLiTDWnZNIF/4hD0eTxx10kOyVplYMnvGiWliJeQDBnsYpVY7I84h
ZkjCdTE9tDxS3zYMK+oK5xIUQN4AybG1BXzO57mYEIU1Y6J8EBq/7Nvy1FmQtl9w
ilbaIIyVxQ7oGWM6coT6bP2oNpQEhcI7/yybc1+rJMOAoP2nsTCblHUVCrtfJA6w
1oS8osCdiOVk4b8NLdSSs2y25ofuXb4rI2HepDk9QM73IXe6KgEepQfK+y8WGqYH
MwGtRSZXS/+eUF340zNxG0Lk0Z43cR7Aq7u1F+O3VTuAmEK/qc518NBQskqMZFJn
YgTOitGVksYbC0VI5yip+4qYoxy8WTaI3OrqZJB5SVrWPFTsshH7Jp8E22bDvRXu
Y/nPWVYyEXETvwCACIRddaJgfqV2fOrl4/xwJiF7IbbbJAik/IDjEO6uoutB2STR
Gpr/uKA2abajZ3yy4cHtPEZmiLZv76E4ex0iLVyYr75pyQwDAj6O19f+EQNjV1D1
nl+dVRI2jkjmGsghJpCsuXeOuf6sZjvwX34pquamEXi0qaEZxqta5FU9fafS2vPF
THcyxkLZVNMMe1bDk0ZeLxnfp+k5uPcCnlhuuOT8pnB0q00kXpgN8WwUFGxA6VMM
LGA4j+0U2MwXAIXLIBARBt723m7MhL3ATexzo+QmcOhyXllW5NJGVQKX0N7K/9xC
eMypxzXTJq8KbHVFXfiwaiHIEeAlT+I3BFvlRRB7u1kfLR7rM6KKuqYE0kua2xOq
mxTU5GIHLEh6Rpzd0ZBQwiIIbWJuVnJDrLu4gP7iLYpt2nvPIcJREKTIWlrrNao9
VQBtSTuJXqndJgpL4BL87/26IM2WIGisuQIaOpTOvCw5QGMkp32BKfF0TAFpfVPR
X3/R+HtQB4MDn4hSAC4vdXuX6Fgg3+Jw0qRaDa8RaBjtq/7Aexmfx4ac1VBeRjJe
ozz5a5pMpErlK//30svk3l0KjvMCsgW+OTz6M7D54k5rLr+KGyCW/S9Cli59i4OP
WbEdthBBS3bXry1dCNA6gDP91nyxhQ93eTo217tKwE8cgbCYKjnkmdu69fiRFGrQ
RI4OaKzpPug9M/KYLo+hLwII8g3XgQEEQaD3rW++k29EQwxufgiJBi687mz6NcFq
ygMhgnN0gJlyF+/mn7Rm7DvDn4JA/cj1NkNVA65ogZ4qUggib5fHv5PpIph88Wvs
KZcIS2Z0uBSYrPoCajk9CUEQvHAXQ6VBK1igQ2Jw6/OmQfIVshdNz0L3AsvwBoBR
tcLKrZ0Mwu2ZTh/+s64WwzoNmZ2bKTqjzS9EIiX+MrJ3fDK2UC5LY+38ESOnOW/X
FTtVcmIq5gaZ3M/MTcjCNaj6/KYv/fdOy6vOBxc+1tNw78TKa9S7v6ZcDk8H9SwT
rWe3sgKmEqLftp21RD1wZdje/oXPv/jBcMRHpzMhZNcaQ6e1AfSFD6uFw35VPHGF
8KxXuEu55fdR3TiHALNUf9Z4g5+VwPyj9rhTQFBLer0ugOFI2siB10gY1xqGm+wR
azoz3hZgZgm79MqlByCQmcMUTfAi+17R8e7iJ6p/4lvmIdCRBbRqAEM3v66iEe3x
41ybKoEVVEwfeFGajKv9xuAFnK2TOrw4OHb7981oVDibii+GHLkcPUxdKmQwaVG7
kRFcxUbS37yJVg5h8kgHDwatsoUTwN5J1fXhn2H60ma3wQa6y7r9eF0xUFh0l4SA
6JzhuDnuXnDL4kb+tF+5CkFErJmSLrZ0fIs9qbsldqjNkJykRC5UeSxxLb3WqtQw
guqt8iZqAvKaKdcErjz/W+YONIB2nEo9bLoEdid2PfifI7/9NgnSWqjDKthEqYJS
lTZHdGPPwK/78ymxMQ8ccnCGiofZZ3LXNrfQe8CDWwjNjTfYaPjEY9uVQwm7MivR
wgZwbeTxl0U32rap+7d5IkZ8LZnOUZHAbHALW0xqvKqM3TwbhQ5IcrSrHWvMRUEq
xSd1zy8KIjTx916u8cYqKq7M6wYRFm3zWhO/kMXDkv/5QuYgpyBDeuqk6xa85xKS
pV6b7KdgsD9r5ciWZcqPt2U3UXmeJu8oG9lutT7DBJ7dOGf2ipta+UfUK+fj6kVc
StLACVcO51cgMyxUuaf0DPAj9wdlgolQHMhKRCsvBKPVjfkDdsbyHVggI027QSyC
0Z6jQiLfRzP5brdFv4VmPQtiX1SL6KP80uiP/2/E1ALQSf8gpfYdv5VK+WbNyoNb
NJXaqbx9PCgi1Ve3gYlTgJdThH7KH1ihd6UUQx8R9qDtzrDR+hDN5SqRpZR5AqYc
7ralxHw3s1WmMigHBhuHLOOJ8X+mdUxSCL7ftcGIJvWz+EBGpUgzz572FqxCmIJp
Q3aAI9lOGaZOtKf4XBPrGQxhgthVpdl0az806ZlcK7V1W0jy3jrR4T4/PXOzFLPm
6ecu27snwujoSoX7Ag55Wg5SQQ4pYwnZHv1pKPoexZVWBXy0bonOAaNyAPe12ZTh
spSd3DoyjJWMQHx140zk90R1DTnlSGy6lQESprDnDeMFSx11DJwt7lXvbU7mMuIx
gSnoL1D9IV+ZSwVEBQNgFQk30qxOThIgmrm/C/O69kGa33ep38y1rvxbPjlUhHIs
jQ6219ja0vNEWic/DR2zLdJSsP0IVlRGQ6IvESNZ+5f/6BHFvaDxgKzKgStC8ins
MNf+52pvU9Y6zzcaBCyNI3BHxjtBS/3cknsSK5qOYXjp1PmR84lrg9IijngoMFs0
/L/e+0onuCPzSVAf9bn4J3tBqCGQkjmoSNvTNiGiZrnQjweObQ0o8ldpvC+FXzNk
k5a2QKg8zm9VY676Mg07ZxmnDNJ4U+c5LVvH4KOcmR5/VPp0s9jJayascFit+c7E
mFnMgQPypo67gTPVlqbNob4Ne1aWNHvsmKQqZVc/XwJbWayN2onWDliG0HgMdxtL
ojlUtIBDsYSJY1ydwS5YQZT7NXEx0o5VGiE8i8kd28O6VNHxqn6QYY1koykfen4u
3zHWCEiPI8b44br3PwMUYEmElC20+ViZY14kOuVcQVn0EXMLr8Hb8ay4/9YTr9QX
ngbO136CP6Z2FVXM/V0oNyjDChMlyKpH0md14SLhiMNmu2JOgKJeMBRHU1LOb8X1
ThTpghY34qwa3krbywp8S7B6CJejPp0hZnTR4UAiYFUP704D6YqgfyljGyjgAZRf
P0LO+cFgdnkTx2kr8N0Ekg13Z1vWWifmyPVnFzvGK0R7jxWauY/bjosh2fCKhl0A
Z+GU9Vs/2r5enO+UU2nttYia2w9VEa71LJRcGsY/yKeuBoJUu35zet4+00c1KjsU
UgSz8cJTfRZiglsMTsKmS/RfxBjidAMS6sxl2pZobPPALfcwZPSmJFyDETLd2Wq0
1nR89a63l9SmuzMAr6tG2wfhFSCf9YcnUPD9R0i5vSuipvSjpfPyesyn1oj29cCM
lfbfIkj6FBeioqH3hjQii12RmFyLVC+NFPSA308ohOQtfH0n0s9QaGMKo0XGZgH5
Fc+9mOcZF2kEaFCHRX43E1G+x7mLEfRKaFBo0RhdzJV/eWvDSsRePmLwhy/t7yFG
wXFspsnuRyP5f1O7XHsgydTNkjFLUvpHvdtBhYlLLkX8M31qF6xIonvLWCxda/F3
n6fxTXa96+TKxmZ8VyXwKWjDw8CI8ChRRUokEYbX8lAjsyf5SbpOZMYJDIo0IuHa
5sGPFv/SVp2JhSMUiMibV9nx1hGszNxDUcBeZQD2QnRczapt0V+oSCQ4aS2YYgfL
WwGRrvl2whTp6yaCSpiIErP63OE0t5uKb+2/PXDn7Y+V4yV98ZLwO6sv2vAkZy0y
qAMt/KINT16dRmj1I9B1GWYxQDCke6rzneL0AxjYHP3FS2PtF3lr3PfUiDcmcWf9
RiGCn06dWIMERtQhSkCNO+nJFXVquTN1LYc4Keu2nkvky8GWMgqQA6r/bV/q9gbu
XvxUp40e5v33QqPFJTxNfTXtGTmOTNyuyWNo2tTBipTZsroivWYoHaU3fX4QGM21
+xNj0X24rIxW4yWMGaAVLbYcNuVBXff1dpV7HQnqBl9K4AMRPk5r7pEv5JHPOZwT
ipFvZN2fEkDBbhpY/2dAkU8RCcgCH09e2Ffnhz3QU9UQeFZA2OYrb84b/APpgeen
FMOWUoG3xejF/31LZuhONRVnd0u9pgwHtPZIIfdke81H3Uk3l8YQZmcLwHkxJf0q
EWz3VeM/kA4BervpqlroSmiaz7tzW8nzNlgg9plJbKhuhH6Weh/wFmbtV3PKUTzq
4lWkjHZKdnLSGoGLrpVEA83L7Y1wG84qK84d3V37D6e3DqqOdmGx0MSDI7eCNIN2
4CMd0gmxBSBoQRX/JX2Z3bMZSuudR6FY1G+mUJOPNKSaYx10PxMmRic+5gjNhYfv
ELLu3V0TbaR6xOnvr/zd8OpHJzlsUQf1ePFZ7NdbW0LzjOxE+2XXlZPt30rJ9FSh
jbhDr/lWaUZ97zXW1qE60YQFXiXCl1oHPsDQjcpXiEewROoLQRUAffFxP6HUXEPo
P0TWwV3dnHmJMtw5R0J0wFI8aVBuPtydRbqH0xwxuCrRD+HvndCYK/nrGGRQ+wGl
UJQ7mNvsvsB+GvtGjNm98AqSKH6gmIrAEz5rG65sZL5cvuwgSRo3bEwhiyxikQTU
TwmxxIidI7laEOpITjpanamuKKGgzl1CJ+LpDvjSUBNKBsVo2efRRZDmCwrInWln
gB8z+fQDMXw5FLOAI1caljcXsEK/kGPRX+in2usTNCP8vxh3XcU47CjdFdkICXNR
PZyA8zAsgyRbPJqUDig2vRkxFdYRde8zszivcBEXvg/LN5Y9esHBYZgDc3uH4/6h
z94ZvAJWGYEXgzFkKhSGuElRoko0p9wL2qlWWvzwshel180FAwoHoIkrlN7ix4DT
ldcEVv0md94bkyhOBU9ncYQEF2pZwG9Rwv5KFGQmBHCZzJB/hVubmC18zF5v4Ktb
FLrBT/hNz/aTYWamSYmUuEAetCIfNUUY+MnKNPwAroQ8tmDgUxiHLj9bCMhIjj27
3PGbgOrgDEG1Z04w6rgfOo56c/aBDx7DbrZ4QORode7CbM2xv3M8zYGau7LkDaBT
I/XxulBhPsqlgfAvnEZjbzopaMpXXUB0TvLS1rJhtKTVjB4yStq9rBvZWDcB06In
goI26a8w+MtPDu6vFVO95tJK89CLBoWdx8F0Th/5ujLU43xyshNAuC8kDmxEkDey
FCE441A+9YKsSjvqCCcKTwZLW4gYLObaNOqpq7eUHsJ9RLbr4TMpHqlvxJ4Vtj87
pkC07cHmp76gHeVrlxuD8sl39YNj3lyOuporrougEW3Yxm9VRVTV5fOyo8eP/6R5
xONqFNBaewuma1eBw+9eBUD8ctOpPdgYC/HxqLb1ArbHQLStCy+JFHmCr6qjE2ek
1JF1AmWXQCw8lptfvo2lYde0Ydls93GC17ulWVO/XDfILqFHYcpMc2xxzODyUv3p
PjwF4ra8YihYGSW+gCQqoO8sZGmlgPaE8GV+2rPg4KptH7ytaYMs6+9njbakukmS
XsCH4SrxaSUe+sgZqE8ky2FGqT/0TDRc69b5KcA/DDnHwDL6Icy+EheO0yJUdfp7
bM8WuulA5Kw6ndsBSW097rXZI1nxW7UmPuWNxDIjFYj262LyKCyWyC8qZQ+F/XoD
mG1BPS466Q4pPjz5TA9o1GqYbXp20Q2r1dinD2rvvimcPbtT+1glyynlJrGtFiLL
EgaWKBESX4V1pPFUduj51Zez0suHNz712c5TGC5TCcJxREVruw8dei8aKt9Ip+Wb
RG/4hRPh7hbA+olVlK/iVcLQWH+tw9AIsDGJqTCvXmNbpiAZTIaVjeZZDuWe+imR
R3cj7wAKhwjHkg9nv7EJ5izdMOq+AWCaYB9wrWvr7h9+Cd0y0VsATJHnJwCR28N4
p1AapEtgDWNvSRxnsKm+fCbiCGdtRXawJ3IkN5Ymh7SyaQFDmv0rsyAggUW0FWgA
TuzaNLyAP2S5hzRz3n1jcp13lbl5ORZAxne6s9K4GOL17f/mYiao22/qp/PwPVLb
uRm8EghuAun1mb6QbWmWYPEmiuqZuHHhR+rTQmkRHb26Z0k7wPYa9VIeROfHsrvt
c32uboJR5dLGaqihhGp9aJgKPtKOeFHyC3LfYOExFxRWDXrTAH1jiTPQybBBmlFu
BSpBRy0w/N2d4/m7222k2ax5EkQctZOJSbZXv4PYQZvW6geNZHMJe2pibBwKxxuA
WAYM+xB+mcFell79vj1T63S1vyPTqVlvqIQzgs1W/2QtsnmrRX0CNZc5iaAwU7dU
VMJfseSC2cvJ13t1jrrHJ6KbZ08Cy7nHfRF6YOTmQYsLTb87Y95fDUcSdOJYZlbh
/4Axf88B26gXgU8l/plxGlR+AfJEMHJ7xWhHamIrVmwYrR7x1bNNw9gcH/EqyDLb
08uAtoeLGx0h6aUXojEFcBPdeJMIk/YIaQ4E4hhwFQeLmF9BcoaTbu1bZaqlx6Yo
hM3TN1Vq2+30uq7Pn78FMCG8kj32NHzrsxpoe1dB+/PTdEmeKbDH/TajFrRc0851
JZyO9U8JDllT9BHlKWscs+dMBZn8PsiIrYLNKC591hSr95MhbPzWWagfo8QqYIgr
jrNveKtHxsMKsohJfhFRHge3fr18VHcXAgVJoZH7UJZiefXZH52e+b6umG1EnrRP
FUS4QlhbXx88j0as2k5RlTvzJIQQics7/3bhuHvE6rQpyCKfOuqYZgWgRMgjUpFs
KyrqKGCAC1Evdzk97qelptcHxQFQz3zjahp+8ckx8pcmT37OqAJAWJgra3QvkBEW
I1bZkdxQ71NCywJuuUevIYRi8OAGb33rsON7fCLfvyhZRPueobh84X5ComIHI0ko
zprSFw+j8029nCQ60wgYdA/IBLYRkxpLfCEMRv07gifjgzf7xYCEWmGEVUEq+vHV
ylrvUo5EFKSsjo9c8buM9rTp71ExV+yVQOyvizOwDi5tQQFXucIBeP5Oa3ThMLOW
5Ra5j8siILLbJKdCJE7J6mziNkxgfgWZtXcyJdtkbB4X8r9wEYwnI6X+qGYmCgzi
41bcUCwPvietCP3QPBjmywDTmS13St2n+TRIAbSZM2G1u8Vz3Iv5wzW3d84OXkap
dw1tFqb0HB12aPp+VIiTMFxKSgb6P7St4TeInbm+otj2BJALvzqGd3s4bjdJIMDY
g1EoV9PNul4gYixLEdE/nuiur7casR/B7AtRbG9twNLhgyTurv2MZiW8wjGa8K8M
Yrp0d7AFbVSosM0cksr88cBehCgs6wsuVxkGazkptionQwd3bFDsl9XT1DoeT1Uc
lHGMiP6XH4VHbZT+kSkoVEszXOJZ8BKrqZZLGi4muSMoGT0U+IQ+24DJg4axkuth
nXMsZJGaoYQN7OZnDs51hF1fPyuUt7jXsbQKUn0+nSvOIghoDKsMerEvKeEFXx6Q
XPZQRoiLGgRBeaZbWAFnNZPhU0WcnyqJE1/bcgztwLYllwoW6CH/Q1k5MxOFQeIj
KTI1VQ79QY98oMizbpaONgsz+S0da9hpPMgKfADnUCtAXCv6IZnFW6AgKhmGA9Hr
6ucoQOa7SyW/1d4GY8Ut23absDd4A1nRzeR6l5GtnfbAhl80LeFm+5GaP5uP8RzV
X5j5NbYryUHdKi2y4zHDyN1XjX2JC++da1BvyU1sN0swivmlHfSik81NiY79QZ8U
nqRxPsy+iMGGEaLNuLtsruSXigJe9dRHEwUt30BWF7sN1VLgZLS0RgiXspxCR9/a
UoctMJPqwqWPObMiiXp4SXNzSPcDPI/hwdxobCfS9S86gNlk73uNFVa9VIWB6/Bu
iy8SYCXCQDuOj147niPZnSJbn5Z3lh03y1RUe1KNfq26GsvwAPkn6NPrQ6BEqCpZ
Rp8+6vUk9p1puo1cjgpum0FI74pk1p9tThrBVVS+29brKZP+Zp/aMAWIRutECIfd
04jGDISEKHZknuCcZe5GVhmSfqSkbrauspP5NYHCckAeTzGgeD5zHezU0waw7oqw
TlXzmihAXrF+FDdMa71/qDeOAEGana+x3XZfOtoO1/NchjuO6wb32cEhg4dZWFJE
uAsbL7rHmlocZ224co+Z/PfOR6J01/3rhnrvXN04T0oc/MkKvi2zSAH1mQ5BEXp0
IuUsMnkkOw3P9lc5AbglgY3TC/haB4b+6+axMJq3B6IImm+fbq4hTR6prooxATlZ
pyOgXnYhGywvkzDtPpTN8U1Ivcap7jxvL39803rPj+WGCMI96PvaEFzWvWAiZbUV
9CvL9s3KqHAuRWYY/AVLhpm2MlQP7O1+f/vGd74PMHPaoUQZVf+pbJqmgM1APNTW
AHtx9BwxT3MkueKIoEacWsCiEeyirrAzPailMEjLTEnAb7bkM7Vgihtbh+cIEUJ2
JqF8IvLfRDbZQuIbQXJxDVN78bTFuMwp1PvC+vz/I9VNitgPfC33U19803/BfD9O
xINsVIXz1dFXmIh2YuSjBmBhHxvKKFS9R7mjk0A41r80gvop4ViNV0p16kP+/hmu
qDqe82kk+Yr8qhSaEYDo6tjXTUbpaqKEPlW7w/ha4c3eNRWd6QhL+UZ23L4GdUEc
Zc6oRggLNyAhdmrWwSJRRg2D58JTrAqP4ss0PVM0FAM3da7zgOozPqyVoE0VAVp7
u/jAd8eUtjB+mumFXr+uuLLTNf0FfiQP0hEJzGOkYeaM/A2ByKLvMRnTBXNIt5HY
cNxeQnwr54fFJp/YvIw5f7ZqTnht8gVvH/aNP5Uumkl3n2HSxKvNpuYG1r30N4fe
sHU5XewCHgktjsqkh2KGudfA6mcdCm3YCeVdisHKY09g9bBvvhy3HI2R9YGTh7Yx
tGAp7MI50EPuKgrtLi16Yo6y8iALufdfMFnHb5F/teG7q1B5avzqdR2A+W+n79Fb
3wwadDT7DlP+qvy1O/bOR0H9W+W8ymrBcBjJBYiBqj7NZM2E46qn86aXE3aRlzFa
Oj88P9qJCC07kYjE80WlcXA0dvIncOaeVqRN+D6EPVYfhPKFdoqGdOdrOJhqTYSU
sN6RCiGv26wqajLSUgJ0Zs4XFsgMorL6ckBVs6OjEV0mFQpsPqQalDb2jKMx+4BN
dmAPhrSYGdZks24rItRW7l7GcAubLvucpNj/1dcWy+VSLuZoq7tUfQb3gHYyIgqM
fqjUonIAyn0k/z5K/OGrqx3tLVzb1pJUrSIq7PT6xQLetzxO9gCjZyvnd3GOEoOV
Mk+xPZLGdkVgLK0uD/dRJHdbSZZ7g4k+qVyH5obxuTtd22CGSzb6g4JAWK0F1Gox
6jXhy88/pSoHgdphyO4hwn1JnMLLzs1hii8ouOGnWf24aTgDDGtWxLaZ2Uxo6gK+
XJL+95AE/tgiXFgGzFgyQaBAM31jA3yvu2Ue301biAUTaBxFtqz8jd1xhdFvYAPE
RBOqBJWjfGCB4QZ2B6VEhmXXpHl1NAHag8cW1aKW0kDxcWB40fhc1QNYwcWgfSUy
k+//ClsPZiwfI6kxUG3fAcN4ZqIoDNnaWEqCHLpux3voLC2aT+gQZ1jjadtZRUFX
BvnHyVOSp9GgmVpY1U3EbUWAWxEFPgYoqPfX9LkWt58d8VXoDUh5zmXyQplbDMcQ
bO3Q0eB9GlF5HviTBQ+j0d/9rLzYcoDnHNOh1XiVgq03YkxQPzcHaQkIsWYoGj2T
3Vr9rWGg2bEUVvOh3xzsdadsPUEgh+jRuZOybqUuhroukrHT8jpx62xMWUZNN0DY
mpPQqmh+TvQ92+gileZScr/0Vai2K/WA9ReBILrbiwPyTvH1pZUWor80AJoxFYhh
ySWLd3p8EJs3UzqTDUiU6qVAItleHATh9YRdX4p5BqRkhkswS5cOo+e6Hfv2nMBJ
hoAJycFYGROBUfDUfjF53UWFLPc1kbT4GpzMWk4ydDYA/laEXMZwSj8hPAu3ix7Y
Ts2FeUM0JbpFN2bLaO7c8CLL9usm3ke2fX4+xLi4wDXdOnEZwImwstKS1vpEUVT4
quJcg74Q5WAhmhfTmHfo4/LaapXKNo/e3fhUzE25aGPFrh54brfve9mWqfOZeed7
VFnGVXHDmaAx+A6nM30vdBQYKSSy94lOHlsTAW0FnIr+YslIFkbukW3baVEHAYKs
Vevd7IFCEpughcKQgz3RvS1Whj03cBNJN2H63DKJPeMTlDMnVF0xTre9EVt4yo+w
Gk1vFudvjVNMvZTB1DWAC1BvYJVdDYKdD/vj9ldDiQoHjtqFHN08Uso/zfDKM7C/
U0d/Y3W+W1B1a0AenqVecrd3RUelnk9SlaDx+psyWiY7k48/ajxhSdEE8hMZPnuT
/mJCKaDxm/VwnB2O2XSahv5BT8Ir2KF58D5Eh/YxecaNX/VQ8eWi3xP4sIF8aBG4
AuE0fqosIaiN09SU/KQKe2jaa8l9i3+nTxi6N9hL6rvfAfs9sjMZMoGS8tAPnntp
nYNM4G1BzOS+e7RWftikKBnLrcT1EjfSuo2jtcfoXqSZhJym5n2x5+OeyBsn6VyD
+V5NEclRvkSGI4zzzApqd13HwE7yTmyvmpjfarrTECpoYEzAaWwhaPigReoJZJLh
Ny5MUlNaAkZFubEnuCrd8bSZzDPzBW81ObTFMc7B8Evrkihi9GVHfYunrSX9wjEP
WZKcpHXjMgoxX27gteLC3Zlj4SCNJwLoIeZJI86K2KX5lKONZGmbmdb6vrabVDYB
wuIOeiGpjYVweEGKPwSw2tnlllhl3a6y+KRVs3r4tzk6EmlsZ8uQkzfC2e5/THr7
prWV0P/+DAq5/iVHU8QCQrD851gm/oUe9zZULZOdqMPv4ywYcb1uK37c4yvVD588
XOup8ATR60BZZkXe1qri3B2zMGP2j9UrfQcESrtK+d2Bz2EZthcUm98i/WpkiO6X
JYSAQdxMsBEzFNPw7/mOrLlbn4shVNdZQRozsnaD7LFn3vEUwA7jR06tk2ST+2w+
FmGSLR4YRQGVxWaD8DxGD/L9zX/ZJcQBPn/Q0JcIt/NZNF9dLXYCyMSE3Xc56vYf
l3d6Gh25QI8tgjK4kOyCI79BzlOYODKlXd9bHy41O99Re5/dKjhTHyLICZj41Wtg
Qa5V6gcHRGA037jqDVjwGkRzKdWGAz3tpXEmVRa0TgmW0tZLVwv1WHXlNJ4PovNh
TI8j2Aq5HJa8AqoDuDRzX5CG/RapgMoDJEUNTgD9i5nQQnddFJqyElwJH0T+ElF8
612CcsmLr25xg+63XsK16jevaMUc1hWbPt/fGFfk2GlrPS8FbTNn5fqj+HZNvYD4
8fHu+15ylkWKgCQFwHJJR7sR8khfRBPv1PjxdlIMIuLGzCxGmgwaxSyQm2Sf9aQT
f/aFlMiOffA4YCjOh68SE+IUz/sk3eakcR3IYXyly5YEwLEnyE674/DxZGJJdcRX
2JFNTUjvQcNsIKOMZCztRXbnpbRgmHQy3RUZ2Z8fH7SuBAYUbw1qjGEG9CaIm2nw
YcL594cqe7dSIXUb5CZX3qn9rd9Dk77pajoMFo6O9v/wsKPnNqSjMjQmmXxjYzeu
drFI7hLiRn3mgwpnjyh85JlH4jm+nQVRlN94bJ/7tm8500w5Vjym76X9UMvU3jZu
tSw/RQMETgr6IW1razEeyA41qoO0l/IRj0KDy5SCHD7ZtgOpi3UpXPhuuX5mu0OY
NanBuVXoW5KlvCrLWQ/r85z/dBo4I6dCxSRzyuBXCfBwRRwOvxtaOhtR3IKFTI4R
YrvIoTNHprdiQUQTfdlHz4JbFVrQc5/UoaJGsheJ2MFzuCezsIW03fFMzenak7R8
c9Vi//R35DBv35afIIhHwQW94vQfTebnGCI5Se4WH3j2ac9x25V3J9htd2RoACKW
GbG02m1yH8IThMlty/GhTUDj9uw0YoNAiL9kBHrb3Ea6qQj9SfsH44Me9sjgbiNw
XgU44oedf1JgeAnueu7+O/lABRfkorg+GC+PSJ1RuC7+3ylOUV/gpuM9w6oNwChv
c3A1MndjmOXDsLF22MyuYGopxdZLpCj6roauEa3DsJoC+KU8NSMg2SrD0V/oEfBG
aycd8gyjB1VsuxOiun1FiYpwTq/d7rkPkTGG6Edpxk2X+BRFYpUcPzS++ixOdsVf
im/7ywGn8YYpasIsOrTjy0QuKvu+VoB7DHwhq5QaLHX9xHYcwB2AXB3pdu3++2ch
oS8E7LgNlxwGjSEikF0LkZjNgd0XcREqk8wQQEiZUBhfIIKcZ/4wnrI3X07D8slH
WNXHDoo6J78BjOXUR94LQimgMOXcRoKTBm/Okrkk/16CZAxKdv7sRpSPpG89aJAA
o5WwlvqkbcRmgvpMC6o6UE4PjE6Nrh1hZXCo9XlTeUC1yeWUTaHZud9U3ZbxcM46
kuWladZYjNIhSNQw0qKYmG/aeRfovncwpl275R6e43D4xVCHAZj2lq99/Q/73i5V
fiSECelH2d1CLO4QwYjuYi3r7JIPF0rlMlkRHPxKVuRx9y6SSHctMwx7dNDCacMq
H0YofllK8eHBXYwsv4NCgdrC9vIW16ABCJsC5Kz9onkCiZCOwlpBqO4Kyn4QuAcH
+OD4p5LThLzxifON8aFlpEM/LbfTsydlyktT9DyQvmojiFEJ+kIzxnkmwS5YpfOA
EI+ZAD+Rj5Ym7xERuERwfFrKEQWF0JWuKibMzUzXHtT9n3WceHVvo2fY99/4tv3A
ecJKAQ1AT6uR9S2qjpq61qyx27gncf7AICnC8eOCCvkAKNLlA3Wbcb5ggf1be0iE
T9xZFTkqp+m0fj6RbOQ9z1BGVj8WbxYNSpS6cCsnjuWclu+DwrIfYS3sqqBsT8vn
bddfNkL8fycUXn4FqhMihMwri73ofNA4y1loyi+efIAKvD1eDA74lAsgZp+EB7IY
7W3Orf7yZkASMZ+p+q1KlRMIxw+jHFydXHjaU5uEb7fT30sYHJEg74U8TZ4OAM1d
It7F0Lqaft6uz7L2ZftTjEUUHHtNkZB5utMEUi2Nle7abHzo3A0kOz7xDxUfKh3f
kqFu85PlLtrlEbtME4Y3s4kctG/VhV9PPV8n1kQnpT6L3MXS3NSYQ8Z/MuTNkdIg
CevOb3yYAJhRqKM0q5NvQwJ1wqgUL5hgqrzpsgj/8bobcdzM/WrhQqCwgZxawz0s
3Wz1ywS8RAe8x8aAXfazvADpFNL4XxsnOxllN39uIKImoH8vFnDMdcvP0IYj9Y+A
JJdTlj/Pxx2d1oXT9X8tnbwBGhp6p54gI17iOkl5bLZObGsKagl+nkYj3fZ9N/XL
XIhk5U0EdJ6GP70zJrD0CYperhcW9K0GE1zNRvvAH+4xTdn0EAg3mjQiEm2CxzyD
ypZ7d9sI2cx9335+/VuQ6+R8asdmRD8/j3pcD2eSXkmuDCFd4tsfTg5kkKrVs5Q+
v3c3cA7o5bdo8885txoD7iibbjHxuyhiXKtBYTxPz2jZprpF6g4/kHeRQdFEdgQ8
WOaGlA2L4hPB9X6lHAwbzzVxtKtojYAnPfJYQxOwqmN2I7Q6Zw3wfaxg35MwELED
69YAxlHeNV+//itZeNeP56PYV27KC6y8z9cE9EzOp5ACDkGCtI9Z6rzpEmCvikjT
rko0GAksFGjg5oYoW0X8+00IBCVwbBMW3ESyetRBXTJKrM1tn4NHbewdqxLmnzDa
SP38Fb8Qcuz91PAxRsKEKcyGWjCyfz0VSozUo++yBDm5I4CSSa7K61X1GBfoM4/8
evZ1+/bwEgSYqQMYEOvcgmr4m12T6WlIpOOithgYOz2WmTmCbEj0wvDdPkfu2D4G
1DAzHyM0pVTBAsXg7smtXqT8v7A9EekTJ+4pRtbo5oEV15rK9G3TZdxh2nsz0FvE
24rxaEyCf8z/IrooBZ3ObIIevA7YkK2xWLQ771w7Stii3Jf/NTHsfERvAAXiwU5b
0fmAJ5v83VoG54auPbq/5KTEf1JnUJVj5yVWLWZW07B2Bl//NY6s9HfdE4Om+fw+
Iox3vrZwQ2Xb0CsOwcMRFZnanOHINtIqswYj6hjYOOjrS0mFJCnh0vuK/DC5sJV8
sE2KEuYziJKN3Rl0X/XXtQIp3z0IOAI81WrIw9C9XbdncF1PXRQk1NusirlXNBdt
30fKNETn9yY6QKbvOE5Uxmo/ZBmI46ZsVoUMS9wi4NTFuU92ItJiunAhQZxgLtAS
6bNzh1qZk2V15uTMUHQmLqhZIvMjpUIg2Ja6KjjvmPQ+rQHsipMVkpJoR9AA3VjY
GsJL2TdKE1YXL+lAViTDdtDmFrvEh22UQ5ylseLHKuZu0+gTq1jWcBGBZBDSZpUl
X7iOcdqx4tfM9dS9a38khA2mld0borkerfa7S8+TpS3asUHa71TMXywsxKDc26CP
f/90ElEjZnmyiouXqR9LoZj3bBCP1XwKSn3gE56kh9cGt7bTubKoMtOD/mhdjplr
Wj022LBjd9sF+oiOLyK39aYi1QAE6mk2loSSSkAzNSf6pLFna9OW61KKPs1WAKCA
9s90bNquOb6kEBA6lY9oO6NXC+Kjxr9awWcqI46R5fsbzDgynoXq93EIEbxrrS7k
3Sz7rwwVyLTqYcKf6zYBeB9cFXc2OzjME2M1O8kTaD2NTPoLRlQY6FKKp6uQWpTV
l5vlaZ6SOHseBFDrbBdKMYVFYf0+2z0Xe7UuKn6qpyKEbUeS6LpVSew7buwW7+Lo
ImvbDpCyiuzq7MKGH0VMJnB7Kuz9fxKr8shfd4OE/Zb5FyczfHTOUAI16oMIUZQT
A4cvuS40P4WpA+R8q30v5QSBiHTMvIBUdh9/DzVECqqR1sqlMvfXtAy3Pz/PZ7LG
KMN6Vz4ZRSrj23FLnMlQIH8cnXF/kkyFr1wqVfHYUVQhclPFBSYSarAbAr8wv4y9
VJ1XGFBGMi2xit0qB5w/Rrqqg4ZAfcZ7EF8Nii1K8dOnBpGLDtxtLNiekabqO5Xa
1OnXi9Vr7SSCkSK9fBYIs3IHsRaO881cScDqjv60bHyE5MMx194d/T5Ok17fWKL9
H5G8ygY07OklMw5bS1y3LSgmFAt7l87Tjq0T2YEnarmioTNAgKyxJc3KVJWm4S/7
6cwIsTy52p++tgh6zWfjxtqTAmNy5ZkAcStNJYM9cBcqrlrDM881HdZ14/TrY6cO
y8rjbTyMpbfXRVO4TfXq4UwFEl96HjU83Z/1Tgdpqr+zLSyzdCMnITq0gx2jazNn
ezJtROEyqSRs2fRhBjZLZUwezpJ0/Rf2DBWi3JyQARQ4/V+Xdb3nxfC2mm7pBWcN
oObHQs0eW8mFPD9w587PKxOCiNc88ldJfZueG8GKAyoJ3fsUYuvOK+WRDxwMYqn4
B82HTXW5pZ43pDsJtKzGUUxFhtnzglElzVMU55RD0svL2wRifvXpzr8wWJtSxh7S
7KpWl1crWbRyUOFyWbh3822wsN/VUY26c4WyQCsTMtK9/T3Nst7g254FjQrmYa3n
z1ZUS0amEswL+EiebdMVbeXtmUF7W0FLTHOMoyt7yutEBSZBUH97DEIJYqCxJYuY
DBvLoiLj7kQg3hOLXclNHavju3SgG5LlqPMqnzOAN1sN2exxsokoex62MWu8X5KP
gg05RjF75IFDxzFW4JRwEh46iHZKUdx31XhQSBwM0nNhpmzYkaFci5LKS+x1GJoJ
Bu0rJJmx8w4ziI32hRwGsvrUZwapQFsq3an9vid34pBU13ute4d7jx5bOEMIaCxJ
+UgiwIfKerbwn5tpQmjlRNGZLPXIJ8aOFbngwkGX6McdjFwu+hGUAYbyhshTeN/b
Qr/WctM0glp6dkPsV7ZWnHYC5EY49vFY0NEHQ7skmtFtl2eQKOzZrrPnubH9UDaB
ejowGk1VOIu9oLB9mDje7ez+o+Oh5libcmM06hcBlvFRrGCikvHDgCt6PTdCkq1Z
DDekmsbgzyXjiMfHencsq+6uATLQBUC9SoacU1dDwsjoQn82TJqMGvgHCCmb26LY
/t1H+lRbjeb8+XkjaaRFdxos0nMv43d6/nE+AmzEYXyBVxItPL8QS/m5dzzd/Brl
YI4wPC56NhWp+fO/1hOlL+x1EKoaSw6o0BEb8DFxRIerozCJuPX/qFb6f1zcOUvj
c97urlHLRIFlqU25Qx7EUfO+VE94OoW1Tyl51XsNyvza8Co1+A21be4dNttkPrQN
cEd5v4ib6LOGT2TxcogFWsiwO4Va8vsROrMWVztERoCoUf1FxstO6jSIbnjY68yT
chdFsvl779v2c5JS7v3RZgywE4vHHXLw1yqptie6I/IsMnjJTGPgdRyevtu2gK6C
pNTwJkC6sYnW3JQNP2lv7iC7sp7rUn2QLSq0oIqczouTHmYgIQyHuVZVNq1pEefL
z5Sas+wpdSju/2JhVkN+JodF98Dvl/niKiApLoG2WbbM7JfOPp+i+pI2fogk6+wL
1I2rLH6MZhaYI1mlPyOZrmi1D/8dXy0k1bQqr5D6wViY5SDMR7V2mvNVnm+r9cSL
OW/anuyw7yrcgxV+R65PqrPcSUA2Kblstyi2e/KXnG9DNW2Fx3GLZXzvKwfD8oPq
ZjizndcokDu6uzlG0KKZWc8qK9UgtJ6QYIHsS0qugU0LfQ9DFkKZZh0lW46dKE21
L4Cr+vdKILubwXeOYT3+B/pCLSKyjwKMOag4KOKWIWyfxO1fv4Ke79QC0ss7blqv
K9X7XItVLgVHaKhe6l3xJnPscORC4LbI+tsuKvYhrhDBuPS3xbMQNEtJuS/9HgDd
2TUpZX677ku8urNYNTx5SqDPJ7voHa3gxtgH32YJoMisOXh7nKd8kcXWZGQU5DMD
8YDl+I+WiVRu48DyzZ6qBMV2VvkAPOYvHMzozkUgBbyjiNPNWhWh0T3Gg2I93bbr
wiKesOfQ5WAI2ZURoom7b0qIPvBIZoa9lcQbbVyiTqmzbWkCmFQLVREM/fy5l9jj
RNb4DyfneQjJaChsQS8Q0CW0YzlUAQFvIG32fVj+IJvKhYRWXmorQdq2WRidvJAB
0gbqm4daBcOscKhit/WtAscjTdWBEyESgxu+p0QC/wf16TQNGDtfUtkTXKRfEs5Q
sd6pu2NV+MshIc96UY89tfIC9yh8Td2sWBSWl9/baKq+s5on2xHpt5o9ZFtL/mV1
UVNUy34qdaMje/RHpwI61DbKiUPK9+H4D/pmYYmFrkmNig41QRKRnEeNWv5CjVy0
xc0XcbDnLgOpSY6mioTZLdX2xVfYpjnYtYi+/slcv9VyRHsHmp0lL18UcB71TYAK
x/4sxHoYgd31QNsCQdxLGUwDg4Lgy1oczCrNvKP5snl1JBcy//HvfdI648chyX9p
oXsgo/E5dPKArCouFqam9HoxI7X29/VD/YnoQWFCywiCFP8ujJN7/E4Ql/+ijyzI
eCx459+qsP/Y4eOooxHbrmhKua+uCX9fj5VgXifsl7dVEdyHI8itk32mifyAzZDA
mKw+UWM+4/igJZ8AOXK0IrswL+vyFa13SU5wspYJ4EtQoh85Bzga0X5CX2gQZntA
7TOIoiimgCKoRS/egFy+NvOdi9FW9t5Knzys0c0pY14MBWdsVPTusoRgXF74meCI
HNp/q4jtJiUvFqATQ6hsMJxfegmrQ+khWDYj8EEBosDIAlHKzpomOHR1+MTWWBdu
eVdIttjHDQcU5zeOl5MZaDWUTvzZDNo7QyoKwA/OCqZ6sKl7/BtObcmo5iD1au0E
Fwd+2FWPljy2vc38oGWnSj8HN2GOyIVZYPLZNQkEKTGRtRajqIXGEwV6TGQYwykq
7lIu3czq21H+4QCytlVeyu3/wZq2Y6g9C7YvKMIHOFlLBaiCX8rzPFobvj+aBMnq
S502WGVN1Tfd95tHH3B2z4hWe90HsWfycjtUTA9mRIsYT+KnaCL9BkwrpjHvuhgN
wGxZSvHBd6grB2L+I5Ukjmp8dTOipc6MvOTzOhB5jBc=
`protect END_PROTECTED
