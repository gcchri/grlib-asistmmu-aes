`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uADga+iTyE9sx/NVqtM7a9pXh1Zu0wJD7xyzAFe2Mq6WkCZCBYNUdZPZ566VyK3R
Tj13cLTTsPiOHjsziYxIP3GgZyMWX7A7j2aDqqQFW9ZkNiVLP6PCP+u1tKOTv20n
WRLZkWGG51cIFtHrcqUVv6aVqayTlNTh5vEN9fxw0h0kNsVViaQ/HpedvxKDbFw8
7Iv6Zc3CT3LiayjImPjBj5NdbKgilfFSO5BC8rwZPMHXQytNI3hYZcG/EFhlK9ad
iYZRES6ax0tFeHehUdi13gKRhBk1+3lOQJmKja9bJCF3XfLO3l6fofCzLS3lT5WK
oXt/BcN2YiRx/7Zbk4FGwgvqZXYBOXr7QmbPxo1ZjpsFGe4I6tIaIrspyBuTeKTZ
4A07UTSLKH1bOxVrhzaus0MyC3SVWvLgKIb2WXPpE4pdEEajmOKco31ziu/C9lqK
2xvWkgo1r/r6kOcuALXTOEvTPitT8ktTsN9FKJAO/zFv66YTX+WvxieUigs+YE2P
om80g8O6andty3KVebwEfoXDvC5eZVj07yxLMl7CPBcF7WIyDhv3jdo1BrlffRtA
EDkEH5osiIkgaVAw5sP6aFiQ/YSSKcbGS6jfRytlDUpgMmKl4TmARhfXQwB5JFMb
fHFGOs7fg1cet/wDdUVC3XsgLJjPtjtqOrevzT4QrXKFjObz55tJ0X0cK6tsLf95
Njgv4+hyDEGK1tzybF1mrpoicFjo5moQQ+xb24JkIZGAOICDGMtOr8hhKLEmwTqe
EZ1Z8JXBnG2r2vqhOdCl2bpDyjZ9XbBu2UBUSWuA1jIVCDUZfA+WGE4EfRok8197
6i4t6qvueZyeW2RMAOxORACAsgd9HmFcvgDzeZwrilNM6I0rfKN7KLMqRq3CNhg/
HZt47IEbXoO/liC/AaIVfw==
`protect END_PROTECTED
