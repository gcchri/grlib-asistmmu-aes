`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AWL0hHed8v57G+nWO/MiWm8Q1Mvkk93Ub+NHnXhdHTUJnEEzaRoGfE3uth003zZj
Q6BOR9qMfpzEty3FPqegERhv8TEd6n1nmkw8SvZxrP3GTTtDcxndXC0hwFYQNZ/J
Y4AEm2hp/t0WF+joJ+I5KTLBv9xe6TckMN2lTju5yryZMmNC4jN46Mx8Ft3NTrTE
H4ACS5LLAem9W2E0ZapCbRh3M5E0fEJQvLA8CwGCJj6v6HnMnbnKmQOfEbv9ppy9
z96bo7GjwQ2xuU87lua1Mv0FpJYRCIgbrv/RuVwcDzvt8zyZtjpMY/gJeAOBKu/a
fQ4+1W+ETBVqwG5w2Pq2e6zndJWkUZUFbReCbTljM6g=
`protect END_PROTECTED
