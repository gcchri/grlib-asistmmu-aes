`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zsbYtFIwjJpND83LCVLB44O1st0mJjB7U+2YwArqnNZjtu2gkPqvuMY0zOYZbNLq
hU0Nv5x4sqZcmh1WOcEnzNgWBRP8SzeqQIqZEdLFN1gjCSrcw/IHcL0gzjg2i/f6
8RHZ8ZD8jTmRePHdY0AMnlOU3k/7FqO8zctkVVKLfAXLRdeQ00yDdA/BzQA5mfvj
UsgXBM/2PhDBzx6XJcRXDG1SfDIhJKS0lDVSXbPuTPfN4y533ZcR3PxkpdMlMIuS
10veHhlI7XVpROhGB7XemNFA0xheFB2BkCujQhpHLr+R5fN7BvwbwgDNtwahfdL6
ZU4Tcq/XSMKHofmSlatunxe9lA+mDbgK5g9PDr1mMupe87jqCP9eCxKZCprWCqPf
8GSkrCnzzTYzNyFagEOUlIwk5TYnzIAdxBhhF21Kqt4thnIR12kBXLT4vAAg9w/6
vn465hP9mZver/5cXBGE8NpB+d9oThOUoNhD9vPcDoIySMb+iM2w93YliyOVUg8c
f6RYOJ1drc1j4GFVo6v5qvZvKQ17l7w75OiZQeK9kvc9eKM690RPM5gRN+S0jGy2
YQW32A+gTJaFCGAxeBUPlgBB/X+ZLXmy2d5OlfwEWF9x279RQeOhPy0urUwhPzOm
9SjiGC+Rtzp79nlIJwyYgg==
`protect END_PROTECTED
