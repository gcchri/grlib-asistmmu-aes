`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kZFTiOpBwaW7RGhSUBwHMiHfQaDOxspoTKviq4ectDO77UthNURbmi7ik6zn+O8e
2biRc8PBJTS+71rNOsTyZ6YZ4a4xXUc3Kayx4JtZ6iIeWTZekU4fP+GO63/b/n1j
bHbQtGBR+6HNi4MykkeU1HKLVQMcMxIBUrZh5/uYlaCv1BRICRk0hgsvVNdrmJy8
HQEE0UzO2rBxjT6aQtvX40oeBNjyCo9LN35R1zeqgOXUYOqmH0qiLKpviW2lXjEi
1IQxJuouPFcBlNxgKBxCCHBiZk1UsWK9fpNx4MjKCbqkYQdChaABDFmLZquLqQhw
wjp4eC2E5RFbu0XaSM8StDw6nbWEujyG/6LosFT0r7x0zN+rpm0JDvWdUF1vI2E2
TV117JOzztN6lUhStf1e6UYvXQwOE33fU7XNA2+fFD6TrLp9HhsiIctSE4hMb80A
eIqRF04/3maPgtBuFq2w+48r198kGiA1M3XnEnY9yVL2Ccdpv8fAP4wHFdbVoxca
HD1l3dYnk2shddim6aL7KelL5Hu5fchdnbywi9o7cHnUC/9Yv18SgamIi+Ai0pmO
oy21jIlDmyBae29RbZwsU/E+M4EKOasjso2l8jxHYlhjnsoAO0Ur0k11DfA2mLjt
0nzndM11DAurYWuf9+8RZTg+WEjqimRETzLdHWNOjayggX0S44SGO5nse+BaOSSL
FlqPApwSK/w0a5umKgHd+Q==
`protect END_PROTECTED
