`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BfKqegRdRuyNxcSOAE+SRCDkyYanHQQwNVERvJi/OZQR4e95EoCPpWVLwkJwdE+J
eQFW8qpDQI7tS0H76ZDEk8R5XVQp8rtalaNyJ4s8UszU60ElDG4RYhkcvUAt3A5x
M+ND/yabr/r2b4B2hqdd2owrT4kzPmJ1YxbFzxkeFgY3nIih+gxFixDIJa4vBeg6
5Z/xlcKAlB0Jo/Yx6aal4/H0NnmSHKMsnZ0Lh3jl+ILad/IjDp3SNksaVd82/vZR
JuQ8QfreSZjFeJcsdNxqd9ym6BXCsqtBTsSm2MwxfPt3QtCrMaVuqzBuVsk/19g1
NgZPeOBnAi3MPo4DTvizSa/uqIUObBkqM3XX2HjYLWs=
`protect END_PROTECTED
