`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gsIpqS7v77aG5iFP7lmfpLHV2VZlhQ7TPFlVQVSF9zV7poDXBiEeZ3KO6F/i6XVq
SlFedoxejY0F5bMHo6NMn2TDUnglVfwtK44V0XEz8BeO6iMcTYCN1zZei97vqZSg
wcowvJhYETkC1X6Xqn70spqGSN7EYD139XozH5wj+eDzz/BBCkbCnZr9pnBB6WnV
sHPrP+xXIByrtsvNRNjf44D3xwz4UuRzLGmPuo542ClBbxrw613kvJYDXs16ECo/
g+uT4z9kC6AG79V5/Kn08NClGnVkUtvcl6v/QmfGuGbfW7uzx78Ri+SkC6e6Fj00
1ykKILF6g5fyakCtftmA+XWYLxZhUq8y3vXkC8UCPX9gDvyZsShhUloZaXJw9yD1
9zWkYMFWmM7Yyrzkrs7q6DCyHB947vfVTQkuEAG//ekQPjSxY/e8O/W04o4Safyr
BGOl6wR6Aa8wnrVkJO/42rsq/LgDhbMFuENs+IvLz5hnLzBBblOW2kDpbXZJCEln
ZHqZdZoMYPU0X5a3G16z/jqowyRDO6V3juOYGaZDcbkXHJ0MaHqmk14deEbv8t9F
6AmJ+HiFVlhbvyaV2f90rKS9MTA3swnpks8UONjueCsCVq8dGXxH2zLEGYqrks4M
DSzJHAUrCnhPxb2QpEiMgLyab1Uca5djvwm7z0/PDdaVXrs/adKqS1j1ahfyrSor
6q4L9S91EyQr5Nl8ui+baE4G7LK6ThDjADCclFIww3y+DLAm26MGocRV7R2lnsFs
e9r7lX2Qw6lg4KAKZrp1M6ZESBd5GH/VqR03ABKOqiQ49bmSbN/bOYYdZG9e32HI
QiwvsCE15o98B6pHwnmsCRtAaa8DtL0Hjll4M+0ieYqBywDl6mD8HC9odDkinPOL
Um9PqG9hVI67iUGwWTKwyrFfLiCZatSEG4wFOPio43CbUngLiO1UL+k3sbsE3vny
KAh4jLPmGIv1DFgvjmGkFDrt7YopbT9A24CpK1XW68zGjtILQXPtPf1na/GQYPv/
jIifA3egSWaow2/Dv1wB2eNQ0RBzxavZrinACQOayHHRvi4O/+L1Y8jvsn7kJi9L
6L+IFIKllULY1Bsn0XSyT61FN55ShuYvE/DZy+Yr8wd2xilPjOlBYQRuo8x+MHBZ
lSnSmJ1La1/CyjGXxG6BO064y720Ybm+acmYSmJ8UQcwiXECiEgs2GY53kvMf+I9
2za5K2pZtFO3LM75fuFOVWaqBZzwWuja5lYOaJBu6JBTf4+BTbcVR+GmGwQbVSvY
JQAQ5aw5fBZ+A8djRPQYpDcLImbl14uqntOw5c/SnZJ+4ReybWh6IAx/tzI2zZCC
no6o75eJ43Q86aTS+kSAcP47u9HXrfBtvY6W9kxPZMA1wMP/VLtngVIvQeN0KIAD
k2yX5quszLMLuZ39FTOszEFueU4VRprPJcSjTviI2Xg3hwa/IGLPsYENK50+YRyM
G+6Hy79lSSuYgOhr/ofSEbVe5drlxR/3b7CTAGlvZOT9kVZkUowXztE52vBiKJiu
e7KQpVTm8Lak9hwfSMdIeUdEtDN3hVCXYpO4JccWNCXNX+31vgruryE3ybuPCD+Z
oySOX+2lbx1ijxr4BhPxLGhhKlICeWoB4GdMBvkLUdNOqK+o72FsVNhAUjC7Kv8Q
nu1YeWTMiEVq7kUhHWJQ5lN04IOg4oURdZuSMCf+4EBE2DsBDXyBT5S7X7TIxEcm
zrsGqGgijHUjVdy+GNDBdpe4qzaOdc+06OgmydOxYnQApIdnxMBfCYDrjjrW6doE
FqRD/zY3JWo59FkefkihE9j1ccxdZITv2jJmNPj8h9q+4E6A3suvWAoE3x7J1p48
Du/GXf46oZqkPJB95FYeRPNlPtTThd/u1RFNzxqYxKlyNBdlDPzt95dLTxDdacgK
CZmXxchBaNFdabdfTVwb8oy53aZKWsngCytDhNYvh2gsM6TdUbqBnYt4/pI9ioSe
BNybCL6wvikVDdpN+SBLvIl9yjA7LMBY5bk2LCPXKmCZhke9yBoBy4n+8s1fmeKO
kQrSNzCr4YoZln4uMCnVd8tYcE4L9m+ab+TUI0OktoC62xx7563TTZhy+55G2vY0
vavOEcH/8KjLCXDV0G5HZ4POCw75b+rrh2itkD/G+wnteExyy3FQC7QYdsW4xRMo
ZYwRFGkvcWVeD0CXmOu7ZvZK6Iv3vzrvLBpvvOzBmIHlmq/6mUY0mqhG9Tck6emV
Jwg9Pn2U1oj4JuuJcxZCkFo2jynOoFfOhainreCFtHBZjQQpeS30Rf3ipvPx3mXU
n7a/OBYqPk83HbuSwMn6/UQ3k+fvc8n2KjiVsvbVydEF3Gi54dfD5DdKTBqZi4gZ
vPntwkXbsR/SXjpTRZOgslqYD46v3P+BFs/nTSDC+m4M7MiBQoTwvJBbrApPa/Ya
/VHtnnLP9OL4UFdZvtg3fHYvQfDDuQ25/vUEFGNyfmGQlKFG88NJ8bAAh7GThclr
EUeg/GMQjld+0VQ3pFqZvS7VTmi5G1sTAGqBwv0Se1bQmzA3w1gnlQ/Y5jj2OG06
eTY8FghCZQaLldubrmP6AGp/Qr6G7YDT2efUfE7iIloNfneSSNsY5hWA3ydl0mbz
s9RT/7mXiwj8w2SC834m3dx4dwOEmOXO7ZqUXKDSL75BN3LIJNQOBMJf7iceiuda
2JAXpe6+jUag/1m2LNRXhqtcZkko3wDOVZociruNma/JH4qTROgd0Y+ci5nQTwxR
DafTGS5LwFAnJvdqZ1iz3JwBk4MZ200SZB9RTh4esP1wMRQ3QyCkZmpZubc8AhK7
asI1+Tb1CXnHoR4ueZLNGgKjACASVkOIZpHIirtTOaWRpmBlAzUAHQ+XuKqvH+ya
+qikJL5ngHifRagSyNpkcFJ+xR0nsjhJr+06seR4C5a7IqZdeAICC2ipXVskACzY
+rB6fs1fL5MSK0LUnHBADaDPaadY/A7EhxQ0lzVb3AVWvmWBW/Zdi+4UienU9laE
XbFXuBYaQ3zLotuXWNM9ctNuFvSvdlWaJsBO2SAt+B+JRl4tEj108O6dAQ//cOVJ
I1R+Nk/CNoddzHvlNVVwuibWF4G2vLv1HRrT2LxlVZtGbwdGVpctU4ajyMTTRQEN
ohJOqv9eGNFFG1CGlCXUmJEPa4d5ItbrssQrKMPhSaE6v0m9Ztd0d8kpE2Uqc3Ia
L83upM2vKcH9vDoJjpvZuu/XQikWyfNoCRt5jDYkYDjnOUG4G5oFMGiQIqhkMWQ6
8eCGT1h7dRmzjv8MuHxnBk/2ae9qmm5GFmJB81GSui8aiEJLdYuuytUCLV6N5Twj
PaHWK2VoWZKF+62Xu9dYLxHclF+lf3DvxLtNF7p6FsBAOW+rbU/dJU8J1xxstlB5
tAX2j9ESDLyirhUwS6h611yQs+WpGM9nufJV5QDgWzxFw4jSBscYPLhBcTkbOVwk
14OLwXUESet66ZLrLsIyaFbctoIudKZwGxoVL8BZHzTvI8s7z9xgfBn8VBiFdwLU
mafmZh9mYdtwgKYd8LTSifLa+0ArAu6tZzAQtNvkANUd1fIGqxWjqj7tnoC39UtR
mS9OAoO+OkD1ijIn04RPSXmVU9grkdo2daSCPI4nHqsQgzVmekPzNLyqJo34W9iz
9ZSgDvHm8zXuxMpj02yNynnvNWMx47TnQKCRI/9xuQ/rY7cugXw2r1BieemvW3uo
vsboDVCKgFGnUSelSg0oYgZ9B0PCHuS0oeuISv1ZNj0w6G5LG4Tzu0ajDkbSkfkB
ODo4HQo156T6jFX4MPz6RpYCBR01NvuoZSrckLvcQXAyfJmTmfjEkP/xsaS4LT28
K/w2oApk4yYGmP5o8LllgI3j+0898QTqFfEMGB1u1bOymnPz2F6RHDzRAkO6USr0
RI7Nj9TnCd8aq9Mg+1qje0bJCgfUTy6UcPxp2tEBx9O6MtuL9LAVrSJizg6qjdLr
Sp77+PyRuj0+91Hxy3M5vy9UAMKuzrQ3LWwPP9amD511/9IsMcbx6jAytJMxxCEn
8Og7FX+oy5JnZQ7bqltQF3CJGkBZm9ZBa5QtIJByk14weoI3BqaqVAoUjfHU2TPR
Nc/6VpqMBAJ1Mj9OPwI6WOojG0HXAs2UnYrq/3615ZJqE5zIw6lvixBGqSRyGNMX
tm0lENxsbrk8Y++ejEiviKR2k/lPVB0Um3p+/6Li0FdLlpAOTcissn91hzPkjADH
kHwmeqd+SdWhyy/pVjiW1zmcO2CmrI2IWcjleIJZGPVcNyU9oSjYGg/x0UGhOkmv
dmFx+lZrWzbnckoh4ZqtpdVlpezwiiSglLB2Vf/ZCoRLvy5iBeudU2ZLagh5wB4h
fWDGW6p3qRMwvUX9/LicZYU41ri7S+gQk4+nYrbJs4oUglCSj7JSIwC2GNP4K4EK
RB9CdTl1hjrF3WWUk8Ynj0Nbl5/f2ZLPUnB3KxG6jF4cmtu2SB/WAl2yhoIxrdbM
TRgFzJBlBeOWvv2ge2F00YxPbJ21BQiWBVWozLmMjfD04AeV1N2MGkHklsT2UHBo
oFw/Y0QGcYFO9cF/Uvi91ywdftUYt+5BFHVGMPyzB2DLFGlwfGff00asS/rlxB/V
ug93azEv+96jIZEf7oxZonQIudFNHnrXop+UcV1GQ9dXJvNXOvGOx0CvG6mP52kA
ZEJaDR0ZwDNOraBvoYSH6aGDdusF9XTDVaPtC234tnsk8TNCc2nSXTxUhSOHb/BG
nhv9LWDY9WLYvSyOxa5i2pKkC2dMXhGQRVnUu7FUDgEZ9VbHLBN34xZzp3mj0Vo9
DFlJOzLCo4BsIdS+WbpJhzB00NBgh7JkKTjYNEmkPxqC4STQlAdpWtJ0/q/4XTX8
21Cnuc8KkskCT0+zQmrL8aqX71Ko8Dhyoi84WUT+b33KS4F+Wl07XayG9Fxsdinu
Roh6HZ6WBVQQTSo0Uolu+Dvef64TP91abMI3TEpaIopcsS9sV7uxA0AzQiKa6CAY
HUkgTdtOvcFoinNGt825gtHgN1UAwPFMe9e6jbZ8QMfH4iCNq2rFZI+h7mi3FpOl
0U8fLfGImgQ/O/AWYT36sOGXUlWhzNAJdvoxjm5heCbQTClfHoa6n1KUj6STqvZ1
KxpcQulmERS04aZ+LARbVZcgSb9Xax642ptINuIQmkOohLKHpbowhaB0rYod7LGz
K+ceCLpYDxSMtUFhlgFrOJfVaDFP26FF72k4QL6wJ9r3Ooxgk12HAxlae+zuQTI/
vL+CMsD7JgWgNQHG+2itxOaLlFuqoI9Jo91xwSFd+5Zw94D1Izd2SrK8OD2pSwwS
0udlyNgAAQHMXiOxxCmXkzM6TVtN9pinFxXmX8eS3eCA0vZ0qqLmpwi+ELR9nfc2
NVY5Of5bO6B809jVKbkLwHOVG85ofkoccReGhDq25HycABfuYjDkh0+ZVnjjKjzI
wQEDYPfLbE9WSrz8WnZ5x9g7WBD2wKasgYrP38P41J/hsYlTNUFaQIV53+Ew1qOr
pca6v73lMZFb31HSaqR3OvRHO69SD6aAojqIM6M1X6yAwcumzvlR47NO051lF4mt
vgrJZPTEJjvxrj6EywNLwJF2TOPAzAOmnmEJK5ykKXHfGb3JXRHE/TxWBJ5mp03g
Nje+bqKmT3PI9ELy3ueULq93wcc/4D6CG1twnMS3rqnCXRWi1rOzbn9EEWZmdFxk
5r+bJFPrEQtNDTM4AfM4F6fWg3IMbIRheXwWjq7wDVbrsmWEOG3UXF57uwIhNM3u
5Mq7fpNlJTg49TmPuYrbZUVCKSbMNjO6rQtdTrLRQ+mTR5mjkRVbwQQNOBPi5ZzM
GL+cVVU24uj1L3R0Qr4at/JLyXOKt4jAkkP/hLSzA4+lLXk8ygYO74BB7lwf5ngc
rxZA9T2MHrCe9SlTRnS/9UYh0in3Cys0PfO/eWMOyR2vyRWvo7YQkqn8zMcjf6i0
/jFS3MK3fhGssPeOuqm7F5Q53Q5WQpLGWTFhf29ytXHbEzBiuEmGqMj2fw95Zno6
HclAl2iPrVICGb+euUQCVwTLIzFULCqMKPJIdIyF4CMcv6rR4hBO44jZTbQcLzeV
GeMQwaiodRzEKA5ogVYG6GUlnQah2/VxHrfaC263o1PoSkrEuTDFc1AqU0h3ZOBt
2nhvCEPlIz/G7okNBeaz/N6N9XnsKsWyyk68zui75EClExgra+UJSfEe0iRruM14
2f9Al5rNKhAERGhLdafwyx2NNDbDnyDS4YkQwWX+44qjEsjfqO2GD1s26bHjyS83
PH6cvrZ9TMDkHrZjJbzFjv+1M6/RroeTIqNKmjBS6gkEKvbjTgtU20tKFQ9BpmjN
ZZQ7rV++VhihtVkmET/+KvfpTnE2VksWzIN4V5sXImoQUHuVP9e9nITBIxOWNg+E
tzAdN/KTozkyjFVDhJCnXXzRM2PXqR/5mCQ89G6Mbvq8uDbFLNBmGrFeQ9CrLtt+
1aV7qm7SxMkZ7FCzK5CWzNxN6VaNqUg26zOpwW2xbz0SXabSkXbSI0RPoqA+VAQ9
bkLSsN+HDoHHsLcenWHLDEChrLMqlfAXzsZpkeqohTAAz7il6Tzc8p6sR2UgljpY
PDsQV6M/M9r0u6JpEJLiUzYjYINq0vnwR0oJXV7lT85zOsSDHnDJLCCoxYgjFkE0
PtRRrc7P9mDB070GwuEV9f2e7LyoBykCgMZvIesLCi2JcTlNOoDG130UwUGOOGC9
rdWqzlKr1j4qyu3vUo6yr4tYJr73k6Ts9koEXAF2ELBBeeQDM18YsBoa4W2ymL3r
vZq1wpkscJ5m1eitL0AdYbun1TjpjLZXyNCeS4WJ0I3Wu48vWW1ru6h1FAryrjXL
JIgbCEw9ifSsqfSYHE1GUE5O1bkT+eYwVmy3L8ZOXVihIKpykBzxBLLzP+toSHrm
xXhXaM5JypGmlhV4wYPh4LhiO7ZfPMY1+yUH5jxKLDaQ2FBAeRfc2W45gjLLJYY2
1liTSZPD1sWnnRQ2TCy1pDkcbw0Gh/SO8/9epfsdvWIbN/Nsin2oMadsimIwvoBZ
1Q4+4miCGYsoEsi7m0FTq56SLSNBgcDlbrBoM2DDaS8CcsgLy9jKYdNOqSsD/Q/U
Mq/h9EA0S3imMWoMxOlqPjygRNnFsEPUniba9ezSSCF+yQy7YVbWt0ZPFAGb99kI
yXi1GWN01zZRYWMS8+g8unKIcEYZjrC9UlAt7FF+ZgTDNEGn2oKAAS1y5SFN+oXe
gRbtqrwBBTxGzNgV2f6TpTu5P2CxUOAH+F11Mt34K5S1TUfZ+oVAHlwZATBX9uey
g1xhVzqy8L4zI1apchfJCSHBkAwSZ9uKDJh8VYDQqUgIV7Z8k5Unqeb7LZFLUNTJ
+9z+bk1n8EBf0JY+KlA0c+qZPj01lwFTRMyUjs9xl4OdlR7XsUFKLAtcnLBiT3NW
KoPQiIZ2eyq9C31uUj3GFTsuamSyw1Fy9gTR35ITNz0jMxDH+XYavLRYvIeh80y+
+YmfegQREo8RC/Y4aPJaRjcpDyFCxh/ywu7zNnQB7ldBKb/qtp4nB+fYPOQ/0q1u
BE0gtd005x7ftAILJbJd1UixTlOASpskhveQ7e4FixYfFkopv7H1+jR4ITMWvmdX
7g5UH8OLNeiKjlASLB3NhmdpkAO8px33JkllG5CyiIko5UY/l63+G1IN/TIQANsb
xAP1dkL2dsHP7Fn4nqhF7+PT/eYGIKJ5CF+RTuLYyQvbNl8WTnQYBZLBtSQUTkEy
9rJHqJ0y4QfYYYAUGEBUCNhT42nmDjqrAspuRTcDMmcXxo2SqHGw8ou4TBn+xyPf
yavNLknvMIBVmiNh92sm4nVDbEobPLmwmUkpv0YnF48C86OUomqiLo2bx1YnypIA
SgRasTMSeBTHN83xySLenfYvpv/fDNmZHyPS5l3L3l4A+CQGGdNvxNh1j3pMSntm
1+IKEBP8tqc8SgxxEocwK7H62vunUpsacVZuYx15AOIV1vhSwb333erKJ1jaOONP
bRbrAwUJ/Z+xsdKMsDEDB5HV1i4094/DApsE7FKBHAeFPaYwD6zT3ZzCc+kPqn+v
1ZPqeKeYloE39z2RjmDp9G4N/6kOKu3zpmX5pdnkARVtn1Upft6fxA7Rql3Wd4f2
gOhJi1U1qwI5jMlwuCywTdPLkgOmz+oef65+MwGvyIVlgwN/mMO2AkcyS8UhUC3G
tVEL+fjYMh++t/3C5tZlgPyJMdwmZ6ZpZULVIkQeBJwLaQGv8zcvPhh0hlcmawwN
nzFgvkTC4tyn0ZqaRS6YiZljmKpZ/GmpX8eDbkNyebILTyGiZ22LziozzHd2LRMI
0DbSR8DcMWSihGhBKAGleu5f8eyTT3A33gBvAk5JLz+f22DDninKP6Ou291WaJ5W
HWXcWU+r3k+S0P/TYxAWv2wIibMbSkXh15pAr72cR3E7XM6imnOwpeC0C3GOWg+B
oqkNtB4mIwITo4HvKNb+Lb+icL6nMIJRWs7SGKVozff+PVA5oPzJaXiIui/Y6BpT
+/o5/FaAxeywERZknFyI24va5on/u41YqfBj1MGSev3lVdt8s32G4GXJ0YG/0m2C
0DItVSha2Yaqbmttirca1gM0YbUEr0aHlj5fdPgYfqo5QMvOOx1/lmKW1M1hIG1N
xoYP7YJ8gf+iBTkOTLqQ77/gfOasfKeKk8KJadqnbQv0ZuWtQNl3CgTc6YNYfRKM
O3WL75hp3IQxm+NKg//wQzh0CH0dNZbsVpu65qAjYNEoaeO4d4DkPih/zsYW1YR1
8/4oY+uEEXmic53MwbxNcJXMQzW2jj6vNdascKJcebjzGwKCr9IhUUgMH+cQ4y9B
MsU49GG/B3KX9iGAd3Sh4IDiyGo7cPWlSCYR2jPaRHhX3B9TwxaNzObcmPC7eGU9
wji5VVT7vmmDLQ+uk6SCLns6DXBdaN7tGz+b1CozbSckBjiatvMsyyu7DJTGmpPu
QGCk2078W9WezcLceLxZc/MCXM1KpT6Sn9fBPuCU5bVxUIuncO0P0+icRoUDGxjW
uP8eN1Aj4q+gwDA1MceeIT0YFZVArzrdXNCDYWRRpR5oqB2RLT31P2s/HNXckPjd
wS1f9y0O3/ebYKMm2ixnxRwbNrUe56yvai4vmAO8sf5JdT4T57Xq+23hi7BLCUit
2cVJc8QIeCi0tLaC/JrP0fuuWazFqylNZ5EaOFJw5cv9Oq72A0nrCj4yd1iIbAxu
Ma7ftx0Q8VLdjKgy/aApC5Xrxxqjk9eEw0bZX+XV+jlnC+4FyEJkDJA+WSQ89pCP
/c3i5VzAyH/lKVhk8pg7ds6TbbgCgoosO9/pQbHseg83eX6WUGfpk4nRb2kdWTWv
ByrJTdXy71y68tzcOCL52TSuZCzJyuZyyIR+aRbWL9mZA6g64IuC8m1cBvIbzSt7
rSYpHe/rAbQCLlK+4lQrQPoqF59sO7dgcNXutCOEoRrm5E8oHU3FwpTPQ0Ad+F/a
NmahUGJ9v9J9icFn/xR/TOTHh3IhhsyW9p456UPBtd5uJ0IomJyckcuznScDj/sQ
6ZX+35msjOHuyVSBynlkahs2aTOLQK2PNQ7LF73E2l+4YBTNqleEC2v+WR6+VNd1
/sfe1m923+JCxA2ZGtYT+jvQR3U8f76mlmY76PRiGJzBHWnEE5FXsfHgIHBusjeM
s2QU5KN22xf0XbJVJ0U1DtUbFBgsdE/2Xvw+1aBbG9E2W0uPHapjwDJhDuQC3EqZ
/0idYAtlV6Bkc4Td4V1KpFSjD7pGfrVBqTu6djmTj+iq75i02OUAgVRzcgAX1UA6
e5o/K9c/cvLudb4a4Rob4IoUkuPyt74PMvSZPmPP0Trd8XKXFGFb7gXUsUmYbeW/
AVanrgqu8ncogmFicp4Y+TzUSsBOStpeVl2OmcvOG6Majbb0vsSrPCSCpi05vhZu
xDQScYufuZbsvx/NaA/2lXYFvergG/DEec6lB4M9RfG2D8HVBdlOdrF8kThGOD5s
/gu+3TdEfeTEZiucvBoKV/mmKzrefZv6XUYJpdAztoCmXS5lvM95BZv7g+79qylq
OCv42IBH4Y3ZoQZWmucux6Gyb1v5bE1mQwfxhfGoZ63igmx4O0OswBWmk2h5e6pi
DKmsAyKQ1Xxu8ZxbLbX1SsheJ3+UhjwXSQSVh7Ndk0f8vyTjOMLyv0ePpp/FZKNT
COeYkpCKcEu7vhcOfluG4pJoqvt6Vwc5oTWaojnuUNjbQqp2YLA+i64nuyv3EQkO
mSU3wY2Gi5AssHdIIwGADGHLnKnVxYq3Ik4kq8sWzsRJ7ULjRsqtBpm39ouT3gKh
mmQjMHhsRYVZLkUBbiIqJ5PRe2Rtkvf4VjSu4Ile1i4fkiI0X/yc9Eovy2kvWE7Q
J9TcZUhbWCvwXV2iFozL2PBBUoC6uxsZsrjgG38D/q1nAqCvO+hJHPkaz2dui4rf
MH/Hq3nKV65swmU7ViF4qMTreE5yYLSmNJ/55ksOQh+8dCK3vHNuSDJHa1aPgqSW
rr3qNe0Yq5jRjIoUj1oHHLMI1Wl22BMbVwy0bpBjzpEl2FMbHAoda1Ocuo4DUjvI
Hr7ev4fwMQJsyH05L7zIQtLWnBBjsjulNYhjk5sTtuqTKMHGwNfVeArZVlIJ8GZ5
1CbzkGnTYBUqeULReqjKFLY/YcGgrtI+RsskBOfXRS1VDGu6bNsNUYjb/kvjvQCf
x67/f8ZmnUuGptyZ8c+HaX3TJc/FDe2Gwbc70sD7ArtoHEVr6o7bXZUtaWRwpjbd
c2/JxAPJru9LHxlZITbCSSoprUnNCJa+7kGk8cD6Fc+gGJRRhEkR/h6lq3YwhxS2
Naa4J07tJ5JfoT3p42cpL66HJqMNyLRQVcDAWJEk1yD6a8+3O18As3P8IyO21xXP
ULB6K+egpOB9vchaOU18aDwZTySnBNGSbdW6IWwqAT2J6mt37lxG7kCyPWOEUDPc
BgnIOwsGh2oq7X/xxiJuvP6ImJ90ibzbUvNvlOzj/eqRNqAifeP0agNkCf8xkV7+
h42GnBTqA32NCFu4qbDpKF8hPXhEagsQ/89oKxEeEyJQZxMVS/J/TrJ0CL+IySoZ
8uUWCKyuH9BRC/X1bu0MWeTf9Wo/3BdS2X6BPVGR4GzU469RVs85GtFn89qttufP
yKDSa75YZiBa476GDqvMAVtNvFPUkSBNMo/8cecwKPCMeLJXwTriu7srD5yQuYJO
++WmyuCISB5JBauNcO3BuXORlOGgRZq1SlmoL3GrBIHmDzUIXCiG2LMAzHdN+/6I
lsCnR+Tyqmf15RX6kEFNHXPFNVxR9qPhhwn62zwK3E2bdFyHJNjPc5UoR3M0UIrh
eCIpKtjkq5lq3AWaAEfwvMsfdwldwhe36gMFI5A+jPgIB3bslGEoPkwnuOkAuaxa
zFyoVdvpOpK4Fo6pBDp3GTZu3j6kxRA40u2OEN2si+XkD5IDbNJquZXE5Uhzx9O7
/smKX9+Td7Zl+vcn2+CMd9vtxq2dJstzsJNd8aL8t29MV7b32c8MijQoIwtyUlwO
dX1+OzDiVCkoqdjy9gufkLv7IPyxeCLhHNxzgI83b7mLEI6zC+im9CCJ1Q30n1/X
+bxkuW55YS5G7PgMTS4vw7iDIa2dhgd3T7QhxC6RNFr6FCEtTO+RZ/788mfuHRSZ
n/XOBrUev5Ywdfq/ioObyvNtZFq7z+axF9M+CbNp2Q7uzuPCo09k6GYvX3u/7cyu
ml+ueoZuua+Wb6UXrI8n6yxpEc8NgWeyU1rSbMoHwE+0rNzWQmxxambwKl7tg0O+
GIZsYA3Ky215r1S8iSgDuCaFWE771b3X7TUkij430zdTlSnEJNFmufiuq/1c0mpX
nctnmv7Rq1gBFsObzXTdTuvOxzmEI5bfEvSLdDkahjOhv8GQc0/exMG0QaN2/YqU
qCVyB9gy6Og/pWtAMbjAjFBFI2Dmta49+Sy0UT636r3yJNsXuhwBmt/rr+Z32QvU
62K4zBE9aC07T+jVVqrbMMEDDs1Te6xtqind3rvgFhxad5LjE/ybo2COokAACkMz
iOM5UroxKwa/13/P774S5eeMkh/cOtnTesrd+I7LdtRtonZxwd7B+AIpyjPO9ae6
kY6qLUB3OVdtBaEAXtgCEKoJi9y0s8GOqT08R2UHNtWc8bcWNr29Ubz6+a/MH6Jn
WMVHTWF/F3xxgA4IvVskLTAa3y/BpZ9itWSfB3YmfBjt6TwB9jI1WcAxhhXJOU4U
eCBO/hw4/XI8CuLNFInHlhc8C4UiYunrkNT0S2dRY0ar8StL+qknz5MNe0kuyT1D
ewaWlYOzZn1WeNaN0Ww9DRP8p3XgmYxXZgu61wakj0Xku9ubYt9pNJuwWPDZ1Z6I
mdPxNBoX0vXBlMro5LTSFoqefBT907ZGvVQmQdEIXtzWiikJeoq6LrYsnms3nGT4
1+YoPiLElkM4ejEotfhA7AS8ClEEzy0WYUJBTUaCFOpX4rwiSmlokPD0f5Vjec7g
DrIGZgCAd9A/+Peb3suMah+8ADU3ahPOk26tnuemG73vCJkLvzST73ph5eJnK6M5
qjNM/KF/rjNhK/NXANDKUVqOOA9Mh7Xm79gNOAJJ5fQ5HHBM4jfqpuZdfCuYTAsY
4UBVTBfiW+SeWzWtulSsPAHNzYmyGy4P/wMcJJeGCTyKYWf5DycrttjkGtRebEa4
uVOvs68VB6KSacbSQHVs/RCE6cuAsH+3hjxEvJaRffoxnCO7XoOwZSJmok5nui55
bpCK4Hz9HEufoajj8tAqyIpQS7uxsavLvSoX8eo/+7FY2zA/Y5PLAsV0J08n/54J
AzAYLv2K9aF7DNBrdUwJBJKV0p+/IFyifEOjimhLtbEXWwxFQNAAyhFPCbFKXNoS
W5EKqtIYnL4lCxPQdpbXqmKubwOXE5qYJBymyJJqfSqzeVZ3oMc5rsjAga2oBN2s
LE63LziueITDqiUM1a+X9uONKa7k0GuzSfBzTfrKglXcgQ2oDTAQmZNC/4Nk9Qhf
8CY5S8tlgfV1U/IxP9ULKX+fKbgo13cQEykPizVcCrE8IaWqPu2DmbQT2VGztJoU
xGfauTQgg40NDEJjV1iLf/2Oepa9Geul4RxV/tI3IN+me/gx8MeBrQewXnEJGiyo
MZGqnVuxAGqXW7SGwLVIuIMaYiE1QtLt5Qc/2OOytpB3RDdNhj7VOZdAslNF4UO2
YSr2YdYyVNmPiYlW87pzC0t/gRAoU8fdi4NscsANfPoLjf9AUzDTrPdxAuW+4uRM
P9WJ5wJQfO/d/SN1mswGBpIVU7wmof4HxXrX1RkDHJHt2AzbSM6jBfblhesym6XH
X0VzBzNJgQoIKw1hgB+p+5dyYtzVFDTnszYzLvk5zDtqHAnxfz9RPZQuk28Msg8g
bP+K7qM7uZegOgN1C4QayxcYnDfo1b8odRIEg+fLPvk2B3IaI2PDxNOBW0xyc4pe
8sL5GszArk2AAcQYKiKVmbhvFFI34N44Ztl7hR7nfVk7xMdWzGCxXFILatVGgJ5p
pwi6mE/0fpBvzuTMVuvB1axKljbiS446JTCsC4B4RNmldTBcgWvHr9R9jmsRGwD/
/7Qhf90G20cv3kqlpH3mJPen2XGm0QTlu5EuOuC51qVUaOqB2ENeRXin8TwCFSMw
QnkDjziiAmgGV5s4PR7BUJF1TzmGzFsioIBIspLa8/kTz/c14vNZESTSqxyg+aAk
Xa+7pEUY0wyCbfaJWtw3zHTNR52dKA+7xj3/eTHJ6kIQwN//mgNIWHTLb3TkC+yY
b57QP1JkMUjAGdfZ1o8A/Tv6z0i6gx8qC+MLbgLOKnBJmT14ugXk6JU99jWjgcdY
56Uy+CGOYSEuzjj1zKDRFzznxnORsPnjVVWFE/AesAebR/vs7qDgytyWG13YYxPO
E7qU28eoDHqyPVzN4Kc0mtKg4IVC7R2QVCy+j9m19hAgazEYzIbgrYMLMNeTuiDV
AlEPmBdgrbVLV2Ep2OE+WkqqPy/Ox3ZtJxs3Xgj7qMnSSbaWzME/mbxHleFudwms
unawqRYLrOKRpqzmvEgsybTks0p5JfvXsrPUYqtjtAh93O2BwtmX2n2032zxCbtO
90u5VmF3dtJECxRgTOWzq91kMwC624dZBvRLs3extvCQ4Il772vZjRt1Dp1y6NEF
2QUxAOMADuz3KaT84TxwDE1bNTXpVlP8LN15JQqyOGHjcrkGwnv+7Rfd3LJLgzkx
aIjptdAL9devNGu3pQkaAC4LlEvzNHR0wAuSu8DesNECTbycUgNV6CScyzE8M49e
sZQC/wRqvGsXDPzNTq+my+5c8Er2U0NBwFKtA4U/owhPg8nweAy4BnYb+GfMo8dm
2icFNjiF+NDjoEzY4APZGfCRK9lDmB/sYaZXyCRJ23sUbZk7V/aOVIBbn8M4g3dQ
Toabn5XpImFkdK5m242ZAHgRNUuWF6sb3pmb9U95vztVoTZAMzBAZYnCOGCCX4+W
xbvKU/QqJ2UvSYClYQC6Qbly5aH3fI+F4+GPvcBpj09Qy+/EockSd5I5gigzT2sR
ktM9CuQsKbTEMxD/AXC65cQkJE6aREZovvGvRWhs92W7xg1ix9yF3n8IBYCv8qBu
tVPzH30VQlx89LUW+iz1rNWnInbtTQyGVNmbALxs/q765gtTcpW45qozwQu8pgMT
hTBBhkroa20sL0h0jkZ+AOQTy2J1WWJU9szI23UDgqpr5ngC239FjY+r8aPnmiyp
u39Mar1jenm/AcUznkKK6lua0TN0FbvzAWI1qwzzK8Ur/DBocoyWZsHiAK9rkKvG
1K08umH99injyOz39X5Vq3yNSpnHVIVIJuYgzvoftSc1k7x/kW5nUOIPxI0alRlG
SExl/3+g/3rEfT1fSYKkoytQ31vR7Q9S0aQgPCq7BOzaKwru6+EbujRhQ4FN52vu
qMRQ+F4et2TIvKjuKaJtlomEXQvRyBu/mrNMzwyPhci/1cR/l9YkYFJXCyI8y7ZH
50h7j+AIXAu/0clMjnZ4mt0nv5bk56z5SpIDRgKy1wbmadl+/uVGdQ6+lTuAxoQ/
RmjByvaP3eX2H2ZbE2hO1Qab9j09+/cYwDZNZkhsLSyOGW949YkQMvuBffNHejcc
UvyHVKUfYj3f1Refz0sI2LUWmQJqtVKfOeF2m4+mJmUyX3MAxc6q0+ntrkqxEko6
k2si+swIyUOC7+IErMylG2oLltLddi6/ICmQzAiwqCk9Ixq2oManfW75VxFpJrdW
aReq12q4ocQ5ICptvEgJMHvQsaK7litAUQ+HBA4U9oxEa+Kpogdy06HruVRt3pEP
1u6nLf7VokaR5mLKtLZq67kmZYAJeiBxH6vq7PczDzdnE6BenPpXxhQSuN8DYkRe
kS0E++PijufvK5auovftiLlBx0ui27CoipS3zdhXqIRR3UWZzD3a3S6h/JIFePqI
6a4kkGVss82F4mX3d1J/XU0EQrJnpgjIYDf7QxlTO35/Zs5+cu3I7/ctRw1oGjR1
RSDlSNIIVEItuRVUvr5dOw823lRbHBb4ozdV75hZW9jsMEdvao5iVwoO02p6+IBr
ej7B14wUN3JGaaMlDL8j89grtS36SX0+jhhPQ2NszrV92adT9QZgUWhzahwwcDd9
xiMJpDXhnA5uTV3zUWoR2OHK8+MeID5qip/+ftfQ2azSy0Z4kSdlhZFZBI5WIFG/
uL2v6wbFjjtINiLzLbawpgX/fIIytw05uQEdKzKtYn51al1U0Af69tkzEyk2QHW+
lYrVr5aBTvxSnYoqIkG1fwOWneX/cwS4SDQTHrxbGz6iviG9F+J3198kBVSlkbwq
ZPHuEv28kKNztIF5x7MmWKs5lyZvBt+fex3tI94rYIYtBRPEj0Bxw5p7L6xU3xdC
EOF9R1REyBgljM/QjnIk7njCJjkByhWwuBkdYf9BQmvjyb0CTKve7GiP2uH1aSuB
CpYy7/Cvpo+dwAd4wWel5TXYKYlFtz5ZIQYRx/RtGl7gBg2qS+P9+h6ocuTQI1NK
9B4wIYD8ELomMhUm1lfpfcpy5H03zvvz0ayMtojCBg/GehL3MgQVjcO4OHPL8llx
+/Cm15hhj6C+3AhoxFlJZo54I8nW4SXiBkSC1vDrRV0ePXG2YJEu6uGIDoCEAqn+
GCHXEVg0Y9Q8zgk/XyDdNcc9OlLS1XFuXPGY/IEtz9n0sBvF1qOebapDdMf1goev
6Y/FuFNGTZePLj154KgD8VFU0TyhwDlVJM2fGOu6dt9aoDpZ/JH//RI5KreJFlCq
oJcpkQVmDWklMp18LlF6JIA1UqHqwj4SM6YmLJCGAR4Azb0DFlnVd3gBWQw6cV0B
6C0InVCqa3213lEqDW1DT+0W5OsyL8q4taVdNgXMlS+SDyRYUhke0JivEmn7GJM4
O8k1XOoQvY3BhZi8BA6roLWWqLGzzVRptqLCmBygVuaK571P9uhweuXUJUsiKmm4
ToH4lNtF87UIHUz7ZxCe5wHwl1hV/qpNnNPSiUAjJtrV+Y95GCejjUaDTwBb7zCi
VWfUzc/CMLSqR3S8lveAOrz4J5TAf9w2fr1b2JyT9aamsFFB9jPmL5QDqghz7RwX
D/aXt10aNq93ZOVMGDEaEptlwSv8KkaqjRS7m7QUIvr+5iqRhgU2e68cVVo9bHKd
MFItm060+UIYLrUAqNteXnRqYO59bJvO6e6gLVQeKvN2pMWUy6p+Gh8wpFqR+kgH
3GpPUQtiwq4APBvY6VKA6BfGRn9xDPc2CjfUIExVR6oG46rolXQLeU22ox6Pbaax
TQu6QsLylKWGzmJNqLggRqQuZMh2XxmFHJF5+U2M15SmSutqQhLVAAmfUOprfKsE
`protect END_PROTECTED
