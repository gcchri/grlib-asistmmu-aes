`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SgraBeXbZ23lo5rUm++kdVTU46ugKF9Nh59fARJZXpLlOxXzJGnSGe5hNLJL7D0X
pL5m+cZs33ikux5euoP/8CdkCfqlet8VYMByi5CAcMxnqVjvaJ+Erb/2pyAbvIT6
fRRQ2pE67ycjYz3k5ZL9s/aSEK4inIehk8NQW6sqiuZrq8Zx9RiMJUtfgRJ+P1CY
za48dCHyH5VgzvSu/9h94K85/BoMfAjV7MmKPa7mJy8HLMlDDUOkORJC5HWYqjf0
7Pbj/92CM9W59S3RiriuVKGm+3Mi64Bf2WuDQd5df42eDKSZh5OxZ90KFy3m6xBp
V4km3JrqVNMvshFtLHPAigzgQhtJFZDdin55q/uRqLfbsybszsX+bmXH/KGv4NgB
WOBBk+iQQAV5ZEDGjmefSXYZ8eK6IP3rnjRXLt2M/RScdNyLGA3PtiuNVMA20Ssa
j6pOtp5n5wCNam5Bp64DPj9HFNCCVepGcgnW+yBVe6/yo3Wm628jd0tU++7cWRKp
VSVsBO7PvOH3sl7lHV2k3aEKUa9MU/U2Sjurrpq7AO4=
`protect END_PROTECTED
