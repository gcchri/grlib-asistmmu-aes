`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NvwHDEkH0IHdyMGlTZk/gEscvE7sRWwbdL8QuckmtInWA9AKATOa9nDj24k5hA2O
TYn6o4PeTVXd5xtxrN8n7b5LgmC42Hi2k8WZmtqkc0gLhjVkemHK+vCMWlnsIsbj
FobMQy98d/HoehQIbbyBrx37QXyXiT09STdjzGUBxerltSmmRyzx62L04Nr+e3wG
5zepnTylih3VxQoo7HbSfIFWH1NrQhJZgUTymA9JS+poY2UzgaJh5ww9FLoLeGT3
JPkaToNLQgtRR+h33mTuOr87rsToT8szilUfCWCaJe66s8pT8HwHuQhhjEGn5xVP
gjK1LMCW7qRISdfPttZ5K9P2SBHeEbht7PoHzYZcMcmHRYRNbLwGSTfZjoFljYwJ
gIv72qaIWE2r/gkIbUc7RJPLktW2ZJShbz89DpdEUEFcEQrd8glopvaLvqZ6VW0u
gc9TYLWJOf9JmUg71JBB0k4+vHHDL7u1iPnBoFgna4RyXXQVtD7IAb6KNzEGbDnN
vCppJaXnxwPynLEktR2BOteqGO+N2IO3JqkzOSbtlojSPV9ZQGJvCBgyEF1Dc25w
g4IryHJWSEfiOVMRHlIj5FiDXSwqBuOoe6bTy4WJ16SW7mVrmoP4DveuQ8s1snz0
FYOTAX7GyvwgJH9HTPbbqQ==
`protect END_PROTECTED
