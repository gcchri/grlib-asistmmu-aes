`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V0QdOtNFE11Eg2KaAnippBj2Thw8kFpZ/FXC59EVV/rrsRaQnL6fcF/B62WH2DQ6
RVo89ZNHWGO1vocN7JyI3kR0FUtwlvjhscX7xr/Wdl1872c6bVPwmjGo3IB3pMwN
U6X3SHCk2OrU8VENqlGM2r1h22Pr/IpDuZtcvhN0VQLtculJDl8vDQhYmxOlImnx
Zo86iS9iTTJJbRPZJxJvteu6kKUaLU5mwudADK7rBsRGn4n1JWbvugqgWFRKMZET
bWXPakx7qKdiFkQCU0UxgLIfUhGe2pkZtiDZwlZF/T9NG+CaJpJ3CPTBnts8OHn/
zkIj8ogcNbpM88hhOs1ibCR9bGoXX7Maoa3GzDPEwfPRaHrKGjiAdJGV9vqpJT0Y
6gQXMKGbgjlL35fuwO2N+HxXA57fZKH7GF5Gex5Tq+S85jmBIm9c3C27Xxl5Tv5X
h3BDmXOfe2hbSoJ//5kZcVVCtH1dxYKw2m3jPC+/y36RXksXpkICWhUd0d/T6F6T
6vaG/zGKNxsYGFakEYHpGGakh6la2RZpF/yW2RbgOwYMCEDZu4Ocrp8F92/WfOiM
qUfLpvXrMS2hrDenb/PkIOOTLHxJ5ujbqSDce9KpKA7K1XKvEeyUH+eq2C4fi2U7
mpToXxAw5Fs8oN8GMcjf46wPXj0EhjngtEMbkvt3U+XJsOqyqbZqsfwMgC76233E
ywmILjwsiA6YSCWOzGRyY/ZalzTmsr3pMHDBmptb70h19QY+eDakv86tOfmYaRa7
oK5T8DwKKWaAjkpjDmDu/g==
`protect END_PROTECTED
