`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T+dl16yQ3Jzz3yCQIct87nDnDWl5Rpqc13lsX8IrwJRawEvgb6r5xb4jofvKxG99
tO6IjLkZUzcbmhizJjgGFxhP62GWLQL71Bs96ARKmQ2rlZRRxqVPj1Hy2xb2MSGQ
dU8Jj/vlKgEzHP96V/6w2kR/o1emMZTRrWLlPDGbBpF9g+Vs0v3xY5nAXlViGS4T
QxlrVVyGjOJaRXvWHEViTBPHbL1fMj3VlrflHbZWfd5bhtgm+X1T2qa5zfdgpKNC
3O6kFoRpqczju0CHZTLIVq27k4MeWls94hd6pTTdPxMAiJuCgV6rLe5dCfj/htWl
epcmd5l3xto2Youmw26c35hpQ0L18VPALknob8Qa7LmST8lnQv2yp4R7scT9vpBQ
Smf0qEjS2t86+u8jSbm/K3AUX6ORN64kivVc4VPOTDJ5JwrrwLW+qtTS1HAia4GX
xlbQqWI4TXYChuRw6ou2Q9F4Il7XeNJnAdOf+xnvYc4teZ5VgEWiy7/eZKL+dhlH
Mq6OxfLlFJSrQJVK7i8MYCGnd6SowR1Zq7VfBow5KI8guHZi+pFqUN3ODoznWIkr
N7Wz6DxfMSdJGwOZAkpVgBYgOLttpuQjhehmEhJi4tODignB37OftSI+c1QN+DDu
Tfkxf4+hgU0NumC/4VndMw==
`protect END_PROTECTED
