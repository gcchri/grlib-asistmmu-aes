`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gNAfsK+v2wFTnnQRst+dbc69jN6YK6wuxWhGIreTh1dqD1ebJ7TJaca7RaLxjH1T
jFydDqfPGWo0Nb9whxruQ+yW7VEOhTR1fgdCaHhPfn+o3+Y9aXRWFDNUCbDB2xEl
KYjX2oTMomyg6XihFlY+wNUSO2YW6RfVipD9cR8G0xGVUisZ4SB6UYZOxXmmTsiT
NgdNcnq/qoGA4eSUAdxJvAUdhKNP9PLwS+9RCylOnI0SMN93Qb62jBruGr+Sdclt
QimwuPdUfVCQO5zZZf05yf7RY3WIE9Ww5WU9zOWTKTnQNhIyPbS9DVQnyOTqJfsG
GYCCf5BAJ4Z0cE3+OZBeU5xIl54lS1wCPSorDvu7WQaBuWYa215+lpP1HTT5TX5s
X4kkOo0NSbhq1D/wgRxux1mvxRKQmxojavpbnCRbecqm0QVuMEgo3TLrpZOxFSGM
vwnDfU2Gi5yH5kr7E64wdqMYZYPSBMnGy9eCVyNtB5+YOwCz7VJIsD94CxF80rt7
v8oCUEXsiq8t/LNisHREy2hB+JyrurtUvWx2F0pMxQaIJi+Rn+tbNliRXqFqJxyI
RGmGhtqOCe//o7sId4M9qK9WJSYsnvnruZ+nvW+D7YjoJ6IpwVxuO8Bnf/OiJa0c
hh06AkCirdUNI+pN02LMQtKBa3IbqxFqCFsF5k//bIA36drZcyzFp1utlZecrxV2
nGPezSuYFT+owQZmYnP66Ax6QZf03srfEbZnd+MQ0NNnn2P1ArGBM1LSYOGiUFTD
KzKK0UBXXKG4d73sinmasvGCYMxQ2qguTwDt2XgOUj/9BbLuwpsXeLU7FHeVjFa+
pdgoqqW/OrU39R1AgChV2Cfy9/SNEG21fCFz3sXeFvCrpgev3CVkTWrIIqFPUvnK
EGwHrI4sGRhoNAw2B1imaiKnrSSGZiL68nZukZGaz1abYAFqdq2wW+QpBSR69lcK
spVv4bH7sOMbpboFWKDW0c7v8ieCETGy6OHRUcpoBZP0nwtm0Yw1NjPjBmv/RJYF
oTDxQgHXfDrciOM976BkWfAZ9nqSE2jqYI/DZWei5GVDLIF4bEn8ImXrzVYtzZv5
31eSipcV0Xppolu881rofQgzh0j8n7rj1F07e2NKrLO/HxSpo0UuWTqWgtpQiVrm
vgsnbVBFP7eeXNCj9c98q4qg0LSHAKzDdLKaPb7YoFoDcy1oRLZLMzkFvi0UEfGx
gpxfy8i0euSQh57hKqYOaAq/6OUNYjZtFp/ikOTQIKWQRiGAKWAks3XS9CiC7KuW
bGy4FOT+MT2ZHcCTsTH6bITK3QjIA8cFfy8TgJYzjnwuAUssu4ipLoHdQKZFZ2ag
Q0tj3zd+nVuBUxDVx6s4fND724S0Y6kGzArvlzePR7XB93KmOLvYzwuvTZG8FPG0
VsJQrY2WRW8W9aZ3piVqSxSns7s2F5tXE3vYDRUEvgfJ6XNg97BqldfpPRpKXXQf
gANdpi49TmoXam+sFqIoRJYNzxUs52WsYie3Lh8rJQI8gSBFi+CynXBKqMU0QF1w
MpqtnBD2zwGlt6k4KIRAKi8izIV7HTtID7RENBiHj0/EdxRg42B0hL+zxjXbwpbo
VfOrmc+FMT4AWlbhOdOx55CsacpawcTmiu6wQknuHDhIw8vGNCSDQfnpN7D9t08j
aN5IItdu2O19DgkpJCGOjdK7DVH691cd00PVAjoqdM7tNnW9RrZ60fgeQe+u3yYr
u+qY/CP9h+vl1d5lJ6hgvExvcdD29XK1rHvo0y3orFn+Ck9w4bbAIF/8CesrGq3S
12W9yyRSjGJuMOsi70mZQtpDcEPHhZQjOc4MOsrYleBYFCcIk1xoQI/HfN4sygrG
Sm0XQBweOdkdg2CH1vctqIjn7ThGl+Wuj+wWvb7NPJ+mJHOW3vBWrh4sfGzpXJlc
6gPRLuL4cCQ9INTIMHPKxtKP1kMyTM9DsxzkDfi1EsMmvXkKIYEhk8w0o4pf4wgY
KpWODnRTpzwpJ+oQkVZlPpAWIpd+x1kaduvfWJhB7TwsHf6N40o0KPjH9XdCnUVj
Uyki3NagUdN/ZFtsIcAjmCQAVaA75ERtNk5QTqDrF/7Zmzg6SxStuu0zP0aeXvIt
0jDSG+NeAQjVPfJXBZMfq/JVkVl4Ey5dG2EYF9Y4kbn9SaUrV0ls0p5RAavCkyRe
9pC/wtWKKyerkQR+SZ99LPV8iFKvbqHpPygtW4ScP8L4k5lc3jQ1hqH6LTHTZbgE
`protect END_PROTECTED
