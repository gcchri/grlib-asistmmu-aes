`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nQ5Gv3WG0GuekOATZOyGK0/YJlSO3SkFUJF3Eg9EDO7w99tBZSSo6CFeWfbDLZB5
L5lQNmatghdE/Nf2Q88q9XC2UJiI8ngeKS0i9CVMaBcPFOKfpThlyy4S1TnTrbgU
5nvUfzjm9605vSouAMy8RQk78/efnKIXwXyN8YpgNR+HxGHfXgqtVXlymAUXhSCI
jDuzEKrq/2CIiDcSCj0os2VFlF8I3ANKnTCBiq+F2fzC4leLsUpaX66rBcHOCjXn
Htgr0IHiH0bMuR6zcr2N9BPlk7ylkeCbSUkrrIKXmXVQN73LZ35WZ2oCeEI/9IW/
4SJRCK0+SRrdPO8ric4zwqmsmZph5UGaHpGchcE4JrNZ2f/h3Sruw41bzOfpq9RD
6OQmPgIcC7HuWIgO1Kf+iyVbbVlE8+RlHA8Zd8LZvEO0yNLkQzabIBNzkFv0PAL2
3gfd1uIUJAuanwRo2AjmtQp0QlGuY6oLbuxedWKAxvhX+8rwbb37oaZFTmUxprUP
pZHQNwg8o3Qn0PZyGYZNimUj49t2njv4sL0zsJklZaak7k0XZb5QlgIDrfCNeovR
dtjnA7UGLDSrkF1LpP4vJSKSJzTbsBUfQoHB0Shg7WxhYe7pmMxswgLDEBaOk1nJ
565Q4dVr9Bsx20zwskRu2Tq1DBsChsxsu9/PA9wubXRq/LYjhux5l24TqLhx4bW8
IzswQUFWaxVXbqRkHCBlzh/fxPX2xvyMBqGOS9owcXh+84z3liZLcrwEOEMwpDC+
URYtvxLJpioFmQwkgCESHaUATvieBLnSVHeSuVU7WJpZCcrxoUYSE8JkMQ4rdNc+
syP/nwwcO8aeY2rgEJulNiWEviXkWAV7JsRQhcrf7DX+LEWjfu8KTCQHN6Go/vCb
79jGr9C4GjPSkjkZeSVUnVM4LagdS5DEBxXS2VBXLu9PlQwxR35FQ/AAzEnqAN41
8I52TrBV19l/Pq4yFM3Wdv51HdmCbE8DX1Qb1HlZajxmkgXd+jqRRPbJ/x0s6GAW
wZRCnE4hvp0T6Jv3bF+k58armSgyGbrG1uIVWtNvNaadJtBQQKYRY9mjYrq/liJY
Vr/pwb1X+YKjzz7Mm7cKrd8e/cBjG8c5LHq46dnR+ZIHXLWSzkETuZNTv6J+Io3H
TxbRP/7qKKWZm2vdvw4qWk8QveFDd7Nb6aFmS3DJ91PWyIEU9C5OJ06EO9KABvXb
AANInaaJ7a9rQxCFl4ODQc/Dz51V/ekSIKnykPqf4/xb2ZRb789TS2xbddSi72/H
M2LZWYDAVpS7CJWlSDxxF7j0Wg/OnB6ErPlcwUUh+D6EeQYOSjQw6WifNaoBY852
9Cvz9kpU2jkrAqR8GPfCHW7PwpdHoJ7AM6s9CS6o4ZpCkdCkpe7DAHc6JVR3HSYQ
WM9nN3xMtWOXM7F97HMNsZ/v/q7nbCb2Zdvqw8a6apKEEcDfpsviLJHwM7ceherL
R3aJFBZVjg2tYkFr+v5wNwJdTZOY6GU7DkjUsO5/Il2g2BhemcE04nHF+j1UjjMn
L1nuInR2aWJ+qJ2g61Qudsxjue5usbqjN4TVv/oO9mqO0SzymCaFJf8PzUTp1A3+
X84QK2cHNx+KTHXupecPCe9wlDBuusD8nqW/n2t6Wl7Kuens8qca/fiJFUjZZajU
L2H83nlM+u15NMCeVnOVS41/l+gg1tgHSWb6goYVicqH3zmbAwp5Qk51Kmt5N4Zp
aL4NmB6bNXDiGbdp3jllnHWH2CoSXy0Fzhjr9zTRiK+8ie8WaH1k9JlpDba+x8QP
mZhz/ymPH7zHj/nf9/GZKo5Lfgk859Ov64y9/1D+gl6v4VVnEVnntnUVY0418UFz
3tg6S+LqtyHZbgsj5lpKUUb/v6O9SFeW16oov0Lir1uF5jLonJdf0K/GLrTAoZGq
YtdZWeuH0RwGeJkkC1DH6aO3Ho7KG6anw/7fYnJ90RwTl3zn+cpJjSMbFZSYfhMv
SbqxtbXmGJ9ZxKmwgSBCk4FpKFVcG+EVQS0gPd5YdwivVkP6ZDfHCYZBYACllAgt
K3NL2JcnvidtpnLH/uYo6yG1WdhcxBnwy/RlvqpzvFTY6vGVpDs9KluJcp5nGG7v
ksjA+rdu6uKzaCsagZKYOZ+vGCA2u4J+5gd2dVtDTPVXisegl1nHsY7iwpfEVHeH
7SjhoW68EMDcxycTn0YY3A==
`protect END_PROTECTED
