`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6DgnEaDWlG5G2oMVx+0bGIJcHT2+Kuegp4Yx3RB+N/iSHX6RPGkMGgSNYHF8LNMq
H7FdIq0ByBRSdHrPyz3RDflNrJ6y2GO1ojqSp0d/VAXygSn5Pen0Tu7Ln4v+iONF
NF7vxFHKkt90mX1Tncdl3U9cu6gMt31xLI1AsZxRp2JJnTmC8JrtLwrio+WxmSkx
gfKx75EF3zwWwyV3JUBokhUk7Uq469qpW6e/XCpJAHuJ3/yKne56aa0yTVX8S9XO
UwQcjxZtstLuetZQ7HTWL/rTJvpAV6r6IrnbyKvSP/b+rsuQvqJEI07PXAgMRpkf
6LOhB+7rfrAAnHd2twMI92No2e1BA7QcXsmb4hZXPhTD72AuKuLa7rZyf+h3C48C
kgNsaPymySfuUxsDHAlIe1KWu38Iz6q9tGCvmKr1MwNH3ZbPziVYtqxCvn9t2KU3
`protect END_PROTECTED
