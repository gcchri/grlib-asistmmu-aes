`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xSrY0X1JCXo/i3s7YiZ9lG7Q9ee7ez0JHJLiOivYdz+m0U6zF3J9qhjm6fjB1bJG
VSoM/S5kPLHdDqgGv+aba3l78qImaKF8uZXgnI6CJ8A6nMDhI+dXJclyGWAl3KOU
4hxA/Nx2Fj27CgVTEyzLfuZYz0OdlKjae86FN2BN297nh1+rfIPSEhYxKD4YxRnQ
2FyW2X3z+px4kO3MuUR5KTUFiQ63agjozhs65ExuX+AJ09J35lU+ZHgS4dTLnLot
ujiMMX+uWuoY1UJUc0sRzrM/qGubOyZWAl9aYNibJ04/04QrRFxKomqoc9VLps3+
`protect END_PROTECTED
