`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ivMcrd7bqQvYk5euikfWwgAKpSUDhXTk+peJ/2lxcvv26PbKJ43zWqUEfQpPirWe
x4YSFwIRUmAm72BGSf6zSakcYQ8VMGPb7hGoww8qcOkMlDNLITX1txdTE2wdmGZK
npWDsJHF5xVxZg5GoNt1sLnMD1YxBRpE0mOp1HZrp76oR7EMWrCQSdANJEnAg7fd
rIP2U9OQHz/N+ffLiIeCMEETcCN48OyHVI51mTdxR01albo5gPpj3XgnnC6gBG/N
Q/AVdamr63FBYMcOjSdH7MA6tNOo+CfQknWmJ2+CWE9a+oSH3AcHoWzCjFfm5U4k
2PaspWlpyMmkN+g4qsxxmQ==
`protect END_PROTECTED
