`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XbnKPW9RCVBkY7Lgoq19xrGLo759ckrc23bP00Pmr6V1jvBO80+Wrrb/KSG2wUaS
fyZzz3PVmw25NBujsvDs/UVnoIC+ve5RGixk4v+yTnmuE/CacMSh4ZTiz744hNuq
1Fzl1J8wT0jb8Pfo8qxLiS1bRtJMn9JWXNAMm48s5hmqnTgMS3RdPIitT3imqLnf
R+yC4Ybz64egKJde+8nm52CUsnZxhY6AuWq4vCoeeKxnB8k8k0o3zpWTa48lfIH9
jl49g0q7aJWymNuZ6Dsn5aEgO8hynuk5Gm4+EIaXeuhLSu3lvS83RyM4zFosKoaM
vf9O9kyy2TFb73xYioSMRgrg9cSc+JM3/cyqXmJm9vNvQCv0OBr503sW7DAYUYx+
+JQtfhAtolR1S6OY0liLhQEnf1lSWq97i5LwPrThto1BMmo65MZ0wrFoHNFoONsj
7Cyou05gyO4YfKwvi1wT/HjTYBTmJCMfg2URYHDn0pMWq73CsvPI8YPBpHgL12Rk
8kozLaom9iBMp4o6tvzUZyFPwo764eeRFubb5imYBS57iU6UUC/Ff8x9G8mSaln4
FzYK/WX5pCg4/ZldHyWseIb9h4Mo2Cm1T6yMBfgmaLe2Igi+Vs40vMiinAOfubaq
`protect END_PROTECTED
