`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D4+JYR84vFTTODpflbAoE6p38g1WPJ/jdD3GtAd5x2/OXq5hPOUDyV5yQl1+mfrE
ez9Qq01X2txVqZLQu2Fu9dHfCCnbZFYshhzgQs3xW2L46Px9HhLMm8C5OlHH9UhX
CtCcAsrnAQ52xOnQ5CXC0iS3QUnMzLLl6VbLXdG2fTpB6ye4kE7LmkOQMSl2Vn1a
ipLQvergJIscVNBrV+fwaMgBevCbPtAp1K7mX9SeDywmtUOQAH4B7p6HfzEm+dk5
zc98/g6yuTtRT+e5YWkwGw==
`protect END_PROTECTED
