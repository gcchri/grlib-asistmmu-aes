`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AvCx3wRIyjFNn8siDCZXzS6hgyUbfNtev85y+KRvhE4e8f1rXVg3gIuozk7Hx1ZO
6fB9Naj0sfZwY/VdjkSrB99lmBfyIUv4ZGntijYWpfSpIO5fW1oYNAka+J6QsrNu
hcZsZjVhCojRpn9iRgTwFmmuiK0FZovfiLInDQY3BUWsBeNLc5xpCjWQwVTyuqRQ
IcLGD0reJD79+giyMnuPCPhMb3nts/AIoY32rf8gajyXJc9jOrKpc83CYLBaRJYp
tHLnALc5LX+7MQS6IbIzazmXfsS8GjLMHKe7u5STpdppSTZGjA958a3eFHd05irk
10HgcVSML9NWzlRzFzdTHDPsBsFBYNCLB7sOzkBvnzsOBecFcaQovVys5Xa9AM/x
GuzW3kr1Ts37vBVbOmKR9waP0WUoWhTZGxO7zRbUZjAe8v+ZwjI/sXBsiG11jgpz
9c0GfgKZRi8dN6GsEz5Z5zEs6iJhdFduPJLONz/564q5KXIb/p2GurMK/r/fBW/x
knGOuwspczBlCkNdcjqeZSGaSDJsToqQ1WC6ipPcUYF2R1gArt2nCEkSq/Yw1iRQ
2bq+d2HnUC2u8Z8TFl04njnpYbVywYOtcjef+Tt1yVg9LArCEzXGohsg0YJlfwND
e8WunqIZOpizE0uguDpLnMvZPvMB0wEHTjNn5Fif1wsWQ8WczdhjwO3jHYaylPYN
GMZDUd0dLQZ1RuBuLmoeJgma5TiW9oS/K8l/OtaHSD2EcmgSeIFOwMDyWaL6WH35
Jy8Sc66RWqd73k0NyIEG6v8/I+cwaEamB0vxb1if/Oz2tr9qD6zFlXv4vMxSLnKt
PmxyV+mCjB3H84KILka2UYudJ4IfBIhT4egLEgRWqRExkOcaxljK8vstVoeTVNhK
1xWGyeCKtVsmJpBATXoGQZMaIQSCujPXCjYUju4fFspvr5YJYiQHY2BbtuZ2Eaz2
aWews8vQ4QMPoHINO/pdLImMzX4xne6tiAbLOZU7IC3j3dHd2HI7YqfH1XXmj2g4
wLgsYsz7/iE6NHZpvRT6hsyKYqaXYXPbcKWBhftmxHfHrnn2hBxIXDHa5IHT0RQR
RWIBfTNGVDxQlUapoDohabtS1G3q1eYSs947eBB+UOdll+JdzpTuPEDEKZEB+Q8j
YGxLPnTmj7B8l6fKFc/f+VC/JjEWSomiZntLUbg/Fc5mH0H7tEebomkVdoJEKnEu
FFpzEBCswrlWgATuaYeDkpR4ABZ9Qv3iVZxFGqiY8cj2ePs0XI1Sudm1QizNoX1V
4FqTXWeeu8HrqC1CeEMrQk4NlQ6dfnTOSxbvOZB247p5OBUjqhCEVsw4b3kZCbIj
l8IKW7c5Nd3jeFn0XYuJOQkFQn62T2KQrKK2oTCBUrUdkWCIFdHlbjXHUfbahwk0
Ou0m4jncXP6gPNebPtxdICKS1+MJOtB7xwXLZMU37jATXcq2I7iNrWgaFtDJjvBt
5y0WKPFis2hUyH7QsmRUDDyWJSANpHf0Ofw66TjZhNc8cOgHruAt+8z0VQveKzGY
E5Hh5CDzim8+Z48ptL12PiCsTzki9laVbWln4xcPux22+KISBe+rvBVrcpZwzRT1
lt66yEHjQVN3HH74S0TL3IuwWfLUF1AGqwcVwi8yap9cVOu3c9vdiSq4CbW4baDp
eXEWrp1qj8y6sNcadj+U4qHCqbDe8Z9fxctLglq1S+RIZ730A8SDiuNj1oD0LZdD
jOVAFkZrN1GACacD6WA7AwMWFpaE6pAmUEuNRIlO1Tr4rKhKUOvsGUanlP4JIghH
xYmmvxl3PA7ovQ9oUvDb/L2nRxjS4lJEFC26jLHbVhIDxzmVXMhFwyyhPXhggmF6
MuaabpgyR9AgrypEBzIZB3xjMJzNv0RBtiFl5NW4Pu/auLc+LSxc4ILc6SJI3RF7
HWALweeY/k64wzXxTxtj1zUUX48rqe2SoG8mUrbb3yYYRscQb9VjF1PHcOA3z0ZL
oxTvpdrnG+V5t1ucBYwKNEs8bt9GIg1IeImOyTvVyB8925hOse29WfrdMhIgeGFW
Tcfyb5+20g7wCR/sd7gZ3pRY+A5VfxqPHwroq2GPdxja7bvboxaJ7+JVvEgrDqsE
iWqFA4OO6FZUWjt03X2QgaIpqgj/oeEnYJppsrVcqxrsr85P3zTx1mtcfxUqFpPJ
Tv8KWXGAwDQfQRbAc1PyFk+FnkB//fFvCwg48FKhOU10rT6dps1Jf0DlYvSO+A7/
wqYEuk3ck2xC3z1uhc4EpZIeRbzzScd/nuSi4OEhuAIbFnBG6QyVl9XlXBvdZfqe
xvMnbH4EzKcSnKPlhtqrcL0LzhNpztYj9BtCBsoiGJCRWnYaNfAYAhtAsX53hrsC
T2yvC11le+enICRwF4urbUeziPVpidKsCmVV41T4x/B5DOHhntN5uuvHNQ1FWCLC
XkxZdStLMTY9MwueKuHXEb94uYP0k6iqKcPEou1nsgJ8CKc9gG5RCYiPG3RGlLP4
+6d/g1OPw6S+Uyu355vfTlbU6m6xxDAvwsKkI8zpS0OIiqmZWN2xI7Z0cjUx9jad
Q3hn4MHhLB2FjU65bgnreltZ5djFPtZ1/eA3JPfcfMzmzldACL4PsQ+BUI7Xghs1
VasYhF5GUzDSyX7vDBulwXSEDPK+vwI32thuyXtWaj9VxF8vXGuBZ7/PwmwvIYQd
4WFNKkvH3jrCI61ZMbdCP6mD/NMzSijy9g/RLYShhxiNOIYa4IcC0WK5E9BADNLX
103LuJgkrFrTMuuDgc5ZGif2Ygp2ma3EDu6epraN3lGanELK9ALP7NYIkObCruon
gz3sU0RcfwfZjkJ1CgRF9zYzH8wQWKgnqcnwAQ2/G5c1Zn7KBTwDAnle0HO0+D3d
G+wMbuLKH+TAjIvqCG0Koy49we/lIdYEHELQiA0uZEokp82LNMJL3uUk/BN/nh8S
/Z0hhB8PBvZ941IrSIhGoda97EcG4JPM92btUIiDr2rzuaIzbQ9uCf/zINrSkLE3
nTtz/tICBgKwOlN2BFRxY2VtGQwrDVdiZ6+t2nF2XU8xd/lsA1P6mtP5ASy7nw2F
kbSJbVRj2AH7sTS6elZ5NpQLbBYa/sI9FeSziBGqHhnkPViMBW/o3cclffsaUPcS
ckxCfFEHaNSR1TKBUMRZpxQBZ+wVPBL++HGxye9E+UsNcTjD9J9KZTeLAE98umiS
BH+1McFBw2Gjh015yfYuHte7YGU2f3VCb1M0+cPRFUZbqE51cvHFIyE4wxv1ZKo5
0P45zg6SDBEykX3CBznW2LsONbavQqcHiVsTRHbAozZ9++6qdqJlOWZRi0/aFr6z
LmKhfmPimXN2fppFvdCnfitaI/CRSjdTBwI0S8KS5I4=
`protect END_PROTECTED
