`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1CDqMLwyFgAs/1c2lxAEO4Bufbp6RUMW6uWGIFBlF1rxjp8u6KpHlV65MUvIP24N
rCSOqylC0naOEAMeFXuI2/8abtr3Gw+FczQrJFmtydNNpyAKTQM814sHFCsIuLGp
QY/+Xrq9cePhNxJEZKIA96I5pgmdRSP9GEE9+CoZWKGRQ8pCvjWjrTrglgNgomIb
TeBz0ShX0kalP6ynKb/a3hStBvQhQtHnIiNdPaZ2N6t0xzjLYrC72wTgyEoEfS4z
094qVT0pI0UxBM6No1Lz0FlteFscGOi/0FtyRc7unSAh7CdO9OBKO8o6s648ifUz
TpCm4CG7r3U5Rd6Wzk9wR9BA4xiqZn6c5uBygYNP2eFLfoDE65pnjgL7nabmN/y1
PCel7KgJhPaSSEEXpXG7FwYryFbviRoWvyTHPXvAcIaExjEgnVagHyuHv1cj1Xtp
inhRAo8JZ/tDyOyLxciVefiLdtUCtSxTd2MB+2l5rEkWJ6gkd1rMJMchv0U9Bgl8
BRocCCgJTEUWdJfE6Evfz+OcaP0y49BvIgRY2yR9Sa0u9+Nst5xQXl1B9TbgfMJS
xlsIL3TmgqEJ7zrHFYTZ6tA3wreHP2MYtYB/K4aBlUZt/m+50zcGfsgCzngeqD9O
4Rba7jKHANI4E8JIXZwuHuwOBNz/qorvSD2Lky5AucGkJZCd8mYptY2hzkhA9S/6
szmxXXII3oMqymLtFBzxRGza2jc+R5RqLGDBC4ztiTrUkrKL+S/ccZJEsXbKBJVC
SEp7aP9BuLwjPe4TlVZjKkbdOd+tfO+BK2S3lCPiWWzh8FCllVAsjgrBKs2IUYHp
i9W3+3jNTtGrlHSFXbu+XIORdDf3nl9tcMmHMQkHYN4JI6Be7IK1tTASyIjjsXrk
0/odx4uudQQe5CDNbIlAtgnsrzVucg7LNe/+GiiQM2BUbzQH+Zl1LiXF/gJ2M+WB
TWilQQEqWagDqj3cOscnneenwuQ+jyC0FaJA3AbidIj3kwWFM6hECUj6afNeMUzF
AyvtfuPn7lzg0qYwKJgXU5XZcSuq9YAC+9gc+g79a1Y6v0s6Sr5xc2b7vh56Ljcc
5faKN5Yvf4DV/CKPekSbxwLvuHqLrGtBNKrftMCbFMkv3cFTLgAYJfJOHGvjsD22
83f4ZdyXz+yWwPMkCdUDk0ubQv7MiVUlDTLLsVR33iNamdKI45N14NUbU7+5N5Zu
`protect END_PROTECTED
