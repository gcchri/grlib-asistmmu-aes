`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+zU0ho2/7eXJVlqOfEXd1giu8gP1mdkeZPTvuxWlpthiogtlNlEeKo2vCOS6Unnk
wmhmah/bDfnCty9TkzcDLjQIoMEsNu72Wf+scJa7wENEOV9Vhr/y+XlFki+pPCZl
oXi3KoGjxJjslFp+5A7AJskRhWH17ZMA/jUjEUfUnG5QNm3jlNd5gsB0C4/ERr85
nexG1GS+gM7GhQy2FO/d9EJh0Riyx/ogA5AhHIhOkpwy4c42X1gVDwKKAOUFnn6i
r1HISH0sUvmYFYXZB/hAuFXdRc0i3BAOC45FKjENCuj9ap2pmQbgIwOq+CfCD+D2
GVTq8uSq9zFothn8Ooefp0Ps7D6qU1BRjVSpSOeuoCkXaWvH+Kh7wIY/ciEhGlIT
h+IKxpUOeyBPHm8/pnmwEEC1O03fkjUyLsgoQcd0paRu9MnlvEjC2LTtDyjq8VTZ
x9b9xspMbAt8aZIxCZzfi8/Eqi69HiMnKge/Av5UDGdFbQiVuJSFdchyWStd61pb
V/+CuiZVyNhVumsxPSsY43i0fl2iusvgm98M7vHihFqWylR5aA/MqWahvpha5hCO
ZqryX3g2IpDcMs/vwnQ7hOzFI/nzd5A4Y812gpZog7+q+ltvLcUMcZak4Lf+FElX
FkA0yyII1DJQhLyy4helCKEnCW7ynH7X8aihXTQXnbneeIUIuz/WSmTng5ur91+V
WUghh60dZh+SFNOV4PLOcoXUBQhkhBOjOkwD5N37wkHBL3Cy4qkafWqQc6Ku2FnB
xaqlBiJEj13Y3gNAdDwPddh1fKNWEIYsXPlsTBJdXYfC5e7vWVdNjm7JfoFb81m8
ndAESMYkhqOLuNv66h4yX3HDUBCOZ9dxZvnfCJgMD6LmGXSEtpze0onNNxtWkxvw
78zTCSLlpP1TwTFDGROB2Bgq5DUSKKMQuHl7HWlrE19MK4nDVjLyBqMCBmvzjFHf
`protect END_PROTECTED
