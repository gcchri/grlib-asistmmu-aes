`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aWE5wRcfXmsK11yzuJcA05lYr60PuEO2zPh5/GVtpFFyov6xM3sx3cCSuGNddoHF
flKdVYQCARsBy8SmfU5M6ZBnADLbfWVFtcEAmTtA/WmfOweBTOSwZVYYw1xT58CC
2Xmy2IDBrd2B5SgJKHCWejQcb3JwQKR3kSAsAX9WW8SpIq/en1iQZ2t6NFrcy/Tq
HrVeLjxtB59wRcTqLB9EdK13mCKq9dn90Bm0dTdAuhh0NovCxz5F9+u8Z32POL/z
3bgX2DJ3kKDZWST7be9TJIZOrOk1qLfHlwAWezE0guQJXIE+SjxpJMLia4FqqApb
AHNHA1DoJWNfguih/hyQRvoH2ucNOU410cM0z6Bx8ntU1c8Dild1JNye+Sx9q92g
QhGMkyONYZcKXSXQCH5i8a19VFoF0ihJbr/WJb46CvdWA2UDnYzDskX7gR407eVy
OyUHvpp5bxfu2pzdxoKVPe52gWSGo/GZeZUd1jMjUvCU+3uuI0jCCB3331ffAev2
leC8hdEAQB5w52sKZmeudyYX9RqjhqROK8d1esUJBZewf0RozFuajJ83ApEQ70cs
M41bbEpp4F7ET9DtWUelpkSLwJjImsZ6b8W2qXRjTfISDhIzR/lvBQKJCmDSQVbl
eOossQbEnRE6osW4NXvgg2qTWsqCgbEnmePVft/12yc3BYd8HtHAYgqSfTsd24Qg
lPP8sXCuwouuBL2f5U1n+gQ7DcT+76Z0DzBVgt1KKC0yfPnbRxxED8xdiSgMStOE
ALSEOxO7cNXJJ1EoXHatsKv02Ymzy1iq7hVCMc0t+7LnyrYGHxTT1EKhV9mt+BX3
nBpwuiWLmQRVc0tyjRRZs7RPKtlKT1ZvzARXYac6jRIBAWK0yVJtrHTahGISgOfm
cddD41BizNAU3QXOWediTUTDeh5L21rVWMW1wiTBjG93yRdaLJKsiZWb/rROHOUb
1AK22r30JxQmxjTizYKX1TrT+qRIp89lcKv+Hp8apn5CQRNrpdvday80/7abr1pR
qL5y6bp3yq9ZIZ9hlCcTzlTC1g507Mo0Q/5GGZ2v2WTC5S4bVv6Jd3jbjyiOlNVU
7MMgECQYZY5QoOCkiOMHuhVfcbLLaCAasR41QWbRui+X+qiK3rFNK9xFb+O61VEn
mn3ZpuIITZ9eE70BPUyXv5zQdruM0QIyqyEkI+pksYBPuse6vCuoVQ4hLwsfGzYI
ul2n89TRtqj+e1wZrPH90OrXo2YWRcewfKED9nqsLTtUBYyU28dX8EaFXeDVlcbg
nj2kiyMsDVMdWpqbeZAvrtPUztqHpa2JxZ8Iye8chIp+NLMaOFT3fjNuh2+//HOH
8wnufF2612ZdfnAL4hJ1rk8YoGLVP/GJ1pX1rDpfdGzpVyZWiDib8hgxy2YPARKS
tuwsupAPaT+LiB7ayDTOgjL1DpWoVHZdYFIKewlBHayBy0No2ip7x+Dw75fYWoEl
ecf2iYZqvnKLnJHIPfePjuSzLTM3nxp+y3n9EAbERiU5Z0KbBBGxbCIKGm6VgZ9P
qW+KylPgwrZ1e0icsSfk1x2AlTOdjuTPwYbeNtrrNOCflRw0hVKds5ns1LBbTWUW
9UYdiewWkGM0dS2ytmpwioC+fhy72JUNxpW0yGdvnUgjNzg2dvMuMMbJsSfvJvDK
OD5eoWO87CtcTLi/Ms55FDtm8N540Nfz58CykolRXzQy+VP0rWI+156vdeaZqLdA
/4f00rw2KGq2i/+o0EXbs6tZhLr8A3pUOzA4qD5NjGG+oqTB0cQJGLXCdZNyNu5i
vxf5nr2VNj3rkepms8u7snCuvlOHaax1Pu1DQFw8q4BpRsBiJZqqDB184cs/MbCx
WB0BBU2C69w55sCMpAixgkYgyazGRMDq08sTNKL7K5HQWWSOi65NDd9fv6FexCM6
FTDJHs4fUlypqNB0ZBwAMAq5hJsMf7ezLW3thAt64FwZz6/hblN+i3KhHTs6wZ8M
ND9YEpKzOFPPAgIzK9n/DlFRX3itFWcjLOlCjuIguoUJsedyWslvSvxR/X8IYXYD
n56kqWHq5fVsJjm68nXZPvBARYBsRTjuQNG5kcH8iK7ldtSDqam0gkz8BeqcC047
FsNf/lAhlY7GHudPgvync0ZkDetfkIrGhm5WzsuheZACoZJ450wEn/RhsOgm5dyq
HLLDeJl4o/pe8joI3HH7LKd1FURHFVuqj0+TEXFf4QrGNDWfPm/rjhjB8uArFEpy
YHlVrBwj+MuPf4ozXxY7DGbs+OldPbNGE6dJ2YAgSt1GWof8PmXgABkuYEnRJvFJ
+pYFnaIPrxEcP0r/ZFUIBReKK+Nw/ZREmI2+uRdRuk2AFIe4bDMZdUpN34FGeqEg
iimVIBuKLLti1GQ052jR/idnrN3uYuvDSMXXdbXL4cpwgFrNmhj1nZhpN5LM0Va3
Gq4KBE56gOdV8ADJXRl84s6SHBqzn2frbgblQo2b01+6fDToUztqWDO0sHbq9f8T
VZ5lIrkqD0smn71n9QyZOrCPBOmefyJyg9/XhoP/feOG5xJMsTZA69Q/O6Jjg1M9
R8EuLu6Zlk7jXoHaoIkXZZ5ceIDjj5ZeNtxgiJohDkU+N0vXU+MzkEPnJfrrcK0A
7Zo7RFOlHMVYYZySL+2Aphq5NHBaAGTvPpeATHXLdEMVAPZjEi4q2GuOXkPb7ytT
kT9TE0UAwwT3FIdi7Vme2EWQzfOTcgNB3l23OguuX+JCTufYbUWsQZYYLtLre/T3
lc8MwXoe/jJINrTKByUoELUctQP6ERvpJ8bYfRENUGKw1MkAX1HevXEKY+HIrpkS
IAV280Xmo6U1Tt2tEdVjRay1pdF48FrZcdZbtLhONrcS3ZEsrZxFcYc1oG8espkN
E76/2cMQwDTyV3d8C5bBitpTFptdcY61REz2ipFSvFbAcm3/8y9TjKO5wd+2UXfO
r2vtwPv9rYRs9VRL6hr8M9Wb5XwQllleqIt2Gln8r3eJGBU9lri+GPx6cmSudhxQ
`protect END_PROTECTED
