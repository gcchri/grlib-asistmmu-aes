`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ovs6f2mSppA+8XcyudTLnNYc2LKShJlMBg69bLN2KMA391TPE6h+WYZLJKgyRo99
8R90Q93EjZTWmZOCT5THKfN6ITIM8e6hWYKDvlgvwNhqWfk2miuwIuYzC+LTmzS8
9nriSp5YCJ1ueNQdpWeGHHBl022nsQwywTfj3aofgwtnazWME0OOQ9AN+xmoYiNN
lUGWaIheSDnxCTlXaW+pnoubk2WqD5YHs0jSuPTZVXseOOrfRhFvcY7M1NOfxLVg
RCwHLNT8vOWKGK2RRxDKemU717RUPSl/CAUdb3pxsc0w9eFtNbExDBQWzKDxl+H6
iKn7W1xPkCPnzGWLdIhIuaRBMCv16AQwqFDJ1Ko/T6JBYVz5amdVzagHFfZnUL9K
Tj8xQwu9Xs19RaTG+iVx0UO5MsTWFFmGtDSkBGjmyfc=
`protect END_PROTECTED
