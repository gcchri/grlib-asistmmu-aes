`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oh4b7eUe0sjL1ODr+jaZW2WyiKLVrRSFlIVRmOH7oY7M4wmkNkwO/v8EigVhEogi
bZe9MVbgetAdK0O6Sx1IA5qpenDFbfDaI/MviJtyeoOmOoxT5Bw+0kxUFPDZp24c
Pl40HTsi6C81zjuWzXwpz87CnOPjv7ij/NNdFDhZ37f88iUCZcy51C7AoeQFb5Tf
l/dSb3q7MZIvOjt819Lpm5tQRFnRxx2tHxm1SLaBT2vBa42S5OGgP5sE485XK/sQ
9AbR5h6Dl/NQ3iUCxvKaHNN1mJJDUW6m9o/HB4625E/khXC+3kI2ALL9Kz8U42aa
/Rtb6wciQc7PBt+r27mFgQYM4YL2sT7R7VLcBOsxKqL23dnBe/4C5Ot62RlSnqeZ
yzkFqxPw0bnURQI0wXumIQOJ4hZDe7HWI9KLrbv04mhftUb5QAMcQ65JqX4U6iZ5
kF49oc3RGlLpyi3yV3BvQe9xGIDf/+tLjh61kb81YUxN4pesjDG3Q+R6AO1kMML+
GB1iaWQFDxlXScrajdoGAp4HHUwzMDuYMWNJY48YW471MACfvLX0gxVTUPnKpvL9
14BX7gLuCHySquGzzoxmmV3KHciaYBVN0m9JbsXTY0gBxNnhVsRMNqTPEMO6zQKC
48Epduiw9Ya0W3yG8SJpRgo6hwMoU8jzjdOmgY6UZZE=
`protect END_PROTECTED
