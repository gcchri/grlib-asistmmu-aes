`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TnJgQqkvrsc01dYjKY/NzgLIGbKPdDJbYZW0vSJ2DYX5989pjLJDX3YT2KcFqDxu
0csXsSt7zbxUDcm2UcEb3Uze0l3akWFJ/ct1VffECZP+BOmnYxgcqa4OUulJrntF
y7NpHnb/LyyJ+pVoJj9pf1xTHWhpo5raZLRc1LksNT5hTD1XdbzPMetLX19VIn0e
zgCHIVhhKxbH97YcQG9fbnzgYQFuNpBmdzx1bmlZzQ4IrrrvrhUNxXNtSeJSZ4m0
nGt3tHNqpGv0yb7ZcDy8XX4dGteIhqx2tFcfm7yZeQ85/TSmzcvwLuLu08rM4osO
p/Bb7brWhEG9CYOW+UhfhUsmJ5UJgnhtTiLPzoGtJf8=
`protect END_PROTECTED
