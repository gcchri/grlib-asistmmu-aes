`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NpzBlN3uOWM4GCRRRaFjpiZpz1vuWrPz0o30UbEpW9kV52c8tbwgDXczGxbps41x
8Dyj9mnh/HxrcMVXmhbQ8mE8ZAyWGEQBUMgkGKvtoSeM7CtdUfFXwHs42E5S2aQN
dXaZVdlVAMpdr2IfpnN+BvlKuKuq7C1ZbnDrBW0K0iBpZ3PySy09E6whlLNpFNBq
k/DSoV2mulJ97XPYoqKVesO7B0wRdzRDNmkwe17T1HK0ZgLOHsIOOR/uL7Z6UTJ9
dALDmniD3skvFRph5TsNwklFotK324eeHpDvFhMBJX+98pwmVsYPt3341nUul/ai
DbFgjq5vV3dF8RIK6Kc0BJIpp1Ap/X+siw3sPtD2qWmcfj/BgGPLNdA4SF1H4vbo
rVTZLlBbqdzQFRCKzKlnQjEm6s87KDWqa3+XJydMgp0AjQNtcg0+U7qGnzhEpLBx
k98KP/K43im1y+isoGovZ4yfYosH/J16kw84ozZxyupnBxaBIgKbHcZaFPfgZpCo
Wpo7g4r9nUm5BXBzbZgBzWZOBYnzFlHceFyHEGEMKwNXw3updGWkP8Hgh+rliYZH
Q3rLsByboOpP7EnwTTLyIbbkaW7PY/HoFbn4suApnHfvu6xQQxvRkjW4Fb9Is7CQ
cwN/aTB+jUir4up+W/b8QMudRFNpKKZKQUR0nZBy/49QzXqysjoXnCWzRsYP93ki
bYPQMaj5kExhvZmOp9aLkw+0Cg5Ehsw3703Eip5caus9JcD7hp8Smj8I5c3cyxRI
DsFMN8S0aA+kel4EjXLrZk1tHhJJ0m0Wxq+h62Bxd2Gap2YH7yog5jYcfXSKdaYM
svgKW9IV5NOR14xBsnh4oAOtub3NLMl56cso71EhoL7S1yCFTripmoPDHdYXsv07
hDvO8tulIRKR37TnSdnN/P21Dm5FMsp7oo1hsnD+Om3zt019YRvEJpSpvTMw6wL/
dqbffrG9NNqwoSjZH1l3GB3FspNG93PdpJ1u0mI3I5A=
`protect END_PROTECTED
