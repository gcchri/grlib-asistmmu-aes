`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QA6OQpMzJ08u3T6WAWhZDWZ2yf9UUSInSp/IIectNSW4aHmucoFT5TQmKiOHwwW0
OSBE3SFnbsSQ6GISMlq5OrvT+LFD2hVJ+yYVZHCQ9eW+tnJGMZI7S+2hAttRzdCA
NguWPJXnHpdGlqsDvsmKb4+BAbJ9W10v7fB25O7Ue1F1B6jWjqPS5FhUGFjkpDtD
hwLb+oIlEGy7ed4r22ETNzF9kfYuoTzvcGI6q3Ia+mhlTykDyaQ7HVb1o64LS1gi
HTnBHvHER/bfwJT9k0CoUQ==
`protect END_PROTECTED
