`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LMXkrw7f2VcxSIHg1IM8rC0exuRfeFIGMTHbb7aCsqfxrRCJUfaSlSwGBiKsY6zX
XqWcSKTvv+GnMDPUyhoU4ppoTC8IYZ5mFJbYenIPJQrpEoVIaTtwyEk8oUWYxRmk
CLC8jekJ9kfumERdMugQ4/kbXOIsP51LQ4tbNFB9w19XgnKI7PpbLw1bF36dh8yn
FNEXGhbTjVduIVaVzQKgT4ocBVd1AsD1uZqKuzKxF/CHRQloZNkGRVfPgjr4xbwu
7Fg89rM7fnAM0fOYWorn4ijwow0clTipt8oaKAqD/OcOH9reYuZMNiaaH6lxUuAh
kt3t6RnJrrE0PkT2RNrZJJpu3XcnG09a3AZNWbDyqYUgqAy+/REdTJfxjPEL2gOP
HM3b2dE8lhg3xjwctOaBw9PJ56DFtfH4ucnuyE/boYjksn8W82l9qudaSsgrAeIJ
+QbkYfJg68LesRzOS9dcdMlHA38130TR72DeDDyUF5Q4f/dFXQwIxp4gz7a34DCg
9ieUJyHFe4md5D7/F9RXjUzPl58cJFndawosIkcsZVujvPkKCxqTGMjufqSMr76z
d9FLbVMkIE+bywaiS9f4yg==
`protect END_PROTECTED
