`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IsQnbQD6a77ZxayWuhYdHOLwiHvNbDdG7eOtQPFC0rFLR/26p7Yrs+as+MNdXYgg
/MCWvu8PYye/yB15xiNioh57rAUBT/yJa/WPqRbnMeSxDArBaK7RbEZ/vp7z9z0f
jDj3vOh5Kp1Y0Zj3meKcM6Cn40PzglGe4iT6QwePQwWRPI5HXceco+Bloqg7760S
6pJBzBEns4njOxNbGSwxlq4CXjn+XWGbSe5LZkrt9Agn36vPl2N/nv4yKN1Diiw8
pk8hdP/3+vPMLQ4fel4w0Kf+bJslHL1QOGNvv/RTJDQ=
`protect END_PROTECTED
