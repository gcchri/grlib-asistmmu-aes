`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qdrbw5kPtPZuezoKVCg6tTgJaz1dbDiIS7I+DJmV6APWQ85+DzuZKBDv/fHvHBV5
sscip/jPkKXrFLHP1yVbyeuu//ktm5Oxbu7kL3NSacfUzZWAEmAxQxDiEevIpsC0
hNkJqYtj1d1FubFHyvWZHsLzbdCMvmpUzANqumeHoSQ5ZERWO/qpLdwdBH8Yfj2w
aLhBu7hVqjsY/7D6CsJ2DbWKOy+DpYdiF41pHujv0YwrJzvnWoBEI3Rl7x81JNre
CoBKB+CMHMsM6bo6oILNBIn+Bu1j4T53P/a9rdynHU5dZ3l54JMkCShBtzTJQN/X
3bJAeux/QmiI8x8ylV4GG/bz9XKXpl1Rg0Fwdx88Ar4JD6OI6SEUjSEwWb/xN5Zs
z+cT77DPwxovG6MTVRTV+386rafHYrFGrcF88tmK6jQ4HkZqCRL65CEe8bQtor4E
fd9VEPx+/e94XfEEm55J7aRzjPskRHRCmjCJlOA308V+0GzpP924ndkAV2n5+cbv
3+ZbP7sgz31M3fsOKN0jDY9nVk/PhNw2S8LXvTFjXcOqTOspD2kS2HJcl8ZdbjeR
0spcKB6SCUBxM/W9fnz5MhFG4qtWO7u2xlMLfzQQkfrWqLq7K8ib0wY1zx6zxKoh
NRnxPK7p1EJOjX25bLOjxY6zSW5eQH+eRYs2aQjbHCux2UayzeF1wmhvCztJhNLb
bv/lvQpVnVjEZzIKRBLW6SIAFjEpAJNdOWFy3eF5/fe7UYC+Nxi7CiM6f6X8GsSV
SuEjPpOnX6JTEppDnl32x9+GcSb6Qhg1xcGF9pLKQE5GIsVvMRI7X4/hoCN/bify
WciGCVhLP0btMVN5yiLIvdwxHIE90/Xt0hohbi8f5UtaQ6CxYbnAXKHN/l7ab8jK
eNwHzqcwPZ7OPYlPU0nn6E6ssGEkDHK3EBcoWftqShBZISYU0rLJFYtQKSBdU8Vu
Hz67yeEN8SQuBtSgHhtKImJjwNeoiakDByz7zLwGKgagvd+o+/YmfV14iQTs320L
AORi6Rg3LXhPIt5qcktcYcV1bXSVe6H20Wotz77mjdDWNVAdipN/lrVMX2EqDWUf
+1EWZu4EHJDHK7biRo7r+LFbPxcmU6fO06VUIwJhLNmqlBM8FLoMujZqjpWWkm8Y
zsMXLqNZ3Pot9Wm3cTZqaQ68+0kPy3lA9u8I+/+e6j4YdwfutT87njj5CrM1RUSn
`protect END_PROTECTED
