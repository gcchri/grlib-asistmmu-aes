`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5gB7AfvB4eoJLer6HdsmgoY0A5pPp56rUHwEHDQ1mn0DjsBPsWgHj0bOD0Vplyn4
2N/pRlMWva2oEDU6nuVsTgsVCveeInMvc6vsuuoBY/mnMjhM0APZPXuywlDQz7J3
a2X8Zb40lM2qxwgk9MBOmrVFh5I7fC5KOA69DyciP0Jit5G5PBpKwv11tsBlKOlI
M4qG/jTc6kEtb5TJqgLXwtqmZVUigrFVXKvwHcRYi5g8s8jg/VMqy5SAxiHl2oBv
leBO5z97m0AwAdHHXaWJU87wrzInY2G2V3PInzZW6tJSmDv4dPoRbD6zGwTt/19y
vO58QEs9VBBjs4vCEWI12Rlkjchy7a67jeHh5kKV4/Y4qC5vDIgaUH5N/KEtjmg3
HtMQPVubjHYNXixDMDJ4ORnE+o7NSSLsQoAdLO7Ib6gorLA0glpaRGkoaqvWsDb5
`protect END_PROTECTED
