`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MIJzPH2N860yrPtHGac7E84A2mOcJQYDpdeeJohqvdUDWIaqCZcYL1lnplhA7ty4
iBRlkEOrDrOJ58klaipNFMAFKMQKvKk0KLUURyJXr47Gjh34vZUtXToT8UhbdT8g
P0rwcKsiA+7DMHo5Xf2DBPZyZHQ6Ae3D6p1iXRyjTE3ib+K6aILvde3yEKi0LjHi
t4LJ+i4d2f6nGCDqzYGGYd1wMr1LFct1t7690kGGKFNqfXgDQuBGyJBP8SFScgnx
QcAvRIp0oxwDGEfcFFRCW/e6tvQmja7Unbay0loLahwiOJplavUtOVcuneZws4Ae
1irBn8fs6mR53w/7jjrT9gxSMSLdFkB0QvCsQkD/mrGxF+VXoAPRQb5aW8fbpsLq
UXtqAoMajHOvVCDc2c66kw==
`protect END_PROTECTED
