`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UDY4kCSJ+gjz3zXdyxYYuC9bbOlcg7UTrhWAQJXblqIX2aZEcxw3hioCDeVmwpab
U9xaFva+3lt2TgHWUGjGDt2taS+7zvDF8/Ur7ZLDUesV75sfnFpDhFDI5zRPr47D
1SuTiEv8nKURrUASN4OV2OqdThRbqamG6Vp3o0QeaLxr1ak9x8EXoAfnrhMGZf5p
FK4tTX0J/kDMWRHvgICg25K6lpByhy87GTQLODM+clOCO0ZLfUF3YD5x3XiDYwks
2Nj4T7GU0aUtrm/rsYwcgWEH6dWqGxKXJ1d50ayjf3O85hT2QMeb5QbSHxXRVnlH
lDHuHubi2F0WzZtHAiBTXQyoX3dgUa2Yjh9lqKUlFa6hWgC6P4+MG5LVuDCU6bTh
sTB9u0hdLgqvSkINRZDe3POICSb7AlkPMw5VfwzyA4xhrNflkl/mrikTGwlBHz8v
5xplJrs0Pr+uXpeShika21F6L8iLRKGTJUguKbV72hrKLO5TFzXr6ZMpFbdXc8mA
cnCLyhR2bGTfdD14C6VvgiMgreJU1gjwCYm+3aWim3sju5iTVuIW7esSBHCF0vkY
Io3GremJpYp1Jx1peCkJeQRbFRKlFqeQBLDQHt4UOkWKV9+50YoGH+jiLeiXGcCD
diLNFuu40+1NP5821aM6sYDMYmXZQ3h68XgnXF1q6NI=
`protect END_PROTECTED
