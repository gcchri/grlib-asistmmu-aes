`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cFkCKyPfo9Li3aSMhnmAKCdDzRNSfzW7pGKBFKr/FlqxgWpBnJNFmefSrr12CoWV
yFBnGUoYJ7p8kIMGMP5tyYWZecmlc85JqY9tzZmSaFidl/EskiX9I02fyWzgsCm4
1ueCYokS92LH1JFsxsIu389E/yKpvc8B47kBrqNDG2/5xucfX964sOzr/neCMBFX
avs1uwtTaz24iN29QrGafvD3nG/9h+/A2X8HAAaHdOB4+Iehd7CvknvH0cD91PSj
1CeGnJvEA2iAJWs2fv70cttyYWfuhllVYIor39XaG+AejutYq2pbMK7imlm7ilAf
NUdxw3nBqdjC16pyK4HmPH3fb9UfQSx5A3d4Oz/8CLachlOBq340Wk7FNGKSN3eI
MrbETPJw2C63eN9OYVpPTW8zXxqkVw32QTPqpg1MMrWTPI6b2kyUURmKZmMQACT1
JVe5i/RqES43iVtdnRHjxpHqQk6hL7gFk1p7EEMs5VFE0PjsoofLIXEGGVjhdJOq
uh5uJmte6oxPPQiOFXr9mcGFmfHooLHbKzJjfS6/hkr08A5u8jlwWhP/MzSl3g6h
s8XRRbRuDEfHVjyB+ZvWjI8pnQgBm5+MmkdAsR1S7yLdm6ENn2H7PKJGwbUVPGXd
CBP7X+G/qWQNCFwUDmDvtdJjKTDBTm1jHw0aUOq/oNmMMC5l0DnztqkhjBXGmF+3
38YgUI1gRppTadJn6kpWZQoOzpCWrEUAZdr/Gft1FXqz43QUwQ9K3eUNjgmkATnv
9yJGGf93Gx+XoUl3mdT1nlF7K+Y1JVcwbicNNkJ6M6APy9K7xXYe4PWWDfUtBChM
4HUb9hC8UDTJF8ePhMGPuRRg8VI67Ik7rirgyKDVN1rfDd44kKPtoJoCM4WrtlLz
G+RgHSjsCBvy1bz5SyIlM059kxPfhpDWswXG/Ywbmzl4OL1UCWbiOrTrskKHI+Jo
u7wnywb7zK6Rjh9rqXCl2B3GH6rXvxTVqfwkoH2YkkdxRlqgY92VBLuMSBA+FHVX
LxbZIZv2SyQFfGSVOT/VT+kq9nm7OeCQFgV/3/1RMU+tmT9vCanHqaWTYccSGQse
NTi7/FuTAWuOHMY9eGLKXgk+4AMjSSCuI5RTmiBjLLkPii5br48lMuBSWEqLsaHY
dVIbalKe9qVxP1S76GhS2OsrLLIG7pAfuYa/QWdCG2RRhX7kjG8gQWbqXwMt0ggg
X3phk49Yc2E0r14M8P63H8qnUxciVqizNL5kE/IP2hQ7gAD0oFPQqvYcr4VvqOuI
ZVwjNO0bErDqsCuSbyMlMQ0RILtP3+0bBenfY2hSwbivvgnIo9LazvCP12REaxHG
weI2FFeScTSpoP6hDpr2gH7eIM3biL0EremAMULiqDkssntfKky9xz56iT+myBqv
XJIj/z8jDWNKdB7KLRTjq4RngzTcZ5AvZln3Ufal/3oHOUnyNdHD/T2+CHO4z4Nb
EnQXyXpXxsZHUKOzRcZX4ojK9H9tPADGfYjlrQlJk3LcYPuLdvglXkxf2hMMmlSw
xOXYl4VSZTcm5zjg5r5zEQDqoLPfGbDRgLNZPER1kRAMPF4pcbZF+feO45op6wqi
kEj8DuWD70yXmMIYVeZwhWY8f07+74Aas3VNTitMtFDbsKmkS0zl9wjMrZVxGxUe
e0BLykpw8RG24V+hqY8UrMPsCIO8g0TFtILR+1JkiJzDSUfCFtMyxo0cmbTilsZp
cleizyvsZvcTMb0XaNlTkgjXPrO/BQPQq63ueLF9ZozIQk/p3heEC1C4gmk6jp0Z
1CQnd7TNJPHuRIREw5YYTVuqM1jSEx9za5XbHN1mCDQzCZr2yvPeiPFFOwmleeCX
qabCFrC5k/rAoiOyw6ijJKhos3WOQEbfPEaLpu0C/AvVuzXK4OwRx7lm3kd+R47l
IwhdCyJbVJry/MNy0+XnGjrCEELtfYxf4N+f+5hniziTu834iYds2NoJYdkC9FAn
g6FCVgrr122xSqIrFRkWuScsGKyvZiay/6IbNH7AQoXTkInX8YktP3yeu0q1HfcA
UzW30Xo9qXrjsLzBe1c9BH0gve3Z0Gi2kbLC70C7+ygTrb5stNJk+G/ryuhIIj5V
mhWIp6hmGIOjqDxqR5fuVEN/swwI4ghV/MgfrsBs3sTRMYf0G1SXYlv+HRvnvoMo
/Fi0vqOmiu+8AngubHRJckryEQ9Rl+3/0h9ZSgy6mgHIOjNKEYJH8JITjASM01Dr
rcQogbaJvRoJkIR8m3FdLZpAiG636W1GHYnk4shlLFEmbzVn7Bo8tUXMoHYOSQ4K
6k9m9HesylMj+/7L30UEzdSXpqpVIgIFj+UXKz1Ju3KT35TEH8jdvungWWzEer27
yl8hVzPDtpkvacmIZcvOm2lxCw2aZ2zjRgDzm77/YtULqs2/BlC8XOrbr3NVRrRP
jyBDTqLcm0E+3TerteZeWg/ZRTlBv6lS6GfcG6LwYav6WNuW3pg0/nzPzeGMB7L+
I0fslpJh16ANdeHTbiooQWmFqqeHQ5a7LyfYf6e9mnqt72aTuAOC2pKEcL9vgkAS
xwJFsXtAkLEh5bGbh4fnmE8qghHqHMMgMwA81eWKMwtdwNuhncvFtS0EUxZWr2ZN
q/72UvAbyKsm9L1vloDATerdywEUseIOCajMUNyYFO4XEWjdK8elQQBxZsNGrgwN
eHZFgBuHypq6vGkoULukEq7mUAAUrBtVFjyjtw1JdaV67CT7+aJY0pmxwOcZuqds
8vn9kZu/0rXIz15l0slWO788CD6SqM+Exfu0GNQrzdeEnbBfSWJu+Sz+r9UIS9OV
nAUFBC0y+3GCWTVN9CHnMNjulzBGBEO2Pf+N6Yal92QtiAzdt8j1+dqkMnrKOCgM
DvLCowmsb3Sd5XUk7/a5HPJuDkoMV+xhH76aP9Ux7v2zj9FjbwhHMVsJaDdImSUh
/UnftaEl7IGs0eczhE5O9Q6DUHgcFK3/tCL10GDgk/rCUVoHdxXosvTcsViHJjga
hQJRLlopzGXd5pt6hkYrNZR8xoCLpBHOATDzR6EP3O+SXm+YbOBSXWJ5p+abiJ64
okxNGtMz7wF04q9ShfX/VlsSmGs82LWJxoBXObSOwQ84Z46YLgTz68B5D7sWuhSd
DtKX726NDDepGK3MzST/pclL/7AHHkNmNpW0CnQUNebi4MpajFkGJWCOqbEcJ3Wo
JOIpqk6hw/J50Ubxn+GpKMS5F+Kn60SVz+r2zGnmS0RPCJPQC457g9bg/AcvEjAy
fIag+W7w0h3unnOYpeyaq0xtVRrQzLqDXAo9Pn0za8KqXkzwQY70cySj/hRwhBlP
Y5TMxn2mJHMbRf0BC3ee1dofIyhuR+qo9ty8TWiyxmXRicNKzX2cdj+BAvnV4vjv
/uLWz4hHUMWOkJg5W+wOd6wC01UdLewpKDDrU7+Z4eRsGSYDvoTQXBENi+LwZuZO
s5xeewRemhw5OEuDj3YkLabFkUUbK2zQv+wfMd4MzPaIbXXZ2/WaZ70wpG1w7WFr
mfFq1xyueACQa5yTpwTNTsDFT3Rle6AN1MDsNiW0iFy2PPIGAYSKOqVGDzDyDrlW
FMj4M/rD7Z+8PWoJnzDN6FJ+rmqHN4W+KwXA6k/p/I79HgbZubdJLlN53dUxRl4z
tLf2ui+9w26G4t4Cz37nozzN0yqiuu6p1+SHqQYEdg/lPcDi/kbB+UX9OPPByWTn
m24mbnvzGyKKTorS760AfGFUmGhmZ6+c0gyNPwrYihF36NZz4VpBOs8+SjP20+s3
CczbVTzkqxBsxMImJaD1BK1igUUl+8tPwOpOb3UEGukYIyZ0oye/UUyhD+AdhEvd
/3XrL7xhx5MczDfPW7iWw97ylSub8z2Mfe+S+LAXcXuim9su5OG5zPoo0Np5BmDS
2r1Q54RT1T79fWGDcWLDi6nhkzKhXSl0DWCC6nIse/sHdl8wnLV1leQ47dSnv+6V
fhGAwPvn9Z3ibsirhnXlXjunleURQKsMN841ph+apYgpYhSYXGF3n2gTd54fkcQT
6xpNya1kJWrGfv5DznrI5iIrdCwRPC9WZKG4ngJWknegChQpVjJ75Hs5REsBWVJC
JsD/5W3AqhvBSl5mNEpLw1G4wfudOEsx0KQs4mNtFq7dBqujzkToR23St0v+VSCt
8GzN6EScJ5Ege+X3TUE0EJ+qW/OX6ltL/5Cr6ls5JQl69aZHZJH42uTdmIqcUCpZ
FBOKEVZrRlT7DhdJ9KQo9HNY7AdqqCOryC6r1uNxALZeyd4OUsJcOJjRRCg0rkPW
3jsBgxRRCk+1Om3aRaKyrAaLEefJqPeG7ohgyxU+csvMa7lmOv4NvQmrwip9qCaE
0sjsTeCNOahwitelF0g6djt2uz9LpsthcPhLie1+rvGsLvCAv6hJW7UVfFjvazSl
tpJClmWVjw8YaROuf48QYr4Id71DHdmUJHvtmSwi07fndyHM37PJhlUE9VZ1Ahj4
SQxR0v4gn13t/bi0eeNC1gr6pn+J+xs6B0yDSYK+Pp14cAtyw48COz7N6Fd9Bodv
x8XTSh3oFEhruCkIub5br9DsjQPRNCdi7N99BCSY4dF/4zH4Fp86kfVq3OhKj4PL
xj7/XHvDp3hUaPmbr9K0P8lZvgeyibMYMooZjdqLxon6emehNFr8WecI3WWUkwLr
9PEPa7QM/r+/CHRdObtEv2dWt9Zcys67q2asI3r5LVTYnhMDKrC+gB5owveik4L6
34nxPIPNZfgUt1E1j8Wsbzyn9i9CzqOIY9i5fEtD46LPfQE2CjQjPYCKEjeaZeRp
wTYdJmpYprHbDvkxyWgwf2jV2rqkwUsEXeajDbln43WfQfiAKx65dAxkuZU6YwPG
GxVjYoxNKdkh2t/Ns5BwZY9AVCODYZDIDOeAKe/P6+6FnGw5ta4RhUTbZnQK+8ps
eURKyMBo9mcJ3yLJ1k2OVtI5vmuUOXWD067l9y5HkRVtjriEEhsH9ewDxpUZaDUR
sljq/mGH648xCaPzC72/kYEdo6FQHMc4zjPYBtJetGBUw68G4puNK7leteSJhAz/
fuB/VD13hB4TA7wzshKGyO50U/vAsx+0qD2ncCYPo2vVsPy28jn1nZKe3OutiqXg
VNRY8f3yXqCqQ5q1mp8eMFrRJb06PqE0d/o4q2K2GGMRRKHIN+kiP0mtnf+Fq7Z7
CvE0dciKyGc1BvrlcwApEcNWB/YUrUperF1IKOeGBQ08Hd7Zko1s+6HK8mVF0Fgk
ofTsReLMKTTE0mQGP6GlLKj0pDQhwAnDtFjiEfvoYncQJXBiZoGbA615j/23KJI1
lSACthmk/pqo8qtoDuC5avk+cgM9wDuPLx2bWYZJU4iklmHxkyxxrJPmXZ1Nn1+E
BlZpJzyj4YOhxTzpf2BOmr4Yb75dL9mMBUckC4sPZEFxUBsLyU6PJOcoxSO86mIl
3OrNR9wWXYRbt0yXm07UtLwNUftkkzexvvnmFLzK3J0B5W9UtnlCEwz7XovJGUhe
Lkxf2K7stQPGylRO7SQ0xOD4MWM/rlOXjXnkM8LGPyY+WEs/bIQIM2dy5FnDX0b9
QsdDShJi/DqqwDg3t+OEcKs418e1aGizwmrDDXVcuTx/OYtwhcAlxLYtB647XAv1
3vl2LDHESDpGkIfqf81qVyw3jjXbNRCJX0qai7dP6aYkR5Q+8q3btBuYbH9dBd1x
DWH9SLIsWolpSMkxcDhfr61ibSAwUEQr6vNJruxVW31btme1S+u8F4EVYZ2EXNsC
97B5DZIsc7Ms4+ColjYg4rwOv1sz++YdX5xvWfLvQ0j1xQLVjgsLRbF8rq2IwJQx
p0ARzIYkkYPW7z5AWeoTXeZutUkzmgMJV6K/pbJtagHcaPTiB3MryW5Qk9UJRjbJ
ALPq8wmhqNToBvCd+37TXfkA582rp3DwXaD9QY7z8bCVp8N6penhkCe6O5csMatp
rV9zUGvMulBcxbfSWekAHFwsGmKpIs2h1TTxdpnxUrRJfoRv6KkeHJLnbBBTHCud
P9OuVMxVlKEXDNwftApRM0FG5WKmWfl8t66P4jAGgYVkABM+ttf+Cv3wS8qOo0PR
tQaco6/SWzWJ2zxFXST/nkSBS7J2cPqiz8dZT8vwvmapKA24sgIj+6abogYEK4hO
HfOhKEzVk2NshJEq2rgrYaWEdUr9NSnCYeIe1Yg0ALrbSGdnftIpYjbMHr/1NKfm
UCLpZDWA+6UIfT3VN1CgsDXZC4qBfzNHXcj8VxhIZtvuunc7WNo2ijruXUycFDKF
rzqKG6kNbaOmaRHcdj8vPrLdyD38LGSG4q4krhnYKGrD4XKGwmwtAegfHcan7BlN
t0s0FtSeMMIY6EeiuZdeHs6AZbqx1NyB2LoWEGenk7oCpag9Qk6ZGEykuAw4KNHJ
EOPv/sJ8VWn00pX2DhWUmceR8YjIC1uiUi8MnC8MJPI4vhQ+R/IpNE1U3rrAC5F1
kavfrmjbZrZrmHsayRrtetZqrI3TY8HE4vv3LD2z/oCbZgaBYndwYkZrKWG6k9Qq
NrRKRVD7GEG4jpSe1WdFZiiUr2n1FOSmIZL0jtEPc3DEJj9mgz6xMpfPkBD6LkCl
0C2+62dFsCcwEF+G9lmxFfzJ89xxoSw2Lw4BjdUfMcvCsGuxVfsFoe2/khPaAtqu
G5rrRakdc374iZzeXNYPsEkK0YOyYXSAVzcsOrQzAo7JaOR3zKu0OcAZehG3tjHr
LM4wEvJToN9HhkdAdzbP2hB3Odu7UUJuRiCc9oVpHqDsYsGbTxgGK85YxbDVngp0
8cMIFzm2SBzgyA1m1bIGfw1gpL1UCh7bBf5GhRmAqRXI7dMl11eqef/AFUfEv6F0
TpQVnxnGJoPtwf3/86Rm1LqpP5nwWYWJDwD6jcDs84NoDotzBW8GZQ7JvZ6kCrUt
P9Hf0MINaFQtIj7WM1yzRDsTXjZc+CdY62z38N2JpDEr7gaCHGwmEZzL7qBh6jdS
Ogtut7uoEFMhGROKP/qswtz3RItmIaxsF6eOoR0pcOm7cU7vunpZ8u+8Esijftqa
O5ByFL2IUAz22dbjk+Orloob1LhZbvLiKIi9pNCelJuV2jkBmWcW1VrOzw7smgQV
OssQLmEiMImN8xTcRzipfwATTD1F0cKiVm465UUMLOWneClXb5C19UqYzXgJX6FZ
GkOfs2iGLGIY26C1L6DNXW4I6r82Q618Xf1t7A7SSOlufHbLH4g00xICsuithoox
1/ZIivVA9nJwd48ukNDb8rXhSaDg6kM28iG9t++UPV30YA0/m/Yn+6aB31Pg+H5+
CXRELWOPj1ZxRM45lkrNsx9NqS2QYcsc3q49MTD6hjPSnHLjm18udWkCqlyciwmz
yJJo0Bc6cLJwceR5Pz4s3u8+5je9+g+RJbvxKeafqnFkD8a0sYOjl2z/dE6L4Pjm
oByyQWy9gcifOA157RSdhMWdpnBxiHdFrdcyhmTOXRJGZZKSuCXI/SfezVnei4cE
d+AXV4rTbBgIX+uvQDoE9z0midZXv6BDcOngTrenOPdheLqFVRJSm042uiHB8jYA
OdU5EDdp8HadRRCNwS3kv3qecbNPrDYi1fuA/QTQmLza4B/uKMV2QqeFMm0ECfXA
xWae+z3KFv+qLe8aVid5W8yrvVLGmZYHY2kRAoyyW0j36XPxg09L7P8vUxSiO0nm
PbMRr2lbxLKHrdGuQz/Lw/yPuRgvgYRo+lIrUpeOgCRrf+BYZt0Br6z8VlRJZgaA
hsWtENm6QJ5U+iA1HKUokmMo6r/mTl2enu7mja8qgEkBQU4s1oE5hStWCAXe/pHt
hMs/5PEZSBCQxogczj6JsO49n166W79ZSlQMMgFqh1eXKhQTZvpVIvem3FP/vW2m
YNVsnHvrip7rpXCedZcVSTbVf+z+iDPSygsD46JJEkz/kwZJdXa5pnqYmQ2RpEeA
HcdQEJ+9JXeQjoYtLa7mtc2aDeB+ngFTnMpE/YP5WNNF8ssrA3YYH6TnvWMZClm1
mgP5RBDu4WKrrqo6YJLox+5F2PKBM5A1Ims0m49aTpT4Eb9p7XCswQgfBDswnX8X
5fxYKJFuLdrQxom2ydrdTboEVSyAz0q4fb5O5jXbx87RQvhROShdhJKA/dspUG8g
6bhEQrBvZ3dBFjpeEAltwg8iBwB+/5n9qlBq2WtgAEOxsMRbPQ06qMimDvKU99fM
ZfRAGDexIiDy18vGzYv5C+w772JXSV6bZy2d2yNsXPRNTpMnEbSmdVAodYzRQyN9
XwJihdMaBuavF4KxffZiVqEGNUz0eh1w+fX3+zVCTnnL251MPTXmNU0N+rj36FKt
8nRwQSDJzk2FSu2vgawNr5/oABa4WZo1yJDRRXLx0CWavUeFMB9DsP8OXMOE2ND3
hnU4Hm4cKL5zUdeD0HcW4y59IIKpdVXawoq2nL3pqau1fs3rNH12qPyhwD29kO3E
biUUYzzFImman3NoYgjru3QcCJwI9wWJjMB7Fru2GAYqBhGq/NP9LDjZG87zJRQt
fBxYT5gtS5q68WZ4ri/fYvJdLsv+enV1521P9HUzeZbW5INa1hO6Uy1d8iQ23+oG
0QpEzTorwhqyr9fhCLXxewBuE1GdvSsGP+XiprdOIUHP4aBoALROgOJYjDSEb0Qk
+u1zOl62exEDoDTUfQlYZ5OtVCYpCEEcdK48z3ukPSRsJWev7gq36fOhkV2+prkY
tHnb3am52X1blDXT2T4SGsEHIWcfSn29lFdElT3QnF9dgKegFIGWOPNcemk1Ol+P
S6GxCgr06NxPHhfFVu3/8CG1dNCAkNJDC0NpyzeFuUquUewHwzvc5fBcXRsSj09J
ulLeaplaZusICadtbU6vf98gLwUIkeaBDlmfFYvpxw36qFupllOi2bdtHcHf8A9s
hmvZ/1VL6F8zJk5Fhbum7b6YzQ+eB2n6o8MyQbRlUzlgJTN7g4eFEbCuPHWaytyq
Qni/0S/Nq2h81gGJp1SaP+O+UzwXJkbWVpIysrV3xlsyuUq0PXq/N3foxhsOIDaA
K8MCbPBo5H68IBgsh8XXeXdFRySYSGDeIols5pL1ydZKJT0iHOyJyFTv7TBumfSe
7Nt6wfVmefWn9Fw/n/94hDzkIf/MUmJVSH5gAI6Hl+caZZIk6a/9/Yh2k4QLAy38
DDnOhwxuTqFct0c0D0Lau505Uq3xA1/qDEHq2woVOP1pLSGXxCsKLTfTJf18MoJ2
XpxqbDF9uP61UJy2Tx6MjhShyGiCJ+K6e1Xg7kGssFT0bUkELC6P5tauLB5k7pQi
0psU7mjur/Io3GsEf4Vnc8Hp4fZwjF0cjqKmRqrj+oe/78unMHkc7QjUH7VH+PtF
WyluJTKIwUUodDx0OeLTvW73YCcvVF+irgZmUyv5HcMoW3T/wa+nFmyIMmJ7UBUO
yMg3mdlxKAHNdk9uVxtU4ZrOWZ35RQ0kuRrVq7+6myJUNZvv0uX7g2fpRwMY0mGF
G7ckRNCxS9GWoAhbonz5DKamgx8azrfbMKzCs83UAPifFlviXzk6jwcLroDin5Qk
R7NnswaPIO5GpOoMWS+aDeJ1Pvz4ujbUy3zKK+7HOGxOCHoP57iqm3C8Gqu+JjFN
6CML0CkJZPRUaht2HSjKwN9xGwqaVaJi0xAupKZoEiUy9zc6MHlh9/Bt7cEvUm3a
jmwuZ3do6mkwXnKuAHVQiQ1mggKwEzec6jyijPedeWVSKKQHm3+OayzktC08N9Zq
uxDzBXbReVm4aGdMmXs4wPx+VZX2QuIiac85WWEwpNDnsfdjiJ+325fDO2Qz/UHk
ooLWQjPNkTdkm7p2cUmMMnUMvEHsdxx2QKqZFbRvRBO3xx3OLN3V8DtGSVxutir0
cCXqFGNxPzfqnFGNcgU9blB6LPDbfI63uj/o+hgz06bVmW+e66QsHhhb728mOfPx
5IEnDa9RXI5AZJwW2BPKvuphGBvk4Hs83O0RUzBRjRJS7BiOEaXhpBjUn87ob679
qeqKmj4C62Xu+b/Hl9Gymq6vDxzUE/z6GEGHr8rJSCAX8/rEojTENJ+PBQaOqe6r
a9BTyKemSVT/8rzlP9i46CAfDRgiOzWKSox9yV+GHvYW/uexfSrzmVk6VKqryxsO
ZuJdgiVivi/NwI4xXGoVPC0kG1jNIwzUfnkaEEacJKku6xo76S0x2T/Oq5kg/pHA
JNe5eVQNI7fNQrP32SH3DUpPCVpQ9IZKPMvfx195KucS1bX3a3dGGRTPP0czpK8X
ItB6QRob4zxTcqmiiCZORPJNshrLpkDN5TpVax5B3QWp9jRl6ob3e6PO+bU1zbtP
`protect END_PROTECTED
