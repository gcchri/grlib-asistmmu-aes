`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CajwwpH7Ik4np2BDq97+LihBDshPSk9hNzi+f938LNmXwOys5jPoEd/0P3Fa5kgr
0gPIBUJRbiE3Ihmz6UeNnr4mfrKDFDyDVKVH53Vj3d6j8m1mwJP7CD2FbGcovQFq
kRsT8EzCPljLDKyC6hsZsGjMkEeKfwhgB1g6FzkFpYjonXMyU5O/pt+eAD6uREIt
56ALLTjimXhxWQSi1T9glr6Pi2Ztro0iSfAHCTpP9x5NWU1PpqzUAB3L9qiTYftJ
XdLVTaA2b7F9D+M4q/kFMyRsNZ1lCZ7u/JxO5k0l7cyl+nO4ClqBSpJfUEwhQYQT
j4IRgiOUPqS6QhfVaCgsG2XJPTxoyqMLbUTUpzYUhv0vOySpTvE6MVE8YmfEKakk
qSyyKVernNWkHdKyS8bJHOw1NXhQI7zHdLkQ0UGvlCS/E47Ev1zDDze4gndFon+z
iYUZlVJDY14ZEoabdMV7zVw88609IOh4rTsrqeRfbESdU9vFOQlHcb/KyogaRUGC
3EOsRnZANPt2YJYlgWTSnkpqtkutH80C8TaJsGvtMf7EEoXiZAfMVLzWXIVdktAM
aTfKLKWuybbNhB4D6OTFCOXxxCBVsecPD4wF+3X4+bLQC95APoXTsGiKAK4nvtPm
qxGyfxmPfX6/z1lhCK2fydK1JDXXd/lRecZtVjbBxfDR+Rlu/7NlunuByjaajuIw
ixdELiCqZzp/4K0lf66vg9uf9syG+5YH6/69vHubOsV46EFxA/menHKJlufhGjQL
eLdx50n3KDFGq4KYWmx9eqoXsEHH6QQWwAkosaGAiSZLxVpObJqYLO+vumHPFnRV
IQBznX0Gi1Ji/GyN5RHigfQgdzD5FUtH1+dbitnmXUbuoT1tK8Gm+ZrM/N7aJUfJ
5hw2yW2GDh1juDqgBNctzdOiXgeWQR52FaNWxHS/kJ6NAYxb0OfT2HTPM21b4cOb
Omi6rcvMY4ifcHnVgWrtsA7nGJsneZiRutqUaWf0kBHtk3paQAmp4Wlvt8Ky1Ho2
TGZPvyMgHYQ4EsfgrFfdOA+H42+bki1FpCZpxzt1fyyT/b1Sg+TDhTmETN2qlGAS
XVAgSre0+TSbkItkZDBLms7WbMcLLrNXUHzZmjjP14B/QUjPDpu/s5bloYxZafo8
wE54k1W68cM1HsqTjLJV4sNJYf03F10No2pqzoHlAum3s9BXkFP6eViu8DZvRcaa
a4es0N7X4RAUOKh1Et3S2dSkA6bXwJtL41caSZyf/avzcuz/bLBZxBK+45aARveY
feZrrT9BuMyhdvq71s4ZJmryWAS7kJLmLYh0IQ2TjdTo/lP3qRFVjFqdXdzgdlTB
TenOExyvZz7HRZW1OJNk8+7fUw4mSwIh5FJqc92Ucb5pAq8yo06HmDtxFLQUKAYX
2RR8vxCvLq3EvJblq9HZ4QBDBf6w1UJameT9frbraGUhmG37itGr+KEKoWjgaiTv
xWF5vlth0W6iuxf1958kdVbBIPdMh0Uyx5d04bcrpR4fbgDWDIKSRNJpDWsWIssx
ORrBr1HJTMQ9TPECkd1UAX7qcQRmn47LkgXPIGJtloAHAoEI8hwWcHlY964tWzMN
I/RzhWlTIuxLaLyHm+La3F5XYeITbZTiua6jQw0RAIdKL26rYq0eORDXtABgalH4
ZPPHxAM57ULdBIbKN09Kg6LgchzDmvnNN/tcWDDJFyp/LX9QFp0mIQLYWJCCwu8o
EtcHb/dgpoluwIvPQNLDxPQx03c0iPXFI4hL9/+X2vpHUr90vL+mOpFJtc2/WHc6
H779yK5AfF6Y7P/1Ti4TVxxFF9LcGWTvO2pMSARNGNx40J4kKsGokic3eQdAhovp
sXjLP0htMBsESrfKEwst8qL8qpAAVZTbtNvUw6tLROSu/al1otRbMUeMTzfC6A+7
Af5wJFsax3uOO2p3DyP/PUv1HbvS5vi6igxL09/TpdPh5g7Gkm7JifXy5CqJ9L/T
gRZX7GVLsjtcdcRljzsw86gNkA8bd0mKlscEOm0DGCIoI/zpOws+AZa+FhhudWta
jmEf3L5Lnsj2i/3HRe+GIIn5sP6yzubOPmmoh3oFtQP5fZz+wts8/GHSCokDg8Vy
A4sQZf/aMAQmqHuKY/8OYj7HQNI0dqbS9UMCvm1ox8PYeU+cImg6w/0OTmYT3Q3K
rnok7SAZ7l5NPzjz7LtFXic/5qcTjxKFYAcIwNgAJ1wkBptrtnp+IQmtU9jyF4XT
dmGcjCD9zEXuEj+UO+l++BRFP4qoJAbeinDxj10FZYS6P6zz+OOm2sey1z/nOGxy
j549QivzartU5DoQJuaoUd/gBujXozXkkmWEDbdHNl66OAUyGSWaLRHy1DzCHCAP
71chcOEYGRiJvoKNqlYuonYjSYKLQVYZIggjYjOi/JzDeOaaqQStdjTgr/CiQVyu
D7yMzK4j29vwcLBcSmf1Kw7+U5kG5l1jFSmXFaTcx/sJRTNDQnXn9PgmV4WroPF9
mXwDgCOfESOmC7hiMTIxhK7zN9GbaUKcVZW77Q4EwJPRFdGeS+nniSopW0RSQhQd
pI1Nve7ZipX8coPHMI3OVUXKZ/Z6RQjZoDYhI3gP0+WFBswUqNO88TxCgGA0TPU6
iAjVHwxn4+OYzhjOeVmzvm3LfGgkDwu3OzVoU+rkdMEhp2ETO8oKY+3cqhr6v4Hp
jD7BNXIVm3jARU3Mf9HGl1I65Ig4SYImXUfsd5tcdizvJfw8PwEWgEHFPzCJj0g5
7n8qUxHxQCBshlKCIGVfGUCpLhrNulwKp08y+StZ4Kc+r3V4ojuPMlhaK6BU4Vi7
p9fU19g+MXOIGAb/SDN11eH10Lx4luhsCAU/nJ/XSTM7pI+ckk10gyOW7Z8Tc+jr
Rl21H/A6XUDa1TgXqDtmiVV8l5hDobC70ufl0Pyk2hVxGKYOrUu03fk/0Z3jljNi
qtC+iuxIxfzsM6iH1UQ7nzrwR7AqOzLcD4AkkDlfEqgTRRfgWYZS/tXm10MLal91
dmbSo9Di6R0FXCIrMrInUHON54suBY1NjXk14ybPY+w8Dt+jLCdw+5AR9UE2qvES
VALTtEtx8Aymm9kJUUVrB0/OrQedAZHrwTRtpe1qxX8xIICYM0FRf1ZkOs/Mw5W0
JobLQpts9F/KDd0EQocWQBf/hnTxf/BdvVkxjrcMaWWToqBaZUGMjH5dFNypoZH3
1AxB75cMaQdVnJGYQOG5oekSB2DiSEGRfEKvazshwjf833JMLjoVI9S3yMaiemAg
pelT+2OIr6gC9vGh/uOG6eGhP+/WUF83su04J4xzJVMSsnQdVub6TZIsAkEnAn7f
JvgOTSheWopjjugwiHablDXpIoGJSyWgkHtkdOU7NqpnS1eXUrOfrVBQ/RkRe/cy
KX93fEm2fqNt8FSAuoVy9nv1xQfT6evadgpAH6HHuP1+DMKPYaCvAPpVyoMMXmGT
T9IUnW40O64vwsM5vAtxgj10usTWlLmnTpqoc8Iq8Lr31lUSBeuiY7Fx3ccjlkS6
Gws7e46zTYPnX9glaM5hSTbJGPnFhClxz+5zk+M4fK1uHwVzFOBlXIErrVg+k4LS
M4xlGDLGXCJfSGp8FObjm3tXwO8VWF5jD//fqX55BHrYUh++8fxGyV9Z9BNHqXUi
V2Y/gn6fzhXaFZXBdu4yHKE6VbtUxJhcBbUBYmrC/Ax/p31yF221u3JkLdhJNAEj
vw5fgKl6+lHDl7DXbEtJDI3dh5fJ+ytuQLtoCCP3K6/mQYN7PGwh4dwJNcuAIw2k
duegcplpd9qIP9QyN2OhixCEOvna1crljzSeolI4uZdPT+Y0U0dSfxRvwmcsUNmP
uFZzAoISWTpthJd6XYGNhdzwDAqSyQJUgJDO3trq6/NP1p9WnTjI3Ujh9JUVx643
PXBU3W6N5+P+pJiO+huw/1gvqhjuva81mVqX8kHeEJqLQ+tN5lF9cdJB3fpfOIyu
1sqsg3uo3i3asr3lkFh3Zi02PbotHlNe9qGKZtwmeaN7AGhPA5URbaM7rF1yJXXL
jS2uPXVJ82ctU7oPh1lEkvTyMrIbfl00p4LnXk488BcrxXtVRqIm0w/OxAr+NH7h
bp9qsHlnMuoz2gqnBCWwUdWPAtRFd780MPciolqwO3XKLtN+KIbLMfVoVdlrFvsn
3ektqgQ2Sf3wJmynROTXfSNPBVmAJGdg0qmW5U4+bTS2cwWoJaZZRs2H6LUdgSjL
SAgBRZf7HWyiipI0cIbGRYF/3aj81MD5gkArPbWbMyWyjlwabaT3B1U1SZADSkKV
kxyZD2V+VcIl6tn8aTGycDGVfaYd/SvvV877LakMabG7LfwXeLPzbJ8Ktgw6uGlR
ySx6eO9KG+t91HJQt+f/1jKFjBYGOVlohcWLNDdf5mzzx0klAvPworyYZjKNnZrn
tBslM+xFbOh1LjN4lws27IFZJ0WZ4WpDciztnz0lpJzmBIZiK8tJCo5X5tcXHIeX
e4q7+Z+aMZFme8gJyLtK+GQBDGHkODvnRJ8v5zIOs2b+BdvRI9X15WzrT6BjuyIj
pdHq3yFP5QXlPMsdvOsL5ZdNsYxoOlqYKg/4PG8OeNPlvBn8cwVMN4yxIBXEP49I
d7HLzYzB/vVeW170BbB2koCyRuNwGNuGkdQmXYktZKEW3A9bBdOc3Cjea35u02+T
VBKixKeZkx0FfeUMspJ2ZQA+x0q2XaBmAJEjIi1br/sab/xz75QUyUsqiXJMYDkP
bBAWtMA7w5I5xu9VFynKb3JO3ux2QZoApyLF7Dbh9Jo4QfVFu6PIsr6y8+rY5V0M
fbYD7z7RIxnARFBPvSc61bP8h2/Z1tGMU+ic8zO1K8GSEext7iiMP21vBzj8165o
WrQwInMJu/ZDyUS7yY0sUw+qOju4n6ZBVs/2EsKlIFJprOnU2qEKgrfi+qGVBFVT
isUDY9kX6r1tnv335BHfpasWa++DGtPdToQdjRgS30ukSnLGmLQ9xPA6kcbOKsDj
TP89X/AivxxitmKZ9sHTDa/pk1DQTNgsljrTVqMtyogd9snqYW+PcntglU66HqTW
sTvjpmv2JJRPcmciF0eBBpUJEgk/diaNoLOGdccsIzcTaogeg2IHO9avDWLYB4gl
SgWVWPWFOl/W12f97E0lbQgNGBqlmQNKetBOahuQIagisxbuMOp7mVIYwsGaAste
6TIyJTIeHbVeA0gEO4pKBB/B2c5naMqgY+ELIjbu00I57XJiDsWKEzTs162nBTFg
b5cB2fNvtDTSnnNPMbYSBFFdL34b/7b7nCMRJ6XUR6GVG+FOwD3eu9ktd+vVWGkt
6RZdvGsKyNtARz98T2EkONmfbF0QWvzRGE7IxguGGBa3fhh1aGb+Pe2rj4wUFbaE
D2IehOmbg3tXhoX9IZeJdBevVdJRoNy+dhB3nz0W5OxLVH1mjCEMV34lengOEV58
B5s+2yiz8JELnIzpn0VfFLSbMU496efIldUiqaJowfDoCTywtG3o273OgbE3pYeI
AwTTTKwjLKEL8Fx+OfcdMIed+EnhsN+YEwPnigdeuX7w46BKknYi9O+sZAjnI9zM
P9jBiT+Lzt+z3TV6svXzT4pjaEPuK/z9REhtPKXOqyZAVJJJKUWQeAnsX7C/N4rV
8+UUPdZ8/Kg3jvLugGwValWWIxYyUIAraFOjJxi8xXHgKMfscT34iQMSvhcKxq+C
bH44jzVrerleP28hsWah2RZTLYjmRdxewmncDayVKeHSCLBXQfsrgU0ddBPRqDVY
fZLnhkMZHXnHnGl9vSPeIoy5pjlaAAob21ehlkwHTZNMtEDba7RYC1YuAwaW1kmH
7QYjadSG81mi5yzHgS8xPFK9R1lIIMHxamMtil1X3SPXfvgrBz9+KMqUYihu4lMU
SP/Qp8cmW4B5xCX+GxKmNUzzzFcgvlJEGqbGF2J0ndK0MWk7sxUO2vf6TfWH5xh5
SmFF1eQeCt4yJXGaV/Fiz8rB6637l52DIaXXAXQUkUo+dJHCq8gpSOt8mwv8489z
NRMbAe+YuNaUkXOVyQdvDqwcdLcFV2fpon4RWHDPFLl2JHudZG8LrdrS5oREXMr/
Jc3R9koYQ7RJ6/uIW+U/dnsRO4pYbBTifsuXdciO2oduPqk48sLzS45s1P3Xf6SN
umJBBtQqYgI0oT7hx0xhemuAKokMZUfmMgIiznXKgk3ytaFdwEsxSCgT33aJfBJA
aVg6fflwNQHsCoNxbVkwj8N3S1aPr/KxvdtiEoPYMrV7Rl3RF68fyfb8ILBTrit+
mFHkt6QzZXLQeiGWwDvlhDX1Lp3Wj6LXqUSP/J1co4sz72TfSd1E674dffQh9xvV
L+bLDVXIN3wPiDOaF6D0/Lsp1zNvjsqPJDadhsfkOVkj9rJTouZO02O5ZAdR9Ao+
ayebuJf+Z5yHIs1ERokHNJIuUW91FoyB62S9WbX7ydVQIJeH236fiFQ+odGhrUSW
YfG4jJH479DKrm3Np359WIh6CeHQDxvRtVw72txN/hR6ZXX/v7sBT1857HevtA35
NlaT+oeEh++Nbuac4bKAkuGkDyN4T5NSBXHga/4HientFmk2s7I10Z5XBHISbQdG
tje6COg3i9VtFRcMOpmktNm//sSrVTFwA8lY0gK7KTs4MO2pKAtlC/rPFQfGsSmN
CiN1GRrMzwIaJBowkVKyLkotOt/3TZH49YdfsqT6UWDM0GNhtA/6mF/TgrlJPxBr
nubdf/x0ONNkVw6aHA3RZr5+4JOvF23gCOSi/UmjxWiX2YMHg3GnrxnRo2UnkfDY
6xYEgMw4As8J/h57oTq0heGzUkm5HWpyxFi4zI7OFd/gE002pkWg583RHtRULbGs
YxueyBSD8K1zr5FLXPBOJRalQwv5jdTdW1zsoKC8hgPcVgej7rPWhCzZ53kENKry
ZCF0mv+WL38iS1GmGVqyBxme7YeAWzTPYqAv5JRGsz7A6SblxinbmR2Qwt8UuG6K
WdsmKCQQ39V17yVFoXalYGhEWkFszu7e6nfQnTxF2hScKmXYJStff+D0vlSIYdRj
a3l+29gIxKpbdFgYFiuo0jkP814t1mvw3xyIdcE8aL247/ktB2h2GdUG9U+X7BWo
/PybESC1pcJq82k0/oJWy56NPh9/VEn7dkTn0X/ucSmQTORHTQ+B8pQYizjtxdMH
xGm0DaB4e8VUWOjx4Oe7y2Gv1qeI5aottO5mQDV1WnW2ao93XcX3lZ1CpJG7msCg
lE6uwBGkm03JyK5Qhkuur4x2G7E+0987vEqfzW6XziBIQY3aIdX6/yZW6MYqHF7O
ejqAk4joOXXDqA485c8t1AuaaY02IAiAyFISVgSAXBprr4ckAiLfBtBFO5iD/JKe
mJ1QTVNPJzg8W9Df1DIdkIXGGX2WVNAEsmPpUhbto2kciAuth7gCPA4sAixfDgZM
hT7Mx8S1eKzRNN8AZZMzODZ/43nscF+rYtvyQ8NQb6nOc9d/MPKdtr+Dl1z2haG1
VGPJTX6BFU+KpAr0Z/JFBVAV8epLBc7EvZDVH9JE8M5GB6b1DnJScD/c3JkqXH06
v8wJEJ4lbGtfKXJjQwiXzWc8XSUlNJYvGwOXUUlAYFO4SqAUlrGGTlDshOgY8awU
tmLdsvu3LeU3FjfhhIGYDsXth6geaBuKniyU0uIp6H2xjQPxI11iZFh1tn7/ribo
AVNwLKImVkkbsLFzmuohTY2eKEl8T6dvx+wYfDDt+5gPZwEKMdqyEcIr8ck3DqB8
RC5rB9xcHmJ8HIqX/g7O1FmNMZIWaSof2A/Buh1JLFI0vVXTtKi+x4D8T87MiV6v
zwfzhNuoBOIYa6i5NtPCT90wHuOqbm10EYc1wDAucSXNpTJT2TDCz/EE0EVpfzxJ
0eN8Y4Gr57nErIKxAP8Uedc6lQoVliAuPIR+M/7lQMAKRELFGcHhEz0K++dDm52A
qT83gHjNemsYHzevX0/yliyyIJCv2UsLPb4GYf1F+ERCDU0YIv8LkD+h071P+yjU
YeN6KTFeqm7hYyisDg3tSk4jlmzWim5akCz+f4oOBwBBtxdyI7JJt4UC8VloRzeh
OBwPQqKf/2VOahfbrIkdoM0X8yXEYfG+oVy6ksC32QPBidAPhW4d8oV3LsveJJDL
V2Bbi7P28lqGpO/eXz9ehS8ZFjPnjIRSX1UKzudnRlF7hDUu/xlugQWo6+WI6Woh
SifcDbePIhX5CzAxvAOk31trLLu36p7CvSl9pSIOG46qiYnF85NhIclKG44OznuM
kWRtQyThZRN+xKp9xnNxDXTgeigUJ8EXyVcDFoAGN9UggRetckYHiPciR0P3Yii9
hjAdYWwmfKFyMvk+fBGGI3IM4d5DAZz8VYgOeJxAsvJslTMMxniCsrIRZ9k2wq0n
BAwOnpQ0yOSIQ+5fN2d4j1mpl0LJ23A7MLx5P/eWrdMBBpgHXuBjgqY718tuEHvW
chRZV8FBqybZ9ZeUfMfEGOwXsiFmAknRaxsUDMaQfTHt7ShEGgaadineZ7Qfa/Av
6GqnQ4f98bltuB4ioIWh7aUnhKRebrsDN/t4eF2vf8IA/W4zxCZ0Gz2jee53fsKo
9kNG1srAfDh98CjGYq4TGsOF5WugjEpA1lOMEE5ArjA3ux67EbDiRgNbv24dsptf
ApqV2dMvNHQXR5gytSBj/ShA/Nko/rRodZV9Brz2NnLK1FSEit5n/X4KW6Gawtu0
K2kaiYz0jjPcW/VWH86M5FvTPAMiE1ExmCoPFnuFF2pwMvc3XDwCmFwoudeCFwno
6hd2GaEdIC9h1Bi2bk9S+vMTz8yYccEoDTcgXCSnkA31ki7BTr5AAnMgJyrJYp0F
7ADrixpzqpZN794OajWDad1C85AK5PUXkprDHKza8nKPEm3/YjTMcAulq8zPEZIo
vZeY1KBukmPPkB4pREG7Wn5bdKZW8A0AzCKS8J/JrDvM0U0AnQXHI8V97isNsIx8
7zPRLNrCoVmBiqTK8ieu2eiCiTx8XmVxZDkZhjobe0IciGGZI3f0RDqTymgXL+2A
dXWvH7PHAzRLKGb/4CgchtC8STqzXpPshavaxeMIOtzH2dBJshw8QBWDGk3Ry1Az
02nJ8grqnSj8QChpAdLcakAuwym5HG4HO2jDnIkFdHeXYR9lDGgjPIN3Os9CqPJW
APjwT9EDHSSlUJTmJjRVE5qh0n33dwsj+v4pkplItv1AJSIbmLuaBm72gCicO2Rl
YWliKwtFF1gHY2zLTb4EfUrmUvxFCVDumjqECNrDNb5gFNxwSgEZZYU9wOwofeoV
U9Ah76GjSd3IXiXYfSG2gfz9r2lbbZ8DajIE/BPRamZwtzNNG+l7OHFjUvU7ehEj
H4UVOe8ReDiQgWJ5RXZSH69Pa6cTJrT6AHXp5rXa3Mv0Ee+8E5uTKRVZ3dEdjQWK
yfrfICJKJMVdSjxtaTnk5OTx1YzRIRG5c2WPMpGW5KagmiM/klgukm1ReTZZPdwq
9YXR6Z7LQONOSJae2gtJdiT2sJh63GYaoLmgCC34u47MjyCly4tBLpTFa+jE4u/6
ecjG3O+Pu5M5UNgL5ZRx9QJQCrJBNxjvKplUhSQAza+8rCQh5mnj7rGGFpSeIh/6
KhgdoQqVBOG6ztaMhODql0bzPHguG1LAhegJViYXviRWlCoJMsW0Jsh/xO07g0z8
tJGPCoL+isAhaoE1aFCththJENVQuFHeKR0mFQR8mdJpB58afkhRa5w+vXZ5OCR2
ug4HkfJ7FkC5kGMtBMjd2fDzsoTopTn9qkcPWCqV76Ld4GGUQS0CrOiSlHQ0Wrre
jGuyml1YlerXciQ5ntGQDi2NXA8X9AokgYH64zCP6YdtDY1YKtWEffxGGdyljYAs
2WFBdsnJk953al8tTMdluWfd8KsYfhBifAjUhsUUzUPVJ7vErxj8hvnXKuynGJd+
EjlR03mOMXR64ID0WSPveD2rNrsNocPR/7da0eQYdxxPQRSdMI6vgFFn1RqsIijT
a9ajhQM+fCpR+fza3PFNyJsUiXdzJ2WHejL9n9WjLEJ8SilJhzxm7eMN99ekKnq/
RYz0RTd7rWuH5QQ8DMg4c1sSLLPpIiRzcHedBb67k09finL749Xg9BzhAfWNYAB/
6eb74A2OH8oE3Wsih56BzePSKb5cETxdm2QM2IwanuCRCLpzpV3BBAn4vl3/c38W
ilmUJW3os/lVXoUiEZqNR+NyquhHTINPe00NMCDXSUqPtTWtqD7Z012sP1skQkeL
95swfnNd2JsEGcQdb4tjGjn7I5sHihpnzXYiL0c4d7ofVyYa3/s6RNUthdMSvSXn
lHWBSIlHQPmfQz+QO/9QSBUx5uxOg7pdrwPupIcnCo8jKfrDNDjVDQcGzVhjAAUO
pn6f0H2U7Y9TFT6cpLTyCvW1+moCLsFoYGFjrivb/jVwkASpUo8Jc0HyX5t4nnot
SW6dOYCpK3h+445UlCvfTq5zkyJfwY/CSywZgcODS5frMUGJTE4uRf2o6lC8H/yI
krRGxbrckXJGT+i/bmzcEdsiMVukQbmBCZRXrsfgYOmdBgNUTevgAUG4VFSW0mZP
n4W9S5kd70Uzf1NomB9XBOmSfSaBHNAODxxKdWCIoxRgZ3V8EoLYGFpAdwzwy6jf
AWVOHs6RBzi+YFjIbbvGyr9wv8JgOBpIrGdO3goUM6/DfV6uCeXwKXCKUx3tiZNv
i35d5vKzjFC9sQcWMC/Wym046StBQfcAIqZcLkmPDsUU7dbLb/yS2yxQZ+fsT2Af
I22AUcuYTBjabUPjDBIvhdQ5friD2wh++DEUsgWhsRqZd5/FC7q/+ac8bxCTjTpb
0Y/ptXO3EqQH12QCv/J4y3gsX2FviZQTB/dtmsxv8nbbLFPXSbWgmzhDXeuNlqVG
lT1WjCjOWNNLI0Qhzdioos3FDwtQcyQOLTDuzdq1sp13UEN4llR1SizfYmPvkbZi
vQKYnH2uLqjAE8nhR1PITlBvhoWkpxAc/bMaZxW+K5kEWdk2dY+Up9/PQ0Qh1Rkb
Bjc/wSNBpKU6pjGl8AsXFypE0JCt9e1n7k4ciuUah0YHH/O/xquy7D+zzhOZLeVx
CHCTFAcpW771dAeFgOy2XvK7ZzLC0orjCxGBgkdzQw1VtNJghC9aMIfErNYi5/a6
TlBzk4l2Lyltf68MGsKgGCYhZuM25kSfv8IAErSFpInW70sAzbH4MEZVf7OiYTb1
+U1UHBsxisCQ9P8JhsTUU4kOjqVfiWLxps8y5OyZLZK33PHQ6Fbh0ZMoNnFj1yXA
RyDcST2KVwOzRvy/PF8DNXfZT+2LMI/5a4nNhVj6P2qV6zyLlDPxTLoEYSbQIQF9
aqsggCckV5cBFOoew8cgQ3sZRx/Fame0nU7+zAYBBGU7mSvcKdP6jEua0RCBNZYP
BVRGvPrRieNV214YqMfVqAvUH6VQ3Xxyv4tKOOkR1GF9EP8eB3ekb8vARxGz9C1k
cTmUAA4ow/iyXzpRSPanGv58ocLZoGDgh1uzIoLjBTSFHeuLtKH1/gENDVcD9JQu
h3Agd535K7epP8U+YBu0BHkSR8YmkPyQ+hSk8mBemPIYptclCxzxFihKJqRkkY+t
p9skDpFRtQRjnrhTJoQvr1A2D0Br1ASEQMhkW/bOsY6UkIkL1kErmTEECEgGcCtm
dahnETmHRFWSsCaX1KkaZ7xOByuSjsEQELN4FAQPO8sxZP7nF85ToEf13k6tryUg
wPr8kycIGoVHbdwUyRNOwQ==
`protect END_PROTECTED
