`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z1xY1WUWfJIyvzRJcxs4/meHjBuETgIjcxRQSiNVsPKUsag6PBX66FcizIuTC8YT
qiAu7UO06eHZUB39kaZyfPj2f2f+EbOAeE6QQ4ezYCw/JG7A+9LEagVVX4LZMoyH
cUImJBU1gcK8Y7F/rqw0U4JxDYPxp0N72b6N8G1peGWeJqvgcq3yFw9Rm1xSrgCR
wjyw19RApegXbzNxPtLwLs8hIpl5A+1T5wybBk7Q7TZ+f3kmT+dwGIPFG6/1Whrw
bpucYPedNNs2Q1BFJZwPwDFTC0zzqw2djUivJW/jJy4PP68/I5R9ArClQezGDb/M
eQ/ND4I9TNcI0Vo26OldNDH5JUP/EHFrQmtVkiKT2AJ5nKo8OuOu4tc9J1hVjgm5
`protect END_PROTECTED
