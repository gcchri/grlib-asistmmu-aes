`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vU4qzoaX6GqayN21amV2kaajEEGmuPut5SlQinRGLZu45HMi/DwZD9papRw7Qml+
sc0usATMAWoDZhQjCue8tCPMXzUWd3dkkyOQdBnQDM0YVb14im5NirpU/slLPkJB
SSx7jinOGOu30V7ckUYHWL3X5J3RTOMVGCJPZx0J4Iv4gG4yOB2rVz4ed4ZEA5Py
ssTlqqNe9twQbtpvKuZJlG8iKhiRAxoIwe0EJw+wj6LL1vgocsXPEqh5fvOWmskk
SkCb7GFqumlfjLqc3J12Ubp7UV4jNVmukKHZWt9tx1hKZ2ZHaq6JuHw+YZg6nFLW
emOG8VrXu79WRu+6KHPUrATopwH2gzIit3TpLYr1Hc9nUk4+KpUr20GpncEj1Ypv
Vaas/fW4fj7nTzwthWUV92RmVYunetXyG6R5uqdX5/mLmJ7h89zfJAxkMqe6wvLy
B6gI3B0SgYhnHXc8/QM5ICeIVMt2kkPUQ9YjEQ1162X7sDEFcpf35zKGzKggPem6
/EDbYQZgFwmtW9zknEohDm71XB24zB/yd3Ewo7bX6KwnqIXvNH2QkKo1ALytWI8s
ubOZuDIX1/DeVWBKhOyI8A8jbg4w1+nNwzy2A7tTCG5ZIQXpikMb9McZOTrxBKWE
ImmyvHUyAJdKRmpytfj/Ww==
`protect END_PROTECTED
