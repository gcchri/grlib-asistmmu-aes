`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dryewhfRYP2tPvi2gAKZTejLWT7THy1mT3vIrejvuSZfa301W2b7daaDPExPYnHV
a0a4MDpCsZO1iE2/gagpJbEseNlhVV4o1h2I0Do8oj8h1LNfEXDNm0tH+rfKWJKx
8GUM4z4hl9UJVFhFg0Hd7w+WDbfCTMI3eYCz1DJxdBghtLo2uIpFg7DDvu4FpZ+Y
xw6VlbvYB3lMlnABc3jcbtilNThdsHlFPJDBTjvJdDzJR4aGipOtz//W6uh1xxYm
ifZrTlwNBEgP8FxT2URT3/PfJBiTvWJlQYWVNVp/h/R3zIGXgXfUqFbBlpSMS1YF
7ejnmpyxwRtcInVu+nJD0TurrZgEAnTQqHR1Q7O+rR55gckQxkpuJdzrUzzICUGW
ywyUaxdn3fnTvM3VxrqfwMGnPveM0YugCwGd2CRRT/K57Y96nIb4ZjpcY+ZJ2+TW
vSOYld0lm0V5UTonMrJa7doqp+5jnWAKeIkX77/jKQXgJu6bBDWM6DJdcuIDXscM
yendT+EFZVxA+quQi4Z+3FQBGTuqsBIWpmDl5S8WJKOWj7odchJn+H3P5mFrDWYB
tuShbr5k1B6dkdffFO7rwJd3wPFsqtfbYuoODkIbUZfIG+up11RiOQ/7oRN3LZUh
sRQP+UKhqEevsnqVDNaCOxH0WyBEdfA28atDuKyux43fPfOqY8SwpixdZ/qL/6sm
cUumbJbQQarMb2h1F/fMtpmTVSMuKonPETGDuIWWTN2U5BlOt2/rZIEz5rbicI2J
cU4iAqCqu1ZSdR1g/myxhg==
`protect END_PROTECTED
