`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TyUeoOgwtaKDij5AhCB8d+Okfv9Q2aeZ1LrECdZaMF2TtnDLujaCAZK2BHegW6eo
NWVqEd9x3uuNIaRMpmy0ryK7zUKd4Im5AP33EtBlt/hPlWlz6Q3XJILxhTaAssON
Z8V0OxdPqtcpDeRAD2hAuQB2DM5xlU2e0Pb95GCb+3a/vrqNYLkdra2mwM8rbbJA
l9VrGgQ7qc4uuVcSk88YBgsfCZ7e5txxH2UgYBOgWAZ6T+FcCybylUWyPgMB7lxV
`protect END_PROTECTED
