`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FaAG5OwJDutjakx7H5pk7QQSpVLxsISnu1yW0MlgqHxzvZaqqaqmxxMtSdTzvhnN
0m3yJlErKp05u04oVGT30GAYH0MSfXXfsrKo9wcL5yYtKytOHwIkhw10PCDuoIiJ
bJUgWTsNEiYS+bqBAUoDTbUhG/iKxzfvsi8CgwwIKYyq456VeLPE7klnzuFcaiDw
jdXI+HYvMIFrYE43mZ+uKiEqvZGCiCbkeWtzm2jqcD3/xoJxEaOuQotFvGgEYdfS
LFqGHYyS4EKctsCzrF+Ehf/ABZyie683njpdvJOCQZplWBB+4ueDp+yKmJb3urg5
zC6uWw+0C7hPtFF2z4Tt+lHc2eQfzwO9d68rwdmY9VkeCFSzpwuFu64HnMcZ73fC
QYTHLkAAz5Ski5AH2uyjMk6+LmenJYCVxme6qJtJRdR7ocJhiDQo/Z9rhb10gX/J
9wwWdtPvXm29hrUvOLofySi4t29LAFjmPawl2MbDc7zYJBuX8MECcEWo3Hpg/r62
KjdkKeFjs80OgqcjwMpPeZbg9itfLNSUee+zjn7JuZjQoTuNIa29LqpD0BLdjrVg
TXAozE6wdTZqRxyc6gkQuP6dSJtuDIutCNezHUdAT/eDSUtVavzmll73Pqt10TKM
w+xy4nRqaBzQk5QqQDwW4Gi1nZD5dj9eZM+ms4EPJZ0qqMs3yJykFfgvl3jsjKmF
puF3JeKSzph0g0E+TjbrbA==
`protect END_PROTECTED
