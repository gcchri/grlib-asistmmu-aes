`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hwQ0MH9SqE6yT7DRzfK+c4lb0GL8cqVif5BzFtD59mncxDD9U85hFCNZlI/d2vdR
xHxkARV2MjkFgJ381VomlcgOInzXWg7A2AoKvcsJjyHfyZrO7ktJIu5OR3wFKaAr
qVMSvFiA8tmOjghp8PXC0SqqqHd9J9sk5T/PVT+Dj+dgquYcSXgiOh6QIouIps6g
s3DEpAULFdnwjfLp9oM+TG8Kr2xQZVQ3L5OJbeJrkdlE2S6ydMCdj/ioH1vQ4QJK
jMPpCS78IZN2GKKxHZHTEvdiArwRQSmDzjFK1uvczxqeP1pLT+qPEqQigA0Dyzpj
xoZylNthfcwS5MHvTHRRcEeU5ETB1PcVhH8bVLARQ79cX9o9LFThvQFsZFaj8YxY
mbpFUPugYcl5LF5yT1LPJFAMuhYItEdQD1zdWqSV//pqv7l8rRxjJTcAzB+zFlu5
KVi1fVkHHeJJTSXDeFlqou/VDegkIJrqQFZZWHhE54sjKCLpgJOdrehXhwqAPfLI
`protect END_PROTECTED
