`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SL046gfzssQeV/uE2kcpK5DXMWH/VXb4wEdS6mHaMEM7EEtwiEHjOrPUluMqPpT3
5fYxPdgA/kzY+Mjwpeev/fDXzCGnqqBMRM4xAhPhhSlcgzvPEkBX/jYO9qG8BLgD
aSbzQ+j5RARSVTFzAAW1t9GgCSLZZRd0qXdPMUD/c1/uanJEyCbChMvWP4uh7QfI
l+BaY5ZvSwWDr4P5qFbbhwKpDZ4jKbJyyfx3sgEAk8x4UccmXrCYnviWOFVuVlH7
ZVDuBthFPn2zUE54R1Rq7P5jbNU9AK/wrVLoSCL2GeI=
`protect END_PROTECTED
