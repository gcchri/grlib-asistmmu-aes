`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qV7G8rd6X02TYrvyJG/0pk83jSi3KoWsZ+y4e82oEx9Q3SSeO0XFPaV9wt9/61xM
3I59GE3p2QNO5D47j90MHNkbZiCPRxprmTOABCw/WcJosSStWCimxpjD/W+7sWeB
4Tv8aTxfyNnAtkWYgEvyn+aMNJ34F+L5pCaECCY1vAvPbCl/1n4/XoFIM0fL8txG
efrKS50p1/dEnh9HxRJlsJrW2/grWukYQ3oWQncP3wVFF27/GgCxoq5lyFYypFqo
6qgclYsCQegBkYjSQ0Uk99QZv0fuEOY7yS7AOUHEWe0WbR3wDwntPBnIgSckhJ9f
K+6elqvrmiTOuhmC8SX4VUFaDya5Xn896efyh7J/BEC//5j2xaB4iU8m8rBQYl+J
qOQVYESLNpHYBg1bGAL8h64paGLfk8u7r/Wlx77LqEkgbRqfgwUT6qZMdCkxSs60
vDr05xlmIkcKUNQhCEjt3AdzR/uL5K3IN+kRBklGZjXPFwCi4h9wG/jYV6oMnM+j
+M/X/f/D3slTeLpnVnUNo/gKcLOHJUaQ/cS93C+gmCX3rRpikzFSqddcDyycPv8I
Tnc7nRABtBRAwClaownAew==
`protect END_PROTECTED
