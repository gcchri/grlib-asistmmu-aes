`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aDt3fVrBrY2zsMxUOGHQt7gd3J/jsp0pYJwgsoy2CuIjQ6OZrcSJx+V6lP4WgPDg
4VxkQZ/KidZccQYZXWgKoru9F7dl8l2W5mNSe8xG5sp0n2OAw6wzaVm8gLz5MQER
i2mGbOEgxbAetLOJPscZ2he5vpR7nJ5k9ZQNVOA7BNWdKqWbMj08guVCJcVHytaB
a7M/8ECdqEoSsvnJhBfNsCLCGv9+ea+QCH/9y9sazw8N83icDAjex0WCf29F+SPX
gPwnbNC65ZPAPYOwS5ntAn0R9iyT6GE2OuVzN32/TSS1mX6tLb+TkxqxEVOLykkV
UOZD/xFONX521Cdol5SpCNKUjKEkbD/l26NKWMck7xl8YWoCJ6AlW3Pg8K54GR0v
31E0cakpeiQliJmpBUn1eop9nUTv2EshtQMJH7uaScUsmSxpkxvwvQU2xFo7CpPB
BHCEM+CEA6UnZYPWkMCKRI05mwCFEHh7qk6sngAa/MviNi2ICf7n1OopoIiNMJXE
nv5zKoqC2e+KKzkNYw20b1aE/a8MRBMaG6CI7m+ZotGMBpXm5bVBI0hAXYHmvn+Z
/YBrouwU3enW0ujNPuxuCXaWd9ahQkwNxDdTkojAyTvxgI3d8D2s8NbL8DIVPiqH
IP31BSu0Kik6rOFc3yqSM4qoF8cKIOEKvxjX3nD9F0FdHcBQpWqI5OJYBmel8RmO
C6QuvahKFFqT9Pj0cjBv6aPmqz+X9Btc1DlQhILNLrkBySLrFO1g/5/83p3sMDNk
wtlq84gr1ZeasMGOThoa/V71jzPYnmeWb/43jet6eMyX2cKg7xp9W96RBNQ8PQaG
K9qUtlB4/s1ocYQuL9ua3yQlREAGJoPdu2HLmFJ8Il5lkD41T4APQVWl4/iEQ0iN
NLibtoxVsuFxfDEYFPNXa2kBWwnNdQ+eq005/TvFMjgq5VGLiR4UTiXiyupCkxp5
AnQ1KQSfzqzgRVhSy/46EFfbHNG43SaMxihF4JJurNRocjvWl1IxA8sJ2krbLDVS
/zX/nE3ykRDBPewBN0aacmZ8Aq3fJfTAkFKw+eJBhCesTsmZ5UvLfhGUblB40w3S
mTToxP0VYdS0NpK428GOb4eWrtK3/mzwgCYGATM6TWECO6BN0CYL3OduFuJz8Va5
hku/9NRleTrCujurIGq16XpqUVc+5BSQP4e33VL0eii/wRJVxKfJnZYhAlgy1F9L
6rD/lQR5JBBKy8x+q4IZqezaXpSZw+0DZoM+dN1uvVewAQDHcccEdK0y43s3dRPQ
hh04hUOCQeoPlSQ8hJeNaoUbVCl+Ud/q02JyrN1sDYjvNSaTmWJEsU2GveWLoR2g
lwnpDkAgNVT4Iojw4u8uKi5T6WGqHPbUl5VPbgRisZHj1SeRh2iD+AZ8KXQmPbDI
TT6qBI6TFyJaX4G9h1jUaBrb318S1iEsX1OXLZRisi66gdYPf3eMxbyJEIxGyt46
sizlPFWIaNrEVcdFukgfiuHGXtS9SyMSolhDGiEHmwPrErDU/hzfFFEnFbm4K/sR
S/kAPIx0v8aRGnBaiE7PDKpMFVZ02viKE7aSL5EcWBOfjXJWFqVA4XkZEUHTCErD
Q26le1v99zEClweIQBiWrDBcEcD34Jq3J5zQzOmsh7jPiC9NZG2C7n4UWmESAWHy
UCimOf384mn/ORArTOR3VvndPFYesLkbisNyt/rnqi3ly0siKfKEZPOvfKLZn2M2
uHuKXfy1mDWEpy5kBDHBanLB/P5gtZn3JO5OnF4t38wQnFZ74X7hqod3s483SeZ1
ES3aCK8NSfFzbEQdeUSV+z+IQcrXpF8mpsPdMOGRL9PWWBXqnlH//GcJKI2CLps+
fibVmgryhncxvK8LZrsjEsDaJHTjos9hpbXOTu3CZ3UtT9II6uVm4fhB/H77FrBZ
y3hhaxCFMdvZm5WC4xR/GvjbGgjoeKqYs/4aCebD/KjNwXY/fvHanWWyD+6F8krh
L6p5+t1DjblBcUPs3F0PV0r0TesHgn/Gzfl50ADa23FOrwrSnHPzRMZWE3fSdokp
A7ey+0jGWMLKzp4GvPcWebQYmMrPnMClsO/MdXlB1qBLdKRZEiuPjKzUgNSwue5s
+kDh7rTCUWxFnTbyUQzH5p49K/5fe8A/ZD43x1DNyFerZN6RmXXoZERppSFxH1LU
zVR5TBPvI9YBDjK76uYHGsCJWdTfVvyXyMOyy2FhTUeAY8I86s/jlAGbdu/FP7Ul
MusSiRmPzHIphtxVA2pM+TwAjwdK0hOwzQnC/2Mm2IbXQAEc80ZjfUBZvJSfbQCF
2dIZKhAWy/dy8KWu2VLWISeKNNUEli+tkvNjMIwu0LM9mpmVJx0Os6hIsQ9RjRn6
ClDiPWTUU0C7GUCcOWHgY+9vitz2XDFTOyiynnx1O0d/fDS7duQEIdwXHj2Ii7FK
X8Td7PVh0T10Sc2rVjrQn1rq2JnTEhnGYsPgQEHcwakljPVUpX+23RXQQP+QHrJN
9E6aodhIdMwUTr1ZP038ckXFgbJIW7ZSuLO0tLLWM2fgekVcrXMgvXRG7xltewFi
8UVI9BtTpggG09LbpjMsjS7XpAWT9X/7zxeAvky8hulOGFnRtuy3a4ATgjoSMmZa
mzYA/yqDbZ1zwbtDvZaZo//dDSAd0CX5uVRssT8rZCxRmISJbJA1iTyK7s+F2n2H
wEzbmpPPkcIvgQmkA58CfhrO240ONufpvh+JXwV8QijnqTBes9RL1NlQ2biCLmnZ
cjYEg8H4V5Tr6Ak5uagZWaYDfQDsHC3x+Z5twIuFoHTTxyS/fV07xBfGGRBt3hV8
q95nOs0gVPTB0DDcfbzoY2ZxQ2qkm51aHeLo5NyRkO6hQVXFrtkmuEQ801fVssOZ
fJ6e1hVXuwubgPQo4jl5oB+7FfhXp+y67j9nYCPWV6Ae6r4167Oq+0ObuJ+DNYkP
+wsg0qqIr+RDpO/tmjcQ2dC1PBG6Xj4Ipdk5lAxiZNc+bYNmhTWmfkuOnPanjUn3
1mVBZCsGwZkDppQ3+kNc1Nry1mksjCsihn1+p0af/KoQJcQYMrXAbSoGF/OU2K8/
kAFdCWwO/ageiOhaLiLRewLptYfB2ogd4Zio/ABj2IpF/AT7nhQG6qCRO/fKHhie
aRyRHrbhexNF8T5nXy7DpqlwurrMXTH/QI235L2RrZVCjfDuUI/LrOSGmNCo7/fT
IuYk2NCTVzTGYUuIFsKEYVdptcsDvdxU9mNDqBqC9md+SqF3P0SFfEfZu61zbgxH
e4ezPVUqNm7YhgnPH9bBpUL1D91hAVG2XzhumK0xdPyro3Qze9qM+ktIZeYZ3nl1
qhzor6z3Ke3ZWNqjq68eJNjFiAuVYrIqO4PnfEWrVYwlN3Y5Q6I3azSb0AedQEWc
+9Uli+t87UmCSOzq1c03FRcsjk6vCIvHTXG2miT4ty3v7NKZaP8UkQf9r00TZEFX
K3ov4DexcMGdK77X2Kkm5FD2Xa/KJJTjBsK9Rz5dRG/rIgtK1g7S62t6W71DHdSe
GI4bT7CFsk6bk4x1cerkbiiCobxLm0arO1B9QU/TUIxuYQv9JHA9gtOP1T+yUb+0
w/GsOe+nkm8lL0LaMwqrfMye6jydx7cJTN03nLnAXbsQEykq2J6/AtfjiaN899KF
iI7KkdzHCmcRREMIZPJaVxUN3zslEEbwNj2fUsmkkDtU6ksi67dWAW2kcAcjLMyt
EA0nzjN7b+RUROWREnax3BJV4nEeOu+4gESogarp0ogWdwGJbKUgCqADN4CjMrbY
yc/OmWJKhvDsVO/1OVRrYquyYLEExY4rOG/DKLRLPaeLtFiEDBa6djWnGbJXHWdh
vNQtPy5MVRjZldDI+u4tjhLEIV3i+DkzIjCNIV3vYXgReEFb5SuRLis9kFyRNdtN
lqTnK/7Q3lQI5Wffy4rct5KTkOHXSz7NJP66WQRSDA5mO/ER7S2O8UuxpnwjRGhQ
oeArvkGC4fuBBS+GPw9kF13tNTenHrdcL8dC0ZUh94TcR/3dqTkM+2igNrNM7NzT
GYqx/ghgw8GxiiG+7AvcpBmXDs+nVGxpRgzR/QfacjIDb+zviMp6AlhAjDWaZ3qY
v04dgZmoPgiosfT02+aYWbpp6PZ8u1B9D/jZwAsFZz5kQ8lFuNuJpO1kEv+AUN9S
YCXWzJpeUhahChdkM4MILzv8l/L89XWI6MaznqFkN9FcmgaDzpGsi3GFAFywjj/n
zTXbjv8M4nb7F+6aZf0luAHK54CmXPSMvcsGA4V1ATHI2E4WRRvSHksjKSvw8FRH
X8gNmIG57x7+zu+j6n5DAFShnP3OzojGET8ovFo5nyRJXKUh5KpQt0AVahK+OmtB
TQWQ7QSmrbUiw92tdr80WzmeQELbJOv0uBGiecjpCKgfal+d+vwfPJ+2OKhgWWe+
qRbsKQtpmkU1D6iNkEzWxV63HgW5Xct5VEN9SX7h/PS+xh//M9DoA/c48ymV9WOZ
+FR0kKFIDaAYtQrXbEGVl3W28smxT5P18c910c2vywRCOn0A4cwxmTZuZcEHxVNe
FLsTqgg1pFtmgjF1SAmooIlPwP+zQsHYl8BkRH5zWoZyAVp+T+0wEbBGlbN+PHH5
7uxsaIRYqkgztyhXkOHyeRM5tPwkQHw69zvG0wWJxlQZc2b7esBKb7Qy492msSbA
K8h2LETXNcpn4rA3wgl3ksho3qyO5nuf4HfLqqt/sm2GxpcGq5DFX9DJ5JtIoMYf
+aPp3HFEA/zy/SK3tiMffwckSov+jRQH4Z4CHeRbtjFz+pwG2gaPNR74YHJgdFKt
qLI0hy4E3M+kgIzWwVI5lieZiA98Kazay8yJrXG+vWZa7IsDgdwVpFeLkeDfJVip
FbilFJEBMEx3pd3hSTKgc+YaSIiVfDY5MSPrd73uwmNtieM5w5sCSMzTF96f8qMC
2i3VcPb5VhvfZaL75ESVopiPHBa7Xm20eN9RbBuKHrVRnfxEwrvlqZlaJNdWh2xc
ywagLoQquZqbxo0InzfA4Emi3FjQ18F1TSG65AkPUG06OxHdqgyyotkNc2SA/0tI
h7pdBCu/BUQyelvxi+zVLbB4If1LxGys/BFA3OmCUcwRWb8l6e7l9s2+o9Ykofv4
HIrA+KHqk9Geo5pTvgBZweL0akYOtPSuV7qpi677iGIw4l3rdx6dGevoc7mF+CQo
xDmUdRy03Efy4dJapSoW9EJd/B7TNTqERf82frDmidds1peifgD3GPqR/hoULAYQ
+Q0Z+HxJMN4NsiK0O+jG+bBHyz5YMQMGdok9MOzkFGzXy0IINh8RwTJPWdtGNDrU
MaPUSh3zJCgCRWY7NYT8ZAwfnSMNWLCun/xm22EdAenYZA3RgI2wuaZijmSKTrnt
dMcJ5ZTCnaW4fBsMvbBIVy/WejIko54K+BMeNR3jpzBxwikazMyjV/Sypt3nf6A4
X8UNt954GaJ3bJOv14okq1W1gj1SbxojAnqZ4nznICoJJshZl4/AAVPEC8qkoyKy
epH2tLy+5UMZuOla+iMgLzf0L9xv8ZnMP7b3Dgay7Uk7BY3q9e0r1pX1FWXHUVYo
XSDkchW1AyMOahuqCuKAmizdghfoocA4358BGxZvbjPyPkyZYQTI2syC3J4dOu6s
Dv+IYsj98FPEwCklg/F099YcAqiZMLkCy9PUr66rbpOoDvDEJaDlPB1JDSLluKqv
VU/WNY47LBTUDAeufSG5H2w1wwoVOyVC3RXpmHgzBJsPIJcwNcdTbab2Cb2eFbxy
onODuhFXL6L+b4eLeBHOGBzoslSwA9LzISIuFlBNrX78Oke3Ef8KOSvUocZMdBDO
klj9kPFxV0rZPIcXMIFplt+rCHA6cHZP45AOGqy6QcErqgSaiZn6xmaDAoveUCGW
/OJEQu3afEZnK/iWOVAC5udSUnj+OOyt5J1YrG4mUplgWOud9jZ+OC5/mWiPC/up
7PP/Nd7Gd4/iQwy6hNNg6RrnDfOmo5pJSO2oYxDI+07p9QuvpZ9qtDk0yk5eWmlO
0bsnUhyQheYWImEq2RsDeDKowhfEqToOwtvsJM2b9BJH3child8mu49aojZ/W/OH
ves/ei6GIq/aMbSAZrIfAX7HRq2Rbp1t4ocLoZfAi06f0TeQNE2W33cfNQbPynSx
wGElyAtDF2eMY6cvpYAesLm3XXpjbmIP3QBlxRhFCzXRUApyVX470udx6rKsveg7
/0AHc2/5SvxFEsdgLdY5B7T8OE9XOwnzrWS/bDj+WzDpZNKB9yXiqjrthS6ASc7H
XLdRLeIxBTmlq2F20BoRriaBiQcGU+sanp1NdHdi7NkJzeGN9slRxXQaBvoz3nTi
GQepKIW6X7qWSOPdHLrtbDBDiHwR25pt/PwE/cl/6e+DLGiz2Og1wU/rdz9bkdaK
/AdZ+0NvYcCRFy8lVHwq44T29U5vlAOXlyY0NlMtzE5dEBoX7c36tUPkr7NcZQdS
l3E6B0UIg4b5DFk3lmIhWTRhimcfdPxwlOzl+/MYjVU2aBZt3C7f8zRLK0OfwtRX
LlFP6AYrzts+iT663z7P9t96sal0YuiiXIjTZK68UW9X2ZD/ItlBSZjftqq0AGhS
e7rAb1SJKnPuMvc5MWlxZ225tj089dY0M6hFINnmKLwwnEkp8+vTijUGgBp9tUAJ
t6NSPrQRYceO0erGgZ26dLp70ywM6omSi//lKMieNGBWxt/eBv0xUP3zWbeMuRvD
S3tzNNUAbWihwEJNzpEe1Ns7353shqcHaxk4q9KrWZ5ODfhfBSlJrmykNZTSlvrY
54J86yJb1tzN/w8RVcW/mfxDtSRp/ZKEsn7ahukTVxTUtv/kjEIkElCyyIGTHpR0
RMhMOWaWcZwazSjbsoKQuTwsZ3tnBWmadbIOmTLmJlDz0z243hmyzpiUHg3pFLY3
TcPQ8XVm5pDbSDcD3U+9mR6wOwp+HBiKgsKWdz1VxczC2KqcxgRhUw0fdxJdszpo
c2Gjo9OIjAEZPCZMktFuO7f9R94nrktIUpXCiXRl/gRZIq2zi5gAPBspa4zNrIlp
oIkLNpKegYEibGI91PjOiMzNIp2X8pPE9/1+MtL+n7WexjeUot3/smnVwYgbKlV6
q6cwVswn+5Mgv6B9inQZInFUOBn7vMBu2s+7etHUvvLhkmXO1qC7YHZjc0gzMGMY
WUcN8JEGEy4iSiureinKZ6nQk2EyZLOsmvBXU+/7xZItF/Kb8CN8xY9BxgR/94rG
32ZE0/toWBqOcqBOA21t6NeMiqVJ75TggFSJ+wm4BUtfDiJQJGPDw+hpl70gSyGc
d/lcxw8/HSkKnGRGBXagY/4cX84JHoNWlXz0nSfv2BaKk+yXBaSvD+Li/OoQFFPr
3p2Et+npu2SjVfmz6U4H314vJ58rYkNQM5W1Xh48zDCDP7wuSp01WSJCxPOMlFPr
+NAN2kF6maaHrCvrGmOdPrEb4KguctSQOy1onRHw+S+/VCm6FNVMGSMgCb/yNaRa
sHJE+Xj5JmLaYzlSpqhfyt+2QYYaUonIuBHQYv8DMzxpT/vxxzKrz+psH84cQFM0
rnkFVv/qOObjlyjTwtiNCZni5/zLbjQLRaRFGjhA69nOpMJOrG/g8waaXEPllH+i
xXhKf0hzCqfP9qdH3lsUXM6knfHyulR48dUO9hVzSiAJGVbMy7MrZGc9tvbMO3QZ
1gsY1VYg1lqgJgoiOYpcScDipNs2f+96s0wEHa8Enx1dbEsdCXQamAuGFL7DJ8gl
LmGZr83nY3/VnF80alZUai0T7Rg7UFVR0BHLlDs/GMbIs6Br91D1zXyH64+CNfk5
qma+EGxs8PxnKowY+VavuovIY9rXBiiBZMF53r4wRkcc+gx8gv3u7B0YjNoMO0rk
x8izFCiRsKyNQdNR17d/pNo17Jqxu5PCYbreB+Ir0Kqkyc/yPRxSquOCffzXb3ru
fuqiLlPXssE9R06MkZl/pQB6ajPxvdJXtSaEZnG8GI9j7uTqSfCUk6TSOYjQiK+U
LAkCqNKr/GOX81kWk28yFkO1kF45I+Fdte4j0/Mz68cQjgyx/ccdCyS0p0fS1xIN
aAcYItlJYZa4Ru9BftRWNGgJOUyOQeO5nTgTf2s6m7iAcFUVosiaIRG40+d6RGsj
5P9VFjUBTXsJZIm2280i3Ezy738rnTBcqPBhMDkAcEg+G0Hd50BBkU2ZS2jCSfs9
T8vBdM1WkSYfj9IXDSmJXMLLN7KMtDvwOAW06uwoeK7xTeWNJSNWHuQuPoTgVVme
6dWs7bPc5A1CaTc0LIRLupbslaMExwtXNXks0lARTLsitzrMzV2jllkCzTjQeKb5
fkKRqpv7HNtposGjmGOwSXJYQnNnYVw41IK84rcYFl9/YACV56AlWlFiArpw0e7k
ijBI3suqjpSpxImphahNYsqY4GIh6Gm0+BmADQsyeU+HmvUemPCnZZxkGxYmM+os
Bq5JmX6l+lwPdirxFWM28h3O1sXuW+79cxzbhDVjMi1KBM6UqgLCQIAz6M8byV58
I5L/77GQ3P/Zt5F/LVeWIH3oLmD+XC0Qlj+VfEjw0/QDoQDiFy6HR8XOU8SkLWng
waXDpN1Eq8HHnhuxk2QECsHJ9DvDqh5HVgPylF+je3n3qRDnl0fZv7Lc4NadP269
edUgVDPIhOnfz4nX2qmEt98n3RXFj3o7U9vSXv4er09ZlfHBBN/HNfX47BuaZVXQ
ZBCShBRGgsiPRIs6o1HNglGForLOJLkimfpSsVjjtZLhwkZljqyDXUOhF0s+S+lK
eO4RLF1pzAgQzWFZbQz2MkXJNX83x01DggAdkCAV5KaD7PZWqbggRK96Uj9ei+Za
ZbFHy4h/3Ox1vT37GliwnJk294qIKSn116b56s700e6qAyU2MzYH/KU0mIXIy7ZL
5FGix7sJEbxb/NvU2PBnY8f8BRbWNmPwVefEbtTIAWariwSnXjeJlAmmvfYDyTB7
GRjFW64hBKxzloCBU4Z9zQ1ZDwT/VhqcGY2BDEVu84NN/hP9fLOabNyj3ZDJ4hV3
UWOPI7kjufYgblK7iCkLvlc0L6OQ6VuetqDJJSxJ9Bpj08yu2o4M8eiDGJopdyen
Q+LsgyRLsk2BHTdBwgqpgcgHmOfGxbsvGmFDCPiAB4FFasRrGXMdQsbycuIaiIzS
lU40/mVi3sP23jloPKT91XZmqPMuBdN4VIanSIpqmzcHaSvNPd4bspoBnO4Qu9d+
T52j0RfxXrvwNNHitAYb3i2NncRDml4jccZH/pl6G2zjDkY7K5Dsd6nwf4ToDnG3
6ej/pdUiSYuW7PD7AhnD//2eyLGyMRHGyWwcB/hbKpbDN1luSVBjdoblpwylBlvK
OK3bqxRKXqkajpYVkvP9XDaUVPshtpMXGkhda5UUCIQ3QRtaMwWzleMh8rkGLAv8
ErFfnQhP/5EI0tujzeBIUJOEtys6s1eGM/o+13Aq2ii6pWnyw0dj2qg6B4PWuveK
CqsndrHHomPQkLzgcCXEcbYaGiuCmudIZIrFL/plsETmJNz6m7/iqTXyHB9dUFST
cTsvd0MUgceCGibc1lahKFFfJIDTqwBKE/jYMIvXd9u75uITIH/xUD1Zc+puXvpW
2ByeimGz4+NedK0GiqpN+zq1HIQSitlLXUj9+pzA+erLezlJ8KKLs9Y07QuwlqYh
2mGLVJnk0IjlDKPbRNEiGfD8/uEQqlwx9L+NGOqx9NqmkVWaFKke8h9MJQnfjkxR
uNP4EqH9IBkRtvijzBKZa1JOxWKQqFEyi5Um334/sCjs+hGPEQ/BU+p3vQg4rxDE
ErjrG4S6CdS+RzrhZBcakcV4AW52uv+NSCFp5bGt/mM1Lc9isqzMBKocjhVew/NI
YlUsv5QB3zaw3lHozYEqtzTPxZKKqx5P4VWGHePxa4DD60u7pnmRFhEFqQ99pWsp
IiCZeQPTuRdmhVp6fRdFEJYyTCY/8Qfz4qHLD8DNHQDyuUHpljUI7MqPPEFSldV7
kAqJ6RG30SE2Wcs9ILnWMrOXYL6MmZSBcEzuoWJ90sZgqszwfaUaFIKB/VAcjzkR
MzyBK7dr62Z3WGjQb6lzQLuNlTUa6getrMxsRUbA18ht/Ay1f2G13c0SIP6Lnmjc
JeXjFih3l8ouZFn38/BFCw==
`protect END_PROTECTED
