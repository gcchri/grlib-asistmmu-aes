`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vxulUndN/F1zZcIY3F9AlRLEyeUYO8e6rb74yDaTICLqGDvvV/wQASK8u1h0MqAf
V5OHMrU+sR3fp8RQMb1sGF+/sEkFZ0B/BoIymfsEjgIapjGarkJntriYwSR3EYwD
PlHpx8FgcIbjugrO8mv4APFjfHCdx2jYKoLvw55BFhWhuTs6jKeXDsSMgnGh+DTa
gI/lHtN5jn39I8hbzb6olwRMcyDsVGudljwF6SE+c4Xhrze8jCfxmzMs9o6FrEnR
RqQsVJBM2cko1gE/RJ6sv5uKZuILAv8QG5KuBN6Y+Y6hBbIvloHncYBg+fkONEEb
6jITa51ZM8dzSInwFxbdpg==
`protect END_PROTECTED
