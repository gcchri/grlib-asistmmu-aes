`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HCb4PV1hQQQ833fwAzb+1DP4OzHaYLeFuleKr9J/1+G3W1pLA8mdzlI8Y9WBzt3e
PSNHJC4Mjd/krP1yQ1NMQM3R3vxpVsWLN3YjJymbuL+w/Ad6bSbN3GK2CXL+KWWY
WRyARcLeFAfp8+nTdNrd3rXwrih/6pqz+PZzE22Ep3LyTcoQ2Xgo398Z3S7K4tbA
AgIy8BTUAhK5zL/Tks48NrkVE01oKgvWn8MSQ9Qpluf8kLrJx2V7IZW1Op2cEZOJ
Q+458BWPxKyNRwQZKdsx96SiTx+VQLHNwMl3zBytGqX1Rhs8Kx56V4tdoqdWFRq0
uxwWIMsxzLjZqOjIfsAPDNIXT/7m4DAIdVG14TLxkJKLIaGEI5ApvIZ1ZIAAT7hh
kI7clAA/OsqJB0y7KS/Bf0uZN1S4NNXUw3d7pMF0+2AzQsxRfaVQVW8JWyZ8MLjd
IVm26lhsb3Ou8J+JYCRtgJDUC2HcvXApBHWzEdPFzbQ=
`protect END_PROTECTED
