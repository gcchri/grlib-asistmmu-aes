`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nJ/XgmcHwvlh2+FSOPRQV5pJMVg3X5oVH87FJfA/ZxlM1r9JVn8Xtrrj0A8vk9zX
14r3miHH43jaPvHWlrn/4xCzYhA2WX2RrbVSy5swC82mfexjQAwkttrDsvRPDtUZ
wbYWTGlm0Rd3tIRMmGwfTtjwOeMpUkpR6aBokkG0ovQ8nfF/hM74N/OJZYXwGTrc
pJbslJ0XoRN36yxbQid6cYLS85Ybqrp7rI5j30qsnMgdK4+ILOv8H5i1BOoErbZA
n9K3whYJYamGopgoSDt0nP6fm+Kr4cjgdTHf+sw/eY0GR7AN5hi0FmWqkypuqBXs
7ZI7Hv2WUzvCE/5OHZLOMYWHq8reD8TYbmIk816RKlstmLNMcVc0NGyc06aoEFhe
jria4V0NLX6wzbnhd+CLYFIzl2FoqSjATAxVxR2hSnhW/gC/PW+XonZIqBJFO6Rk
0pSkypSIbGmYN+ZjwBl0z92hN359LHPvr4gtNkKbWtNfhUk1mZ3vePY5pC2f+qAh
ga70TyRlZ/PjGpBOpb/+aXh+p5lVEYtVllE8c9H96MzxQLDeg9ph5RxqFwlgJPMK
9FzSRhO+WC6l5DN2XYcNolFHksKjyYKjbZ24UaTq7r+Py9Bchbeo/q4fYX14AmPO
5mB2CQF3AOt6QqHtEY11yxQuagN9BpAR/68zSHRkvUSQbPHAo0j8xwneikZUPNCX
q1YfINo+UazrQSk28+RYF7Hxy4R3DIjX+E5Gh2oDjWUaS0LHJc1t8E2iXWnrg/3+
xIu+c4+XqkCHcr68yNWIbWTLjXorWfWg1QMUL8gYNW2U8TjztCoKHRsC/6FhvXGv
2bmirHSIEdCf9lKMCNRW00av3TDknWgYxNg4mDU7JC0755yhdPKY3+fNCekK5W2a
nJLlICtpoAO0mgMruL48QslRRtGyii/tEb/FNhszYP2TvUB+fZzSCCyEP1kuCir7
VcWxLyLT1ivLd2YyziRoTyL/7/gnTeR9OALsJUqhG/xL7owhdkmxQssIAl/8ii1C
8NGaYu78YAieuKso5a9wkoV/Rt93C/WrZ5oydlwqZhdzYf9jsm3+fCzpXgyfFvCo
lG70SLDRL2TjQJfxrkNOKCG70jW2taRDwLm8U3ieGeB/9tDj+rxih4S599aOwhh/
5X47Gy1lpfyWxvDApqhINCOYFiL2gpWH4Pyo1DrwvjBvQUsRSX0oViPz0AknlcHj
Pev0T7sC8b/w+LkUngug48d3RgvWhSC9xdnoqeNbPUd1fuF+AwkyTNyosBX9T+Un
dzaP3eZiQIII5a6esVT5xNM5KpLt8JgPFJcqyZNR3ZSVLPN2Jscb0e3e8DaNLfa6
8zTROhMpCf852ig0oW789jJwI8H5VARvcTDNrDmnwGXi08IGaJH9dYm4Tt9n0aUQ
y3KsVRSkbasgLiYuw3qEWQ56AnShDF4/b+BoYHclL+c7g/+FFkNhZnSUYtsOFARJ
WjUuBbJSBGsXB9xOIu5rAmJYNJn2KEt4SD7Kk0CSnpsUO9+kPvzv8mlX3aZkEbE6
g4G6g9nS/XlSQsCb2GtyceG0avFyv6Z6NXOWkRfCwgU9arEejoFKLpn+TM8mOkQP
ImRR0w1F7q1SZB+TfCewvgZRGyEyCSAAR8YibCsSyo6tXsHTckMOp7uvROHZilZN
aDWp4VKgH0xmXYiGycaZeu42Ef6UlzhQ6pQAvu11m1O+Mr05a7X9S78aAee22CVu
ppAQ6xLHdSUNM237wzhfRpBwsMGqJhwSvqd+h1Iw+jdE9MRl6OqhZgcBa+eVmgfV
NkqrLAf4gcsuZFAIGcTnQ3X3Td/mCsXH6x5EaaT4JO1G9CiOrvRpSREQ8hSCIjb1
dHYOT9+VnOSk/I9sc3UmDieOI0LaEHr0SdLxmF5efNKKBh9ZTnmS18q64vqKXQoO
imom1XlqRcPVp4ELgvTwTelQwpy0PWbyVhDawWmtodr+pIYhJKdCpWa0StNNcYCI
5pp0ehICOq2AyhFhP7Z8uPcHC3QF4T2xXu+RA5fRJTp8tH4imz095Z0FNRtYWAXS
AnXtP5GYfjLXhMLUiwpZfwp+Xanr7kOKzWGCXSkpLEEq7Iw2vghzFLT6gUzXse+D
qeYFiF+PsZHN/OSP/x1/qa52hKdAjV0FgX7D1OaPuPk38xlcVq55JvdntyznDlzi
OtUn+FZPc7uAo8DPDtPhNvIsrzoaFRVV+R6Xk2NGBYjZ2Kgubi4Kuh6+mZuA4A2n
RYddMJIEM/y1O1C9eQDlOi9xMwiMnrZkpESApQ/+3+AYUaRfkMOWUJZuGJWtYpDY
FutccoSThuwB8g38pPzgsUj3Tk8ig3CUD4pTb4iQ3Cw=
`protect END_PROTECTED
