`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4FhcLvOzwtevsSCUMErD9MaRm09ANlwbNTDz4SU6LE9nqDAydhmiL6OJXGIvghPi
qdzGd5dz8dNwefoJ7Slcf6UUWHCKpoGLajjJFMHiHO+MHpqmBdVZUR1+0K0d7yrw
yMfY7HcIVJGdlks/4MPx0jGD/If07MDS+9qO4z73QFnU65HAWE61k1VgGUdv+e1j
aUWwhtfCisQXmPx3S11F8Eb2vANiKoziXg8jrWMOZ2rgbKYydUHU5lpc1pERaacl
UU7cSQsqpB6KEwTIy6itnFEH0mQp0opcGtliluDJkLHQ/v2rVGzJ0fm5APCOS8Ky
7sO2GmspPPhBoDiAOiDtyO2mqvmW3dN25uiUdBa2oJuLKFRUTWvVR0ZM1QW5uhWd
dKC72kUu2B03YY5DlYXYrokCx3JJRS6+k3Nw/dnroDXfnXOy0RcxbS7XBxn69oVt
Cu0WI8Gt1KqpnwVHWLvI3y1IXStacNfT2FEWWgCRoaVINuorPwA9wLyGn5g/kXvd
uCbY30M9BZV781zit4ooATRKFl5H/V9cQ1a8fNNhmtY+k1urpTkskY6TlXiFlRtZ
5K8iOEfignT3ZvYW6EKQsT/lGgEG8M0hpTjE4KYCgDahy10EsAcOz8Zw/hi0lDH1
UsF5gA8mLIlQXyGxETPqI2u0t62HiI2l1nGl0aaBTbM=
`protect END_PROTECTED
