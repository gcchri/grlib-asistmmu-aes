`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
36G2PkAMVdhJPTlp/A1INZNDOGmzczz9HT60npe5uwKsPHdhRecYFjEhI/HZhBdA
2bfCBggGU+skevQ01p8aBN6GKiUNC5f5Wi7xyYQORY8vkONlszkYTPF/f05cDHPM
nHKLqXO7nK0p6doH9Gq6kUn/yUHQSkhlA5Cr+HRzbEpMTCpu6FUc5KXU0/48U1Ic
iKP2ZJvZtexTiYP3jPaKffPQ66JUcF8xTmgDLD25jMYd0oaWu0tAtiKRzUntOqIp
TWq/MZjUPVPgaRprgH56WltqVnWLS6fF6Q55l6FvvKUPMyCQyvATX6KasUaL8CfS
8qjYh2ZkrIZnqKObgn2QWr0ea+x9RHEqNB6pWIZZHbii1ijI31oOkTXHjSy6cP5w
1NWytCA6awUmtyUPz4drNpVFLIZz/JILSBlc4a+WKM+6mzqAVWj2iwoGZHa0EAwm
9zAVJQ6ZwFPEcVnCsZzKCo57mzFS7SF91qJ3ZZ6hdsMukgqCOhGn8RRgcCQZWKO1
/Stk8NqlDe74g3YqJYn51NyLm2WSWDChnB4838+smgIBeZE99Ewn+WgMhFaNrILv
aVdKkYLLsZmhJzmvPZbOPfrG9lQ9uh1kVurc4ZQCPco=
`protect END_PROTECTED
