`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cBZvLnBLV/lxtB3I5dtz60gwwt2j7J7i6DVJ6DNNWyzjbMSSUI7A2WfoSfGRTBe0
/DYl6RSH/xLAbzIsoO4KG8CiIxHSxxf/O7lBOHRCggZVF0QFhQ2qNHT1CfkUj1aK
6S3MjYBMoWHpsjcJcP1AkrxQ3Xcxg5IuYdkBspW2/+JzOgVlT+GuJl7bANpGO7w6
D8HufWh0bpzBvmiGdg6nDcKD/qFinnQC8+WtlMgJHB8a2kRuytQ2dYCPVSDnPK7B
bRQ43PbWF/zBi7xUBtykUKNqd/kNE8JRkDF10JAgVK0iua1mSs/BEycfP5u+/VWv
dfp7ssRkhQUpHEu2NODibpYCg81xsEGr0f2pPw7LhDZIYKb7l4OMICGZcojdDA9g
nmTquB+joAgO8jDGN017AR9t2oH0sVDjc88E2Q7cdBiwLvgw9735XJCP0HJHIGTj
PhY+a3b1BE1uzSgULhXQcEKxBAtgsIixXzLf7qWPwvWyqvb7xBED0HAsm6yd8smQ
mvgHTTT+eylfxLLMEMz+oSh3oHzYMVGk+n+cIYPw9/UTjU6bI82ljqGaCtXuGjab
j8eekXTmN5prjjyBTZRqM3vlFhLuKA5OYuH6pYG5yEy74B2lsMsPEVAcKGcW0pt+
C9GgCRprh9bcQuOa0yz9+xMHGvJAO4ASNPg8iSlIYsV2G5mrNFwQFsvQVOruU4Ie
TKdLlpNv5Qx5/8TSXMo614bHPSwLGmPrjCw33Lz8d3U/cj8eSElJ8Lk0qsL+WPFR
VgaMbYSFqt51Tl/T6TkERmf7S/9nt6W/TC93SeuDdeCySJ5NOH/Ms223Pk65ZZmX
BAnDm8GygG9xdmlv1Zwf07h4jMIDadnwlB69pudrrdWKyjLpH6h6HXWB7mPCkMNM
uG7NVJSRd5lQ0rOIXOgfhEFPjS3rl0BIaljyww2AesoYR3OKyVdceG1qpTTfnK/x
/wwhSFWGEXVTBCuJVe1jOktbqrUALOJ1nJtDCpKgqJ/+zucIYgbbXaD141OOtwlj
Im3UrC0kR8A3M+PuwmpHd/NSPmtRL44E8K8sccPyjojO8E6t4IEL5TaPTucvQD3x
alWbskFs7bWaVTGZQAOcWSzqPyH+j6TitrQ3MkOmkdwDINLVT2sC6wbLH/lwLD4z
LHzo0WHiA/8deDsYgX4l5LN6TEQoMOTJbT4ClGQIgPOfRf6V2IYOlTKsFesnmivg
H2wi6d30rS0S71F4KMy6VOxsZlt1d33LaWtP96kyUC2CfrgmOghcJpKpqaakuoU3
2VfZgUeXBD8qQlr4oUntNX0ouOAXClnwEsS49o608OJ5DTyJPu6CWqnRKk5YOsHV
+ah+aA+rJhQRdXwx0G6MLJAncc3AUpp3+V0GPjDzqC9l3fgshuipwKRC6dHtCI67
OLmnpBX2EIlBd2exBlDP3/8xOnbmtsYFM1xc/PHI9QdZQ9QS84RgYNl/jJtTU69X
44+UF5uL2b81ubuZ59hyaA9jz5srfkaVbMnpYJRMpHwCApTT4n50SjNXTsRBVNA4
4f2vIk7SLkicQjSmh/xTe/Kr3wmvPjAtrLNF4matJKuw4EdKi53ZyIU9SZi84NWI
aF181F+1hTcu9Ib4H8Dc5ptVO6f5v71KlV23zY7rfb+uVpN4fQ0IFm3hKgbB+cWP
M9lLmYmMa5gn71FZZ1the/nm9Nrl+2AH0sIibnzmZZ0UwTA7zKCl/h/7YFQwa7FH
FaW+qMD7hRpv/0gA902BNPHqM0VZcsAGK1PN5LrQlzUACko2lSBU51Vp7037D+HC
TXJC15p7W7me0eTJ/z8ON1eu2PekGuMB0dYIRsoaP/It/QC3tIR/jT/Cgfvi2Psb
LA/TDjM6QSz1KgxkUmSz8QMTjZsMe6gKx/GGoxSmoTDJ39sfa/FHc6R/Vak28F2R
6gMaRwly1yhwnVigQkxBYp9RYseL6BwcNTKpmKgn1HBIIblBAUv1CvkzyA5qL2R/
Pb1clLPn6DBrnT44yX/vvPy34n4fdZcvU3opbOXpx0k=
`protect END_PROTECTED
