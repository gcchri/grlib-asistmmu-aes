`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0DwEppVggUrnIxv5X6C/6wpHXw80bUBTGoMXJYKPp1on+O8686ZdK3LkoKLJWRdT
synMsCU5cwtzCWpA9RdMu5ZDj8kyi0sjdVxOn1sCQI4q1ARWZqAmTiOt3CeEWjr5
Ti34UbL6wmGECWtRiJKja9uCqUxsgo3hC7xtzzbYLkAnaU5w8DqgV1okk0XOPBRG
yRLc0Yvzel9zn8W0pF1jF7QlLO96k2etd2XGqNupDQOEmT5SoaLCEiGpPVCaPw5H
6MOL/xAz06ym2U+kbEv5m/DiJyQZkYafltE+ixG0R7ZefsjkjkWv8MMf/iAli82a
Y1mozskUq5RjDmIYYtdSWNHZUUPYN/mEuyAZU81hEY4dgTfwS0NZkHVL4EHKWNTT
fN5ynmGYqk9et2BtmNj81bg2drJEbBR0dSf5RXsI7NoU0oj6DRC8kQcgZApuXXAo
cohOQ4hRPM5+FaNQmVRWcS8AkyzebTbzIfIcNW1wM2Utg+J/1Ao2N4mM0hMXcGzT
D2mMnFaApJuj0tO/CVNha3Ec/gWOOr/0O6T6g/IcSNekgDYrAlLYs1A7wa+jycVf
R31REWdE6fnRvqg0LERgRAxKs61cvNB9qQjDyezWdhe/BIZtvJ4fCqi7SA/kuIIy
/YTmZxf6P6+iOfbbm2iczUjVQ4FY0rVfukIbu8QNPpDIVjo29lGkLf/FChTOd1d/
YIZDACRPalunwiazsKG7dzBE2w0pEhpJvnJipMM2jLBUZfnknVN+dD8iag43N0jv
iiGdneF0eRNgA7Klg4xkbl/MK+Q4T1Mjbrw3p8wkjBXEGNR+40ykEoNiXPht4RxM
r0JeaIUiLS1k1K3yIEwOOl6m7x1kBzPsF6X0JkfjcIRuTG+ldj6JDfuf5YNZH5YX
Wfk879W0gpqXf6yIj5nyXtkyezYhHz5vXLPla+nU6Nzo5VoSwGfxRM3/OEPGjeN5
XgzN/e/0g1g1EbFEfe+FVp8+5Bkt05V4/Q8XkLwwdw678B1QpHqNY0v3OZHHRsAr
xpd7KW3C1UD2TwsQX6atWPubHxojcJ8qqjTLQdeEkSnH9/vAUx9SzfWa6DNi83tv
ILqhDp8j9L3CT53wtBb+LJhBiVFWUXy5rHHB3Pj00l7Z4KJY2FdGRKaYNbnpUeCG
AXeFMbqBIvmCL06tb2K0KLjYQ0m5Yd9LGh0FFO1cTTDI6k8W9D2GJgectrrKSA+k
EZL4nEN2jGBiNj8d9Fs91Cas0HdClFurOn5gF5XmPMzsLUgAarO8l25UcdZmqCUy
eVGHEpua9CJ/yheggQhfqLDrZ9xDxMrVsXer4XvG7yyETtxrE06ZY3QVPoNyrEDv
43ZJpLD+y+fME6mpSVtIRvwUB8/5y7d85irXmzbAaiznc9r0AYV9ZEeUZsbl0WjP
JwyLlebqgnBG4xJUe3Wagubw2hfO3+nf7L98Bo9XpVXtF2yPeQZ43cEJPjJAoSxH
jUJqdJEX7WJXsOovcalfQPdiQ59zzpbhU01D2TWDlSs2qdmII5fgMunrSGPc0DLz
jDHPqUI5puvYZ9S/6o+e1rhQ3Ybl6hYZ4bybT4lTsfmWYgBN8jaORE/g92TsP6y4
AhhQogLa9wDx8XMbH27LKGOAkZIjD2SobKCEoaD5a6BP+f6lbtRr9QF+hqyKrQy9
tU5JmCfWfmsfPQJPnUnCoh4XhMNeuKm1vz9ZIxerpGy9gh0NztY/QfrwVzVdBn6+
I+2EMn7bqJkv2t4PyudVDfxdR1nltVP1Q6zCxa1tw6lXUIVGsYWx2e7B3E8RfAVD
QxdrVK5g6+brTQOEJFfj1Vwh62qMokWmzIaSZq9wkECQMirLw494uh9cw1g4X08T
PbRMDEvBlYoLM5bBoqHxoGPV1cxv05fWnDqyNPeT8gmgs45HIONhqzGti8+Kk9Q7
AEEpcDfdVizB+6WcjMs+Er9+pqXxNe4KC7X2WCNgZds9QgDRwOCgkzxdimLXWb4c
NrBNOYcXyMGw5mVePayGLaYVVthPsuvHSZCjlR2DiH+EwAUOoDWk0HfbDGXtXY8M
La0OUT2zxEJ5pFvrLrv7K2BmYnqkg6oa020rtBSNlxmjFC5GoSLMpfC4/3J4mH6K
nbFo/wXNowERQ+wXGjtI7MmGowc4BAG3UIneyOa62zj/m/X1nVUnccB+pp8bbH2j
gSdvI1m4BEK598110F1cugSVmH2flvvZqFO3eYibD6C+5tjcZS9SsYG8vbiNPBAY
izYMJcsr1SpCciyPreicU0p+VrLD/ucQHm/v5vPc4Jmr31qnPDreD6XvR4x/me5T
1p+lKT2OKBJI17ujq7jHVHh5w7FtEiIoyEEyMyOCz/+sm7vhIJVGwyO9j+uoq+m4
5wlCC0q9vnIMTlU+ef1hh9QsfXINnQEu02c/jZWWqhYcerEredSb4YE7fK6WMFdN
HxMEPxDpK0FXBKih7/9v6w69kXTWAsMpccB8VW5uQF2Ovooq1dbA+PLAVdFMAkxN
HENZpVHJ7XbdKnsHrlUGgeHll45qEUhSO5OwhFnKqOSK445oWTZJWdaXx1Kyt7wV
BTE8OQ523HT+UfiBkGBb7x4R9VJxxaFasrzm3GKD1TFDB9BxrGlkO5ZipHLXz+tS
UiwCD8jEXkNbuV5fDWJy0Y17V8d0syhG+Pu9WICtaY3Ir6umfzLAMmN7/ggv/AtT
y01Fz5ApPStbjyxg6bSe0vKtGdANnvRO97iOBqtcXWiHgLWYZ9kS3ovaOum/DcSQ
1HpJtaJ5d5ZCNKCeK8kUe7fYE5Fhfp77ZRZnRhB40L023gDBgcQRPLXntOrNcwww
bQSMugVvNbanCbPtNRahbS9Tb8Cb7mFJBcwNcmzCGRLsh/xkik/ctg+IKQTbC6vt
UFyjyFQmZP6CB9twU2MCmNS7Mc1LaJbCuStPdBd5vC1oK9SQjPga1Un4UaXFaIRR
LXvUGFD6qTe5OmqRbvzGjhlJqNd+MWHXl8ub+0eIz9cIoNoOnQuoM6FQMLRovIzS
f4jVOv2W58VzrFvv9bJTLJYz06wD5AIZPTjS0dOicnN063tiPI72KYW3z/+KYkM3
Fp52EGreA8DtW/1CqPcgBhEWilpVMs9g96Vo/zHRN2Xl5JGZQnY1RvyQx33r+Efr
zGqo47YUkqAb/mOQTGiUtrZ3Qjz4BbAxDYpleGxK//nG/eX9H/LQqwdbSMpnKtrz
VszlJYbtuvVNob4TJqIW1q24s8iOUkWys4q1ESLfzg30uhxZwc+Ta4AQI8uG/NL7
K47/hu/hOymgZS7Llku0eLji+VFnRnAG/WJSsPF5U3n1F1eTuWMgb2idcgY5GiNZ
Z/D01f0EJ/lK/FOSfMdtzQ==
`protect END_PROTECTED
