`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pOry/FEIWk/Qrc2OWwTHuSG+mgJjzFowWkW10SHs32EC+A+8UTyWMJ/SGKz7JB8A
oqrayzCN9Zl7aOGRxZl8uWRRxDCgqZNyx/oZ/jSAAkwZPU4Hkn3IVuk7lmRoYXBw
t9c2oYdv2IjUDpP6FBxliCwlXGPWNV3BDdOSyAfWrqmHdJE6wjg16tRPcWp25wwt
cmozeag5ZqxjkXEZg2yYolURFWZ5RkXwGTuiq387Dg0X3jN8QtNhvGB8ONTM6Qhb
xdwJqlhAVZjj9AUzgL3obEfsL3aSHBHlLk5MxosbhdPjrFZRWaIVRIdhm+e4cIP4
P0ErieSmCsvJBfDI7nX0vvTH3GRxaa9jGwiEblxzxC/SaVDmO5FY0MX4w0Ht34eA
N6NteSAStoKhtBYCruFfYOAv3oOr5AMUp94SiduwitiL1GqPkA2WFrNQZ66RndL/
kjtV8soh5f6l1+elwwTf9UZKnjyWLaGwMXEOUuYywYTzWlPpJ5BLCsDsIZ4o3QZP
uL35CN/iJi1G/HvpmtChQ0j11gR7YlFyaTXf1ajl62Kdd9XxxTw235uFzgb3K6Us
oaX1iv6SboBQNWXcqi0fjh6CF3Hl3qoDbMv+TUwDByK5I4i0yZSHziqEiBmOHERM
vfcTxtI8po9y8ZOgAraqrQ==
`protect END_PROTECTED
