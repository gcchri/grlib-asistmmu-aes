`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OTn84RscCsu9InL5TUNBm/P73r0qZdP+KYqeVBZZdJv2q6E5gd6sAoK8NtP0GP5j
+3gOPMrtBXZpc6UOMZhW8GpqEjZWOGZ7AlaU3p3HQ/S+oIy1MFDyJ2Owzt5/TQRu
E0KAJW8xu04rWcjITHgDPxTcpPhofDz/2istdxBTGKEysy8p/q8ZAYUXFf2ND0Ym
7svhYnIGfy+WNvdkvQQJn6DnDBC2dHNFoGCdlF1HO3MX63z4YnDKgJciMYNMlYE7
pmSNODfCLsYz9h2YYvPRBDF6YaGoIQwqdr+bnlCP1RIP5OMTesqmMJeHQKII0in/
7m+c7D2pPQ8eRQcI+KEbIA==
`protect END_PROTECTED
