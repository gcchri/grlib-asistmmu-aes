`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nCcVoZPsiCI1BNa1YbnoWWUW3WM7NiEOyov+Hmix3iRPCOghqWUzGZg9Vc+rVxHc
QkJCOd2RPpeIWp+e5t4JBxqYHaafQERzXOckGxR0suDRvMq4pzWheC69THIopeZ/
CFp0c/v0f0kQ45lgDr1KarN9aUvAMFwVwOerWObxhVHrACzxcNOkwLQpATu4zFjC
iXAHg4GzdgRxEDQd68sNel0araMROPM9R5AT88P4EEVck/PoriXoXmm3MB4v7ONu
jPaNcYifRKcOTHnzwDMJ9qki9g0asUNW3TGofxCtUac4K0sidmreIJHvnGM20e6b
vp7JIFh9YdxFmci/fuWRIZ54wNoxe5v9zWLOxc0lU7znuvzam6Ozm0qM6B088N9m
4VrWd2RE5UpBrLNiMvsPx22I3irv9bk274GPW8u1MrZQCSmiiTDogK+adQygDcs2
7CRHOTKO8s4jkk3YXp4EnLd8djE6xJ2FUQ5Gl7VnOwRzEkKtWMLWvsWdAvwKN3Z1
r5TdpM1TcrCzbe/4/ItwbFgTRikXAQ4io7CUaFlz01LwL5Ouzq+noQVgrSvU+Tep
xXwv8SGpv096f+EwkNpp9g==
`protect END_PROTECTED
