`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fRfKV4PpQTEu5wwKnshUu3OCM+4ALNXV4OKFnCgVNv/bFz34bJXgVtptg8CSTLPo
4qW3CmjWonWzW3CFFnPjCJxP/IhdXryiQPOUsgh2l6SBHyG+xZXeiZ5cvlcCqOrw
e+jPljlrtSO/DcQ1plRqGq7Bzz5nLn60sqXixnTSGVODN+WR/SBlHN1Yc3vnQxYG
Rd8GqDwKbxHwly5bTXo5L2KAqR5j/NJtaU/5jKpxoj2UhOgssVzRvn68ZZYk40am
PBiXeCfY/A/k2IXgYOOo2JY4gqS/cMdvBYJEk8ial1pQBCeFAqC+wXHBYFbNMDB0
wvIcK7EJkw40dU3FvdcUkWd5uiqUvVs95CssNxr6uQBwRgH/nU0S57qYQnrLYjb9
uK7xoGXA60KH1IxVv7URvQ==
`protect END_PROTECTED
