`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kpqK+i03MvpZDv5Wr/+TGZvYo+2QpLlLRVUoVeJ434Tn0yGKi6eU6SsPvF0FB+5R
vRAGoSdc8pX9rCf5g8TTOBtfqKR3iiNLH007t/Oi7aKxVHbIJr6QMDT/uC5NMGQX
2dHMiL63fpLinno0UGi+A/P4RiwHTJcYa1rvhBoQk/Ek8LU4H0CF4TRUxACwiQ+x
48yB6SH41loqM7ANXyYn2ThhyJx7QvZDA1fTNX73WPEpuKu7vnDhLXMojNbVUM3u
FAKnimWvAR6cUzTrdH0Cv5Vy9pBYmfZutDtb0gqWa2ZCYBHrWGNyWn+voh/EJUAg
otVDRUT8DWcEUZh6+EQRvn18ZtTmBAcYUTwRhv1+1PPIWCAsSTTFbAW1c2Gklk1v
oEVHJMoYh9cpnpYCiS6mYgIXHfF1cZ9YTGfa/FfvaKIJhl39vnMWdXdFGx7GuUb6
MwKiKBK4BTujzZov2TDAE7p0JpVgigCPBrTn5o7E2HTsblGeZfMSMl/zt1bqVA8t
6cD0AmY6wppihpCpAYn2u27l+cCLHohIDvEo2tTS/z+8SuC7PkUDJtQPfEH224kM
HKDkv6yHypQ0J9mDjn0TscNBRF3kefR1ACMZy6/0me/m4k3+RrI1Ya0UiRcvkizJ
YVbkieiNnWI0jpVVDNbY0RDcFwQvZ1vemK6VmS9nfRxOXWEfT5dVRzlFtqo1aUo9
wbhrl399dG74rKgIppVuh/FDsP3Y3Qg6fPv51akX/X/Zb1VD3C+29i4yg+oJs7qS
ZwcoldPPHegfBXurrih0ODkqvwErQu7sc4H5WRVdM2JUPLNajl8n9DEf8TbEqm/K
hzuo8awTLDZMdRleNE7H7KKtKsGWUUufzCQJtFzchasounp18OASUgh2zUIFa5aE
X242yyYAWflXA05zRYc2t6PrQpTB6ME8+ewVIuAPMfoWT3KsoAec/DsxXxXI/svN
EnudJxrdhhL6UZ2o7i2l3F+VRE/CWpN9RECNCK4fYJdLfSdzKeaWV7FEP6Z98sUB
W+sIjCSswIoyX6BPLDPWeVlby/Wkj7yAxhgXSOcrC+9YX4f/eBQMjPhGHNF/zhoy
psr8B6jfpbQsHCHeNDIf6UF0mM2/yFQbsRRXY/623PzcVg7Pnnr4nL8AaqTFPOPC
70LFIqSDp10U2mJG+hQ/A68cUr46gOQdZt+uzn+b0Ys5CD90Ku22f/Ef/gLA7gEi
53vP3yVbHyVXUggtFRjvUwFcutmycbSd5SKIGhxxRkvGrGP4gfQmLdlqWvX9pXzF
LPORpOgTAl/tgPv22y1+Hv9uxI34a8BC2cYuI8u0fWUWSDml+sUw3pMplmm0FTx5
34PzPr657NM4XE2zrf10ac7CBkZTZF2PkytP4PnGyJGlJPxob6kX0eWNROiNVLcv
3O0F/WARzdsUaOw5zrVguz1evg9gTbDj/mdD5GCxXChh4MZcoVNk54engxQWx4ot
iO88orH4Rc8roTZ+ZBv45t6jagDiiIlCnZ5Y9cmsqFnNerszul5stY2hG1hT1mWD
K26LCPqLZBohKRihNL3LJfgundwDPEl9VUBSuxuUAwnLWcpHxkNWRmrPCmHv9SV7
U354av+ZR50qHdDVWyEFNMo9/q1m5LgqUmZ2kJdkXh9mM784f0YAuzh5TMzJiOSP
yl/35UKoevtw+wVvb54tWlvwwVXeiZhfyChbkSwVpEpwow4ANM5zZDJbUo7JU0DJ
X0JIkOFFzI+AE97CUPldCMi4mcxpTCKN/RsSLFWm866vsnI5H/hvNWiN5rniZtuH
rDXoEWxsNi0jTZGiLnHMAb38suObD38BR1+wNaRO8jKPIScwjBUQFIKLQyrvzhz5
Txi8sK64sTN3ZljxjZk6vUJEJt6ffA5GPRlu9ykZYZ1D2Xo30vnKNPXC6dwp5Nce
C7l5RgbeKS5Vzjt0XfjEE8aLcKfnVaRpnCoh+aZgkfWTXczXQsPblVzDwdzWnuRL
+A2cFDnQKNjGJFptBe+QaEHbnvCBZTl2uqy8s0qf24AK/SVLF/JeuNWaUx2YV5CN
XD77VipBuYGRZXgLeigpXYUxZWhC7RUr8Y2uboSVSjjsDT2NIZkuEGaA/LzQUHgg
MIRFreNjAU9p5G7RloZLwkWNJ/tS8XqCkC6E1kJeP5cBlc9/xHcZe0Zq/gye0Z84
pTKShHRLvA6jPFFZ8mQqsZTupP/M5HPZHOhAeMD9M+HLRL6D2Man2EPnSGkqOEWk
AX1YlmLjktXhPpypzM6MWsfSvR8dwwLlfRyvnnYvSXNvASi6sdtLa0NQXiewaPm8
0Cenb4Y36MWCxSGilGk1cyq5+m76jrHsIBz0xkYXRrTNMP5aMXfRaD2V0qNJWsPD
mZTlGVKqBDEOxvjAyARl2GiESAbG2YhY/N1Pf3cF6rPHyo7QgfGlEFD3lPsykfBv
OniC+xW6hmgTARTIiPD7nD2g9uju2s52ubmOU4oWc+cnwYWlOFQYbpEnDy5L1Uf9
IrnSL6zbyngevdhjddVhLS/oGQba1M7M7aj3r0U+iKyM64onQE2HAZikHOMwqaK0
51ax6GJ9fl1T+BjFSPThDHRrfwe3jUYZJwczLpavUvGd5AB0EY5CHr7w2j1vJwjF
VNiwvButyTP7epjHW98ctm30W5H8KZiVsFG3Zl4GcPJVkghjEF8iQuLIJ7q+L6DO
wlDwJmRdeur9hJL6glvT0Hpkv3yAJjjy64RWcjzrTODQdhtJqHAS+o1h2mhFKEIa
ey0V4WNWJ4gV1SvBmcRBgDUj7iUOE+cOHW3qHUDFr6mPnvcDFNf5UBx6ftp4j7Ns
ZuK+HFBv+UCoMNxG6MV53+McAEAmZsTwj7OkEOTj0q3wUVCW5jGBk/QbVUWqm3Z/
5pli/BxUUA+K1o6f6IALaS+OdbsdpSNsfMcZypL877bsfvR2S44HFVadSqi7rq0i
FNB2m1v560L0wrS1xk/nQVgbcZxPqwlk//5KjfTUPG5GeHNPAO6AOKwvH9UxGGKq
YNBaJJvCypaa/YC4mchZoeuMKj3XTf483+CRT3V4unNdzmGH+WaHYe9phLGR7mPQ
zF6rK/8JqzjlLbMFs5PZEWHs9ebkh3UiU4IsceHu09w7/y5emdwqDt3AXDSNBYDZ
SOochiSalPL7U9YL5FiBC9VJyiScnRLGtA3ZphmKBuORdA8kMq12xZ7tRvI3iLlg
o/uAy1qp6jABEZqxZup0QjVnRNPDMLmB7qQ+cSY+8WO8IpyToLcrZmUsgQBmgz9O
2fwII7zqmkgA5hrsnNDuNirGSPsvSVmOi+MrkhhMRcuKN90Bf3nOaYwwQYjUhxjn
mYSZsu/Dln0ea1BV5+NrB8vytaK7E7PqHwbhCkek/+Ves22ZoIl+qGcGUFeWopNk
j/ayjOUxhowf+R62RCZ7pmg0wP7YKcgmC4lwojFJJMb7/Btcd8hhJQyYgfIQgzYl
ZHOGrapqH2zrMypPGR0g13Z6Bn0oUn98Z4bUjP9aNpe2vp+CalQeN17NOXKViLke
7wrVGcrA4wm98al/Qkn9693x4qbeeMqGNfFbpi13SDFFHc8mfRi/tKojODBMwAte
Z7cEms0TPGY3wLTl3XVpFTvDxlsFMw5QgjvroGL4PIXF0VGv5xLUFZLePky+fd6O
OqhY5SgHrDpa3JJ/uoo4P7dJPXTqkBA/ZbyVdkH43Dy3rluJiYl6rAMcKJhRsPjg
8nCMt5Nr5a/vQHZPCAeZ/y1CzPUJWKQKwHEKm5W47xnH51ULeveiN+u8aejgG6Vw
JaCWrGEMMrniEtL44HnLX+lQY/o5yOfvuqpSsHN0kwy+xbmaGolZdprWePdu6v+7
ESN4cqqcpztn/vB83CDuTlQB5jLISdoHtEHDhEV1+p4MQZyOapiA6BjDdlSM48WN
MpQfiCUeHQZBXQjo+W3FsPGG3Jcn4G9TEUu5psgOrMdIh5MvjhUlK3BNfi2PI42R
lU69E1Y7r1ZwOazikrkZ0wKllLUQSZqNNNPrFbOHuUTy4AHV9izn+KqQVIH5tmm9
IXO+ILHwJ7lfoIetn9VIF29ui85LBoXNkXBJJkxPln7wKCqimVY6/ighA5Hoo5Wq
3RPI5UpGUYJF5Pq11MwDHlKgCB+Sgg/6FbRsca6ooGmIdx2BWyr7MNcnTaYwbLIA
XkMzeG2x0faLtXtjJYnLvvweFrK9nMWlAkIzTeH3urbuFZ6aAdWESTWf8Tw6ODnT
gJJYn2gLROTvtTclJL3ZpnQPQzLVgk66VbRXNaTRNC6hahSj8GXuEz7n5dt7mH2H
jTF+SvNx3WYbxPUF2mYzK8JJqSFgVHTY4DLyxzF8fcpVJacb3lvJ6myoaDCEIkkK
5M+uA4ZNG9XLghoXYjLJbTPJe1dyfHfRtfQWUVflUm+pFg1DtpAm42uYPIy9vkiW
X0MSbTuTMLUhmpBWSgaX5yEbEhyW4xaYpkRmTvFbPcdBS9yYWRVAepQQCtuIcMzV
o9gf5ywLblJPDPCcjayXj+Ds4Khj5B4ST01AgK1/r270gkg0SPFkJa+EOM6UNOM4
QDHD5KiIcVwq+d/7JF9Iulk8NzcLVsaoXurI2waRRTnjcmNzJrvQZkcYUMX2C2Qe
A7Q6dMt65DNPEaOFb1KQ0IkQOd0+gU5M9Vtag1pUFKvNTleAJXqSkUPw5kvLYwVA
il/GjHD/Xrx96CBUOSouipKD95zJJGG1wGlK5GRTMWoDCS3yyS1xDBIRhTTrXowX
fjZeFZ5b1eZAsUDEyHshx5DgnBtoB002m12NAbkKi8B13xv4KxDjAaRmnoj9FdSK
8RrPrJeESZnkjpU1Cmbp4oPXkPvgeJKAD3068t/eaL8BkofVfTEiqSKfJap1S/ll
14f4FXsnJhmzEegiO09nW7WeNCjvhesC8qsIz178Ap/wASQ24ojePX1gpsBTc94r
EtXOfsLM66S7w6ckU4oY1bt1h7TlfLeKVubGoTpbqkea88c5+0kRBuBAPzMjAQDk
y7Bb9ni7n9GLFwzbjWKTMfIF+ZXMvo4c/8b5nMGItiZ8+QOUQIMItvjJfFPrIomM
BTNmcEKc7+H3W1BmBrZ4hEo0+lU1zXvvVCU4aV7cA3Ti+IHz1cb5juoKHeY5GdSN
ARDuHAkYBxGbGxy8oo8usXtgYFJaEMpT5zZRqxTYR7gWZEdb0XbdTalH9a8ElUm4
IzlBNyIfrjdpJu1UU8F1p1AcVP55RWVhkWIefCA9dGt0LIuppGrQFIFUOCVlqzS9
oLR1d51UhqLHVIeIbfwykfnQ6BqC5W5K7SU8ASvmUn+ufqnhQ1f/pxQ5sd8mtViK
otcYGKYm5kXDLbJpJeQmMWpjU+tyFwDxrq8lnVFAYFFHzMsy5qUssAyCaPC0JZ6K
LFtFEfsgmEziyoPqCNlKVk1yn8wH7v6YGfCA64sHlBTB9WSjWVwMRp0CkABeo/+U
PgYFyM6l3iBIRhydow4oz4mIqnyrAPlHClDxUyatW6HESTFjm/KqohMRkDnXJx9f
nbTXL1fAQwYAGCt3uJlkiG9whRtf71xTwt3i8kvt+Ky3RYRZKkvenfgRuQnU3lU8
xWkC8MpHodrAE6usVlwLzCvHXQ595cgBg3N+YwovZOLG9a7soIopqpL8HEUG5QUF
9j+VS+NvanBMFX+XFkBWOIeR90O8KBHVIMRCz1s9Lgl6leSrpkvBC9erEzKEn1Xe
WtihuOdrcGoUCnF4/8k65GZ/LjAbhCQEwXeJjVXW/iyF+R+dLTJAUyRnQN3D/+cd
Ya6nQzeul+P7FCvou+s/RLopWv/uphDXOK4IAInx37AGBw6/3WwEkbL3F2XYqj7Q
lpA7YhHh2Mo6Ia4J5X5ee84OTCtaWH0kRmYeDrGxfj94rO/1PfHKZi1HPgZrk5RB
vi8rj2NzUE2i7wxHRGlnBZpwTDgDQZuYpEbooSFZ4XUKk1uLD1yNuJJ3jG+WnIIh
1D9w19wn5zU56/Ouxhqu4L0FaY3CMJq3SYqBy8zlZwsFRFyNZgJycp97yHo5yCMW
W+gSRypDOU/0hBpDuZ9dJ7EjLZBKxsIUFziSSCPDzlGvRCXc1+5PKVlV5dFcV9yb
DXETxA4S43Swa6abzA5TECyXp/tH7uz0vdp+3piLxmNMyXdg8sAbfKVzCiWKyEBm
nB0kTmnBvAwHq0GSSOyEBwokXLwiYVRWCWp5oYCgDVc6/R9rkPKzNhbrP4intRRW
dhRetlV6NKLIwc13aMl9S7P7yUYeKGXF1AaQI4OhJcbzk0MzSQSomvpQL5wHs6RP
l52db2zZE3eh1Qd44MjbUHO+ictFuKkrQ5Ontj3gKJ/RZk6PUqwbQdPTNd8Pw6XN
Kuh+s1Klx6KW5kPm6zQJgvqB0jNhrTsCgcvUNLfMi9hlJi3IgmOhmgVEyz1p/A/w
EGA3An0yVPE9b3lDLIp0ZQ6fgsCG1fM+pKTr5qDBVu6W8OVRLvqKuvmO2Jcu+FbO
ck0/yfHgcGmoKl+ii5MbxcT/KexZu1ksTRNlfo2i/8stoliE5SJB0j5XvLCkTvFc
L64YnLDqyq7V3yg8QbsQ0mpIxFGz5FXNFJtlebM/meUNUdeOXWnreUyb8Z5r7XDS
EJT2s2h+ZfF4/eWYk/UUwaFiTr/l0O/+v1pmX7oGau84h7A7bzCFqdllmLo2Wf60
NsEXH7COTL03fF0ehxQ9/4rQ5yODwMgM5OqDpB2cERE+yR/oVfL549Nc1J3yUhmS
3SI8EPiQdhwPcZ/DIUl8ryJTn4DvBg2NxHEDp5/5Yz1RfLsnt/VqStZaJv6Ar57g
MHGdgWlWlc2bGC28PvTatsKI/wl1D7VJfFSilSFuZooMSLtGV+GCiLd9QGP/79dU
neX027WCvuYhW15nl+mw1DnV6+8VdaLM5lAspAD1pnESe3cMwuJqWPK3YRZbYKK3
CdZlLcWnydtVKQpITN/HInkX5yWjfDdwNDmDT/jMqSHltX5VIoTqAJXftVHGdO48
OW8AspfAaDaiD7GlLUYeKrjR8N/0KdNhIGwYiEKijcTlAQWc8nPMj2MjkDPhxUSE
iPGvNLYPAoiQIyy9yYGUGyEFlUAccva/j+p5ytEoYpcaja6r2R7g/E+TeDV8K9N7
GKdZcDzwELwSFMetcWGqG4dXB5hK1RuT8m5BKehW7x27pB6+fElUZRHQzX//D4/2
icf2Gg2QHxDonV38WsjIA7xEFc82/AqjpTK/EJNQcfL/E332q6iEzMZ7t2ksgl9A
qUe+dJfRoDg26PvE6py+/ER377wY8vVjblnyf7fmN5p/yBpXQUioW2Gf33HnBtJz
ehMC+crn5knYwfaHTe/luyBglJbfqbP3HNeCGwK+umXU4kYYTjkyB7e9gAbWxm9/
SuTS6aX20EzjNIODpKmbuIJpfLxyiXz0JKVP4yN+hCB5wHHcuiw4dq002Y349Jnp
zXH5DfFGzzQVSSks71I6n+UVq82QCXb5imXlMQ/GdA2Eez3qupDdMmwpaUn/hMIp
F+ZpTtp9RYG8m6oQ2lN9cP2DiH376Tt3EecoRCjz+8fHkTdYAmD9S6PAN48Lih7E
lRVsjfrmbgq3hv5fgWdVqgHeL8/agpSXhGmIOmCjvaZVbhW27ZfCE9GbDIi/lSk4
fafCDZnl7rz+3SrEZtWKwY8hrep+femYH8T4HIF89LZSmiEsn0oajyS1X+hMxyWZ
uFlAoJhGuoHbea+Lg4ibLFVrGrMlfG1Qp+K1cgS5BzggWhfYIAXMZjnM3UYv0CQn
KL0tjBtPmLHwiEUEI14nb9pDV021p7AA40FOye/MFI3jVoPhMrxOAqJUq9rjOsl8
Rzn9gYk5n9ElL7iyyGzPtdfTimAoUF/x2f9RO0dLo+A8vWGkJVdwxmMYhXebUPrl
Rf+kEGKZhrd1DvMRP3aL2lo7uuSAzg4+8oE6fj8M8AAiGnm6wexddunVBrkMdUlQ
vg/je3EjvjGWEpuoZ1J0pddnEKtYYnOkErb0/bqhLbaiqTASvGy2mwlkQYbcG5TI
L1m/u4y1H/dTydn6DPRqXpMSZ2os3tovY7WIH0MLRjueW1Mymfkk8i7XVCdJLV9T
nCkZGPvKuFtrrBf6qclfyCGAU9V3SJ6Ac5PK7tJqOS1bZ5HtLh+0diENoEPgdbra
P/VELJxWO5xA+NltDBa3gBMWBAvHPIqwQDp+KVod0B5FBJKl8KQZycYYfuJK2Vmk
azpKO5SuL8yTCmr3Vzemxn5GgxllyxPvUlPPiEDhMv6hAuPly3tx7GCl2uh8VW07
MIb3YugyAItQmJguCRfEUeLnzxn4ZDZs6Pzh1SRGXbGtm2DAUhYBUEarxuv9iqnP
YC3/YnsHmsnPEhuFYjCQxi4XJc6hGihlQmA66c/FiFZc1jqaVRTwia36J1RHqyZI
geN1XlJXXZeOv6zwob5GyQoDiPZANury1kg64ovchbpBEmaXxyEq/YNzIV6db6sQ
a0sDTbSBHUL0wjTfEFxcqXSihx22fBlGRbQhgmn3usWB8Vru8K13bIHD3IQlIxbD
ne7K0OK7jqhHGjZVxoy5bZFSyaHwABeK80iTCbNxXu3HpAJ4A1Ovn5VkJs2BlKot
Or14tK8jvOmdavU/RwjUacY9MQNidzjzwv1b+kNaEM4pLGMkLhf96jhL3RUMaLoX
Ch4lwU6EPggUSwjaIpkRkdSpMx/og+sVqT5btCpO52sEM8+9rPJJAq6dPJqkeJfR
w+P8KFXDJ8PBwmv5QGdVKuMUdPtQzgkmxPhlDS3v46Ek8kglHkLjUG71QGomuGL2
jHH+g6Gkp2JTR//8k4eQ3lgnepJh3ndvFI18awxY2U2Ji94L9EExotQ9VY7ssg5o
ooXicnmGXIhsw0tX4UjmFYxVgaxS2gCtofCKKL8TAcIrxN9mutlmKyY+wqjMDn4+
vtnWoYsydYL7UUpaspC9zv+FqBgG7ByCkiYSmKYLgfp6xuLCrEQ1+QxdUscbBdZZ
RugIGl+mPUvriih90nwU+KVJkRMhvBdvC8xLQZW19eF0Yqg8M6oMclzEF9KrxqH3
SG9+kU8H8a5cJYaiDbQiOMUGJRGp3w8T0VcNKCwNGbBaPUyejl5FUJNrVtrfZUEC
umD8R/N6SUuTJqlJST8KIusGzaoQPZfnbTEfrrV/3xLIRh2zYx8xzZ/KNmM/seK5
IQcBV0EjF75LvbKYb25dgtUDGnxWy0D7DgWktaFvoNEJPvdC8yFVQZ1P12hQ5f3T
x7ri5NTwiGm5gqy+QO6WviQePoTREtPFQjwPFehJDrwYM4iC8Utmq3r6CIpn+3qO
zxu6kd71ENoRl/9YwnyNbc0S6QMNu8JaKc+7aPNgb8iF/ay0W9rbTfLJtQOaXzrS
6WZ4f7J8vR+cKduvG+VJ2w1YaJ+lklLdEsA/BcEz4omC8fen/8eq+lca5+MxwHAn
vAN0KQQf/dPD2HoYFcU02lPOwjGQAcfWrG7XsKMl41SMYM9vyaU2Q9Kfx5QvtE7/
SdOplWY0diPnjvxqPMPST507cGm931e5tJHc5G7i4QhS7+lZyEKhZI/OQLE0sHub
udhrmKkNsbJISZS71k6tEu4hm7nG0aeoZWhVZ6oIWl00ezO8JI1aRUeh1xBNmfxk
2fRTkf8rXnUDT8WaQTJaqe/WcNbty9bHuZK27XycsWsZ6O2WHNH/QrYmmSie1Gxb
So6mXKbPdAzr38pOO0wyD7JHjnoCh6vFyf+tfz+NdaOwd0JjjE20g9S4BJbnneb2
NKSI769FYj3qEj4tZk50mXzHYOWEzIPxDlBiYILqJvgoXss56qGD773c57pMqKle
resvKOlSHjaE5DnM1dVZiY859q0yudCs/xco+uIT0A3o1bJq7IIvemeAkvAqvWPB
oPp2c1yj4XWzukMAGFm64rajqICxcAFR3bINpwQtQ8h3TMId4Y6EFTqkefZKnU4+
mphyp7LEqG6AhUZ/0M11XcwGdmpNGpxvCs8DFkIXlI+ccVbE9sFEJJjwLOSMmZ0a
Z3JuRcJsExcZZpghc9bp4+Bwiu5o0tCM8xSQHyybYJFqSPXUzanHJ2Q8ezEXMNUR
sQLqZ/rwps8F3eil0n3Lidlt+9cOMrnG1Xq2XSoESKrbqnEirL1BMFXe/HQvogDz
ISg1P/AbYxRH4UERhILHdQ10f637pXiILsyf0MkVt4oL4MIyZ3nKj1KGu7UQ5Czp
nKs4tCOP8wK/MxSx7vjOU45TaFPXLOy4zYqmeE/s9I5PXr7toop6++tT/OP0cDoZ
FS0uzkH1yWpyH6bEmlsh3YLqP7M5PVmY1ht0Gpz9BhWstBxk8seuaNb3MIj/ZHi9
8Y+GIiD3SecadgEoEjWerKZ3LUFqgNUrrOSDYjkNzA7HYOaJYFRQzO7qxdP5lZXg
6t0UWkca5UZsYfQ+47osITdffYxmMeKdmSy8P+7jSiXdMFPtWQINxIKUU1WyuVDS
AIGBIPrJKdkz2OgkSpNiYdAu5lOa/9NDmuwK8qI5XBM8DNYrsbAkAacsPMAtiNMK
SI516Au8HPZNreAbhg8EUZNYnciIHPA+/isfSuAXVDoTqjEerlrRupNX+rpoqJ8x
FCapMkz6Bu1B7/Eq175bV2lzrMqQBcmC1BiPecJyyhgebA7daWIUtcFi4GQKqDa1
oDf1PzY4N+w48OvP1882+HLiakcDvzIdddkJXDiLpGsxwfUIZM8ImqYLNG3Vy7E0
zZ4DUcv/ej64QXdn8bImFIpm/4o4wll5TMaU4cnsO3QILcRS+eWsdLlF92kx9AQj
ZDp1L6XinDAd7bTvsRANQjS6BlBUsYAVFBb4OcsojQHDIL1EwLJnQMuJGTQ9o2t8
nUsytZvczE0sYvyN+1XcMFf/6Zt+2OWevyRgqnLX2HnqAIkqpUQ/z78smjZhFxCa
OoUP8FHHyOem3ICJJfv7eEGCi6tc68Z2OVBPLX4zTINnJAHa51XBEVGdV5WWGMrU
xQ6oAMcsg5aPal/07AYXFY/CR0Ypva58t/8k24q0Wn/XIbulKxn9dICi6VwkMfC7
2rBG1CDl6kcdULyhHlqYz4rP8ZsgC7BOcTPllU/lOG8jY8SRnXLDGNBe6KW2HViB
713egSH14PSgb6TzC3QmFMq/cBHAH33unUZxwnY3ogWS7CDoF1fSjZ2/sf+w1MH9
Wt/4foPtAHDg4wO1gqNy2zy31dXDrDAgXNGaojACax/DnsqlzAndxUCOOui3XTOb
XejpJFwnrxbnt+24cuSk2hofBhRUOMhcBW7bQ2mR92ZLbmE4N8V83eIQUjbfa3bW
53lGOD2E8y9gkwzTfQhwpkT9/9aEo0qSE03VyJVc8cq5LtvzgM+ub6Doiyv+ufX6
O8ZBIPpBiu72G5ivdlsHxU1z7XI2kZCqMPyHSLRgbGo4HCcQR5o43JGYZjZzMVq5
a01n4i71vYCYVSDnKigdLG4GIisPLY2Jb3S3o+iOV4+4z2/Sd1KGHnBPsBQLcJBZ
m32NflGfqAz7B925tVg8Nzzhk2en2ev3/1mZtvwTM+FVQ/9VKbxuoiaYj215cwQk
wvX+uBg3SVF+94zBEMnIv7JLmu1EKNrI+NUgKM5ybzllICH+SK2Tc2b0prK6t72m
2buQOp/dhPeapQ1gKPqPANymBATm7gMJmoCYdc9bfYv7SdYoqq+xdsqK+NYAbwbb
lMC4FQY1as6Ou5cKEkSeicMgiykaDWRkBnbv8v1ahAob9AtcfmqsU78kOalshxeH
NOnhydqgzdWp0SeTuUif6edVFmcNl91S51mD9FzwmxVndK7StR7GMe4BMirvwrKX
VhdH467zr+ex4dnV+ZAEoqOgeGUAFWKcCFykZ+Q2bLVdf8W44SFkFHzAV5aGEtWD
teMliqdiph/bPtQFALvrfHpYJVuRjRrE1THfro9Me6k30dQN1wEMtfTmaRNf1RO+
3wtXwYogZ/3NCF6Ml0wf+WeQg78nBz4gA7opdJfxWrtDnrQQXlTB3IjrbNxY/ESC
yS0yiBq4M3HbzVHaVeRcKR5cdl03r/W5BPXDmQ0Qr2L5srPzmmoO5RGPOH+Kev+X
g3WXpJkUDmAUwZF4qt8aK4CgrTCY2u7uY2bvqwOfnQqpy+cypbEEl5JjY42ff6CD
QJsATic1Xq49c8lLr+fe3fwPsVARVmiK8+ZtTgwdttQWIFZcddLGDbaf3WaZKztl
akrA1gY095hu52Ec3I63l/cS+dgHkQvUfolit0tozVrsGEumcNu4oQtwVt6vT2lK
m5foN1Si6n+Vx+mse+rjgbZ+j38wHJXG0H1EW/t4F9QLdbHp79j0f7GKWXQw5Hxq
pxKkVavSSVWQCSoICjWlSX6WY+rx2AuAonCHHSExGgaGd1UDlDYoHZvWOZQdzgt3
WlkKjBEHtl6EzzjE5nra+cTgkLBtrbF9I8FBdXWMsovQOeSJ509fRzj1WDSqzoKR
3LMb9Z2IPnM9H+jnbErvmEoadQ/0O49BzmUXSjUJm6duGZ6iLFCuFRAz9IpP2QNF
x+VJ1XOwkF3FgRxBhC8plycgzsgMQkimwSwyWA3HkSQ/8cMSUDu82mXPXAxpYGkj
/8eqkox55QcgNM6jGPKSce+lVeEFvXaNXktKeDH7Cnm5k04G6PKMCkpg4s06TJS7
6VoB3JtSA3t1DJFfc5rWgMXSiAwipMgt5UP3GQJfUGOCp7kq2kwWA/EsuMjpzuFJ
Z/vwFSVqGkmII17hl4wQon6MrBBr4Z2du/81EWyQyL93bF+vMPnpXpHcMpRXMmg0
rvDXEyPXFPBT0h6t+XWtAJpbCAlmhDKiQf4PfyXlGxA8WWX/r+/9hCmO7CO3s0eG
IPTQM6Vf/XLlAOia2Cp+Mod4xmydubw7pJqwb4kGmkYtkXglnasQIXndlV5VuU8e
Pbh2+bdC2oFCR1uF0E0d/sEsPsYyc7H1G0Z0ItEEa8IJAaHNeH+EprEGBwvKBPr2
9xC6E+PJMuESybI+tOjBwzVhxItOcS/++Cs/e2Xyw06BqL8kkzhT9ZL7Ac7dv9d6
PZq5sgr4GGgh4B2BFpuB/uY4dsnwLfQ2+w6eyeNdiV+ZQCeKnrwA7u8C4BZ5r+ao
0/KXbpdxeWghznfHmXt7I/tr0ZlhHlBBKrkKihPBriO0gh6w+YwQDEAqI8Y04v0v
IYrQu0xwk6s9svG/WYBoZhhPpJPYd7UFIuD6zIF9L0JVIzpGIpWqryblRKKe96Ho
X3VL4qV0xV4vqYscn2flg+xoaSJjSfibCHWODFw+XhN7+iOohDd9cbJHKzsaZXKp
j/N0UI3rfxzEYaSrK9t5hfXchqtsdKnv7pDirHqRkqORf1LyZy2cL04Pzj607Xy9
3xi3dQDXfH2ItHZNrj14s86tCNtdtWRpwJW3X8xKsBJGY6NHANOcTMaHp8YqIGlW
xR2AAYU6UDSuBJYkANpsXWo7HVaJPlwRKAQiFTmXRDiNBZxz08q7gW60Qqune7S5
t1p3FTYP5UkmSaz1JKj0To91MRcBILGzHVw5Q5Dn/pHosuax0Ct4P9PmT/+bqUhr
E2Miv3dDKbgH4M+kHmLB652Z70Vu2xNNAEiNxLtTGpBoyqtyt6yTxVIW7BX/21m7
/GoW51Fgx909kLMZdfrCOW8DNCqcPF/WIwrlKEt89bMxkxDEvG4szhOtRTe2WJfu
zPqi5VpqbLBpdTsFA/ZvLQ0y7JnKCmTK+n/XBWAgMkyag1HA1PKEsjOjFeLI/xlQ
AWSsNX14l1IQ7SEdDBSRuO5aL67VVRrSv58Kapqk5C7RssK4aDADA1yxJ3YVErJB
1dMhqeaP86mAnMACwvnaBikS9Mf/J/ojgs4OeAz2fkstggv8sWFJfklkht2HGmWZ
ALXveEahCqyDek0iYcVtrGI90GcKqzge5skydLgji8s8ZhRp5YPuj+LwY9fjVeEh
6sKsnPmFl0Gnc7kzTIhIZTEtHLTMUhML+ZYhkMwPxIc=
`protect END_PROTECTED
