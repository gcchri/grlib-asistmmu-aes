`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xIDn2cgEHu8klA7Xe7MU/C2qh3rByruw4SxJL8FemmVRBWosljxGI1GIhZLyuP0f
5pKEtSdQKzKptkrCgHE4hFBiabDV2vgW+6uRbl/EvpViQAfYCQyYFkY4j75iivMK
DAiHjlxIvDtk5qPL2CD/MZ67Gj/3OUUSCOW+DixLapqCxMnRm/dGGqbMme8TPG96
zCUWTysfMRG8YcRQ3A8O8yVWpYWhIvgxZgwHqrlK5P9wI21tHIKWzYO4pA2zzfic
BLgRzgOVtMe204XLPqPOKyRQs5u/lvHKFVmv/HE1Onevgh7ygzw4MJ/uKGCOYGDe
6Ex7CQ8zvGPPX4v5fyLAw/0J7m7WWvwLWw0VfBeOTaua/YcIoo/HVo6ZPY0QPozq
14V7e6OlTk50KZpqo0+3vp/c9rbbbNoCDF+KQtSXbbYPXfJzMJDr+t7YejwUK2EF
SeDgBrbPSUGps63h7ZGny8wjpc1/8Ovzl3QCMAXcYaZl/ZFKtZ2veaeBWggf8gik
ogmwRQ1GDBDG3UkcOADsmw==
`protect END_PROTECTED
