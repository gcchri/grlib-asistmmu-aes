`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9LPhDykhHM5xCPkkkQ0MM/3rpADSYOBGHWdhlsVr3cBabiVtpC5/59PcSyjeBve
WWYgJI+yG7wNYmC9m95dWdUYlIutHdz8jK84xrNMCcT3iqnqNAjFXtd66EjRc5q3
qeBHIKcDxYxXrMvd2TAUZJlX3oJr8BO7eam2mGv+TyaMgbP6sSIaCWDvWSXO+k5V
HCTHx80d4tvDghVgqbmTvenHbjCYITCK4SS0wlBXjpksOgGBYEB4xQA9cz+yC2qE
wpMKXmtCIW1dGbqVaZXb2KMGgPhyHrR1c3LQsVGvHREJ+RN5ubNmiZnxWiwTMP1f
oBVvpw7NflsNN86DnFWi5WZOK9N7bpu67OEq3aHYxWrdcCPMnBCIwmBXAnKPd9bs
Lr3IS54flMMXp6fzw1+z1rKA916++JrrZ4BRziPvvSuNTB0wj7Lw7qNLttkUJiFP
32BVZtxNALXJ7JSOBuaZOfhO5m3CSS2fydsXwief8byjDIe9TG+okmgb/p03F+Q/
TdyMq2z91PBeaeURJH0o/fd4QhBN9gxg/0TIvA2NIgOW0zLeYkLYXPDSyMgCMlMh
dT9UpCYNVEfWSJpVygm9r2gvNZR6xue22DWYz3blFQ0bV7KfpSpOfCQVUDG7AAdn
YZdL0JgS1O+GzZiMbLZWb+/xpewUXdfzR5omsvCtuQFN4RoAe+8g2hofwJcn4puD
ecdpIFOboDeuuM8b6Xn++7/Yj/ekQyL2cNkmZINYXaLANX+hOXnFB16nttqwu3ea
gfSULy51/MNWgMAhNmKOhAQihPTAJAkyFKCGK3yRopGOBfq+wmt7nZQrlK4cVefY
TThrFqjvm5xk6b7g0xH9KAQ6PzoZZh4pA1dOI1Th/o9qSpUG24HZCIOiqwEeJLOV
UnM2gF6UBTjoJ/x4l46rMpcTG1XqnfY3T+nMFQOAJrxCa7YeuViMsKBR5xK/eoHC
DEXXyw/X/r8xd+/8F3IHZhz6Tf8F0E7fAXfJXCKnyHcK0N5sxT/e7XZRaQu99IC3
2IM4p47fNSFAsOTHyO9Y3LcYlwUOkwh3Dy5UWnlAscNOKWwDE5KYgW+phM5vmBiI
DjqpqvmSXZHY8E78bNak2Xl3VtZEBhLXGO20Zg6jQKjueSSYP4RwQ2BbBPVnNbDV
mP7nbKzwJ2+WZap3N8ym9qfTj3G/SMoyp3eVgF6GVqHd4APaDbYLJAqavJfrBiLJ
A4APlurOlilDzO+Lgyjpf7030nd39Wbqu5wy+UaAXRVehZ/Uyf5zUt7N4QwtS2EU
gkWOPQijsKYNjl16i/Gn6NqgTJBja+XKtz6w5pca1975D0r3ETXvitOvzHIF92oM
KdK52YlFaDelYa6zJjVzgjoBCny4PdGWlDoU4ei0wCAGpbRkbxfLiiY+MJYiSvgE
sIY9x5XcnTCgfLBhxxc/O0Pj/IO5i6bcPcjXxLlZjqz9FjEgQigwTsDks8GNLnNr
gWfvn4wIeZ7jSeS/RHgJKx4tFNKMa3L+csroiIDHz4loaFp6xYITE/Ii9PfkEEQI
/aPNLCDWyK050k2UJi6CMP7HG3D0KCV3YvJlPyrjM+bSMtjQxDtuMLjeEpoQmVcE
+gN5WF9w6nfXCbiOP+4X5uiwfkjc7LfXowfvNlyQgyoqjdIIH/cSkaO2BP0nhFNJ
IupzEQLyfzJXCKHI3CvQddsE+C5WbCu2ORMC/FKMclEVYLg2zIUZ5Lkl1C7jep4K
gg0MbtKTQNvD1ZRVtvO2ncgAFAD5f2j344OsE9EjMt87E0VFpkW51zKepKaSeIVk
UTUNne6BEIsT87qnT7SLx64AGpnGkLDk8nlVjLMhAE+vBA6txAaGz+5uC1YtQx22
THQM7XmRDeFQgyNpGQqM27C3h6g0F9YuxotP2Asq7RSrY8pOj/pfcWpyUbPl+LQr
paiqNTWb7AiAcY40s+rXfhCgetRYBDU/xQfvfK2vSDCKu2CwT5tTX/T51Ly6uncT
faqDQCAP/w/4ftuoaoXYyJ1aYhqxCGJ6uNRZJZyOj6NIuveii9HVszBkn+sGlV8d
YvvPzFdksW2NfalPoHdkjiSFRLnvDnfmkxDM0FHhhOQWqb4R2hH9hFL3K9YPmd3N
6GCJHiJe0av7L4ghbz0b5rEDdW65602V/wAtPVCuxPzLDnf02z6621eSKOJ+0hfB
gaF8oyJgI2F3mHoJqG8cPpsz82q9LPfazufEu+sP4oyX01EsCMjD6+1Tjl8s0KZq
6QjD3Evz3l+bXVQHzwu+oDWyvXU75KLzBZoKlDpsiyWeM3Lx+8Ky2SS+DElqTGxJ
MbsFKTzfMn6ybvfqpuBSTqB56jqPLCk44ng8W88yJg5bL1NMWtjzxHADlBrZo3lc
56SR7rxoPPAQ2ErxVGiSwJDEv0wjZJKPyNV2L/zRLzsEX/o3skSp9U5yHgux1tew
050keE7FvpP/RsM5+7h9KNUd2xU1/PP367xf4eyYMrIcMVGwDHfOMHLuo1OBnKtQ
523h3+rNUuwD2tXFOkYIoojJHHN7mXWLq35lkR+vQQ2UEsHS3FiTLI4k8xTefn94
sh9M8Dfx8nmJqJK8eO6mo9o4kal3OjIxK7UIbqLZElHrJ2U7KeYUHGcLW9a/BoRM
Ct5/3tlvh1tjubWgkOrh5RTKUl9j94byIhGu2++QpFIRkyX932k6rZZukkYhR+Yf
JrpuEOsjy+aL194gm+RNAB18iduKGZvExtlhR1PGAMvQ+pDHIKk87INdqu1OqjB6
AfVh/4VRyl13llCR1h35G9wGp4V9cDt5yjliPb3LHeGH3ebc92CiQ1V5iF/3aPlV
9OJ58Wyy63un7E/XgXFQhwwxdIdRftzh4cvW9DmlA32G3z0gl49ng/Os6WbSjvll
OuPlFAxehEfJYoUvAQxojuKKABkZqcMfVphks6rV5iUsYSjqnr05agPet53PqhHA
yXKdMjijO7zgl5G6bcHqrVi+skR8wh0hImcao04NbrURrMDkVSpmsyVwVsUoT3GI
qY+AVj9L0xFshZvAepFdVgPHUc2MqxT79Tf1KnBlhtVXh6ZKHeRvlnGXXrPpX9EW
fmSTKHR5Nv2A33sSwbI85j99WcuBpE5uHcwN9WQNNjDR8tRCKADUtK0MHf/TdvUS
L+82b2V40ZMBM7H4BzHICF5mrsxzP2as1/1ZvHI8LVtPwSI9fmiKTjTdv/TEJfAr
cFO/WFLbKUdbn4aS2xJQGzkQAxo6sicKKC9Cx4vdatmq8Xylg+oB+l4v3pTBVG4i
ex1lYw3EsfL6cwRDlLYJxwJBdXBSUYLD8BHnZ+kHO/75vyiUhW9Go0NX5LExbplA
AR+p54zrnIRM3JjdQW7YMByD/TIequn6XOiIJ1wqCW3Sk7bn9jTS5qxEocnnhE2M
fnAFI2uAp6nGfEUXdybdY1ECekCOELRNf8EZ0VcpVZ+LOlooa2QgJTZoFu4beTqb
pz4wcAMGip93ziPyZM0oljXl2uKnhvurkbx63SAErVy3/1M75ipQCA8hSFOPzYgg
c2eNLKMK18x//O3btBRb3eDMCARX4TbA6lObhZo9TkotyokGsu4xBOcxOeFJC7AG
BkEKuLic4NVfWMcoQ6rcjvQDizXQIgNNEzXXQbW0PR8ByEbAzUcd7rgtKA9on7bY
r1vUz2gii45Vt0AtPhSOxQsnEJbh8CIqgwkRjZCBOCjGt/ejV4B76vD5bE7A50lc
Zi1jMWIP+m1Y72pFZk8cnuMKz3eZrELteBlEscUJ+lA4TVxdA6jacbZlRH8yKZmT
5b4BA1LYltIypWgmcv5UKhz9fVN2QnreMylu+hF3jiLb+GbqfL7VJFtGOOAY3Edl
FJW3nbu7y1KCba1PDYMHE2azm5C3EfFyLcpQC+TqErhwSmo/u5EYKTpvRJlxslDN
AB1wq3VnUUalJLT4oVaXShwCpYHQFp6enB/LPUit/IAPEpdtHGyvZ+MRfTsCllLl
Xqfv7UWgs5GkDTi0TKWfmtk/zaFJHHmV+efwns6cF21SaiQVemicq5WJsaKdX6Ho
utv5nWNGH0sS2Hz4oY4Y/MyboU3GhIm+soYzlOjo1mmG5pP5pUbX3HKXe72IsOBa
+K2x8NA48VFocR1ibJJx8vbDDcWMXKbIzAB2L8zsghAxmmoLYgZIhny/6/r2a7cf
S72b9ohUcaaOVLYsIfOqNQrf253wuoTKfqJFbTZzqV9IfnfrNasB9CTYz6hbFI4y
rhjG1FjQS7gHjbwmxzzhp9mi4/bh+BDOP63im4QHIZbKcgMrGc9+7WZH4nhV1iKd
8+H5QgdGmPbmuKCybA1G06ureqcglGGdSkc2Ig97qJLQ0418Mb65eueatjhok0sR
Jg+1paaefl38pUpAtCH3UNNkI7zCdptuLDQoA2xAaiWQcNJOudNnXFU/TgFY/5DE
+IT533Z0qlzitb55cTOYFuPDW3i2FSuDESbnhIx9ZpoBf8iA0bHZ+O7tpD1kAD6b
hDIun/LMWlmkcnACXsFhxU6+IRRfmjtX8UeP7nfMF6A+L+7+cxR4Ci7iWQYOJ5IZ
U2i9Mok5snTLNCUhD0MzPLrUh9ykw4zi4GLbVayAQcNSNUDZgbhBXZgJ3pb/ag4K
eyD6DEXYN8JMTa1JL8ELWtt9zAiQ0dSA5qp+v8xEF7sbU+96xLhUCbiEk/kYFtkd
tEv598mLQeLUwTD8Jwm2ffcKivbk85w6Pa+m7bHV7YhyTJlit3WFoHIFiQeKGisb
4ZAwGX32aNJ2Y3tbPglRuByKn25ruSavPYONknqVr9HKt3RXj7ujaRZbMUcJX0A8
B2F4xy/vtzczrrhW+aRSaiUTCPtzwlPWKHF0AcH7w7Hd/JOpnORszi0ANPB6l0rs
7PymzqjRDjGcuoKDWXcYF9nAlO4teV5s/qTcE3F30wiHCqUZRiJxbvhm0eImUVgY
/jfXE3Md5fwYhKLJBOlMNlXxlgaooDisUQPebt2nKjqEndIEobop0+NqvunZ/dcC
Nw16IcG4c46DrNw/Z6+CkxywSVFiK6QKKtSUBrsGlUi/KGj+06k8ZacZVsNrNHDH
8Fx0EuxN/C5fvSshMG/MahQoLDAgY0F8mCFWMC353R8M4N/htlSGpeD17Y/nNEk5
yVWK7ANwjPPD7bVy6AJhCYd5Uu97NWQd+ymp/ahCzAb+Rp/VzSmjV5FfsFov+w8f
do4QqLmHgJyBt7xABQtG7xAJLu/lUWItFjkuZANxj+JXuOUE6IdSRb42oOT1hSDj
8+fl+2+azEye6/HB+e2EvggBC0VYcXoqLXtL0pC3VZsFhLJIFmIBNwl+ZcSF+CEh
7Pxhoi64tvHxaGud6HyK4MZJwyUIT91ak2huVvC2V91usi1e/teYqayJEmP2Khz0
1VpxsaasQSHHwN87BHVChC4yh9I8kl6oSknIZQoqFmVu5vdm5620ngHraExL766E
zCcIIvfOp4XomcdILay3gRKwRHUZLNoScT087P2knyG8OngTbUwlDvj3aMPqQblb
EnoFTuLllHovkOS2HDnl8Alpvzr9MgBRbm0FHfjDtfbCY975uumXjuYk2TEMd98N
daJpG3XNc5lHTG8mt4/tyB9/R93ACks3Qchy5GTQic5dOQk2aMNgqHiOTCeiQHrO
LYqpgs4JC+DY9wupgrGX2I4811ZvzBIq0MamuZtJY3ywxCcbxQtK9MpiI8VCEekq
+FiRcJ54PqQ7zZlyG9o46ioeVKGc1qeFGcwiqRGHwwiS9Zd0+qqON+fsYica0E1x
/PZ4LX84mkJp4hbaP1gZPxOBAF8UxFx/KvvTvMiot1Nx/iZ/QCGUN8IlhgMMj4Jo
WqwFCBAZveo+ON/J0oHda5paXK8syhQZVdw0nEZZIAYjBUYfU+ruINsBCiVWH6xb
Tw4hXilnJkNZ8HOEqcJlejZrG+Fe80FS86WXEZJxj4Egfhn0GbDUgd37l+em8WMR
8ZzdyUEg1UmJ9mletiPylHRl5nW/ANJdDAQmJK6GV5XpKmbY7RV5wjscmPBHlB+j
poQxokPkxFbx2OjWQ4+DmSmeg3M6/RZanOyI7aTQRXlKuwYyyIqBLCQu4JZOfgQr
gTCuWRRmVVnY7cKI1y3Irhv30qdd9Gfhy1QTveo/sV786cs2ff3evI8ZCQqBdaFF
FuFUSCUo4tFst28T+YRZ6+Hx/4g8TzrIg/l4/Lb2PxYYJSkx63OsHVQ4v3mnUGTg
8tBPOKxPR19UF4hh8ijbhnHekm3SQnawqFsXXi+eeDv7qaVAU7107bngCembxn1d
Ed37eIg4C+OEJMvqf8ZgWsIIcyl1fOdBoXyILF6B0iw5fglfUWTeYvQtdl0GKqI9
5M++dknOKRvndR6wK/vVvWb/nMuRYQ44dCjjjiYSaQnsGpygPgz5v80omdG1m3zZ
AMMk7aEAJ0KCGYBEBLhGpV/eL8KHKoWbn0ycJMayM2L/SRNlQk7YnO2CZdL2ukEz
pU3Lec44c2Lrx77GkRjT0lh4vZUJM5lenz9clPRwTSDJKf0HErOzWOtXMSgGCa3w
jaqHtXuGRik1Ho1rBu1VOrwmXh+HReLN8fvjSVLFAJQ=
`protect END_PROTECTED
