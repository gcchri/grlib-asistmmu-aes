`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C52I9f7oYC/jiK8e4oerMB/fHVC9Vx2O39a5G1YsrSCuEZmsHwbx+fPRm8f1lsSH
c5//VWqRLz+Vwev5fYjwbSIK8dEdTqEC6EKmJkKnYdC0YHdJiX4/aT5dCkO6ifdw
1vzMaxlloypmI6qnddswojkEeWhZx1Je7xgLsy1PSryOnDSjmIGmdOTRKS3afjiK
hmToFYU6kzHEXiainCQ+XW2rrtZecg9RprepwlNX6bCVICxd4l+Mqq6lWQ8pCSCa
qAgfaNIbIPyH9L8LPMk2nipq1paGFvaUcLQVe82vopwySSXClxZPQYCsvTrRenVL
fQOpgjc5vFCPL4US/l5z20t6D3EF1CN4egFIjpf1S7dWCBN5iHMkhhBd714887/D
fTEfqYBqng1N0MoD6VUN6/OoGMZown5MZH7blVuXKpnJXRi6Lq9aDY3Dv9OsNCH7
O6hCZoA86fMVkstq9OqzFSppjehr7V0IAw5UQW8+XKVyjnEHtNsASt17gVqxSUR4
WYl1yXyS0GVuWTpK4Z2/MURzYn2tYxBUXIUcsyhXR6JvROudOCpcqoC1cfBarmlT
91XRYTOxKZJ0cxw5ZKwXYdMLikGx7fW2Oso30R0jGbKEbNXIZgkb/xRQgUVjeO1W
jqeLJpFfz9TV6IWvi2dR8SCzQxEASxxLBE0M558Yg3QTO1+YdWXY2dC+ggM3QCqm
KY9KZYxVs6YA6FJ0hUJGlf9RDpvopIWssmu9ljc3C8B5uqO34QTZHuiqCuin+n9p
WtMNrm3wzWyOUvndaEfGsaUywDPk5iXUzg0s5K3jJfG0Yt/WAWyze3bqL6dRH5Wn
bACcwT5s+3EtBu0vDnv7PcqTca/opMTueZCmYe6rND0fFm0Q3EZCVaCIfwMQ/JLd
XnUlMQOqgpqKNyKIwkJ9zejQjs1HfOTd8KwyljoAXmKOSWAmJ5g1tlWHMt/QZnRm
EHmpVze2Rgx0MtaAFGZMwF5PWGOD8i1/Jrg4Yek5AW9Jlz+JqLPPIDfImetuKR6T
XT9xDPjDQVVcAcoBN+EOvJEsrHsFGQlGANe+AOXTkVolep3sRSr3A9mEqVjF7cga
7bzqSSHNyXwr2HvHyVgvSqfKaobl3yfgQHnihxehPjY/pC2Th30KySipYte7KTuA
`protect END_PROTECTED
