`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZhHJLs+NaTMF3RUeOUzki7U8TpVqKlLY6VSu0FvJdc611aSAuuSFMm8QQmBjWGKW
uPZdxjOnZ1Xxx/T8fBOqCMSqIuZetav18isgTcysTyVJGNNmxdxdK9+f2V1jP3uB
7KPYJz1eVlNm19fbASjxrV70bSaoI5FSuxdgMBZYd1PnuV4KRyUE+qYIbJ/llkDN
6Ow1tU8aZ5OnseMNEL3hr001GUMRC3LyBnPavz6G5NAuRHqBiTx9DfYYodfjoc8a
vc84d0o7ReaHY/+8mPvJf8zQez0QVhBalH5RqQ/nFZ4IdmGhXu4vIOIcxdDBBnIA
AeUs9Z4M/bMOTN1VfX97pDw8Who3qseJqsjtsLqHk7sB3KnmAsCfojx7ygle/kHe
uHO5ej6y7V30SQVjltoU17ZgG9PmlWa0VzidUlyWuLYqE+OfVF0U7rVtmfbv+FSZ
8v2RvVa9iO5xaWlFEldQuL1TU2gXyNB1qv3b4LAGAv8=
`protect END_PROTECTED
