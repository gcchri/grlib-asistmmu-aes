`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oiopWqqQ1JdF5N0gKQ6M+7LzuZq4lAHsm/9qK/b/PFzmblbngq6gT7H+enQp/Y90
GDDQYdRaq4KRLNr2T5w+GsCRy03ha3BoPw0N8aHSPDT58chJtOtrRukrPnjI2SCG
dE16dlq+K6PNxuYpLzb6+Ho5QCAN6wNA3chCcGg9EDo77PKW87ruGkOVoVMkljDz
yZwblzFI2dVbWunsnHwYsiLG1pCetc/jj6wQeKAoBxGA/rzpqRCeTfbrbuh+nKlT
pOWrxR7Qm1grz/AMpTHvPzP4H9ZwhRmbWjtcxdP1JYUyb1Qjrpab9m1IztP5KrbF
si6LfzwkrA2ZMOex3hf5kLqMMswQkHl1nFdHR2hqlAu1/JsG6IQJ2YYa3BkEN1jj
J2igJQZjGFHU2slOf/YhgkdMUOk7eJpuk4SzLQxDaCI2jVdGPo5tMP118GYPP2eD
eNjhuWvGHHmjCZWy7vLXGg==
`protect END_PROTECTED
