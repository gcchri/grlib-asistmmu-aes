`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EI/Tj5TwLAzpxrqMWv5Jugc6acDMZiSGChsl+Uf1rmbILNPIWn9JoOncP2+qtad/
lBSDDBaqhg23BhgtBGk66bBDTXEpcF5qvMVha0ml6kk7BbYs26wfpHOaFaqtc34P
5lcH7iE+MsHHCzyZewC8zte6eNYWJQg+FRh3BF7WCdWNgyMixkTinUzkruCvFW0s
a2MLElCmblgYvJnJdNYTNX9Tzt5it7X5QyQPZnyGxwESmXJ/zpmztS0jDjLUQ/23
MX5OmClcvBgDh2kEeb/qP69RJE4DsnmnnB+pYSyn5/gZGnp363dz0bWurChZolml
ydVBZ8r+4Qk3NSA4PNFDZDJp05kCef5pRpsTC8W2ZVkqsDjqDzZhRQO9jBVPMNyG
`protect END_PROTECTED
