`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PfH/X0ZLJQFGZL1PPP8Xlez2CyN2hxklfUg5o9F1nk9WmLKJaOP45Ji8BBg5504N
i1pAD0rEePJGiKb7eBH08fMesay+iDKoPDf5lYHe3Fbc5spaxvhC9yxbyCnac7cq
plilhDaixw6i3rY/GZ4bTblCGazetiVEw+tBb/I1FZAYODpHnuhPJOeRDiXhtMZy
dBLaWCxO54aDcXDShf/Lz2uHiTmOppaSSGoRS29qq/PtIEKxY8nRV8V51SxvJsVT
6InEwpETZmjSLCaFvy7VXV/1BVxnrC5pp1VJtcEEOeaRAOPmxrgsGMWAArs8z35v
mxlzXZTUcykg4Oa1r4ljaZU5fzPmQ4/JM7eP+Z8PrpWqtNOHjifJDTFztywTKJjL
/hwMVDNK7uhHLLBsFnIe2Q1dhxGijD4WructuJ7DMnsBPhZgZCsUstmvz0HNX38V
DdExo6UGj5snJTRvAoxpE/TnoIOm0B0qXoKobQ06qOMNs0Jqwsqnxwuonfxm4o3f
`protect END_PROTECTED
