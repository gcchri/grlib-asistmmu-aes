`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JUkRvyalutHoQZKOTSyzNb8wmK5+EuZczqyQYPfZnKBj4x7KWw8YxRrnpTHNpiE+
CrLQWRYaCRaro3bJlGzp1nQ++Na4pKOOenVTSvMsIWR2EFs3WSZ7xjKOmhQ6JdiK
bW4fru8bxgUUf2r1Q3cmQE61F2LkJAjKXMgwezKYAJg+5HITEV5qAZVpqTimo0BP
6GinTZMWezPYYmRMLUV2v0rMMRMaGTMggC3uVLzxIXDlGj7WlbTkibjhncKTBBc0
JAuT7/6sgsE0ueuyV53ysx+eYr9rzDRYsb5OHj0XqtFxAkoUr6/cpRxqoEgFArof
2aNJYX+zIJqNScbb/uiw6uPaCv+kT6Gq4pUyQ7dqOlD1KESqiGwpueyeokZiRcRT
cIn2jSb7xacqiC/O4HrfvG40tp1rFr5I81UIWhJlHumbXeRRlVbGZIc5duYwn/M9
ex7TlDTiEZSfPQWuF43F44lcKfClD9QJWnkeeqqTd9s/4B+VifBlgHrsL/8bdpy9
yfJ/cP1T8tSCI9ZZkPhJf9Fw5lqVKG1k48DdM6tLUByk7lVd1wRN6n1EBI9/n5D9
nLfyTRxb7gkFk78bUGoMOf4YbogO2U/E2UN9iohqOsHvmPIVZti4kTsKZUNixTOu
LplxGhZ3fh1+xeW567ZYwUAG2Gh5KBJjcYMKTpU5hEOkuHxqqhLofrBFIMb2x3hl
dHZzaaAtq1FZ9cF4TuKbj6a9ae3sodySLMV3SVgzv+fXJL2MumcapXujP6mtMu2c
rJ2Dk8+FhRNjWjeswGJ9ATUMYT7ckDHm9+dikKszrGT3H0q5irqZGdBHoq+tTScc
`protect END_PROTECTED
