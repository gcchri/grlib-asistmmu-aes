`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K5HEv37ruZ/cBh3rVPoY0R1RbWAh6KbVAczMIbzGBj4GOF3UCUhooD6UTDnYnhup
m/QjVc16eiE9PGIdaLgtDzfKf7df3BuUrUbHErFxJIz1XZDNUNZgPgnqD1J/53W3
sM6YEHp2rCIYyJGA2ySzkhnauyOI2EPXPJo2xqxrSaNvw7eteotW7iKfZ7kS51d8
h6V3W9qGf2CT7J3OFVDw3qjmwbI/PMSy7mWRRb9nFLoWI/yrn9jByIdeBggT6DbF
aj5s32WAyJMmz1hQsJgo/ejadaAZ/j2sqJ73dms696mNJbAMsfjeASgeLLsGr9MO
+f8s2U3xq0A3y6jJgSB6pBZVn4Y3e9cAUKs3lluow9ctVYZRgLgqoi1RZJw0LOEF
I3ohepCJPD5Vw8+10if/VL+q5WJUeRotf7v71LYje0Ul1656lnx7K9Rha1ybHlht
oYSEN9azDPZ+2xBRxWxTEvMk+rPskCBWc267QuLI4x41Yd9He3iAXKP/JweqKVNL
s4ke4pN1OIZPvlSMs3AiqtUsHfB6iMokwueuBlSlaUiz8xWVGxx8C7GzZvTzB7hg
DjyLjmE8PpRDkP4f6FnqMQ==
`protect END_PROTECTED
