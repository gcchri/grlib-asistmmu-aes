`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NR4NxZwPbS4B7xe4W1B5KyPVAHnbiXdbbT5/b6RhltkKk+ZuUTZsK3wDWYB8u2fU
QhTHlsIJ9BX2o1gl6CBmmyK9jcQq6wda2oDExKTAlGOpwCDDH0oejH4oQN/zuzu5
OM/GrooqLMNnyTXn/V6+HbFz3D4ulR5LJJ9k25kqgfdpcP/8sUneFly3gRNxegNr
IuuSOm1cY3CJPdhYuLgGKTpiJkvXDaZwb+QaEO3BkzZTI7JlOJeeUWNwfoQWijg3
`protect END_PROTECTED
