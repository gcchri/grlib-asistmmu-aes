`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oNGg8vL74yCX4n94L4ZCQln0lSuHJ6W/bs7s7CvABgkuO+LZxIApVfmhX5uWi3p1
TXi5a2BYI8NvVT6jogJaR+fiyveUVvC8X9NGF5kkyV6GWl2Pj/LF1kksJiur2ofL
uAJGSiXN4cj807iwA4mHvfno6F6ORH5CsKzAHlpJDcmXQ8fKAh8lH8AiFSEMqjeV
J12dgvLMQyj2gFnQl8Jkl1ePeETb0CuplpkAZn02wqDEoWHu09UiroDp1nsa0TSE
3/5nkCV45ntzPocWmE6L9wm2T/mH7BzqSGeI5qxIm9c7elBXwJyxeFWHqOGzRF5R
`protect END_PROTECTED
