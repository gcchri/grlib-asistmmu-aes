`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DKFEQTF0YlGVsmjP8H4UpCaN9G6ikbu9Xe3DqtMsAheLd+/dViJz0gfB3MnKHkxI
OYm7PD2dfZ23SscPQcf7z5KKxKRNvvsxmDSvgu/ms+9e+2kL7t6x4MeAFxZ2t7sT
dU9yyycoTLwjQxRoMd5gCZ/zuJWEa186puq2Gh7qOntDt9sM8X915Bwj64+QuMeU
eumXEqosADZqpFMmlzn7d4Eq9EaZ+8n8lUuWUPO8BDPgtIyIqjJ1oxxQ6geKRZeS
GlbJ91tw1fh676QHnsq6cYmdeQJpYEwr8KPRt/3qsvQ=
`protect END_PROTECTED
