`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f8KMJdEMg7kIa3rtsyD8vP9KaBhTVMDy8PoVxPGTRL9n/SkUQNWPPEAz19XKaRcd
6bHkkynPFgJZPB35PeodspfIcT6nqmU3qgYLWkPJTHILpKHzUwc+ZZhPr+82P6Ks
hqSfn6VkJbD+5nzESqnGbFRoCBhEDK7FAqaoJyjr5rv9IWHvglws/N+mt4ihQZgc
zEuc+noBR8MrEi7TtpjF2kzn45eAqv4ld0YfYf8zpC0IQFJXgP+nF5Yg5MJKseOn
2sSwxOG/Jxt7+gSkFci7N0nA5jB929n8oopyaLelWl/P8ps7HGQ8XXvwmKump6fp
xYp3j2kmguB9tyyEyi8rEzQT3HwQBah7KMOH3Cvl7wOAGhQs29tz9uZz8ZQD7/2F
RftTlQk1pDGCg0XXDRUimmV0PrLrIXNEUbXFt0vCV2m7N1tvleV9IUD3AGVINz0L
I0pI1zk63y8fN6srEPGHqc9C/Ed0FzdgQS6IFwCyYypv7NGD0Edqx/a6oqNltgZZ
HmP8BzaAsW1qtnLjNh/TfcisEas7TOeblD6llpiiA+xrQ15skehtv7c58gWkh6w6
ZZQOQNft7hOLXWiIaBL10ZYkqVr1KoaYr4VMJp9C3kC9bz2KedXBXHbFy5DdIJ+7
yYbQN/tMFyrXPB6fAWAvFWL0aEspRVfh7UZuTqkWt+AAtpF9/o2klWQmhM6L9dLM
KPHlHGEng8D5os18eqJwkAh2uPVn8+oW32+YrMMXOkLB4nLPDEOixrrNvDtgeJu/
DuUvKpNNEREyhcEPIUJ7O9xBSnOZUadRk0OYCvFnLxWEldMHa9Li+kwJtDqbUb0+
poR86Rpj2owrEcfEAmUzqEM9AYCR6M9ILfdok61HChWpkVNbQWnCgXjOw7jUcvze
0d+ESaGBmvlY+byTnIeV0LbxC9HrKcXTxVEjvrImx+eyAPILSBgJsaXRtUA0mWnU
n1jVjOj5CF7ImF50SYoRbjDjH+TovDtQJML2eXiwMsrzRjtUM6AgVUaN6OecA0rr
x8GHRqRb+75ZBLneW/xoGFIKVFqFqdAXcaZ09VQoSSdbAYoHIFHw4sZuKhiEMbp+
5U3G+D2tUu9NCUK2ajQ6goy+LZVA+RQ74/I5sRzfzb3C19/p4q0R+CQHH2XddV54
1i3tS04QZb1tyGp0Flk71HBNrfMv1GMGbrsEgNSKdBRcjEf0wP/pGZf0Ga9N49hr
BFIzEYi0YCCw6Tup6ezMv++ip3nEyuatXs0oO2PhHCxN/M6QDepH/sjHdfijED2I
WopS6UBMKlKOPA0eVKW5mC3Yjy1KMnTMR5up23cVhh2td/VKNmRZRzvjGdJzv/BP
bTgh5/G+QgFJNGi9unUrLw+asEoqQ1wGrOlLgkGohi6KZvwWr+mAO4GRd2hgFVyV
ezGJhRrrmF+C/XEkmFc6qYQQaGJIqkgv/o08pD7+R3XfCcDgi5LAkXH86fdRI2sj
Y5vMY95dNKj2JZnzd5oTmS2oKjqFHPJ+SncJCTr4p7tvQVujAcpVx2IzWF2AA6/A
wqxlbbkH10WhZuoQSd0TxIs5B3RxKSG0Tmc/vDcKaYqUvBy9m1PsQPBm8cUDe7HF
J6ovnDlSg87mBLArH9oyrQC7fTMTonElE4wip3AAinabxK5l6ettu9WGcPg1BGnW
689wewPol21yHrPG+tsjSN2F8PKBGqaj5W/Ph6O2CsxQq1hXkov+O1iQNAk4CX3L
vMVlxMKGm22p72tDBi3eYRZtJPOuV/lfEK868JMYV2i356fup5xt5nTSlgxBT2+Z
9btPo7oIDQALV7OYQF8h+61OUVQmFuXclY4anxoZ3Q9o7Af+W3S4Byd8derUGXti
v3OwyQnPpY4gWl04GZO29nEuAon9oejQyID7lVgwfU0hOsKCHc5hdqDvJ5sWnU9W
eYgDLEc5NboDCrSbJCMlL/2A2qPAbaQaUTYJKAFoY61C7Vevh9CClyewFSqRshYt
LXCnuJNoYUplYW+3BZGHtd7vZAUTqBxiBfwhDImjLzmJ94JWpGZCUoOGTROwjf7p
xMarJ9xOzU+b6eqTrtS5qBZO/ycaOslkFtx/nhsEVZgDkNVhSzYSDSW/3qLrx2gw
Y+I3s4HwJFiC/QGFagByGLh5NgG1r3bGfDsMiAuhuS9mm2M4jTmoLluFHQUf3mr7
swH6ny/qyFwYFRtY9L1CeGGN33Iv7J8p0JWUCf1m2M2e9bk9c4V/EpeNXNXxfBUn
HE3uvUF0gLgOR4VItD+mC3Sn15Fmp7QsGvGHCvYiLH5MtbbAEO8ZHmOGwkBWLb3m
4+vY1jc3lbmztqUzFtGBMVl363L7WlPVdlz8VAPd7D0tAJiA8BkFhBr9k1Kxex8q
6/T8JmKA32NcjRZg/9poE9WweziKNPL2xQvyMHvGvt394sN6AcPBkivOiG7YaBJG
Slu2ynvz8egGraTtOQ8wXuiOb+s1XvvJRJAxadvUMCH6Cl/Mtj415jwnNxsw6hkl
ejhp4er+KRMjNSBfTE8h4K52C9gyJr2WGKIvSRIhz8iYxwW9YUwqREe8gonL0000
b9T5EWOVAsI0yRfiIE2zoIVxoNG4k497c4bty034H97kgxVX6TTXj4r5qQcvX3F/
Jy4Cey/xQq8/D1ahiZyvvpNHpCvNY8qcfI+2WbJuibw7mz+KFK/H1tsFJ22SdhRy
SoVEvjMR4gDd7+BlKXVMAONfo65KZI0KM94JHgrjPWj62PKDMd0G9iumqQkyge/T
VLEN8cQRxAWXgR2Yvy0ZxUYTKYpmfgxJf8pLlOmDThoI4IIPCxbf1odPl+dw9XH9
tkeF7BmRmkqLJvCntdPkcTq2p4Mt0nqvn+FMx3zKRptPIx6xMUwWvlnFgvvasK18
uB8nTKt3SwZ0BvQ74jdtPVLbMAB4qlnQlsxv0X26TveSjecxqlxmw38K/mV/kRWJ
76i01i6oyXtqu2WNT4NqhrYtAJP8pz2TtuwXBKN5dWjmIZNvLQ1EugtEFV8G4u5/
pAAD5+oOn0XapjEtwtQb0mLniTexFxbUb6vI/9A8NJJ1BuTrknTrr89abb581hiJ
VBgXVTv2lMkue38M5tkek5SDFJB4+LMiBKbwXfKlPnnkHYNCRU2cKGqXb3bqGlDB
hXeH/S25xCOj03CRQ67eOR3AxFtIl+55tqdPMiR6cgXy2UrXRDv0X7iM20AHEBwT
r5jtQaeanBEgUYjxotiWPTw/m4GiFuuqIEUsQWfgODLTrLDLiPCYSb0j1xdta9/Q
Le5qM0J8x4/ow8tc+uk56fNEXrbMwU5WQYdeIAauyOn2xIRRXmYCzuBiOWGhE3mq
+A+nPVO7yrg36OtF5ZyZ+w0MDDm9F6Pyxn/hIC9/UYSZIqyHZUeWwJr6wDvcL3ti
jt60vPF5Zh77fN4+6Q/KyOzr4B2GOmiqD41crZvk5UB0vNDmPcusIi6tPS0OaaxI
d/VVz39jlN9mLHKezBmPTSPqjAQOTX8H8UWzafvUBKvAudGjAWLVx/rZ0tdrMzFC
BGBmbnGDVTjvxMdE+wimin+4qZc/QSJ9HSgDU1ZOSerjHAYPV43eYd9tviR/ZF4n
gXcB+DXDHqyU3uqMh2YRWbZcez/Dwe2u64U/XeiMvmt4pfnSvsk5IM8R0oCIf5Vf
J+6aWkLi6iKlMnfH8jyAlYBP/3IO2VkITDTcORRg8TbIaOF5UkZAQOGaYCiOI4Vh
fu4ZP1YM2Sg5UDpB2hzk/9yldVsaQrpi4CAH6fpy/o61MlvX+nEc35LH8nDNXxMp
2JHaVoFCtgCZGpQ1SDB2iE7FoURbWbILaowJp1Qox24TUuNp42+tyaMIa2bCHrGr
I3cnXn5R41zsP/lEcSgpE+BQQzihq4GflsY10oqrcsKsApvuOtzPMZySpPKrglsN
b6S1E2J6P2vaNJ6NrTn9xEm5Su/9EjI701wMa4zPPFNap4HCj7pJMz0B0k+2VNR4
60CyZyjTF4L0r6zeFb7ghjs3iC96jhFFCWYcRdLnFJ3entwzBlt469WGvr6uygjC
XfE4C20HhYWE5EO6j/QDKkskXoaQVBwv21+0Q/0TvcIR+yTYqgG3DDm3ybf9hPbd
Dg6Vg0euno0klLIXJjgI2NeV/07VzgpuDp8c8A1I6+rKkz0AD8ut/BZFEoVLoAXI
wlRTsL3CjeKp09BNFOhy9RDbfiGnw0hAGd6h3OIrgciX8eN1MqDihxE3T9O5XsiR
EPDW7Z0p/mL6LHfslZOyNFNoU1u8Er7eUWkTO7mVZPwul//frV6k7q5oxOq3EA67
1CnkkZRsrN6f4ArXXdjph01PEwhfncS5h2PwFD7pXPbdBfRy06sz2/T2qFWepU28
bQ6CdsQbcJAY1ReY4upx1zKW1oMRFY8BtIIzvdpAtLasHfPCW4YLA8/KjgiEEl8G
0WbIUi9QKKQIyqOB6q6hdrT3Ho4rx8vgssoMZ38C+VZSMn8gOHEIf5qIVtDaO11D
i6pBHuBwNP3xFldK1eaJQhBwVGidntZv311kv6H0GhhZ+WchMNo9asjaYhTCxnLg
NFfOkWY/EcQ+xSqF5m9bBUQsk+d4HM0DBcYChtO0rlWYcLTm94rgxX7X3WDi2B8R
bByqVwGFSsaLEwdTCfgcURPKIY/jCR/j907CDNrqhEAUjs1yZY8LfYl0o3WUfkJr
O6o8SSZjMv0x1sngf6V3eOh0PzgkqXPVwTbWFIyZ6OZM/ZX8qbkQN55+sq5+PQyT
bJK7FlQjmc26wZlsEXv/HaWZl/wCVDqMJdBNlRr82BcG5OEp+zIsMoQQifuBTWgZ
yhNJgkVr/4a+46ngySRruKtWnucvmbsmuuJbskJIuiQBX6fhstOLkCAWLW4vYdkq
77Y60M7WPDcmKjoGXOpfHVEI5Hsb/rnBLWbC9t22DFrObW918rIlnPDKexExJkH8
OnB89w1Hb+7lg1QQ1pomCUjKqP81VRnVpUrGTICzkD6dWe81hcnw4Dus9ZMRId3q
qfHIm43ubbu7Di2H3IkCeLMtlgc6c4BAmLgMzJ+UzWXs51YqVCy2JUu0N3SFrF3r
rOTp1iO9AZZueOLuA83+605R/XeDCaFNWROEhcgKkteN5bATgEjCCk+93lw4L0xc
FkPPt54tEMcYmDy4lP8wiGuqKExTSpmo2hU63uV8e9VuVRNvejIiqWlOdqqXyWO7
LcFXNINfIH7SBTB0fitUxQkf+bzHuqPKq0zsVUpcyQ/hpHqJoDfQtN4nGWZ+Kr6E
w+vftUXZV69ZMDDIaiAGIC3AvaHFB2FPIqYM/jSjrQei8mUz53Q0o6TTsCanvR2s
B3fCbM03VT/6PU7kWGD+iwgfZM62vGbc5q+NScaBzYiR4psCwfHfH6y7m+EcwUdt
BsCxKYOmScogeDzs6TuNOlqTjdYW2x+KOejm/fpM0pMpNS1dvTx80Atha4vdBBXV
kVgP1fImh/zZAGr6ub56W1/PGBxxPz1lA6TwigP0E+2kvxutKZCgr1MRrIR9xsTX
a1+a6gVDxG8t2x+7d5XO14KQQCtYwIVATOIhcc5HZx3f7+I9sLd1uXKPVufWCf45
w4qiASRauTjMQzKo0xoFu/Jl+zV6YvwEDJBJ71FbD2nlmhKiTf9MHh1rTraYa17n
oSguRqGp8v+cBtfeOU4DFL1uro7f+1V+N82yrGtQJ7C20nTitBz90DCJQpHB7Srb
4nxleLFTzpiE+qqcImVBTJC/EZIcAuvHPFEIikcjqcdtIaTiXUtZml6XENuLt+in
6xS3hhhXBjVhRPApaaZSwx9xY7Vu15E3/z2G0/EXsV5JO6w+s9WworkWRZlcq0cK
J7hujUEsyiwF538vl2dVE5tbCmx5Q9KzEUsrjNgPQHwr+Yg4Qw3vb00P4Z5DOqdP
Nam4v/WnA7Gweb6bJD1B4KwdK/Gs5u67BFE1rBKqt9zi82GaS0hp7VaVa7PnWLj2
+W5CdiveAMxWYpDX+t7o7FCgjf0L4YtVwBtbhyK1CS3P5YhiDDJqg+CYWb9E8+AL
v7wdxaFS6QjbhjMsR9SVzCpFjV3ZAdlEvZ3q62Vtss5QXTfkxzV6sCUPgsXhIIpJ
F+c6a2lrMYzx6Kivy2ZwBM2+MeZmzwObTLt5cLkdjLyVpUoSaHsezBxzbFp+krPC
+AXv8eAIvhw6rETfo8n2tRiai8b781HKxdeVMqBEZ62C8cqjpazeuOOxD274dtnw
9Nc51hS6CfJ/8O6zyARULmqyw6F4+/3r3xRfaSmuAqY/5u+1S2UbAUVa1KyTknIv
JJCVsfpv+8cQe+jG+WsQAXkew2gcVKky/fygo8cmCNcQoppsKvnk//jLw8MECbE9
M3agD1dlsq7ZiZLM4CB5XbZ0X04O3k716byjnlGCwkf6ZzCpbyC3N6gMRdDlbUdb
RKb7eJqJv5NJ6HSifRt2zso/GlEepp/8UUWxJVTbtWPvMDTVIo1zg0JZTfJABCER
aROcEiLgYVW638w8NvJ0mcj7dfSofOjafDS9gEv5o58eA4ZYJI2s2peS52xetpf7
uAnKVCZLXrqCuVZfhaBMVyoByonC7IkPBrUMkuKf6J1546ohOgcaR63mS+Cz4LHl
YsKEalRG1FIHPpi8iDbKeVFHcG+ogl/mp6HBGElAaGkuT0f98GuMJIPhHdsPuyzL
02DB/PtxHRjRIK6NxtGhrVQcWHbubDhN3edyYUINjmrJTotI1THOCwvDhDqzLMbC
oyhZSRlTDT9aX2JMDkxgohkGPTUiaoiEigEMhaFSW360aUv34EgfHbON+KKAs7G2
5zCOX4mf06fTSE2GV9eKpH0K/2h7Vp7vQDNadj3Lqdhh0KrOLedFv1voiOZGkSjx
pXk1XgjvV7DeFazbaqIM+Pg70zwr2BFdkBL/jqcQBhvWfhHwhDL9Vx05zx3aAKet
Nc1QMV7ifqJJjo8MuMpsY+o5MYiqXjIXXDU/lEj5PMnE6zS7VaLnNntAVqRMNAl9
Az1XAHGBgVRFQltp2mXhCeVI5lXdSaQGitkKaOpdEpvCumjOiUq6iZ4p2BNxmAdi
ppZy6cE00kFysGEpLrGDwSdG1zNMQqP3OKgn3Vsxd6PgA04XR0gUqzb9l9kwAOLM
E47RGyZ8vHf8nCyqYa7WIPlyMyFHcgwFGLozkNaOMGJn6QK5pvLS1GLKiV5z/IvW
n77XHo0e987reLZRdNtQ4FrH45VEJ1wNW/K8DAwF+rQBldPpzqyOE8SQnP7ySXtb
bUvhifOnLntGEvMEU7DEnRJ8srgq9xlbqiIICCsujlsnkoltKfLeYAkXPEjGkkec
gdv+Uo8SBrfvs++o0MefoNT9Q9E9kmgxYId96U9l0droJtpJF2KusU5PhAuxfpw/
rBnKSoylYiEOIOFQo4XiK6niCH/8WVzOI+oLF2nXcDwOrryUixocN3FZ+3Rhbvua
uKvj535S4V2OxRQPaq+DvGkIGEbdGEQJgNMDE4ymKH7m8faNkeenhptkcXJwVSw0
68NWY5VeKnCm+oC6fhsfyvtcgXtghoxnNqSH/Jhfg+zAlgAVzsSn4Yhy7RuE+nO6
+OPJjSAVIThOdTbc066pCWfclMvfvRFqQUc7CHG44FxZCY+PfLhGQdms0DLMIosm
uMwVkLlyn7j5TI9+zlnQhE33OAl9ek3SHYELjIrMV21q3BhQUOYnEo6MOqRAfGV5
amMuiHD4nziSWaMFqx2u7uIj0FCs+KfaqWH4PVzGXV+FtwqwVDR3+rkXN0NxAO/b
3kyGEteEwU9qQzNqb6oeWB7MWb5nfpM2PeLU1I1BcSwaKGtnrWYojb2QHtAftMr3
k+9zsFv5BlPnQwsF6bRwWtqrhokJD0f0S6sv39mhTMhJE3IDaAQlmzPkiYku7bmd
adwo8M3C2jEJX1vr7d5AkCMKLjchi96YPv7zIkzQxa3o/4zVwNmnQCqyzDgzIH/F
T/eZ01N3DpO2/XXsRF/SDUfM7522QIxkEQhijT4Jod0AAQ7G0dt+d8KSBTDtoKI0
xP1gc2IEClC9nU8cKZQx29zH9sLW/YpJdsNgrtzbpXsRYmbr5dRNh+R/ocyF1HiW
o+D57X7K0AIJrJq5bMrLW1I1v6nTRUcHp+e4YwQxV6/htukB4oXbNPzLP8A4kf0i
ekWZKxfPuaY+RKFSv917d8Dw04SL2RTUCnzgG6GN0fPCZKw3cg/3jnbBMQZnNg1R
lvVmSigvQntjyHPpZJe+DbyrvYTFe6EvbM0noiBRDWJfsDqTGfX8YGCdlyzRvGl+
ZD/lcyJnCxCgDZjmrHSWTMt+8ygvUNWh5HWhDa+ZmpONcJg0oZOrKfm5Z50KICHW
41iK2lrPVSlrMEDjROvBNZH9isQLdqhwAUbbJv6+gnX5+NgYrzcqf+DNCDf8c4Rx
PtwxZDs8N21O9E36izNYfluPKFrRX1Ec6ypDzP5+e31R9wv5jUPuRMcdWsuYQBVd
1UYJiedGlPrXmKT4oP02UvSUO74mwRMmrwrShltdN3F0Pd4q7U5FauZ8tiJRYhiC
opc9oVgmGAeCP6JBeArlsd1r76LLeE01Exn4YxCCci9bxHyTPdvJwGEvSrO80Wil
qIR0hmRrsRTaDd7NrONCwj3qciS1mzg9LWzXkXysDwXZ16vl9EjafoMUM4R7r/Jx
SQjxQ4f42wPoh9zk1rirMCDc1MxFksLZP07iLIO6MNPxGS49mq3Pj+aNXzaaCjLQ
Z9ceeqdYJc4kW0z1VjWXDVqdTgG5VZ1Pia8lCJmtUdnzrNih3Jvz0DkUkxwQvXrq
i19c06S2PGbQm/HOQ2duMGt3KP7wLGnYbp5zL8KjqVFxFJgpXw05Y7AW4i1gWsLx
+bQGb9gmo7kmjvTVNS0lj6d7HNHzZZ0/NgZCT+VONqPUoLtrDYmlvBS4OalMRmkZ
heUn85eq5sUWQ0AXFKB5GhnV3aJdP4yWDWrW0CStsLbbolxs/d/9DJh/ntuas/DI
Bwej9bheTgnrdI5yKumzwhEaJEh1bhWm9BdLIVRgNqeQv4rH4S5gz2/AMFJG/+lC
Ht14dL9qendmsLaQdv311LYVl8GGxcTzwADwjrmFZbwc9B27htr/16knryoB2hpq
9rVlwNBuDq1nwLpGcOFJ0BUZJcCDvFp0zNJBSCPOoccbdaSDORWOlmjNYRo/9kYh
QrA8I9I/blEJT2Vr/qA1zvybCc08q7FZmDzXZSJdNkNsI3eGp9/YaC8zqLu8tsrf
TlWzeZUkgP8QwhYOoXv2kqUeqhDlH5I0o/P3Vd6kWmnZvnPrmeV5C8+Tvn3o0P0O
gw4BTgdL8pR5YPsvS8uKYfXe26VrkJRVu+TX2QrCZA/CCFoIqg9ztCt66bNFYphZ
VdgdnTFPO7bmSUeyi1jeq5z0qrhmwDGX69B67QZGwfM7m4GDhkX4Rdo9SItgUMJr
7BJhpeaKYrWd7DvpEi+mQ7SkHV0bg1io1mapnOKF5GFRdW8uWHOYu+pY3cytQqgZ
i4jnY77pihg8W6yeypxo0RV05JLCrES0+2apDFd9mXsCLLu65EoeXAEE/W7FPrG3
Z/p5bvaEUK9hL99/7hdXV68SEmfE2gbbMJ0yqKFBYcuphNAoBZfEhSxEJwpdQL9v
OGcG+PGmYwMVT5RiGwwSdnYZzgfFKH8iaBVQPoW+kXv/sVpajWu97hZmOk+50L3t
Hvg4leEBxXuDWyhFLw7H5K9S3NpejWtoEBHawZahfMm3fUC46lzZpACymhrrouhT
X+vmlCgxmnue4mst+qjuusTaaIKYvR91YLETzdPZxlTCtfV65KwdVwhMLbUAggnm
yePHZdfyZ1FwiEbDhvm25zvw3y4RC/ebEL/HV9D7U2XafaWeD/iDgYYWSqqLw9zx
VMwTK6AjswllAEJ+Vx9TLnDY89kCymwz+ag4P4Hf4wYxsUaiID/JasOcZfqxEBcB
5jTBGtkMTPK46Cixn01R+mtpsbsKS/I49DouyI9qthvbDNyb2wMnmaWzwK73PAXG
Kr8o2K6Hq+jWaM8nyJCW0+n5fDSZi8kTu2Mc44DTkJ1+cwDYBx6oP53BSTVrFLbm
oSw75ner7vxRETfJSQHbIVbLj82ntlJDGN1iNr41mHVr/9KrC7QjT27+JtZgEih3
x6RixqjrNl7WODpvJY95wTWmt8eVh7MkxSDq0x3jJiqZ5FxW+V8NJCRX4THUtrFU
QJDJTVg7Srn0+1CNqLPO+JxnwXPFnKAJFqZZFasPU0j3IQgxLBPRY/rOxaOq5ive
vvFT9e6duWica4wJqoKB52god26QPd46WEvJ2TWBb7YAWZCqkVsppMNwgyyfvy9j
a1tnaXooqHQBXZnUYPOVx+KR/n12RKFzjWUMxqOPjkH8q8LSlh8MCoBCMY7bblmh
7CmKJWW0GkLjmFz/skDytNj7wIM6jEN2KmJcRo7XfsA7jbF5TzOmnZ3Lw/izZtUT
op/5nqes3H1tKdD5PxNa38HrtpDVrMhdca78U1CeqLAgm50RhRnes+JIISI0uzAl
2xrpsx7P8pyU2IxwtDdhRv3AhLTlZA/zGr8OC6BX6a5OIxrNpkyq0yJViVcQG0vC
MwQm2eVJZEOAf/KGm0TH8BDs6lTz82dUyJwF0b1XPfxOUVoPtLYwly0/9qAxLRqV
0I9HV4Tf1fH5wQixAAn9Lh6HwXG9U6oXcL5JAhNuDn9ENtg3O/nWxSnSNidVTU69
y9f7TJJztYxZVY+Pr02cQdjqzfUsPQUnosDgukBwWLSu6Dp8ftPkrtNT31xSbCr2
k4mAX5VI4aWioOlKd3KmC3kbR7cxnrOmmhPLDyFUMYoZQIKwIW73Dq/OjTRfPcPe
M9jumvks84gAKjBys1DIvGym0v/+maUjFwWCztcQH6htQBvnX0YsrmjrbSlOtWnN
gkjrig4pI1gJfhpTSSkj0b7GTCWASYK1+O7UbjsBXxMKkzazqA1UlLGLn8VYPIzO
1s8/EJFh2LzTTK2+QfaRCDzsNaUPrP/59TMdZYZbjT2nGp8NgCxneQo7qmI9CiLT
E+Y0ccx0d8GQJ1OEyEDXaQ0H1hYOPk4f64X8HK52SjRzulIWBxMURKJLp3dH2z+V
sx9zAOQNZyoeehTGeQwD9j/8nhpROVzd6KhP+lDIx25laSSqknkt/we8YgBNZgX8
lSW6L0fHHxW1jHeSugsxzBfQGq4ut+XHESyRl/LNzcPvVFhSl5jYJT86+As+vQS/
/kAE0zg5cxNtm7/zdcpVWqfB4UB0mGxbQQ6Tz9KTra4BOTlO6gEoyM0IG3B6CORl
Xqzl74G5f8N6G1XNLSn65XxGin7JkMn0iEFxZme/73E0g6w9FIPcMdnjen4IxaDF
EcGSKJw9oiscn3tT8MI1Em1F9p2OGiuK6/ILS+evypZw/eMpBROByACBlw5Bq6gq
7Hb7wr7h9zVmz/iLG57KuPCFaSLuZWwZhAxOYn5lQXIPfXTwKSRUhDUY6YO4JZm+
wihwf3BgJQsJd8Tu+maJwzA7uWAGUgS6rv7apcKI5sV+N8kqFYPoI+OgISAMCt29
RY5YOiTQ7yo7h4rDfoc1PnNaEs5uvUSIKBS8T9GyFWhZi7Zbw1JrYYgxrDXFrWGX
KjqagOpxKB9t2+sfc87qefiHHiv87ruZeuzVcdcolxrZkNVLUqs5XpiqQhRQ8Goh
v8Bn9Jj2ACgHmkSu0JHZFpqfkt5/KOhbZKIY3al2rfhL9R3JwEDuh2pyIROkOaXG
xn0/VCLuGnzQ4h62QzIHEncgvEeiA56+d3sRNygs1He0Vn/n2ohVog4egZPIciir
KX0J/Xi2mioMAe1qjW+PTIV/88MrA8UCTZvKj3KBhqnPH03Tug28mWTs5yU0bTgw
FYe8fiEEMy9o8nP6IbOs18lJn1IYKES8sC0rLzzAFpJLk94hl9uZ+2NdxVmewg+W
+s/0QM2dUHUGVoffSsM2KQ1D3RDyhSsDn+80orc7dJMIkAoC9AqjfjLex+TDL8Nt
wT9PuITAjo1vJ+KgWV7uTKdcmbbO/tLjyclLCDI1TBs0g4ShriA5D1wMxQZ3ykJR
2JeqjgLVJoVHUz12K+2BHfVrd6OQxDvKKKVJJEXc5wQkvustrofhhdho/k47QX2h
XjoJ0UHlINWYAIwiJfqelcBq/kJe0TsEqioGPdEgeZAY+4jnnVSQSldCPsBgz0Gz
LyctFRhNNeZZX9BCXohZ7EScvRp0+toTgGDWpvtYrGn2GjQyWp6d6PEu+U6LawOC
laEWac4LJGdqd+CmhQdPWQ2aeRSC+ra/WEwyC/O65LwWhXWXtBsfjJQlviWA2w/D
CCDRQgAy15+rtmV/ld599Xvwu496yhEn8mpwhhuMgxJXNy3SDAvEstzTTFSrfuBB
j0HOsBoKZ5Dd3e3LmC4r4Zaqw4vYe46LCqGhhAmeVgJjkK4j1HfEDI+Rj//dLyne
ehxBKJGFxx5cujY1AX0gT67fsvny0poADEIBiFChhf0bSTzvJYSgovqARx9pyGuC
6eyaQEhdHGICkc606RS6NwVq0jVoALhzMSM20OBsZKZQL5I7gMbNfNLl9XQzWbq1
KVZdsmgN76mMdUARi+u2LcCYBQdbxJryWtLJiBiLPVl9hw8v4zLguf1sxwIE13VD
/gjA+KPJyrSCXaY8x+9xGM7G4LYFgmEhL6j2L4ju56YtXk5grF72vk4Oa7jAlwH7
vRWtSJMzo+DAoJfHY/NGpRRQylsWXkGYqW9vvsXN7myy9c6MNQ5dWYYyMOHtljMu
FDSRg6YTPVaDP/VWCnPBmXuJ2VRWqegTNP8SdjUTyVOs100Rpibu5DbFzK82YriJ
F7asSm+rsOrPyx7/tG+nfU5Cp9aFHTqY7yQ1p4kZ8SqbQQYHXawU7tXA/AR9Ow7y
s+Klz9nsqVPXHHf3UhcQ699M3sF3rop5y3sJ5bINZRlNNDOHOz2X9o1y2INvco1Q
sedSifFZY4LHsfT6cmATxn58C7RoG4hUIdMwhiKCYuJNexG5tTuQIl1N2z/7oVmc
JetWHTk+vc8IVi0ArdVMCYBohjdpA513kyfi3pb2IwX0sdj30EuqC32IQqHHZg9m
WYChJR39GM5n8beFDYfk0IYKOQLmcAf6onbQ4tqbMdEzZPhxV+OtgIeYzTQOZuq/
h1zc+PGBG3oFk5NwHwOUHM6SxAzMMh8hLWImUuEIsOvr88c9EJRGMHe7uKgY4ryp
v2XDFcEUvOuqnBlkoknyz0e3dNQbnwc5Z3Gnm9z48ar5YR79RO1cFonnGDFpoz+r
S9jU/bfiZpnP/adIEA2xIWObIKrE8kd243DcFo47DDpXfKi6yJWAmLsgJItEB0fT
S2cUjoScY21o3z5H4hL83AjxX+lfbGZz4hRN4G2nnvn7NHIoKCw6cDSOvNsd+U2m
9nwTr1UVbdBqR5dER0mUYliKl+JLAHPyR56H2Vqw5e/jiQ1yV4rDJ5mQPJDHkldl
Ezl3kRLWfNCPLoPLSkE2/vAe0i5SVX4pLh9Z2GQ6RDJdh3LFm+PLsYsCzL95ZoWd
alQfKkTmEmZ+Ict0Yswnd3uX3TxRNygxjX1WKeEI1iVKvgNSuHT+sfhfUvH1Jom4
ikStNQ0Gz3WwShfxDaFuuPCKA0K7guX0m6YWrkS7uZKSriEn3oKw5jYtOVD/nhwG
kEF5q9hgrjXy7X8+VUeT70n0V8oKzxqA6tULiqLH35gIib2ggN5+lIRv0g4h5yFl
gNGzs0I55fQlgAM//3tzbKXV81N80PkrPEJcvJA8G55Nz2EC9Qkq0WAkV5LJ1RhC
/8xpU1/vdYNSwFnb4Cj3NsQtQUwtHakFu+b4uAiYFit0cB66edHrQd798Wba9Ho1
+PEUBsIPcwwvC6jsEC7VZyepMXDTSvxUiNR8f1SQWZfAM3i0Vgf64fXA9BkvPVNV
vkUlGykSr2MVoF+JfwHKbGQdJc+JoffmGuT/nrsZdamUpwQ8KShf50312NGHzUQS
HpunjLF5tAZBQxd1JQ60bz9P6+WE+u838UBCy87fYrDOxkQDco2/mCmkSGABYg/p
1lrDq0Wjl2drS7H/NHTVdudKHOn7+5L2Ki7zVU0/i4Er+Ko8lnN6mrJLWSbzwE1w
+FcDoZtJkCAPmuDOJ3PqRRCqpp6soOOMyg88r3w0LVn98RZtqTvVUlb68FW4uDo7
gBmtoBgIwVqAobdpSssAKVOu7qTMFyszC6jhFQbJFm97OAWulHxO2xv9YIYeG6b3
qqAhKGdf80dSsldLQ+EPmTOqVzBDH0uph2KksGn2f0h7R4WKRsyb6KH2i6qpsLwu
7UCsTVI+qkS4wTTUs6Rt2O1lEhcLzTHmpWLAnawmAuWd+IxmZKz1YiNlzMLMGbm7
lTfWSg3LAoiaLxQ7bdgWsCch95ReJVdzh54lcxIfdBlRn777n6Ytug4z5VKUn5mR
8Lv+lCZAdfIut0DH/7xLGSrR/dMbGyYkH3yrPlXLYHTBnEiCFGdgbZ9NAc5Ncn7K
D9fz/duaNg6mxhE3+68rPYfPaFtpMqc+Wjp6G4AuGMh9wNFJnNmvSD9lI73SsgXV
oOvIAXjqiKAE31HtXBrsEuU+HXxOWI1o2bTrqT+Z7rGkZvOXTb0fQDO6vAd29i+L
l1o4yraUfBOauYZLMJLown3zCatEGdECqLINmbenYnvQh2FYwKoo8srR5Ql9nAPQ
5QTCi/OYwxXaVOYgyLwR9L3Su7JpBSv+kEvkn0dGhPWPH3RRGpSqJFYaistOelWA
9Splp+LoyWxriFp2Q7XpKD4sAfVvEECRdEUXrUsqUnF3+buRhlBlDgBGp6uHV6JM
FTpiqhOzu9L0fAOgOya43v8rkXGFvJROU76+7iKaxWB1RPMjZeSBq3RRgqROXNpf
FyETFZgKEr4fXTmu/o2+z+9MkYGgTldZZtFW7siRboaYJk8ut3WPIz4OlLtW+/Nh
+6JBeF15itf1hIUVxxG/sD2qXrdh2tPbgnJNmWqICvM+KgtR3p4/8ce4smJ4nBdX
W7g2IuFcHFN7qgzS42Hz3rePY4hjPRe8/w18Cz8V1KwzjtgLSOlGOECopDLWTB9r
zk8zMfiKCEdpKmlGha5rSET6oiuMhCtx4d6L11kY2vMr/D+c5ecRYXg2OGIKW9Dy
qDdXZ3v3YYXQcNYPzE3klU+q+O8MaSIKNuvCBjxwVaW65h1eQzItsyClr6IP3fjA
KVaf+mYvV+EhoKMwtQf1NT9qCiBFQkwbbtfxoDD4Q7XLli7qxMBZzQAtwvIsz/6R
PiNa4fGPAGdcFn7XsMYdtHqZ3RuUd/kD20utsf6NIQzjzgNyB9vBRWzwNT+3Q6bb
ThVoHalEvrFKWL9dXksspiJc732N5H5HlTzZSDGKQDOwHppsntj/T0Ju4AT3vnC4
8hdx9f84qlqfMqQnEIwL76l68UJK5Q5ESA52nvl3MoPDADgA9z1smmAWDq7uREUX
a08lOmS8aIyCW8htKaEKoKEWbqjcupURiZjcXHemkel0U0t7QDSqixyKXGWJlimw
TQ3HdU4R2cwkAOODIT6fZlPFPFRbvpE2Z/8Fqt8sMg9tImNk/DVS+kPW0Kz154tl
BCqV98qz+MiOAdTDbLsrwgonAEwpVBL2n1Myc48JwUGfzws5lLk1ta8E+vy0Hr8J
EKlMAwaCu+8WwBLvNj7jEV/v80qECp+qHzZSLu83xpBqGLc88ZpUxMF5QLh8tfx+
nDHux9spYT+n2YJudrqJpNJHhALm0Ub20VZBGt2dlzFCk9/qUFjh4fMhr+LCLRhz
aLPgw6LD5p6UJo2WLuXmdvwZP3YmjENmqd3ReFqGxZG91vNuF9aukuswe1vsiWW1
yESJ72sUL4n2vZdeBEDNhtY5yLb5pQpQCAS0eqrdmrMOZCIcHLS+yQo/sPZ7iKLq
gsn4y7/yiDryjnvGS9RAK3xa8pM4zLqd437b7iTJkZosG0lccFL2m/rOLhsqF/eQ
k2r7FsoLGNmVg/PEVHnp+hsMkbNk/LJhF6DWKYLFlrVSzXXT0HKanzn2B0yFgXGH
JH0pBY+NgpFBe31ac36SSEleN9KMpx6KXelPWV6DKM1sf2LXYRi5D2/tBnzhfcyW
WEMXQ+i7WKkvtmzn71jn1Flk1jjF6Km5ejfBD9F0l/ErkAixDqLc1K9fbXeCOLjk
24r+uk/X0PMK+GWnDDfsvcHSXLr26aAkJmvSU2D7wb0JcUAjW4g6uTJzmtUEdQay
S2Mx7sFTBsRwR41qT9UFFB0JzDRGz/JqNMK328R/9LxU63yTvHDK6ArzPlQTuMFn
yAobqcFDWV+KwtO3j82tXBaIOK2XXhcNU0qPhMCX6YM8RkjQRSqmXNA/kuyDa+tv
HS7P3JJEJH0whyfjKRdz8Q2ABjPuqJvFyFutp7cEK7W/YcL4lS/DHMQYyZF2GXgQ
qtWIkSR201K7JzpIRmXao2+gvrXpKBTFFqgpm2YW8RJGvNVeAuLUAV0K+dJnAhiS
w5+7dUMCTBBdiDe7kdkV3Ssk9zUH+gvcxwrNB/OhNre6op9kMBkFKRgWW4CCaKp0
5X6IwAjAwOae3ZUYIHbEiFeOigZX5LPwbDZDSiQoZCKKvGPdrbMVfgaKeR4unO8O
pqXugQrlf0nyLGNcoN1MFzc4PyHvxsEvRHB+0pQeH9pD9HuS/7ZoEXjUsPE9liMI
ajUVFXl4Q2MezScZFMNXOA2kfha2aDr1X0/TVw2LnN/tgXX3v6QDtJ4FEy6Z+tkO
DDAujDR9SKkMkBNYrxhG4a2JQ/6PCIPLYNR9KjXZ6LdowV5kr9wxaRMcOYmjtIUR
lJuIwDYeflPSP4RSQzBwST+t1k56cHNSfeNIEMU9utbcJxf935eYEWWc1KVxW6wP
DZWhaDGw3Q2AwzWJOndKtPEeCwy+6E4jYdgRzSTNfN/YrcrKIdS8qkvZ7ibpi2Ah
ILx0zCHh79q841p+U1mUMR56ejV7folg8o4oZCrxlOXzR0rIRZKvcd58DqToOuVA
aeQxFVwFNHNKXWStWEcqvWSio5ubckrZgCrMeiuFlK3Ca77C5seXm7mrv2qb5Fkg
zfyxhp1cIqoQEr5UOQzQjtRVHFwj1e35PfJOJq+hHljeRJEu8sBu3+YdU5++ID+X
tYIOs7CRuODLM8Ohi5DJ4bOATORbcveP+1YSvOuQsZeU3e0PxBFxRkBnIeDnLEQz
d2obShr38yReTfvzn1oeIzZ6d7MSmzydtfQeD7O2FT86Olr7z+LJ7Lew1w++vz38
c1Q9SaIyWuCvrrjwKZlf3DE91vjTTD24VuT0daFIJvJpg65NPbSs4tPfjbBxeoxm
7pSvK2GVeIMupcBBd2hrD8fba2GY3aOrVuxO2GfSZvLE2Qf/jFWQebxH08QT5nLr
0J2GPI5TR+IEUqiM0QX9bhBzAEV279SjcTyVeidanaHBaOszhrohJsQGQfsK21LP
lYhHROZWxlyh119qW+RsFdnFRTFxIYnXGh6i2ydvcfq0rcWg2AsV47rKjq84LGNp
FH+ShlJBXcPDCt+NpzpbljZvbZ3qhydEWZ/kbK4AVKAclM5hafSEOyRtm4AYys5U
an2l2ayg5nk9Ku1olFPuXFngTsCno8zCUAZ3mItW4ouAy9W7nyTY1UtzD2FIreNF
5hp0UsoiOZsO10EGSJIuLG6g+ZQvuh2O2hLnmqPLnzpOcCAYhVO5fagqD/ndYs4z
0742MJSv5o8xf7FcuudUbl6YtEeAxR3usg3WHKa7Va1XyBmwotNEBaKuewq4STlG
Zfp19QyHJvLuuKI2mWy0kWqUi3MOV3Ux30dZFt+7EyxPOBkpZmCcwYLJ+4wxpOSW
qC/nUNm2VkvBEkuiws4KxqJQ9pecbEpvAGQa7CKzOiCktzNPFDpnpV9/TvwZbyc6
wW9k69ASrNodtxKi2Bvim/ZooG2n3wC8pgBcIdICEPdQGVKT+LipASGtzZF4cg1t
eJwfA/Nbq1MifT294Ou4vc5B0BeTrEJOzmNPOYgGIqL5lvPIq10jAMQO5yAE0gv3
uWibMgqJelb2zHoYZMfpax3NDhWnoeoE5cdVc5UUK60v41qqvW25L1FLbJef7C8w
JhJy9iFeunie4ZFZR8+3BgKZwL9QXA4QdIYdc6LKTRl/9howbwEwRK/T6rpBAF4I
WIqFwsN516MfeqtxrG+VRw1NCaUZwy7WV+h4yBIGQPxw/6fc0ef1/EOfgsuCTZnP
fVuYoLzHkVrz2SFoMpiRmf7RG6LPiKNpFv8GqYryiolmMTSkZvmxVHx3ggDKX1IO
MIFujdNV3871bprwerOBFDIt42Wv3IrTt8mLXUd6UxOOgi3/iBg7WhzdUMa0QHCw
RDKjAN3TwLff9dXdmzIaVn5u/HKeDdUVym01NDSzAZ3cBdGfNvXQJ1N3rquWeXP8
6EJrwR0n5GkRAA78U1UtpfQ/QzNH9clleuW6N+w3bWqe1eOfOR8Z1RNQhenBAbTK
yw9tMl3qq1T9yKnzzb6SFUgccgqHRHWdBX2Nc2FtB+4pv5dX3fB4m97jEpDAM4fO
y7gnRbcuJU/QLVYbymQJ0cKrj9BQk3Ibh6VxuE1SLg3g3lFh/WCj0aXktySAGlHR
7PybhFpbXr+EQY8w8svkOuIk3UN9tBmoTQA0OmPDqHF3B57LekqVorKaDS4LdnJH
robFzG1/uRH+IoSeq+kCXVOPxJefHSSaU45H+LKygKZvUuxWPBrlxOveWgtPow89
s9K/dAK+oydKCnQ6jhqXxzMg2TVK6Cu5RTwfq41iF36O1SruLPwbS6Kq5BZYoBto
oy7Yz5ncHxcoo3Wf51cTn7GY/7dxiS05I8i8O0fb37eum0crwEuS34zfaZyloxhR
nonjV15SMMEkiR2fjFkERED7rHYMJiDuloyXRK++TaVaSfll06ijhy0JCA/iCb4v
O3Rk50V/XRlUV61Zxpb9cWNvTpINAHchfpPiJ6P4reUwk4CUcqX2HpAF16OUYAho
IQT09sn65h5TokAZqbmNFjWJGoB8N9iiscVV33P05sibEViQzQzWIEE7tjsMvf2L
0KAWB+FYLx/JPxOeb2JnBeJv/00LYyIPVnsj4ae0WVgZEqTnPP2+6eFIZ5H/c2pI
6s+INfDFzdne0CNs5iq0Mi+IVR0anOZjg5YhM32S8+vNyX5GCTfUXa8teTrSqriW
1K/tO+dmtazWkvFUNuIFZy4a5HI3Nwm8bBe+cSxuAa9xPvrUIZP5dAVQu4BWYfc3
MvvFn1iIXkoy8yDXd2smCwylNA60pSEmlB/cCQPU6Fmf9dYvgBsRTfA+5x68/y2n
uD1of3Xn/daQJnfxO2x73cbStXKFyKkC2sH02K8GiUZjuftWe63IarNlJzLjL4uc
EMWzG6zpz+3g5ICXcq28ntkSDKxGWwxVY7sFQhaQZmYN4gg5kQRN+x/BkYeHUyjw
3HpMi5HB98JAmXUy8k0AZlw1OxHVci9zx7re7kWXvVzfn7m9bNty/Y7RFNIUOxCJ
75P6GhKMqQiAoIebpfG9fzlRT2Dzod0FmNiQ77IesILe7KOvu2PF2eTAJPecCsky
d1T3EZe5jGEKU/otJMLhdAfXkd9noeDpfrTIr9/7ziczCzmwak8uZ4gkRDigVpmQ
GLwkUHpkzm8Ktx4Zbz9V9m6aV2b3QgMSrz+zY3WghbGF4n7MRUyUt82EEUw1y7Hc
DDhhxL1ESF28EDAfSPcha0ISjZQKtRW9XReOga2mAFhDF0BBy+RUlVCojO8tfal+
NhfA29gpBrfzB8O1vHTYIBOU7aZFFIDEOTKwyoQklhsW1FIHVyrYeSyRk3J3vmzJ
3UDvCqDQ9UCN3r9bHSfI5xToT0V8VAowLAaRWMGLCbdsq9toHUc2v4+z3sDlK/Xh
vFZ0BohlCB/6BorUuWZV69jaXYXn1lOCD0f7jxYFJlxYE1iQm8O6X5F8pZXMHqZf
yVnQbgdciHVRIADWmeSJ7Irh3nrwWthfdVNtFlTm994ENxuL79xnuLp0sbIC5LJH
/xOUHyoVNJi4jZoDKiMcPCnrOSyGB2egYCLhPsymZW0ZbQdnEHpTt4dIR3w7e+xM
Nqly0wx1S4mRVZXrolGXeLdhc4Xymkg4WBLPmdoFeXn9oVarADGK4R8VYt362Djh
IoBDJyNZua6P7fo5iY0uqzVfDf0CAlq2HQ0RGWQBRrmAmlGV3ZJm+h1AM/7XbFiL
ouoZe8nE+Vy2ioA2Va+BBQsd7rxc0u/C6ZtkSLqq0nhv0tXyjKLINh5G/I2rFQhl
trBPdBmlBgQz1mKDN7M9lRavQd4/3IJLXyN0ujyKSLJh8fBCsjWOqCWZSpl68ysp
oqEW4qHkn8Hion5e8dXA7q/iyvtAQP8HjgIwKQXG38wVbLummTzL3qDUGdnTj5wp
KSNf3JJcebVo/BHnx7p6qpBckGaFoNABjyKaxQLi+eZ/MdLttceOIR2DU7/GE4vO
XFS9xgXuKd8eVUPhZFPy+Vn6YATZjuTbH4RLMJs54eOVcPZHC34WqIG9mAu2zAIb
oXc8CBazzRxhb2CPMSlktTX9OeunP/pec2wzBTSp6NghYt65E9cFCye+0serzESA
q6jDkQ5wHrGV3lA488dm7Gk2h9EgBJx6n06eygSbrfAJQw5UsYdPzTXDUNlwI5Ff
7Tx+DWaYE5Rd3Lk8QKor6spMm9TZltp2jX2PalBYPjg5Swql5lXS6YlwZkMXIhcj
uuOOKhVns0LPxwu5Rr46FbPkXhfX7aRnZyugVqu/y/DPR5dHof7fc4Vw5GzbHvYk
iDGQHgXSt+T/l2nMKQCW7JjubNpabkV9V6PwgKxitWlQQBI05Jcz3Dqh+MtKLMgR
5kpk1ctLGmSRcMratqv7INn9jI9byQC22JClTvn7mDVRDUp3rNWepB1Xqf/4NYo1
eE6xYgMISiQngs7bNupTsDI/EJolye/gUP54C5cA+ekpUxNczEGPArbqgrjSpsTL
GBs4yz6k3GgDQll8gOup3xHDs4HGHLk8CuF/0PmvHlkNgECdwycx+3cJkAxTd7Kn
T7kc4OigVZwPpd1u83GoEDzu7pAx9Jy++5H7ElGCxQYHQRjT3/njkHqEj0hG0apl
sLBDwz7a8enrnsu+NyfdBxsoIoBeB8M0KrflaPLw6fXAXLNNECf8fPj8XgC3OpgV
CZMTdhu74qnA/5pSNFSBoO+ABrTzMLTyVmyJrJhsYkypy0CfVZpAJdZCqEHKRhvK
b2yW7z39730hVe0gI0TJElqdWenRR1lYSMI/mg5HQFKeXvHEs+5LsO/7hjyxzl1o
7veIK8C/KjXCcCqpgTMmkc19aQ1VigxPPxp0QYSLR9s7D0cHC/8J+QuckLxrg9Pt
6zt05qNY8JlZVSyuED5yX/SmEAvT2ITlvGd7aMixjKuuBb/Th8Ut4d8EQ4220CNP
xbu9m3i6WSxbDl21L+wy4OLovpjCB1b4bTuE1x8RbydN3BznJ1yfG4ruqJYmrMi+
Zl3OUN8Mqo+d3TA1fPQhpOM3CzynjT24QNr1MNgZ0mMO8MEsPHIOhfFYOYQ0AABn
Jnsmo1YtkQNdt20TTl79S/EUuJGAWy6CMrpYQxbxMfId4WgTWR+jLupkXnkWbOEm
GU99hq169V374Mt1sYNBZ2LIlh7xpgLU1osT3IGcL8M2prElclMxTCbWLMiRA37u
tMjXQLDjhKrKf88NddTflOZ/+ritioJNm22x//IqsRGur4/gVaEOwGvCnn656Krg
B2BPt2o6exaUHwmBvSfaxnAaRggtSxaCTiyowe9mevkqkunvUo4h772Hc2MRnJ/d
iaxrDMMEfCVBXFDX1XnPJGjNsZuZSft9VXb7bV7lbhX01lNEN0iCut+a3JTBMyQm
RwmHPTvb2EqELT9gHhgZndG/f2KStq0TgHqgQDJI3CBYF2uUd+MvbGzcPVFjX+fK
wazX7xboxZN3O+E6kKNyaIBa9Re2h0iehE/BcYUgtz81KzP6QMtNDZI9Wkx34ljr
QV9ZeDHsXNv/rRHxdM32qWPsSMP70rbhyCS+dtX1uZkWgzEBw2QB4BcZKdNdIQDm
7umapl9TrT6hjSAlD+ym5ujS80PMxs/wpkNOep6JAMyDCvohskIazPmL+PMHNdy+
BNMYIYs42GITwVJfnLIXVZNumCnC7DoyrijJhP13KGXyrQ6lNDbHRgdOyFo3uIXG
EJvHU69xEs5hZ3Oew0naKxBp6JwSZExQXPXxVM5Rp4a5Z2aZzvvcEKjmPxTraamD
JkScfNrbcm7r4mgqGJZTr8YXb11oXLCmURBmpAXjLvNzsx+mlvHB/+jmOKm6HqrO
Nb5XAh8a6D/APL998tGm3H9uiS90Xd3VamQ2C6u/WIXtLVE2VwK5++CCCf7BRjPZ
csGoKzCVqyWQOcEWtzYTyMibPkVSSgokmOKt5Zs9rb3qrdMPrhU11WqgUjMLP7o5
1Kf1BLABhwaPuTuESFAOqaFV0uAWp57HrY9TJr06Bp1Yz4gnxcT/HsTUK0f2prZ3
EyTa/UEcZD42khrxgtTex0a8+NcbuzkhOpbcCehHwMIh7zWu6y70Nj3KtBkFuITF
hDj4FBFW0/KxsnmBLqHRlfNT1lgPG++VZKLGHPg8MM10ZFAfCTM8mQ9WGs732AhR
z3DhOMe2e/4mHzHC75tcu5c7CHu10IDhc/BLmzmHmAah0Y0L01vfe0RLAtz4OsNU
7QvAaXrqofYE/d3KYNLeYp4LG+0SjCSBSoubtgZ+u5K6dcH6a4G3QbRVpDHGzgbj
YJlA3+FK/FAN4WxG8ZoBcAJz+eDJThKC77FYCAApZqMW8nJN7g0mhqLZiYMkpYhQ
Vkhkm4ewS0WZSFIqLDX7YheDD6DlzOcPHRY47GzKImo9buG7NVXaDh5dILCrGDqy
PVFJwPQc+/3SwFug90ugjArXS8Ks+Wc+87G5rW1QSNDML9XhPXlflwYpbAYAVrEb
vSR4YBhbCEdJGl5Jh5TiIPXqill29lKItfvPEeBf4j3cVx3FS45SOeQNl4xBDscf
xGF4kOGKutIlsGTYd5JdUpFy8QTYcbNbDS0e8Z6Edp/0R7CHA4DTzcmiE01fkLMs
osk0YT9/uxT1Tt9rBC9Om7kfENEMr9UkgIouCkeFabyUmShLLLb95fkdo1xQzXmc
ScBJg4/DRXSwuKOKkgBjRpxycfCNxPybM7It/oq8xl57NvLxhzBhqBkBmmBK8zT7
HNXkt6sa3/a1YZ9KL/KO0B9ZHOrxoH1pWASqc62rru0Vi5o6nB36b8zEHgu+3KKV
xQ2gR3O8/XQ87ThmbaPQtUlfKDbgy3FzcYvZB7PSa0sNu+I4RWv1jxnwO12+1lCN
bGr/NrJ3uHKQ2x802c315QA49IxLbimBGO3V/hmkP9B6PFxwa9PKdJsh7tlT5HhI
/+72e89mKePYY8QkS3j+yjETJSMj0Q+9aYH3Y8B4uG92sKOQjvGFCIkibXPAhZ/r
sSJ2jIyhM7nV4P2s7dSSAq745bN8p/hnNm5HX9Yo2+2YnQzu0Y7TOL8TbIMAAo/6
PAaHSY3nFMd+t9PQ2rLRzUeCTWfog9hOVG2jSjcEwJHTQ3lwPH3DQ6YfHjJEswQe
AN4/BBhX7YXfJSeI67zNx2hvmirLcGTuttKjbSLogK2Moh5o0F1bljrxKj19EiS6
uX8LPm3i3qZj2bvqETh6lQD0WqZ4kT2RMvOU9hPTC/3fZuYftlYMkNL8hem0NVjl
QyXasHjHsYLb/tXQYgyTEjPpjE4oDsb2Wu291ikYbCE5pF3IbE8uVT5DVdpruFi/
jd3sfvjkoKkXsu5UKult7o517RCg0W+L6Ee90Hc9U4LQg04PHGsqVTNR7UsuhiQO
R2KnlFHj2d5x8XYihhfqABflu4G0szOXHAUsYoLmTQFyQAXq010vA+jQKZ4KA1Wy
s6OLae2kbgyYCreaSovKcD1jBg6vSHjDKJDZEZIIknqXBF6TqkzXnXmqI5PXpZho
1sbv2ddf9y8wPgHvJp/xMrZ8oQU1v93Q1zrCLACYrV80MBT0vLCbxqBD9by51t+s
4zxW1l3DyAs2BIpHNu3LgxcTZ5Ewk/lKY/iOdAyc7qcftRMh5zsK+0HoL17v2RZp
6KKzT6HCratjK0yLWFvVL8CQtjLNfSGQxJCRc1hqvapDo8ZluuhNDtCibwe6uqBN
M3tmXlTTXg8qx4jA1sax9KHZo/F/QJO9vXdAdvsXWwONqrW9aCy5ReD1ryscd//L
11L2O48NSAIeYUjQVzyw74OYzq9TT9Htexmf65sbPZGSzZaoJNNQAmI96KgMqBY4
foUvL0cGVsrlE0yDb1gDJ0lDLe7uk2T3CJNSjydeP49TKwnCW8sYbzQG/G776jV7
4LX7n/sv5m7r4VPRjMw1FZqUFCsopmU7wW/STxTFty54UaDh3MWE24cY5IKR6iAU
7V2rEVRrFhLMx0Q2cpk6F2Y/QgrDd7HfprcxHKUihvehJX6+/Lg5k6NtRAEaT7DN
MlJ4AZlOFmvATDTuz+QsOS7dVVQZljXdMYqrsG0+CChdgKxBZ6zS5lAGWo637F0u
MMhEn98f2yCD+/jVJUfgJqtyUsQrvlZdiCN/XCSMdHwMbg+2FMyQwmDRUy44wJpY
pcFSBCAdqbdUGnx+AAXac3WakQpX6KVy+IBtN5P35UsFLWHLeApIzfB1m4kwWcrK
zy/8ywwM5DzIuAhmxr4R9B+v+qjgA9lZM17H48GII9bfCehe3H62Vl9KiKlgYD56
SfrzqsHRm502Hp/43Q12hPvRRrjfh7yutMHYLwokNLubpoI6ndWyZJLXgRDc4Fb+
aMO3Psz/KCJvF3rPXSIbM1acOanMobd2bhSpGa+rxGLPovh61HWA3R5qym2XVsmx
wtXi09H29NtRwlQk/b6pZEAewQfp8G7d6bd8HlWnwFSJ8y4CFRtvBX3SKH2d9id9
KbUwWjXT+qHlUd6WEHFYWbWE0EziZLtUqAj5tjvYteYRbAoae58sCOtWTHsWwVXt
AAjWx1vE0ehT61Jvl/AkWqBduZUX8ZDVzCnH2Yloe6j++Uwl6mlbPxpieFcftFgz
E2v8bvYvqrd8kLvpkWzYgQqa2ecNPCLvfKIfic9vEY+h4TbPRlFF1e8Ma+kB8xQK
I9TGiMEbQwuoTz0v0wVCBgXSQu69affVsb8PbigptYWbvwtmerFnxxmsi4znkHjg
mDHjSN/tDfHhi5vWK58cKfE39eY12o6IYusUKscGry385uExDx9tGysNBgZM/9Mb
mL55NAC3UFS6lJFiZapmEuFDTdkLETww4o8ZbTlY/7M9A+rBrnAkg+E1THiTKo71
ZTRYf1MQP3ZpbaJG8yBMx02mM5CY+Dwio1nE/tg/qcHrk/jDVqWmRzxSxA19+wDY
BrpoA3qJgs6CYQJfdzBYqaggn9Yys3Fd02ZH9WCOYhAvvAp+8PNtwAQMW8wUq2nm
HMZ5p+BOoWYlrDBKNWFs8wjq5+u+FGnOuOlO3OdKgqsZE/889MgFpk4LG3Zjh1ja
lW0Gt1+HqbfRa68cQeYvPxu+Y95aBVZrBxiujGJPxElq/dA/p0nKnSJUK9LxuNAq
P2jsykkcYpBhplpG8vJy9Zy02vtZ9WEvyonLwU+0LFbcWy0aOOk4/sL7I29jfdmz
AIUEidbuYJrUgMyyBdnyDE8P0rCJ06v/8hbcn4/v+7DyjDhmRDZhLLQ/vW3bPyM6
ebuu7xOWfFZEhcpkkLPLuBhINWeadSxihCozsGKq9DTNfrPN/BCHCTzeFYEY4/8G
mCd+P3lt3Bxt+tt4n3iHrfEraoIS+Bu/0gtsRIsMezjubQxVPXxNoC0Ns2z0ohbO
cKlmfkjO9mCEO/rG0x4CotckEFyOjrT3tCyy/2vRuOaPXeDYySiKBxWooGN3OpzE
ID/PxoHfnWr6Q9qs4J7aBGsULhwlA2O8dgb8aXs4tcIw1YqsuaV4wUU4qYJBAAPh
MmXExlWDoSlCI3OaSnrvYiprHkoUdl5qZjOWB8O/LGjiZ825D6mGITVp9GkBk/w1
17WNDuQFffEJVkEWechADdOIB/wjNdrvphi92FSmarrPdjSApOefdvocD8jM21++
85PadC5VP4S8+d8Hb90DuJltQPvJbBNlNS8nou82z1Ccvci+W1L8HIwobKtMIDm8
GDiSUyokolB0Fvzm+wQc6OIhI0QV+sfQLzPj1ismcrV6ssEo0lgIexEIaf9Ac6sC
56uoalw6gi3lyJLgoQbYU+sMod8DnnvQtwKsxZYbG2xAM2cvwBcpZZ3G9vsSOlPx
BglQXJ5U3/NJJZjHb0UVZ2XZf0rG688XbZTaUEfVqjTu4NuGqxxR81b8nMrBUGRC
YmB7Zn/1wz0QRKQeHc11nmAxhv+H/CQj6QadjD/A3C4cqVHlXpK74R3DnR3E6AYB
sqOlufdIit9bdhjCSX1uQTNHbbJFQ2AXMHxsiqfaHED9Rnam4a7JvbUYNVudJWaL
+NnMx/a+M1kzOWkOppE22AIxRazdJMiaBbTUWwDsp0hR/T+Bb8dZ+gnT94bUCrWu
5vVZK8QqxRpb0NVXx/0qIykDcJH3JumCM1vW30U7fcaz7fE6Zwa2S6y14awf98eS
xYGsyj5DAIZNl2hyCmSS705GQzQWWupj6LUaU9jSgAJxSVEMYb9rU7NO6hLhWKyC
mBSsG/mQw74IWqT3Qsky4ldSbyI6BC/4PR+DtuSHdhREItbu2i2vkfpD1tLVyjlY
MYjNUYlA2TyBW0PI6GkUjdEWjYWWuesh17AMcgI8an5OGV3RT2NQ5XM1GFz8HoFH
NMGIXdWRJ7iAkajPGRfEz+RQlWm6tZKhlJ2hbGkIOAnV4/6WE6uGquY7/u8akAce
LAjn+Xu1K0AzSK3j6HvmDLaYcJszR8w6QJKKfsmMSefDrPi7Cq7jh8had0BNcz3o
fPAiiG4kXv3pbnR9Tc4Dlcmtzbixo04KLSI7/4+3MJaGebp2orRJsLtKjmS1GEgM
DlDZF/WpMR5DAWEXkH5oGcJIWPERwaddd5WDpda3Cv3iRdN5MwPL7a/KYT+9Cdjg
RDRyJ8Bh2mlKM1uv2I0j3ubCqWFmUahCDxHUyRQL9lm2S/dcK4lqVVxrxQ4Qgahp
u3Ctta8J4VL0FsuzlSGky/burriHNcdV77ycNSi8O4XqEU8BEcp/ASH21RpoqVUs
kk5E1OKMKCzj9XFk/h9fIFuvNMqPqgPV0T5VgOsL6nyJsIOOmECFqmYWhFPnWd9B
MUAPu6lb8DH8dtPIObze//wApXsUtfJUlCf90q/et5J4SEZj7kCTkTzQ6FMcAItg
IL/NdZD8+tja69Rvjm5t7vepeCmHQtXvs2BIsK1p2NPR3aPGTOUVfZOglB9XjjZp
caoIr6jVPUn45hTRoGZi7UQ9iTVrfvsvUWfUHwrD95DOgwkmAciHLb+HFAZAViDV
UYNT7DADiJP2fFT1PZ9wnAAxZ+3zOS7Y979Pu0VuE0zgExOuqjQB+jd7sK/k+MxN
mrcK3+NW/dMk2klP1pUH3nr41Wd4YeV2xCigt7aGpvX4WXhK5qMqgEXrUhsA8d8y
8PQnzMqPlSZeLLBOLlrZjQuhdPnK5JMkE+AwAjfGE91A5sJuVtvXfYGl6ri3phd9
M7cnxNe9rGXfedJNjAxizqB0E8mPnWXyW05ctWq5gO0Wu0YJYYjSP+hI/0sF5U6v
xe2Kdtef3RYOGs8nrT9MYUDGYIzspq9ta5L2WhF0qphA7E+paILQsI7qJSXuhB1W
bjrRG8GKVkk0pjpzz1UElzwgoFbv1RONxJhYhMTu/K6i/HKpjrS6ml4so2sqABfD
t/od4pMYWKwHKzNnDydaTv5M/56FGckR+nDn3Zzoatjh8Jk7A+bVxgAuMNzbOqbL
B7WBjLbrESVDJfwi9VabGumEdUw1UJdXeebkYbkANOtX0TsqW5/ys+bVVHRI2KPO
D1DoPFXVxYhR79aPbepHMxu05zH7Y67gIkgAZnQe116W3FKmNSwq5jla6hQEZ+Nl
iiaxeIMmUu1mmyxqKHRCA9GaTTxLmBqQL4mzcpJubT1r0vOvN8YIbVVaDwjOWfNK
S0XpkWJMAtszaUed4KGODSeYE2tacRBAsrfw4jpVlLxQfqH1YFLt1sQUz9/9OAJM
6L3NH/HQ5yLXrdMWH2kmvnEAv0rlq1MxfFs7r3ZY4trx36q6E7dtPoIxx3c4Tikv
mKZPXrSxL3oj9Ib6q68JmVSiue6oTcwqkkNMCSXaudAxbpfamN+8AwggOleWqjpU
zCCrY+PcKx3SbQESIAZSUztrLEVyXhQLutUHWPjsp++sTdFS7lKRt0whb2EYOg0H
OKiOHgUFjgrS8AERUbQdPgo+JpAEzEkpcHLdYzQoM7HD9zUnghh4dzrBzqnZHwsd
w+b4wbe0qjmGf4Jw7wz+wQfgUjVH7srucMA0JSCDf1pE6IU65jz6ZUeQcgQZeCxy
sy3HvCpvsqOv23d1FH772HrwZTpzsjZZ1c+RMSzVQO1TIsAIPbRUv64+z02qx7O2
qsy854Ani7r/t7VQxGdHDEB6Fz0ufdNYb07rK7+q/BfqE0Zprjn8J1oblApJugi6
U3kDNSAFTtGuLvbbLVgXqQNKjZj/LLbeanuLH8oSbY7HQ+jCaIkLOJC9ZnhWTHi8
krEplP4vzS4XBmgFcSBwdmB+6FoOExyYBOCdu1WXlDnSiq8x+eZAa8RQ0xd2EFJJ
ZzE1atutmWSaPqiuNdbCuBLnIn4tF90VIXzvaLG6dXpAj4U4FquQlsGGI67qPmZ8
/TmlQhpXkmgdJ4PWhpGR5NFzQ/pcDyRtbVzJpj4JNiayzBPXwoQRBfzkE4ng3Z15
pdorwr1xibwzOC29DcZbeoWwmDf/NmtsjvfiEmjxWOWDE2kq6roeU9sTlSaEUI5A
YPKBT8ZoCHao31OMqEScsyQ+2K40L3AU7e5rI0Zkc/4f8ZR/sX5M4vDm59tk4Jt/
IVnYSgFi3waae4Qx6H9gwGEj4igLw7IHwlnRqiCGcAnmKYKOvQDxSDiEJEnAmgOq
1plqnaFYkxAeNBRV5fgSWa7vZsCK6ceM7OEgJZhkqup91oCJ4pjj0Q1eMZqbQC4O
oofguSGW5I8si6VtrSoo8GzPDfkONyYeuVwgXnshYeAi7PdM/svsR+Iu7+OXOdxk
7cifysQ8f70G4LoALAE0Cz59qFFUy0KvjCXapR/JUqa/VtAky8Ezik+1zyjrVVie
VXcBQg5vr99SGbockt0sTNbUheYT/M3QvaI+HEM1tEgER0qJAFH5RVPoZWKxuMdO
FkpsWysyCUCCLD7PniUUNVGg8IQy66frL9maCGusyMaOd4w60AYWV1mIH4oFTU1E
oRexSFzmvcTQioHKoo50VcMM+hMTfibnYalShqAzNc30vXsxe9yk7A9zPKdw3iE0
ZkFxE0qEWiuQTylgHt7r1dZXc/S+wfvWCGxLTvH9elW2han25r8LKYhxQq2DGgK1
/oohHMeXKPfCQvl1neGbTt7VWmskNlNIV+OU7Q5xwkR3txzQz4h3IWAXB0NlXvgr
mJ8XEHlJRb4aiQ47YkthumXxO41OuBo164QnkO05KpV4XUlaT7mIolWH1stZ0ARR
IHn+Ov/cBatgKuAfbgw47nAImS1kYreFUtuHVaYKtAvm0J5nOhBwBzqlDoMQBbYW
d0P7eygHzcDbLGnbm/qHnjGpvK0PhNM0Qq/fYjorJCQXRg+l2VKgP2txppNrlim8
znM6Gu9wbnHm5LhkjUsDcog1M6qF3RWVnmXLtmHYWDhBhwy6sbSfa59bEYIUV2kx
f8t0WoSnXAK4B3DReBwglV5yDSIkosf+tpm+11B4H2x7SwB18ZZ9FrnW+lYACiRF
cxVAykzjXaXyGPsRiGzHyNoAR0lAcjUcZrEaR4N5EAomZh6yHj9MVcxRU86Dl9TG
UHEFsHdnMaZDLRL5n7hUoUkCUt+PVjB3DTNW1XFDIrgP5ssfQfPgKK8rt9bn1g+L
f+R8VYXkrFLYUO466Fl19Mbs5eubK75PMvPACC0jmt/0LQeKdPSonR6+BKNJUnnB
UQF4cswkKMFYzuq5j91Ttf1gL9XZVH9JD8G4V+BLyyQlM4ueZDHRQMF0ZOJNR2pZ
JrYIlUgr5T6PSIKESIAVObTh0+nMKraVQ/IJYMYvyWqjJuHEP4YefGwTQDWcbuuR
ip24k73YXH9qbQL8y7OA5k/srzXVJZ+ZYQ7m8b7G1xaNth7zUw32brbkgq6FcfBJ
eDcIkUDONKjclkBaECOiC5UumuUBQ3I1IQJJ0ijOyKNUOTDeQFlBjaWRfvtRreqY
4z5Nj9Ty8SJMPobFr+ybWCYi6gqBoFXmqzZCU5/ZhWOW/D9jgqsRnVwBgVuo5ilu
vF6eVIyeRPpvAbHB/9aliBqJTmA3Cks8DIxeMu8Q4+brfeRkbKmgqXeTAMkYIylk
/a00UDl3kjKHH7UCVyIhHGHUYmx0K+r/Ys1bFY5JYAYIGUR5PqLuUbKWoAXDUPGr
DCMEMyBn3bb8N2aADL8qL4LKJWPJWQhIyap7tODVhN1rq3Ci5cAI7mgVIc+2kv3z
GvFTNh3V4uo+HSXU5o3hcUVkGnpi2qL43J3j2hFWBhQ7spigVNvInQLHKgXMvnXg
2IaebfLavSpHv2pKHpGJcgQ0G1ZtbaNHxT5tzB2KfwZ3ASzDhXftdeHrMkoDLGS0
REaPYf9UoaELHlbDZiN6Y7ftq/dCHbIfxrm0AFdXEPypajU1UDbLrKdde6LC0LoR
k/qrT7p8RcOOdz4tH/1rrijcthd/+SqH0N9GlcMR8Zi4JctLQDSs6+g6uHET1rX6
tA9bJBPKAoHxI1yubrCsE9dsfVERFmR4irxuAA0BQj12OVlfC7v9dKRHdYnMxFiw
/tN5hbG3cNpPc98nkl7O8cqTGEyeyMeA56u5EAqdLN/WVDAXLHi6RAoIP+vdDVWO
4/cfAJ0glbVakAsnFxiIWMkJK2UlTLOIw1brZ4on4KlXb1+gpjz8Dq3pBtAgYdrB
4Jp4YnDJ/SG5wto4wvBWNSce9X4FsfbNSLzN233yX0MFyWPfHx2bMGKa2rxA7+jb
5LfvIczCrrw1oa+/CtnkMmRslWsp4RP8IeU3uEPNWeU0asIIFy5+DOrbj+IDOyeR
MLCIriZRIDQUYfA/ARDKT9yOCNf7z9q0vF/PcQkr8ewqFR5Gjs/GYyBzPo4OEaKr
feVSijeDhoNrLo2UX72ecWlJnO/ZFEPx7qLRVq1snXcrWpSuM/kSjoIOfgXHbKXt
vR06kX7I9khV6aeYRB5BWhalEkwsA0eXE3SwQg9QBOVtWdCtdPI9ijrVLGpNQEgW
UAU9lqmcRb2swt9pQihLkTrwChXnx+hOc1es0Sb2ck3Fd2nrkOhBzQvDCo7jFoRv
grkh2ROceSGifay3kEdMn2SwY1myd2GuRx4qJyvMP2S+MLBW1Kn3JknBCv7Rh7Xv
PPUg9Fqm9QoO0CI9WL9lyoea1BsLK+3CUMQ84L0GuE/vaAYdzrlAY4oP8tYxLlB/
uGRon/E4KFcjf10FhBUjlQhDzp6yzsJwjphjIESVY0kBu6bvZZ9fWV5tDFZCKxyC
sc7ihR8Lun+md6gm2Isj1AR3pv5YjJfwKvRfqWN6xjT/rkAJ0TOQVLlzICCxjs7y
5kt0HP4TuNBcMShgzXk+S+Qx1VE6vxHA4kwDdwT1J5vhUH9GYX/7qbNdQnbpvByi
l5MWPPEmeP6/T0CJj0xG3rmPUQG2gaYx2i6/XI/tOKsN6i6guWPBwagne2ZSJqc5
/2gOVbpixCKkaFjpP6sfMh0R7VV372bl2tU5VckfDsvZL+SD0mPiCsIzNsSYFjeF
9QjtvZkCh6A4ETfHCWJ0KpY8KMxnlMNkU1IWl7x+IDSGNSdR6/ST5XF2vpLhpDdq
NLSfBhjNH5notJN3Ffb04Mqh2Iufor2kszL8xkNZtDUj8L4j8wud0UG7uY0ypSjJ
hufTAX0uF/SzAw+fYCTO6yKrJRGQy6/BgHcHjJHWwQGhJJXCtkFpyUnYkv8Kwiji
Q0zyleyStzMYG5uUTTEwJvRWnvutMyoyNRtfJaFVin2dyGBosTp6/MhmmmMoENua
2BqwSdPaePGBUQSBWRM9ULvVuLK5p91HCEqqgxFdkSGFKfjSN3f/1RuINPOSrZK2
gW2dXk7rgubpQRA8rQAht3EH2G1bBjNLENDADeU1JCwTRdaz+zgowQu/PRtjiP65
Ev0fEF6hJMFWs3Uj3R4O29eCOIm0CW17Do6Ugfuk/b4yRKTFLNTDUrc1g7MZ+3ps
hnQ7GbdbrW64aAXS6udv2CQpvUu3PADADDgEYQOb/yFIlfvXep0+IEsbLdnCX4BL
m4e1139RZLIgSFULyme18tl/eX4dSYRG/WlF4umOvNd1v75QJsnKqacbY9T672La
5cDgLAcgCBZwIiNPz06URWy5wd3gcaSksWcw3hLlug5stk4bDx/4dg/Gl6GOA7tG
fM88OhZlE3QoV2tTsZCuEbWOWBiwQbBPxYRf6AcX0hoDh7X8wgnVnSMpfEfBQ32x
VRHm2+2iIaScXQdFfjyLp/QLAeSQnqz7ysuY03ol9tHkDk3cu9xasyLoJSn9IZKA
9K6xJIZERfQ3YXn5UtIZrJ9v+ddI32iZ1w14L/AxChMrMhYjOweZhdSsv5hIXDib
GlATJOZzDeNURhWfhJ/Vh6xl5JhQTulknjri8yuM4XibkA90Xkp61fJUewk/xX/Y
1iAJvLu6N1gj3Kv6Xtqs/Y19ZP+Lye9z8trXNGLsuZhPSeduLLoY33eNRA6aPXI7
+HE0tvC8nn4gK0kjDjSpkzpLH5FeX8EMyJAqaB0e/nbk25wMg9Xq1xtnAUvLJq/j
KVgpm0peQzgOgQfIvT+PHI+RiqDB47g1plh+pwBqkfIYKTHeeXZcgMjx3xIeoRDs
wtwzDEqhCWEhhPQMiCdrJSvbXMVSUuvHH/+gJcZrcad3rNZr9sUaEXtJUtyaOcVR
C7a8bHUDYyiOiQnJQZOZA3Vo0G0Am5JYJ64/k0kYbhKuxPl8huQoEKCNTOK5GSsY
3V78aLLBr3JPaNXHZCXLlyGs46HfMLd2yLF9bbfK/bnX67FePtRn2uYR4ySzp18n
7gup3AV9kfoms1fw+R5GArzOsNDQ37CAkLEHM/G4Y97UfsISLkcmSsPXUzn+Nww/
XTqrXvcZt+/nWnEujPQ0D2xd7rPwK9G8MBTRtu588POF6dhegZzzPAiZHEbkXRe9
Njf1wJtOIsvZz9B6JZxJOpvl4CJqrDHiyvw3GM08oTExv7hH6sI6QFIVkob84ztM
f2/AXccH1z+YujECAIAVTjoE2RsG8P2fyktba8+iCzHfsyxd7FggH4cfbC1q12NJ
+XRfuWDEnw78+SyJuTbk/wFrFBIUDva5C1blczJet1RF2/w4XHQick3HrKkcCDrL
jOjMcF/Y/0DRYh9kgjHJL2MTJSkS8V58I4EqbRFka4DVbbSO3oTTVvMPj5F7hI9j
/6HYxxmO9KbokKpDf+ZMry6gCEk7K8+NeEHfKYBR9vP8gms5dbdsYLMVrEsU5Ff0
VCQIykOf5MajG99+gyFEgqgrLFddlvxQOvLTsl2+kOc/bYVwLjn9U2SecTfPAdPf
xn66N8XbNVgyTqwuLjEKy1LE2UCpwTZ/pCfTKAQVrwhoqDBTNR8ulkpkA4P1EN+w
SPmtN/Z/37gWM/46Ul1VaaBD/J89eFN2A7PI0CV5qCgtyc0hpiHtTJg2Aq9h7ytw
F7GxUJlxyaUv+t2qfRTHWjTjEe+e/oHdZZ9jAbiL5MACZjseV3XU/XXumkRpk68q
4XqprSRlYrvDtFJC7vmXmq3lCEV3DyUHvjkNc4E3vcka1xjqngZybzhHCUST1wpa
/CC6Nv7PiiBjEI0O1czFNenfj1t036YGMlFtVeAlUjWLrJI3apqqD2cZ/lVm0935
TIpma3aT2rvHS/Ac0noYTZ3rnwtqnPCaAv2rHYU3u4UX9G7aqC9PhmMdqOoO5MEX
C/ZZtBybvTXsGRNQaT/XoTOkXCggCiSuanInLMrXNMYgZ4L/UmAlycWDTOZBpIbu
BOOomSxsd4ijTmjcTrkV0kcLuFWYi2QW1S2t/5ikrbhUWG00Am0lT3PlEyw1B0Iw
mLgMLZmq0PvJlQFwIYWJeGh7pETn8ZETv+Q/oqKdWy62XMfnP6CpQKP1jHuCXdrz
0wcA+l97iHWcDwxJxGimNamfWab8dlcZes+KcVTAoLS/g71fOwAxqWPJU0hdnamk
pZDX1/D14oUvNUQIabt56+t9HxeYFOknRXNl38c9/5s5mCQWtpNoi53X+jn+Hk+V
mSyj7hwiJkENNpFb3tWRGpbquF0gJySxZv7dBcJic+6jm1BTSU4it7V3gD28WVwO
9xDDBSEFJiNc1fSvSkMa30FwkyaHL6qJHRU9Eg8HtwdkJlcjMC52DqnYyT1NUeaO
XJzdSPGlRrM4SjTaU21iGoLgSwVKiB4q5VtMVMWlvPxYNh1jwt4m1aklqoYTVeu/
MVk69FUlEZvPnS3/o6qXy5/DvwCaTmuF4sxTr7slqfbTF3UB4o/nVfO7VppAiw1e
k1yWmtS47qPry+x2Noo4vorJbFOaEuS4CZH0jRJjY9bEzWZoYLyv7W9SmWjRCn5Z
slKChTShsdNQQfptugxIOq9WHJJOxdWdCGBH5jVoYpLvZ633PiCCJYZfCoa8C8VW
E8YdpyjEszNEIz8VkumQYq5XIEk2KbCnM/LwZdoVSxYmdhACA7IiV2/CnWV4oD23
yF2jMeu1I7E4DEFJPxIESeQEHIF30iMoFzTFZHqzLBVRoLgcYkWFQDKqh0ihNZdq
f33tx5Y4/N5R1jbk/eJ7RkqLNa5V9a1NF+8uLH4M/SpuJgEBM3DGmD/Tf46GIuls
4B3hmEFn2oMYQqZ/gTC5fOgGXi1b8HUYSPc6T1UInRb9K6eykRz8wSvd/2lOAORJ
0q4H74F5aKFR22wwjFT98j8si+QziVCWqdCEsxLbVIlQPHMBq7NE0TVz+d3+IgrX
OyUEoMf6Ml7ikT6fHtqK5N1alKcLV5GVI9AEYcHxvELAgIhfNa8l2i20Q4QO3Tys
ncCYGYj+Dhs81WIeP8qi1GBeWNiLJ7GnhDbBzutrT1fe5paobg21vbzxOcUb6dg1
kki0h6qUCuEh7LUojZofgH7KoTEMasNgbsQBpQ2an1FEUaQHRC77Zt8Ug/xfAAZx
aP57XDtyyyJ5RkczX0iamcyLjs6qEpgAHry+sVBFJ9zotIhpLk3Tu3OnnUIbPOdF
XkNOpt9V87aZqOPz4f4S2+TwaJ9OOqNV0ZOKfhXlC8ArG7le9r2XIF/G3JVnanWX
bIr9cmyZmLmCv7GKTpiwrqNkfHjLkIIs7GoCPfLsXjtz36CKo2AT8RG22s9WV+YP
hBhvfnwjOrz4hKHW8yrdeU/TEvGpXAW53g8woRQNBgMEaJbXX7TpQ8MtcRPc7iDK
L4y3hayckDo8qaWLURBVaomKNCbOjmGUzFtGtEE3WFSrDgwLYLPyKdjmumknwyYK
dkm18bbXsQNqcy70p2eIPMzlmp2S8Yud6QoKU/C07RHIhDEhGnTW6zqMa2umpFpn
Fi54Cr3Q34QtLdKoCnUcjUpg/saJHo/IZJC0peqqCtgPna/mtTEMLYx+sBHzP+zR
dYvrUMTLkGvf6gzd259ZnvSmjKWO2KgW7dp7XhWylm1RKdG+PVY0Ykb1Zs3xxZKx
IAX3TkAjN9TudVKUEwPmjisKworp+TvGcPzpvOYTmTCCD4n2Loe14pxPKydyZ7TQ
tQybn3xBPV/ntFGrJyHmKcu4Iie69HlcnATcGxks4g/ULEDT2fql3qOKmBUx0L7r
mejvUDFbKibGFCpL5bP2t4+SAMhCXpUa4eqElf6cg/jlwntYqzf5OBJFN6khBZQz
oOvx4q8ucTxK+CPvpbARnlXC/1+OjvodoYdqaeZoSWjyOK4ruVNGM7dbzvlGnwGR
s1P9Lj24SlAyWI7DFPiLZHvKmtCofvu+iF8BshWpCnrJJqF9WppNkW0dD1Y9fd4H
8LbhxJrZoL7uX/Q0dSYcCpLEWgnQ93O3xWzjczsVC/2rV9rsl/PIYm4aJ6wWq6bG
I1VM6YwrwcZvBWuXzy+egAE9cmqvcEgrfgOk5KkuAYkGrm3AqW8azVuac6kNMk0j
4FdXgEeIES1ULEzPz3J7NPML3C32scYqzIXkSzazTa6EEFA6/WqxKPE+8woZgd4e
yGr846NKxOHrGPImWjDCYRdCfNmhenNIpKJ9zJFt/7Ses90yqR69caMCotapdqqo
SeJPB4W2iBy1qEJ//tLbs+gCEEXsXPqZPaivXMH39nP6a+K6KbLqg6hrobsGkDB2
Ro0UAxBf3EovyWzBre9haVTkxFiTqDtTl4pYPpn4sX/vlWyhgkYwegcAFBvfAh81
zNXUHhUkxJJvMTYqeNhxhyUislC2CCmYXGlnPkZo3y0KXRWmbageLviRszCZ/cBO
3im8QXb01GIcrvADVnOk5ynS8q3zq76Rd6IOZl/e+bZTEG1/gRopgP//9iLw7z2q
LE3k9xlPK1THtqBmeqC7IkLBggu/UrAUuiObDYSQZEpPITnmkze59ZCDJBC94Col
98B1y9gDkI3CjeGYTtme+MYtJX2cSB4Jla2s5KLXn53ZwhY4LsBnkeavXGwe4nTr
a9iXfsdiGxxTZNRuybytCxmYigGXagt9AMyrBrJ2ETR5sylKgemwpf3G2wHpofqZ
rvCY7tkuuIMWiho3r+p5grgdH9RFw5UQ4Mn5he+WDddzQUF90GXmwwsVu58sz/AD
wBENztRXnT+4a1JrU+4B5k8pYGzZjvg/lLAXT/CXMfQ+HftNZQsjJTbENKpSb2Ny
uYyxvJitCDvD0x8phrk3YwEoZmALNEPtQh1laCYddwXySMqRXWLLzBA00+tWP8pn
3fCw/woyqwQEclZjczTk2B1uC9fAIEa40gQVoK/yOFNWAmON6VRhQKWgQesXpS28
YvGDC6oZaBIRE1lT9Ild0TXGwwBaJiv9Wj1YFl73Lf5MYZbgxHqnF3rkZYTug0Cu
JNWtU0u0+SOstQsRtzNFAIa5Swt3vdA28JyWq+GjKij3rS+yWW6e7EKM/zLQoEEC
aqaEcczMTcnv/tCRT3qg6khyVIs25emWAPRy0AMBps6adkbdw9OsqpKrTKrnqwWA
qRMMLMCQAVLwPnUDLnhVGs4JhBBo13gbhWsRF8384iyM+Hcn1wJA3WtjhJVcgasR
lUcZQp4k/iPtVjb38QfO95mVcQ2HJvakMYyBlyXVIHU96aaZ16N6mlLxbMp4hba9
lhMIXUs+/92En1cUQDTByJkWddaPDpkALGS4u8X3+5TaeiITyNCE0IK2yRewEgBD
E3veCjw8oIIUk/9Uj++vPcylcOQ67/s+lkI2m8MD80FDWPqs6Fu6DM+RhcWYqCTs
CNQ6oFeQpsRO5NXuUSgG3n5nDOkGYeCQyWIvOM458vyIJmUVI78yr1yXfPGPw77D
5D0gEW7YOeXv6j1J4BBPS3pytv9ZxnyTzHmhxYRr9sYRkshI/sklli/c+hBln/WV
ToM2KW1Ir6vfDdrbbB8zAIHCjQOYLH2PRFlKU2xSOsy9X/R900uoaQoWAsaxrV73
TDD7m3UGhMaElzzb4JhSFu1pDyKOScwhJ9jjcjMH3fSUq6ifF7oFkamrZDKpjVBK
QRyJUrh3fQxTYGION1FSH2lFsC7kODMi2kLLF/E/4XTTLbZr6lNKvCCt3/Evp4x+
Ejc3KX3iyCcrk6zW0TFHSX6DmeENPo3854exo9uGCfCFcf1wFGkNo67sSpl6yD/b
1s6sM0wHdt7AQyvUyxmQ5DSFjCgj1eqvk7RvvvPxiM7Q0ZZGEcYiggGufvApKvHf
wt7ycZr164gA83dSTGAFRJAojIOIW9/8WaNpoBqBS0jy1hKp11eq3/noPn12TCJf
TfHP2RYTNX/sDr0jyX2y35hjA9/IOtH0zdct6Apm2lRFAbkk+xD9FpKQrAp7SFmc
DJ1IqIcB5v8Kv1oy3QbaUKXaij7zFvJ71Q83M+7PhcEWrLADo6UMLQjz9fpEoaU5
fMjTXwbRN7IYDhXZNGvANN7rPrHuG2Groc1pGU/f+WcleZ+ijH4Ol9KJRvxIVRcE
hFfZsiSPXgg17qZTaKXA8YvNNsGG8MYxQjsAOLjtUs9VxucmwVk666VPP4Vi+tBq
DTL3I2CP96RG7op9f1+PRIgtFy5FJvfyPX/jo76yYkDaIDUp4p+zQNCTIi+OyqL4
F3Tc4E6haqusqI0D8XrNdUObusV6LaM9g3Y2IE5KMa3RI94EDOWZq7mJtWFwPd+K
buwubXCM5r3SJ8/we9clGPrMAWFB8i0e7yOnCckY5oGN1QSJcHlNPc4xtpen0XY6
9ZADMrtas3UTc4RUBqrlyoUq8pMqErExn1pRvy0DGB1DLx1FWj9q6U+su4Vc6xMi
9oDkE8I94qvHCLq5zWArsG8kuWAK4JUl8o/NyyLdc5j9pZowH80Ngcz17dzK0NV5
g9JNugzK/La0fNWAow5dlTf/xdfRy7i7U92nI5k/H3hSkfwfwxoGoIKreVZBLQPV
++2TgDrwpZEJ/FK7xlXCeID/XYjmd3pvPB+Jp9YJmlsDr5cnouAsyzEJOvkq3NxE
jWGEfCU3fxx6DRuSobh2NFm717UxQRV52M7EVHEA7zxVvqexftuiO2hq3cY0LUB7
Wo+79tp+USmC8OcF4TT+FFjPk8K7Dl5hqdXdcXx+oT4WEzHDS/39LmoTodlJ5dly
AT54eA6bqrC17yYHi67GluL6WSRGCJ9OkoVXHb2aRo3gtvj4uVMYzsa8ZM66ANV7
bt9iVPyRokhDwvhDB2X4xVuHRegqw9GlbIXSruY94DgGid1PQ1elsy2cWFUoXvsw
d5KQueY3fiC/6xpZLdqclHIT0HwvGOFLQKdmAzK3i2YzX7zlFI2kk6sXs9+aNLte
opPPNUPCEyLz9pdjGnS49tNN5S3XQW0KDv9X8cQybDmhsH7ygXJ0kaV3oc0pB3hn
5UPGm/K/iVQkjlGYDlQXran0EkQWii0qcyDmgDhSRNQLAl6nUS3hQtiqlwReXHt4
`protect END_PROTECTED
