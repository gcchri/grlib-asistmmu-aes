`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uP5v6U1H3UHTcipUfVECHCdKNaMKYbJXYOptBXewwkjCihejCFrkS9tEIKCbjwLq
aaGG6y1Cv/MHz0qwsvfL0x5c3Sbfpk+gAhaDh+Lx58Jz3/c2pV0e0p1Ijx5CXwIF
74w00/2N8ytbDFDXTaRplGgj4Z+VixvHGddVLVbEThqzAlCrCtkATA08MRXgrBFJ
4YohTrEzKZBWQdpOsi0Ht6SslqGBVEprv6+YJ0TtBPQtNh2COcOzJoJYGDw0xoiV
BkAPADauMp27V5sOgaFxexDCvU6hvFqNsrfIUI4kcEoCYMGt9atCXiPZtyWHyDef
jYFCMFl1WV2pR3BHValGWNZaO0YRLEdTxzLhcddr2eIB07XCEluTrS/WycL+uXOn
WROH8hVw8Q/ZkV131HDmnVn2tzD/Eu+EfrAvEiPF+4CrIagmpnGCkdM33kx8LRPh
BBNnkxq0WUWzy1X2+WQ9HrWFcXNXRVNvLIseam3vdNKMdHCksNEmz5RjdOuOI46W
tThNCHpIg6A3YHdVB0w56aj2aloR0VsvjDdltksCg+Z7Rl8fBQ9DNuX3s19SMuEa
U19AoPebp4AZBiw2Rfj4S0afLyP0r5GyPlQJT9pTNuxqFyMc74khqIa08/bR/jwo
PsoFlLH514IX1PO68F1oDdlrIUp+AemixQucaHpqW4dapiJJ7opnLSUqPWGLC31I
ZlC7hymn4vgC11gbB/fCUhuQPObDdRJiic+BsTBT2obZNMUNKl9eJPN5u9AgUCcP
GPPi2h+40Y0Xct25X5sjAEqIgjME+DaKYdj+3gyT5c92L4nRg+sOloTHHB6Uy+QX
cPBbwobC7+ITen9PucM3d/Qtwi0k0gRwBqPDrUDeDhJcYyZ7kZEDzWMHqlO5f69B
Xy9ekqKzjuuoe1mfGLjIrwn1W8U1JxzJWPulou6sfoMkp1n2EP9JNqgUSY/oJKxo
SyHswbeNx4McIaNAahSlqv5WjOkY7CQWtwxgizo67dobu6Rlde+848343LUK2dl1
Ukg+I080ERmToD0ejtP374gtrqTp9lcYLxddeW7dvj5t50ZoYZLV4/NTMxL42qGf
xQg7z/TFv4aCjlGNpOn+Bf2FtPceMl9/ULIE2cAD1OcTsJ+/Pq4Sw+FccTTgh8Yq
LZL1Odi38LGybsbzS0sqyvju6PIP1E793PilmOKJYaR6YkvLEy2AnOwlbsi1kRR2
Q21KYY9ZlRgG4u1oMsWmePH6imY7MoLw9rvJPmnvL2vrvvzfwhxyIDNnlX48eaqA
q1w+CvYxA1z/hBR9XWRkdOcBnDZYigQDt+8oizxRMhZvTvLkiH+w419BOgelQZnS
P58+k+KR0qfaKtmL8jRQ4RuiB73AAskjoIwh6D+GmWRaOLLlNMq3V15iCALXVZwI
vqhH5+oeGZy753wEL/Jys3Y3ume/8x/hvF+fFc4hs500lsixWlmKX5+YXa7GsLFm
p5yttE14dlAIMXsOYrdj1zIvcFAU5H3UDKPQmHNGsjoiwqTFGZftc8FteMKnhvDb
esJ/K03gmdMAfmgxaLRpftGouqhJZNob2eQW7Pm2IETegFVgyi74qkl9lVVIfhsD
JMZeBj2QENkdqXghm6xnN6r7xUVC6DDEfmXoJ40kVLY9FLvqRse4WLE7WbPNcqwQ
AFPmY9tJO/Jx8tsRvzYWCQKCyVOLSJlPajBN4sPzxxZpfU/hLwqH6O19kjud8dGd
6cgKK+wtwe3dG2tZosJqdiiz+/I+EydRwcAhsI3BjDDBJdjaAYJ4vHI24aPQTBK+
KsALq/C40o2iKTq/ciWeVNLfMbXankZtwKJuzmcI+GzGzQBWVAMSYZcnk0gmzih/
3HMAII9dKQt6jaogShjtEVHogVrOOIUiUODt9gblpUnxOWXZ5SsbfnDfqDVzTK00
AaScj4obMp8plrqAeg2a2xPcQYPhTK5vVl6EECLCwun6DfgkcRkLKrpXMXz5+AQY
tgtDWaS63Fh0qoHQLn8e1Bdi1x7cgGp+Nz8c0nKRD6OPExSvoUMs173sNhSjSCAp
GKDUPjW+CA7TtErR3sUTyjeUinIp4680kzRrZcmAlHwAP3evQb7hxZ7sOWXnLbmW
L/lcD8a8BXEqRpzg5ncKiBa3Gmv7K434iuMq11+KiZG//XsT6J4TfJR8kYnONQUo
lP7eWpAZOjvXOnRHNnkqeR2QmYzSjhmFuHFtJki8sPi7JhZcJBziaDHnyfK9iONY
J5IeudCkhj+Z5IhRWCD11wnhPLepC4WDI/zvqE5TT/YvMKXbwb6KpnWqRHwSRFaP
LVozdvWC8J4wks1Io3CUajDxbR6xYTIR19+GlOuF0skkcNA+GoGvyDwtgUvjoIri
KbBkE1d4OHMZFb5HGd3RaqamYWk/m37KL6yceinVMDNFK62+5A6BHlQiZBzM+cAD
+gOQYac868e5imlQ/JcW1sDkU2Tq9f/Ifd2F8LYK0Ob1oKH34U+m2Uk5+ASHSa3+
xJZzbBXTTH2cv8Np/XhAWqLP5HLXLuhwOhg0rXFS8MWKU+ISualmVKJ0l3+2ltg4
c5Dg8ma9om+U2FnxVequ4SKlS7JHtNSn60g/ky/qPOxDVNtWpcHkia3xT6JEpqln
jVzsw1nsQnBMBH8cBZaXx+aZNqntrR7h58v+PP5OtLjEewtFSwXdwxV8L3xOmpI+
P+T4ulBTysm3JDEZGZT2OpI12m9/d7wl7F4Bsh7wOcfkfZcZKJfLazZhSgeP3jSj
cUkJAevvN/RtnylbFa3gK1hQ3eNDeNiIjmBAPLSkKrMobUz4JStsp0dFuT8e79MA
s8LNNLicyu3mTex5G4G6KHU5riTHNhjv65JqmQ7ICHSYBu1Uzr0VfSdM+dzHC2vw
wBlxpPMh32tcGwIULjcaYFXRu7gF703XiKT30MSo3Leg8FHtxu0prNEIuqKsgVZS
WpTTFRgsDWkoDyoPQSQxrCjdzAhT7Oc6ZRHG5ex9b5ZQJHHBeXcWcKbHfDyyYenp
QyCXQol4R3G/M7atqF+kW2+0pwPqTotIk8dB5emgckCTRs7Im/pvkhLy+fk4qic5
yB6mbhW5yL7F7iBhYhDrjoaWdpvFCfSh9Y0HF30zrE4PnKPfwC3ey1Wogbk7kx3O
1ySxSNL515QkNfLPy4XMTAmeZutoDXKEcFbmHs2/daZ94MwNu0zGCNDOPVS96pqc
xGE/7pKrSnaoE5P4NTsIPWoF8wxZljSz36euVjfAjnxf8wJokNqD/PU4e0jGujPc
Ll6kKvuPbt1Y4Tvptiw4hQ==
`protect END_PROTECTED
