`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FUambXeAgzWAySmMyLSb+QmCqVihqKvVaL6hK5HWSO0nI9zm7mOs97j2Qsr1Ilx+
HmU+TOgDk44Pg3ar0NUX96mws3nFKo4Zm5myndlJdXxvZ1JN/6Re1SZH8YzDxz1T
r+Ww3XOjVXGiqu7K9tSld+dnxnMStWVn07MalahNFfEk7eCT8WmkbeTZ7jZkXmeQ
qPcckgxnXDmlZXmfnHp6BpXkVKKurRUWUA5sBSnXcthCZ8Iuxp+duZi58rKCOPtH
3I5vY3xMNAgRkHoXxz9L3ZH1vdq7d04C43iMqITuEUv3vzRNvDMnBHaC1TI5VWo7
fjuQ57wBKitKHzeo2dvi6NCr7no5Y95Gzlyw4iMru2vXb8iJDbBQZrmomBPzOtgt
oO3oGa9BY7c2exViGUy5D6itUP3ZcJyMZOfWZ37srAak0NVjg2tN42LAXT0fjb4R
GTq+MDoo1nwU3bUgSIItM9Ebq7Ygk586TitPJu5eVY/RTOyWHWPor5x6Wkwlw0lF
MgtH1VMTE4tu+Q6xZjKVeA==
`protect END_PROTECTED
