`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7m+jhcpL0osETvqAB9VXZZlyfac/K5BYz06ZEO/rY/3Uf11+ATC4/V5242I/OmY0
EGEabgg+4llxwTp7rUiPtoXM1fS55hOeVjsIgni2JawImTP4RZ6dOBb54JAshedj
7ifZqLnH8YuzQKZWedV0tSpxAws2dPqstdikkFuvsXc7sOTuRHBSVZvtUC7uO7b3
ZtOg9j67KAyXx4x37029iFBa2PxT5WuuPGnaU6YdpeRoEgjrl+IYRclCKqoTlx0w
/015KQ8aCSSY+f3+wvXuidXNjMUimVRTcsWsgL/yfXYgEoyJ78ZNoO8zmFsn3ka8
nFrlfs7hsTWczm1/ZPacFUblJfMb8Km+fjY3x8mV9IaZBhzHdfAUv2VE/AJMUgC+
wz0xuEgWnefWXJYYzpY41jVdwNdUrnLg/wfkB1kUgFkqOaVwjs2rnXgfx5cddEmT
nyhgiTJmZRRt9mFE095sGaF8DywatYZK1+VF28JyUD2aiNBVUB22MrVYu8v6otaq
SQ7nxbP8BQnz4GF7+90GimJRk4qc2bt3frCXkaPzYBu9VKGY63HyL14ArmvxUk6h
tKKdr5FcxNlxf2QMAFG87FGEYMBOVRzE0gFyGmeqpnMXNpKIcJXb9U+C7nCXNU4/
GZnaL2YMHT0c4mSkJR88MQCiwOp+9As+z4bnLpgP19UwprP+UfiASyywkgLf9oJ1
IxfLH3VHXbFVytKKBIHueALi2MFZkcxTKJOBKOESuHI=
`protect END_PROTECTED
