`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q/pJKCbOUw+xSis38yacoIxjVouBoOXW1cNyqwPo7eoainZvSC7c4AGxPbKLe+GR
hO9yVk5xt9x2X5b3rK/14zoUdoeZVMEfUH0xYIQiZFSXMha5+IQig/ue4PC4zhUR
ObQzede3vTbF2KZi6PxmorxfonqSelzi+peidW2Q08dx3y5vYWfgooJk6vD4bOsu
z/dRNebbeNHv4Ru3NanQzjbrUtjDlD/aumQ0ZqkNMAvNRd9NXAkMvUSP8KCFaZZk
E7JPhOQ3ywzxQ4GbJyiaAzduJWB9iNHQkIM2jMyF+Ec+FvRfPHZR3WdJlt/51FSX
sriemQGGauqnpfV5DbilOFNFZEvR22icguXhewnGSzUs7E5H11naE7zn8y/WvrSX
B5sBa77mDNI5lxDBG74h9xjM5IGt/yRVD8G5xOR5okc6C/UPBzEsi1CegZipvXzm
`protect END_PROTECTED
