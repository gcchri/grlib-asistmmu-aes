`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XHY71yZ8wdZ5wL/IZ9karySSUyKnXWoEAGAC1CJBOtEfW9G117AX0BuCzRvMWB5u
rKJodODZ9ITpJuk521FT72JUbwqRjjvVi5peLjQcr++Xa7YzeT2V3GwkBka41O5p
TSgLDnLzEswn6Z3JIgu3ob1mM/QCkFc8tNigv+3QNgD/f+QtvsA2YCFPnjS4se4S
tQ3QqWTm+HWYvLI0vBZEMpI23yWlFBw2QSR3KGc6NrdS5IA+VSDL/iB2ytKs2skX
iQpN/DYkO8sK+T3IW+E80525NLgaw4bUHlG0teYzlDUgEd1IQBUD2eXP+mTlwCou
5m62L+iPT3PiE2+ce9soSnlgRtuj05lbIkkCneWQfVM32/MigGHCBW7cZ4NSDw7S
PIpG+IsHO8jlbGhrk/RMWc/7rUkk9ax55MdsRDjYXOtBphNLKaZ4he0uGuhYYBXV
KEa9l3lfgAU5h+tJbkLEmr7YRjEFll/rnQnTPDrXZ4jwvJJZHo+GQb77BsJLWdsl
oHsDJpDP8AERrAXJYmm09KjYyELeU/LAFki/y4bsNfAE7suz5EY2LDddCICt9dS4
b0+2LklEqoBYnkKwZ7cgFzTCl6C2xW3nN468Ug2dYradOsL95bBvtx0GO82IkG0H
IB+duFbcAvkEjyTOG+X+SqxZG2HE9hgBTGWWGq9w6htA45CZHChXpJlshH9WqR73
pLxtDHD1kOYvvm9NFxJB9DmRQFFbSlwWqmeLchEM0N1HqJzq91AHl84TcHjiX4Ia
vpcM1uLLl+gy4PxFpw8/fbb/MnhhYRXZyZm0bO4jps/2AVK0HH27uoC1aOoQTttm
+9orI1oTAy+wIWCjvBBAE8hR1qcggtRc8ETf+6vDN8pxjj95+Z2l7qHtI4aJNKbY
aSW+aCo7rcVm7JI8DYiKXweR+ru1bZKekp6s2hZvLugeTrMBLhy7SuBGRwuyBJRP
5V3UXz1cyJJqwfSVRAG/AZ9bouBMMoWXYwRZ7K9yoh1ROCjQewOc7cbbOfkoBNsm
ufm+MFIe4avbyyMiunyKaKkFxTFOtxwB5hNXs+ziH9N523OJ3wOxzmgsrZUWF+pD
5NoeIpuo8gJvRu/JhKPKz+MtSSfw6uXAtjwHOWuC69Z5OWiRHc0wNRQdtas6xZzn
L0tYf0KSdy83KFUM6dVrYMiBKaEy4KiZmEyK+pBFKDAZ5LdsSuKxupax0mXIkzFH
vFDsOWO2ga1g7XoF3BmManCW721Y8sND4vUZzKM4FZZD/TEDX93oqIxCZJNljXjE
kqZGd7s1B0i30gPoulY5L6/tu0Pz8RAq9ERbK1ESI36cWsl70g7TSSfLJy2cf0zp
JS+5ft/Oo3xiflCk6HD+Wz3S0ZV8zwghkXO28JA/AQB0BC2JdVidTnFntaHNg78v
velwMF6ID4W8cbgSRDLOB0wQe0mS6DXAIhcZ3n86QDK6ZaYWSrJVp4Sg/y4bix+J
XS5iZbnEBPCcrGh4eKYfdKnlmsNcl78aM0Gc5Vt9N7+kZhaYlULwDKuuKWse4jD1
r4suXNgYoO/oLvSJL3k/0Z/q3pqNp/AtUeHpH4TWF7US2eZN5glqEn8gSwMV7i2k
WGN5U70vCRmD7Tae+sIbwRheP95JfynQX/x/ihATrPYW7cyt1RQWW8iPkLIE8XUD
9KQ0nOL4yXsnG9fl7NO2jKJDqCmd16sADc+yXY6+YNxY6IbBieBXNrent8ClBO2f
ugHleQTD9mJog9NgL5nfk8b3NCbMaEWxrPuKHK3VdwqzFNVh3oBDlUbcl1AwkMT2
TDAvx4UsGj68BIN/tSkdKREv8RGJV/u6XC/0uHwYaGEcEpHpYhGkgED0uxewZUX/
WB37O8q8Sp5feKehlG9MyOJfw6Aktte/SzSd3YwVoX13cgvOaKMX0eCsLC00alTc
yhCsGYi25YJ/b4jVUUG2edGBDE0LaYGNe5trL2e2pBya2eUke0vK0lpAp4Dy43Ar
MekHdKxldFNTyOH3aopuLLm9ZvWdoPSG1SlvdR6R3GP3UH4XVGOENIGjibZ66XZZ
JWl7nkYdGD1wdL79w//ve9Z9kajZOnUZjhkGxl1CgPZb3rILLXaoPHyaD2q8s6hv
Pspj/rkfiLLRjIFKiqF7kKFguSe5v/rw8Dq59It14oil5yFJXeK4QJUC5B038r87
z7l3shWKoaE+uaDuqH7G89cBe4GaFXRzUP3ivPFdmBu+7zG9xly/JWqUmDSyGGJf
4CONg8KNVrd+KdmxCiI8aq9Y1WPiyx+eK7ac+sGk6B03i78aQGjS2BYxAwDMfK3H
PLPSpL4kniGK7gEMKADGJ0sOq9Ng7cZ8J1UKp+MUh2IZ9u8yunZqAYySaYy2acio
ve427q6UgL0dZYMBf5Wwgu7PWEq9yVRUTBI7IUrCUN/tA1hxAHDAc2qubRl02GBt
FHMtDYkKALVl41l+kWuGBb2Bcv2MO2WF/oy0rQ04+GTFJxYmiOWWaHjEbG0v9zpx
RFXcgNpsxAxJopYQu87YFktk39bmCz1LYaP8VpBKSdlT2/qyQsRxeRJNzvlenH/a
SlzXOgAht0N71N3X+7HW4Lc1pzuJ1ehixl3R4mMmUMCQXHfbW1fKF7Hryrv/Af1U
287yWQjwgaIhsaYwjlUjjsBi6gLqAJR9V8jvbbHQRjOA0VhINLuvviGnm67GStco
C+njN5y5KxXQENS1Bm9xkKFeS8nxoc/oX3k0vnOLJZ3rBwjT049xsqAGAIA8cTlA
AGXRTriBx8M4IAgYIvjsGpUrrsUeElCh8vSEiUnRerOpPnXeJccYMGJiKPTkXGUa
urE1bQOqU2F+KEY4sfdlLOZ95N6xXHS/cw1jGObf/yZmgH+42faDV8k0uRDktqjU
W+YgViTaVMJQaQFKn6iKRQJg9vJjRdtHo3s3l0fGYaqKTGUOLBbfelqlP3twhbAa
WS+k6eRUovGRbacMEgxundB+epjOEb620FjmCcFIGXJX9Xl/i3q5g44tMznoJLrp
AMzs4O8BlN4+5QtUACJXRtFyJulgkeAIXLaaVwHMWkB/rsnHxyLl818X8U+XKL+d
8vEixr6dv8d8EJUUbW8EdnQVRFl2HtdcFq9cxsSj0rsEvRvFal+kOgYNwVjBlmyA
ViC351f5pLDaX7x6KIm19Yncl1hNGdvjdeS5A9MW2zDLwsuyhni7HHGcYBUXdS6e
vPkMBq+MW30rog074TlhkYK34cGU4/GdedC7C6DuIMN0VulmcYAV/yv/SBynMH7r
3R1Dm9WpeAmJvurU15P0cLzNSiBkdZWPY49n2/jGQkoy1hbctfEqNnvuwZT/kzFn
15oVclxUPBDaOZfo4+BKrArFzp73SofETCDBL8vSTWssTIrbu+I8LSIL0bIIwD1C
HKt5kZUvSFkLwyolftS7pD3uu4ScaavlBj00LhAwSG0c1RBKkooTUqHVphjhqXV8
bkkl4m7Jhei9sZaF/W1zsZlEZ+Af59wdKaHrFnMOhtOtW0a44JyeY7Iv1AV64fIl
k05WLFTPFhafQjOulQW8x/m5Vk2SL61BXFQPAiqR3B2aE99nakYHP6qcZqBQusVd
p8Big6T4mS76gFRrPpOEEor9bjtlBV33TGr5ac4C2WBaob2H0M8B+L+0CVwJG4jO
4ZvFMj3YtgXJz5EkKQKp9oQ9YJRZzG2MVF6rNjc+ymhcrWgct3A2D1Y+nppe7GS1
E5MQrE72wBORuV5hJb/p/4T+TafZMty4F6MGDgHnLCRh7se+esEq9MqrBjQlGTIa
MGbXuOksymYQG5EDzSGe28NHPA6in52WsondJENP9qb7klhxbetXPeUQC0ymYLgg
yBcK4dWXD0rd8wb0E/AUPClYLlFEM1fL/W6Pkq6jVWSVj3F6zWKpE5VXFzvoWN+s
RmVvDZGI8z2TcMooC+vp8wfIvUX2cwABMekr8osPqt1PRJQCy2l/PUE5/X8ALvpy
DAbKegG5Ib00/aDrKt2MI5TM3n9o3xoiLVMZIbHX3AaRSyxRbHb2xaosFALNzcbk
xTt1EmgaZ8/ZAHP4c+ji7odPkkZF/mqIvuJ9EtMK4P1cotL2Q+z8vQmQN5wKDJ1x
h9PxvhYtt2bbp/Roy3OxFgyoDNu3/d4HzEl1EsTfog/xmffvsBINV5NPSeoooXaw
YfEhEcpk0TU8VKzI8dNjmb8r+/0DxwPEEgNJ6fm1M6krN9APgk9AD6Ldqm7UxY+d
Pr8TynvqvkjA2nPH+fHr8KZSSLPfGkOvqD3QKjcxBzzZO1tWgMeKLJXCbr3IY/zE
OgnS801S1cS2NQn18Hh9nQjqwRWD1imCbgjax0b+GVptHdGJTP2+yrSr+gRNoYtd
hsEqy5kuBbrgh56RMiFZ3n7poVizEnqZ4Aj+RhyqTPTRnlbFvRKqQuUnjH05JsDT
+sIJbN9wocNkYYNxnPDfzEhLwrtaFOldXbqrPfJBo5ge569cppb+AP41kVTZLDqS
aL1WGM5JrluVk4tAfsV+3Q0uZa97fMaOGVDUW/CpttSns6xa7kLLnw2a2j0QGjic
PYbyvD9O+Uo3z1NIeUHDg+WUGhZItr4cZA2OdpJFkYhCGkePqu5GQk8eEBz8I6zj
xkjWxx1XBGb8UXZqq3dvMlet/1UzByIemlj/5afPGKk3vgne8NCGcCRNOd/UZosD
+LLgNgv8KdrMZGeUE8mGBiRDXTa19ZLKg/8pN6ydA+5uwS/QIvqyNjvDMOauvI63
dzuv5D6ontn2Ynks/DAOY6cZJ5uoGutwtwlk4912GUPY6Ct81D7i6p3rGVwY92yA
yZ+0k4wEX1Vj+BOYol63ZWQZTpTWbcVV8hta/3FT3lqAsfn2V/cktwPGMUAfj6Ov
4TTlwZDaaXWJV2IC92mgSBLVHhKhTvUZhyqS1sSBfuXYNPJmVx50N/zIrqKvDhEN
qo3fsJBUSSU12bW0qG64bbaQv/DX+fLFmMdMPuZfCQu7yc2F2qSJzSY3dEDLUTCk
wc8P0mtnXTatS8sHpQllxSUj+hTTe3cGsoyoIJ8apAjFNFa38q2agHXgmDie2qFR
Ipv65KnI6hHnSgDZ4304YBPfrywn37b66t2D7q22TuXeQ+W7bw+BA1w9qyZHyrFj
`protect END_PROTECTED
