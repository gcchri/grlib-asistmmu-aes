`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ctnt5luu90K26OmdKXyXQIZBaDCCHFhI2ethsyUH+Qr9UFQWUx7NeO8hZq7XQkRq
bE5OqQKziJPYOt8aLpdtt+2bkVB2VfcV6EoZSYGyZELjxpsrAo808UiJklEE0yvR
8lkfdmUUCjFFZyZ3l/TyJKf1PFCuUM4jo4MRhPYd1y9wbz2lAMjvZJmf8KvFqpIx
+Bhu9oIdBIoDNcsLdFoTOMDnULfMJXEolhVnsUx5DslZJqaANXG4kH8YUf+Og1fq
57Ad4g0+EYFX/4qwQuZ65j01TjcLvvdcc8qaIHiPUGyt/Oo/In+gtJ9Xm2/Vn0vn
45o9ZTw79MzyEfDx7dlQ91lY8TSuui/gsea4HLX6o/SKSVfNZ+59qrKmD2p0Cbxu
aMbBQOy83HObM7YmMuAnN5IoZE++KLeCvxtNB/osOd93UK0vJKq0eOzYUCdVw4My
k3p+UC/lRkJ7AEK8yKWOsd4aI+1AVreKDrz/4izh0Eu0eMKpq707Bv0rBd6vFSeo
a60evvlb7r+Yz52PQKLFTGSBmy+sXoJ36u1NKs6aSdUOhL+G0zkxVfXvCAt7LA6Y
xpDOYO6ZgfaYYAAt8eIfZ1BmyqZ8mwm2+/ildfwnPhs=
`protect END_PROTECTED
