`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6+6xQ465blS72oog0VyAaDE+d/iytcy+Ae1szII5dTEpZUxr632f/bXoliMFweyP
d2S4BjF76mW5TQfcdDqJC6wfn0pKQHQTv0O+nswRHb14Voy4hWe2yPyDyWx6hclK
K/Y6RUqhmVXgKTaL3b+fr3n/zqojvUJyZWBxaY0MYQ/QrAQEZU/jVqX/25LyxDGC
luYG9sNH5bMgM97P2ZoZGaCbC+kjRcSMbBz/uJXvJPiNVQ8oHAbcKN3BOsVSJV/1
ZYkkOeNOd/XpjcTrLzhZsUk2lnOIA3r1Fxq+6CXaAa70qzTgTwIb068saJvmEtDn
jvbVu69N9nUGRD8yMV5XWqS1uWiDUofHZ9WelXgUND+rLHXQSgXCPE9VkauPXkGd
nI7RySfbn8AWSxQawkQdOBKOe5VdVVKrwmCCprBksMt1S90fznDOFzktGhfX+gPA
7pEFGj+8lMkm4Z2RTOTAXqE9i6RaDlPiTXzxz1rmYexjVTQQSdDwp4UC6ELvYLPE
cZkER3/6vZVAtH1uovuI3T+6n990xdsWf20sqOy8iHXMrLvcFO8osQBdKCk3Zt3p
aftoyPOnoFTnW20KMIUUmpaPkzC4E16OsY05WAqGyY8q0ifdpNahQ5G/RboJG/Lt
gHW7E3Rl1D/f8L0eUjXERmVoMitVYnOUZU+5tga0CGOCTzz38hr139IN63H++VeW
Yx4ipC1M2qCPaN4gSc2V6GSryf0UX/vTKDi/+uABl6Fd58+UX3NTavkJ7WEfe0CS
7UMt6QiaUZWZmAj/CvXmXtMbyMb2HJYHBnw0JyfuAJF24lGDC+osnV1yUrIbStS7
ya0+SM677NIumMeqItZpUCY0rkRfAzfDyWL90VBQl5z06uSftooGfKk/qO8YIhB+
x6bXT9Ftd6CiKwuQ+/FNCaBPEjDNLlACfvQbIaY9wT82nB6BEmD5Qh0s7wx6Uxy5
KO6vMq6P0fI6u/YXpXyLQQ6NBPA8Mvk8liQVVL1uUMN8hekeEYT6tzj1103JHdHF
yqd+ABDRYLyolXZO+OPyA5NkZwz9QveB2ZP7ShPHBTo=
`protect END_PROTECTED
