`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PdPPSsuKGZoNiWcYP+GxU4VE+wXUsdJXsxwAsnnYoPOSBmvD3WC++ONmHJzM8wb6
L7s94LkPiavFk6Gok1q3JzPPhXw/VGZ0XQ+KcLtfiReJqx8GPskHFIU74XTeMYGA
lHNn/sbjcBjg997VH6pl+JkO9YT3rues7HsDLJbKz0g8VDd/fFVYY11axJ/87HH5
mhCN9mCD/WqTxJGqVAhpSshe9Est30POlgvzBOcCVIHVa1OEmR9gqR0Lr+jsShvn
QFr04EoMjmWaTD8rmPvwwoJv29UU38TObZv1xla4wvs7yLTf9jF6x/MfUIDBhmG6
69MPrLeJ/iV2iBizX6utCbgJB9ajyM1c4W0fMXOpCqizaY+dpZbHmlMQ20Zpm6FV
MhD5R/p71cTohkEVa+hRKXFYDIoDQc54vTl1zyc0emJHVXqGaTwLlC1JmNEQuciQ
4ZJ+wfh+a9Ces2/nyx5/Gx7BhDjVR55fHFe0Co204Umt0P99SmCk86ZBfqhBN2Wo
`protect END_PROTECTED
