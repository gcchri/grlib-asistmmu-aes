`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AXAaejSDK745sz2A2mJua3P7WiPTxTWSOUpYH+I0juPAdkqJfgNQg3omXZ2Rg3bD
F/4VdPNXSq6hr23d+lSM9w0erki5mQ0yBKi2VrvBkjYzA4T1dVGV53njdJLi+/48
lrdd6LqP4vZiermH0BbNgilyUrmyhss/6etkRE0Hs4NjPOLyV3vYe6/v3+ccMZwX
hnfbfq3BfsMAdA66aab0yxMbfGmJJXiG1u/OaQlXMGL7TlmwtNE0NcaznQEq+v1D
Z0a3KTrLLIXv4xHMSK/Gkhx+5/Oz2mH6Jl7EUSy4LNCzIavoUFvgnqljkfdzZNRG
+b/uWUvmbnavZzD+AXIgdKHCk/Jstf2UEI08LL/KXWoN5Zjg581vTjC9GxX8ARy4
iDk2a4sabGqIq5+P2aUHtCxG8/uD1Ig5Mn6X3eE4Nq4=
`protect END_PROTECTED
