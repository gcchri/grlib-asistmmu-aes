`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gs6ivLuBl52/u8EdvLaeEqDd7ehOCfucj1JbNRMvqCHGw3aJrwDml/tkvbjEDxeH
5U7M+54PFTGuINbQ6FskrNpiS/n/YVqhgN2vxbiqy2naTD2kINlVoBC1mnRKr9L9
QGB2mFDdnqTjdzn1azWgAYVujqPsLuIud7tJIVtv+HA62qAlkyWDwuy3yXtGU0+h
dGTLc0AEDkMjfJF1OCzhcn+wIVtIRV4aBCtz1skYrsee6fSg8T2EqxDDvuzvawWA
sJl+cXyntafjRv49I8HoaX+XSBLvUTZqEwoLvpmOIGVphQYFppZGRt8ZmmjmUHfc
TC4ipz7VZE5HKYzbTz3tlEYmo7E55U0JwkvfzMANL1T4U6ztzh+voRTiU/Kwjv9y
kRUdx1e0qLuKPRvkjyrFQgJkW2wzFdUt3tg3MZTgDEAa5TqfDOyrkH3vzh7t5GgY
psf77pnDHsEOfMDb8jKj3VVhRnshEd57oZ85LWKCHx5fkZrDht9j3CG9YHWddSzL
xaUtXcUKpCpD9o+6kxxY1ghfsoflBv3MZ7xXUKFtZ6pkozwOclh2ME41by8+stJH
`protect END_PROTECTED
