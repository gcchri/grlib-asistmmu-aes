`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VUJTbqE5vF1r5IkCfwGnkizMykeODmhIIPDroiv0z5WZDWqmxJJrd+kDpKtdta61
yBsZwXWZaqQtXKHZiMWL3LZND0Jadnq54jKB1Zr32fW8Q84ABPvJsYr1kmtgj3er
1LplQHTP3uMU8HwtMD2MLBG7bbxWLISZl/GV0HlDkAg0krK0vw4BfcLINM8hXwAe
tJkq25rE3xPwsq/2ePJTkvfXTzOZPqYRBy/TaC4A/t8nqk1nL0knkOOZc601mF1d
Xky6FEH55mMD5Oo1OJncCrWKOT+cLcl9bAMB79UJ8qlq4yBqVSJgrMxz3PB7hctG
zD2oWhqnp+b56TOF8ti5c0mz0uG2oqTpZbu0fb6kz9QhgSsv/SB/Krf/9LpRqrXN
0DIyvQmv6PNK7vBrK2VPamjuYTY+HI9/qmxpgiwiixSah31zkRiWkAKlXYM2yh5L
`protect END_PROTECTED
