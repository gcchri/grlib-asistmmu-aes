`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u738/h4uL/AA7ePHYJoNJYB6V6bHZPHTIlg2uHIcbIJOQp6KKak47PR58boIY3sh
HMeRUki5doT3uwBDi0shYes2POX+2LQwgQ5jElBu3QFifjagQW2/X2Cg6PBouOAA
QWYCFV3k7aRrkwEivYxFZviDC0Irx/95//90XNdl5q1Alb50wylbjhxoST6E3QbY
k7zTP4Zukj4rwOkwjRSYbztXT2o2KeGOmACHt8HdskXhrgdgENha6v73xlUaJ5TY
6yJ5/4z/iLtEPQHZcxW1j/a0DRsI4TPqeQR/C/LJWeq5+Gw+44uSIAslsOHU/rU+
`protect END_PROTECTED
