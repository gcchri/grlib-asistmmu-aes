`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QqxlpCrLou6Uh2XRhcEqEMDmc3MCrdsV/7b47mtS27fRAgUf6TpDg4//to5LREPS
gdV0Qda//TY+XPiDXiEBYPH9tSFWxFsfuGjZrEBMPWJBOX2Q2I7D2XXzvfrXvcAU
YLzZOYCK2jzhHU2ARU6a4VazFroSrdpB4tGdBXCp1sGi/qr6dqLa954TGpjYdpnZ
AsTiKEK+pAfj5pjJ1gs1K1mDdR2qcirVbSUhhrQyAcy8GyI1ZwVjb5nQyUvhDhfL
ck1AxLyvt0OhzTkEwBL2Jl8moO8ctvB0TgsrSaL/vTnIGK7qIewUrPqMZP07QcL9
8Q8J2jk6PPB1WcNITVXQjPzSNsBcSOOgDdXKkeYX5MhPbwQfYy+fFmEjDM95KWAa
TI07DJcmkGivRoCpg5oc9a4XnfpwJDZxaz0mEqEGQ4Y5S8dfUWL6gjNK5vWJHBKo
dEunjnaLTLVuF18Nqb7DECc+l9F6hY6vMQKiYsAN1XNTcR3kzuVaIaCZZktDN4vD
`protect END_PROTECTED
