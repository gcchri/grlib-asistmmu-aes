`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hN3z0KiEbznNIbsqG15pnkOz9b4kzjNGgYU+/QbvGNcD50H+XJOLSYKOOXd/qJw5
N/Toy/nBF8EuOLTbtLYhFmpR380dqCIBG4wwY3Cm0MTzjSOSi39zhJc02jeDpt4E
vi24kRHN+93lz4a1aqwVzdDQQ9wSVRJ3ZOUyF+dsdWpKhE2yBPnZgp/HGar5oQHl
YGwSXhdoYS7FdYSUnqKwSnn+0TxeqP7rvgDAYs+RnJ8p0LWIleIS7LpoDdc4YgRK
PXTMdv5oULg7lSn5Dzg/2UFIRm2BvGK6TG8WjF0eB2ngG+OPL36t/8JfAO3vrrnp
DJW4pc5IXkGiMpRSX8q6x/NQAq9BRp47UA3Kj+O6DUfhJq8pSUrc7B4Z6C2jibVq
L0LlEMgmaEcykIV5xgpcJVh3wjZLhdEsCyj8h0mMMz8sviHbNpzxK0/EN4Va9ozm
V+qf3GUI3w2fBFRc2PnPrBevmwxYbr5d9CAL4zUK6Qwsu/L2eU0qCbfGs84PTZN4
Ckrw6I8tXzU5cMXOSk8ZPBv2u1zmbWO4wAuJgnVj5Fv1J9l08CqypFLVUrAXZus+
HzNXYhwwMaxzdN2mxRbhjg==
`protect END_PROTECTED
