`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T/jiWt8CLGvRhAteuIrMx9TNWTcqL9AhSonykHcxCiZuqDmlUZ18JkDe/iqzMFkb
ih0Logo53TyLZktQ8vNuKAz0dsoTwLYR151mDgl5h8ESa9ymDejjVm54OL22janR
TuboSdxgLf/fhcmxioQ34F0otAD0POL5zwiMcGzg2YjhaJU2nHYPE8sgXmLmat6X
KA4Xyd1jR6yI4rE3rVdV6hS4nx0uW3ErL2q92dzgyDtOqOT3hCLRHYRzAKibsGO/
XUE1BHHXW+AaSz5BarEUKpooQk1GTE7lSGDTRCVjxcFNmf78Dn4xX0IKyYCSJtLF
D7ACu2rBCzsdVcUHh3Odc1Ppl2vSmCRIe7NCihtVSd0WYOqOTWyvSiXBGhLtgdoI
akOY1qSCjJymp2nIaUS76LKb2m+tQ9c8+w+ReDUL4KR8krYBSKD/iJzM9EH/p9Kd
eJVlPTHbIvYb/xD0VFc9TokggvoD9oM9GL47a90TP5qTLc4ei8otQmhGtRN+d+SY
Feg/ZUqdAPbYtDIZYVJcSdKtWQj8shH+ydwhnBX2CmySLW9VlF8sAdocXMvPbh2V
PPjk86Xpne7991PL7RoZQztyey++/dIFsEC4QkLTjc6wT0U+OyIETGMw8cA9aBB6
/gdqpI9njqiSYHKKYJN76+w3aekfevxgdRV8KmgeVpPzwIQsE8R138FLBTsPEyDP
mXV2DNyx7L3oe5XO/pcuqJJP6P0zLSg/7DaHSgQCXDgnz/OzG2ulZgNv8jHejelP
cynursPlUv2KjcGetZXz8WsqavGNJI8QIePDlnw4yz/I/Bvj+GmymTGtYUGLTGZP
pmtzXefDGLaRX2Sy38TjoNiWdXI1l+YYLz+vgWnZYksS7IDhEsiBmpjUefGLOo3K
c/NgVEDBssiAVPcy3DE8ITRA8pxU4NVWchCcJS+3Ki0=
`protect END_PROTECTED
