`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rzcPJSr22hGUQHgCQXOh+jgSV4XCcuXK/Z8Pp5j5n+eK05B0HUY1Zzb6oM5YciJg
JQavdkpwMELa4fLjiIzMdviC9QJ34ZHDXwwfM3F3U3GQdNVN+TdNeuVWPr1lOveE
ju0fcfJAjyWlqQpTUeBSvARerl08Q6a1l4ZaOvZPG4rpRUDFFCCWbpfsc8ujppSU
Bx8jyhCLxoVtW2ER+rMGgDiuqVKXLocSVKG/6j24525YypEGH3gMhgKyJJXYTLsh
SZ/u0GWDq1wmMh333IbG/7MjuCwbXM3hZ7vC1x/u+fDYqNXHkYeSHlsus7+TwvoN
3AGlc+Nwm1etgSFtwXsEZ4k2pEaq8fiZru7vPiDNSPWkUiQcwHvQOoPDm4NxWN9D
2GmTLEdk3uy7HVKX50llGdUlcfsIAUzEHMdWnd4NnsNFQrNEXcngITiNf1YbFDSZ
qdQwhfYcvwLZ4t5tLXzwTU0+hC3B2/OuQ7vLAew8D2STOMlw6ShBHjdCuuEgwNxK
1uA/GhBzzoMSdacwV1Z+iHE7OYQFOCncXpx0fj6VDvVGAvz+PjcOLQ6X0iJoiSUw
IEkZVYIJdD/b/hO+I+7wqlBy+U3nvtpV2y3kcNUrjlphG47mKJSCAGMe01mSuIqb
ghcfz7mJ1P++U9LfBBDb3A==
`protect END_PROTECTED
