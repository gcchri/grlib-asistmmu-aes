`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zjWujBiiaRuq0VrDYdxNriJS5sIEoNKhT5IGeMX2lbc8xtSJinsnaTHRZkyivXeB
6v8TgYd5d1a7bUlJAWP9qN99SSupW0cEr24S1RQmjXlprkZhTnVQ286v3dcSSQLZ
ENg/BAXJRy1kp2q2OgI9E4g+ZlrHCeGx4fF5OWJ4VGvILsWTSipFoDheO+lCYQFA
RhRX7KYcfK1d+TOxyFrvIFFOC4Mp1uh4QkrzUTiqCRVAwjX/tiu5GAueF8Nuumnu
JDctqq6S4upx8ycAIOEg6Gnl+hcSDpuPxLz2mHdweIWmqguK1ftbgOI0qIcgweUg
kWxG5TsYxK6FsFiUF1WZYbB8qwceu2L16D/sFpSgYpiVeNAbbEHHprU/GJsWByVh
f28UDmCxzVCjl0ZGBlaXWp2BZAdlQkbFIrPs1RjYDlfOBk5xupNGyAuj2cwzoPyv
`protect END_PROTECTED
