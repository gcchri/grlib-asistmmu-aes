`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HZ7MgyGxZwOdRkHmMUqwc7Q9WBnoBcZnyKBN9sse2xnoaVV/UXfhXo6hmsWTJRMr
atvRDeyjbAFbQ1CPaVs9johRG5boFVnh1O6BgEgJ79OE89EV3t1rJaTWRuFJnQNs
Tl2HTNxhYDkNnbKVyZ6BijRmsi+FGLYRjrS8EDtU22r+3T6Mpvskl7qbXha2zZRR
ddHTcHQQrxL3g1k9Nov8c+mmjlVuKSFSCNeBQm2K4Pjul+xIx3wsxtdtAsCDhuXO
V1yvhqauNeDPSXdwUdxSqUrsyakweaEyQj4SvXcbS+c/53pmGonhVH3VCmRU9Dtj
UU96mbjod0ct1lTnRm6Pj9yYwxJzVtPxiSbwcLiEnPScbKCIIpEQc0unyZ6tY1CJ
HhuvexuytrzMWjQE3sSDkg==
`protect END_PROTECTED
