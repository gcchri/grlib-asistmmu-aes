`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
26eMF2mXZHi/z5SWPym/+/H5TsG+mvwzB/yaXJ3WqJxgprbFmM/Lkpz28xzbZHJM
Em/2ne9A4+3lh1BQrdxYJT2PamRPcjLnITQ1ivv97z9JuK4dUg5SdTHPCA688R39
WkRQAG3Z+r/hFAwRC9jn+Pi8Fkeb8m9fk9/+qifP5SkgFrA/mhuRhOxVXDFYjW5v
sCe5ljGd3huk+pqzbCI2C+nmPpfXBmnIaITLBGaRPacvcEYD4iJgpko9MnvO+VOC
iNvLbtbDo6EFOjNxh20bYFo6Zd6wW+xtDUsqAnT0fyGe5mpJOd8lu2LmjZqMoPfd
ZEeVUi16npHz4+oNmWWWFs0iblqYKCsg3Wtu37deZOfgqBb0iAm7S5sHvQEONE9o
e8MDcJSCtjUBa4QbeEQp0SSnmsSzzMBlDNrQJV/x6WpjeRh16mh2JsFDhaKcYA7O
y9rw4yxxqM1/fAj2FBka1behEHpT7k+XKtDWDwh0mMcdg0M8fY1J+xPyxVh4D+1D
`protect END_PROTECTED
