`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
87Ci4687EsM8RAmnxqz6RzOx0LiLewWAG+vZxGUZ5v8O9sFG2SNhQLmH6tE9k+yE
Ma6xlIuGmaqArQD7NAbeibNuWbJLl/3vWJJGiDaSFP41ATjdNROeMozwthQ2DuQn
4cqszger2RH+9A/qDFP1dM/9BaMhKzUhNmB1y5ti5I/VIUF/O/dckbKoHU+CDNTK
rvJ/KY+ZD+3tcmxSJBFU3V3MRmhOMORXt8/Ohg2tv+mHl4EvCTGbGgUSOr+JDMZe
rYP7P9NkxFqTNbUJWZctdaTuL5gLOowa/10bFPzGOcgX9xzWUJdflL+YXLVW77ay
6SEGBb3XXDsNdmVr6/FVEbR06jnJ5a28mkpO9nUQrzaiN3OKFTi8ViOGn4pe1aHR
sKeKmaVCBUOI8LrGVx9luSF4UU5bhpeHG7MZO1Tu+jg8/IknjI46pl8A0DG4JtJG
SThHuGgiepf1o9FMeaIbR2StgxKcZcy2kB2nY3odjVxJmFg+P9qwKpNTYpZeRXXh
`protect END_PROTECTED
