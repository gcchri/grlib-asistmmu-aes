`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zcx4AhmEfo+ZnnLpAy0zlcXP4h/C1Otu1p4dmT4VMb6xx2zt5kB0ZmhUwYcsMaca
O20+6PHDkPG7lkX3GD591L6heZgXFibBtNKbIVp+VoZgAi20lb0jKKsTLeKn83Jm
EDI2UQtO9Z0pOoi1b41LY/jVQ31FJZ1KPQnmMUFYY9c6qUiYYVHWKLiOtq3Bm/os
RYwCklL4645APET0DqdxVyY0jBhhHWmdtXmo6gIZPzchDssLXtWORyXUMkMQzEqf
rSgxT+k30irywvouDY6Sqx4yBSIAzk7wSkV4WPt0zUkqYB6vLSol0N4qrnDe3aXI
ZTKSVPSLmILseWypnTQLauPth8C7xUd/m164YOQxC/uUvY3jjDDPtPJN9zsxMzIG
+oCC7D3VcuLIi86O83QE/C1l0L/NsQCHPpAhPJn0DUqHDLTEpfKbE5Btq7da47L0
hQzCQ3xKnrPbr2OyPCC50NJFayZi8NqoHUTueM5RcOYWsXe5gp7mOzF71Mh6sfm8
C1NNZ4BBgyZCEFUo5upfZu/Qz++y44OURijeTOamuM50VxlD6J8HMCWTOL7q4x4c
3SEIyKqAV7UxcK1NlYE7cGz2fNgAClDCdng30cMDQRh1KIqiFblPhEjoPdwQfAz2
45gR4VFuhh5+ATjsdPsEdM7YodY5GUuTWa6I8dF2qLU=
`protect END_PROTECTED
