`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vxuWsm9oTOrC6m64i37x1l9+wV9X1PZ9TrbRwk+69RPVaOUwNOxi60Oy/VvRGeMm
m7VNhZ9F53sgabHpNayFgyWlMTMvd6D3onXBzzoxny8PmGTh1F1wa/n7eidG01bI
08QfkhSR3t4kdzcenTkht6YTlAK0R15MQ4tXIj1hbA0ea+tca1M1WQdELBC+9J3x
2iHDC6yutCbOVGg62wwdc01JKge7RGwzGEiHBlLOkueiG28xJm2wIO0J7dAR82J7
OG/mFyNa3StBC/y7gvLvHvjVc33ETfstn26Ol+CvTbmeem7UjZzxGKOzlOgverVh
TQ34ptsr1hGSjZgXR/1jAx+N2bbLnAXujFFlyRWtWaC0MST73mK7ZSKgNhz3eqfi
MUZPnG2g67khGNjtoCtbK+7Ctl0Tt1Ck0d/xWJENaU+IydOcbsbE4i6lq5vEyEiQ
nWXsfRhmy3V35TzSCXT51Nn91uEf0RIXyR15i7760fUGoU3W+YXhMJj3S8e9jyUa
9mISf9GTvDWSPJofeQ13qGk5No2txCaDqfZmdaqbFEOTGicBCAqk+fQMyA/xq+S5
m7NoIGLtMfa0GtzktNU1rSf7d8V8jKpBZhbngPJfbRqDSHF/ljCHkenZF4WGstHC
jpsrtuyk0kSpsRqXVcSAqG/Lz7LSGYKgRmjcm/PvlpIFnKMCGrXR4ERyis0zUlVn
SwFdfiGjR2cevzDqW+jKAnltzZDJ8jA15CVC75ie00RmFvV5+bu9MS0ISDWFM1ny
+loLh9Ub6LwCspXApB7daFxw0QFiUGexwjZtiDxEX4Mwy+OhMUu7C//APbdA+ZQO
yK1yycSf2Z59fetWIWmSuDKJ8dZ3fWwNcGIdsVlO7VpnpnS5V53VuEi+FslSI2Ri
nsHZ0IiHJd1X/kHEAHuwTp85GPSmXqWpcjZACJ3AscCX5TEz6NZPamVbdPDRkrgo
IdRytU0tVpqDwfEpcoIggK+LK56eC7c576SAw8KNJvdVLLAbwNfTd+pdYdyg9Ln4
7NQW4syaeeb85iueXpJ0A6uL2Nk3uUOAmA9xz/50A/U8fILgKYyoB9VdTa84frLQ
CtNClExNpSXAsNmpgvxeGFLNpspLJyCjhTAoAzASxQl/Jm7xg56RwimcGASn7t1O
W2oLp0bRWMMB3ckPogFo3J0Mn8UCV7jf7EbWy1QT72obGw/5vlnzVCTFhi2LGFSi
EUOF1F6F7FVpz1yp2uH1SWqAnDX4DGi/5Le3HNFJOJtDtGZp13YLIIH5WlDPjiny
dJ66ndS7mxLMcpkt7AxX0HBspNe6coN2QoBzd+eco729pvyfCDa53bQeiQRMAC+h
1WhYLBwk7TBfICbyLYmoMCE/6XVrt667A0GZrcSoeXGgbxsg/RkhkOd4ajNapf6J
+AbFvksautLMgeBdR5Wu/XKEvG25Yt6s5QyX1ZJ2C5vWiCI90OzasVwyaXmQOPgQ
/irWgzQYaASIQWq+Co1+/01lbz96mSRFnJrNnUnETbbMzFKI1Dkxxn+hEiPAp1Yp
mHjdNopjhdk90oHOgHK/Amhf0Hps0uKfJgWcBYth4FOxT+kp3MiIrzryWoWDb3hj
0Noxbfg414xyG3ZeQ4EtcBD8hedBj5lt48LgkyRz2PVzd970XLuCICQXyVvBcs7r
gVCMsxgtpSlMnsCaHxlHMbYZYYk/LDhmQI3TyjBPx7Tewhm1v5bMbWNsXKijwnZb
WdD3guoCvA0HzDiCweQFyof/d47/zwqodhgairPYxTS5afMBxJUclmVyV3Vet9nT
MsxBzl5o22f2V2uMO+ZF52RcI8ILkOIpkuSwWlI7x5YUxWNSMhBuOnZ5DVOlhhBC
WgGleS3P5KzHHXaO/VXDM/2arBaVvaFgx2rIGVgqPaEL+9vJKVilhBQr/ljF9N2I
mXwwQL+0ZyksuoXb+TzXQMT3Q6KGjmY48n4xFRKKwSIWZnAh3f/fTqPY88hWCj8n
fwowzHdtLWUIGr6l+4GMEok+Db+HhTluJB3AMvFA4WCS1+QsR/gtmGENd7lR7EIH
q+QN9g5trv1j1X/JmyIF8vIRlDJ21Yz5gCP0SERwt/ARS3Au30y1INk4aGGDtETx
xzI4WBK/LJ6ZK6Im8bFE+zZIvxLYO5Ybtg3AT9KaRHMUvzdRANmoGmj9a0fM5Hr8
NBNpAOqPY/slUfSQMm443/ODsy4kmwehnG11kNHq+3gnpY1b/Ip7Dy29I3KMv5Ep
zAjlWsy2xFzMPaK6X5FAc2eZRIw3BoyH+laKZcbNeaPh0Eyw1y9u6P7jaNk79o7v
9POKtxN1jM9dDLrQGXr2ukVPr3gvKWUL6JtFrYwohxHaTsgcKWNv7k1fD1BdhIJ1
eFTKoPgNXVulegrqwMdWEXV1jXJYHa+E1OYIbBbVmzebhrYQ99v93KQZjvBuyRUg
VwXthTZw+SQ/neOT07lCHZ1tqm5NbYf/0ipOjTPeNpBwyVBbv7eqv1jP1iA/TA0E
yUqV2DOTKB5HbLm6ZPFKY/QbMsuYEUx0G9B6xnbabLfNo/LlDpjzhFSL9ujXRTZT
DHH/YoKM75UXysgGSUWhbWCK4CChyDjisrjNRYG++FI3OnOXlv9YNMUHMu10R8T8
46CSompvJ7airHHRcBsJqUJERZ9LUSHQuXIKSpr2PntqPoth2iRL2PwatDJvLveU
OybdBJlf6AyIWsbgXdAtYa27AeM8W0jU0MAIP67eREnL/Xi3dCnI+ffDNuWRNNc7
LTBds0hcTnwagOrKcNjd5aXlhB7lD13HJk/Ai6h3jWoo8XOB1TTluyyddqgjGITk
AaRbyX34N7ScBpP2pm1hr6vX8qCnbSTpr/n5WdZLOystWYP7xYbeqALpLmUYp2W4
NvY9VVDYXTrmlOJKe2geQKzHV7Cv5d+YJvyyEdkXT00GF2KiXElfoFqc6cJnh26a
srqlRRz2me2LWB9VE5XgFJLwHvR6VRMTRjZdE5OzZ331GdXoT5jcC4lVEsAROGJs
/K3C489N3tZCBp1j9Pb0FZTYLF2R1I9BRGEkTvW8wDk5D+ACIQ3IjCWpXw29D88w
2U6mEtR8/jMFOzEM8gOJWSsAjKk9iidLhZ4vjR8PdxYVVB4mT5gNVRMZo99mZ1rD
dixMFrzBYIAHRFB5S+wj/WlabNaVLj5/IczNdwvAIMlt0mkO8x5U5plWJqZ2q61b
4UanCLCWpJm3ttKFmZMQUidZaBSth9xJy1nYp9TYH7QaysdppesoQ4ikGkCVqAva
j6qEJe9ouQU03pSv+2jnCOGm2zXg6IJjfGcwG9O3J3oNip73EuBvfYnBe+ECGgWH
AJo7WJ4olHvJ9H2t/ZFUo/haV1citB1PS0/1ERwZRJqEN9Frv8RMcv33wQYDlQLn
JQ+Avj0D8QGWKumLSwzF30ymiXFHAyYlMK11he1eMbXPyzBLZLWAaP2rl9YcaCV3
67+sbIKszvT1M76j5Fh9YY3/vSPsX7bFJoqniQPqSsCcmV0hBBOTho7B8Os2A6m6
Tg6J9p7euEemqQJklcfvsX1nMF+Uph7BpigV4qIQM9UbTPE81ZEQmTb7ajQvP23k
HDad24JmtIUzPmFbDAnyqa/T8QX1auzJT2w6zmS5mTgkBgva8TFFR2AMYhIWl5He
Y7MUdBYSHIQnIBXsVUtsktzTgcqr2sc7X3qVz6Fhnu168VmdbVxODC+a6k7ohNs0
qgEjr8eJnRBGMV7ZdCPHUegSmAzHx9TWgfNqkNJG9Q4qRrmZqc+3zOMgG0Yz20Rg
0qDopOa16431KfNevgCSR63oH1U/6TbZesLi2R5uMCLT55mAewExZSXEr4wHHyC9
TcRbNxsAKQ4q4dGWrIr6jjm/9zfzrdcFa6ifeCxaJQCUhVfWJgzJ3eksTTPf1uLD
h/8VahOXw/iSQ3kzn9XhIPGA6HG2KuoR5SqwIVILRmvaAI9scn2sdZ7VJ2UJ9GEC
bVHpnTD3CspEv+gs+4t4yT/CzveXPF273h2S62VK5qxbTjx2p86VIFfgPzoAld+n
DxRIBIc3uOdcXn3siyjWg3uirKj2lYPkOTm3L+XL3Z+nFFv69O6w/rdwCsXONSWJ
1W1m2wypMu7T37EKP+aDo9H8mhdx1k6xOXQ1NHK1VbC22QaxNNHpt3vMRcaFLRgk
A/vPlSlLczF1xfpn7dknFDGSaprW3Gtj8k3RLWTOIplvK779z20gBaFHSjlSk187
G0zYBHhw33QT14HiFQlYq5XC4VXWQxitmzElykSQp/reH2WE0dWHydftJo77LFi/
xXf/dccBU2s+Yky5pRHt0AHN95x2Iza7JVnM6bNciRoSAHl4Rov9rfP3NO28TMr7
uAN2W5xCE+hRuhESV9Z5yA2fQseMwQZjN5OElXxA6elryBJvWX6Wq5qpUUllwuY5
qq3+59q9guzY3D0n9nJqRP/cjK96Asi8ojPvXwJFYnY8LJDI2UuC7NGEnuuw0FPn
yjEnfGQFEjEqERLzLidK6RAjBgZ0rUDR/8KncaOl4xbRyKNVyndP3jRWSM2pwmAI
3LjYk34rla/S2LgTSRMJ8wNllJrIUAc3NnjHHNflWn+9mzE5S1h32hzrIoanMCcC
TriQk/lOhWRkYPy2iAdlE5O6xxui/qJ2cgKSSBS3jj+dqIxjyrrJDvJqOb8g1I6V
DnRSzdFHBUu1CpcZB31mGcQ/oeJhWzMTM1bmPk1JANq2hYPiOu3a5CjUGkoWlS7I
zgt10isRKI7GQiytUtYx//dMB64hnjGDmiz1PSs7vO+UFLTmbzXHj9Ep1SYAYgEP
zRsjGjOk46JUpSIAp97RqMr4xxwrZow9jKJtBelGmFdPsgaF6P6GlWOT3pjNeO66
JAOQSlZmMaMvz8minXUSb4zWIFTbtlwV5ZJcJxmJ3i+gS0lUjjSaYsgauFEiknv1
Rc2Z/KfijzZsuvEzQjTp5TohG+Bx21kKR1EWc8gjF8FGpJLI8klPduIfat1IpUkF
tS4d1LnEXmmAm+QWbRXdY86pbcfNCEh0RQObBePLLziNGXXDrQbK4URRc2RqacC8
3WquYWyR0SY722JTqKh1b1KZ6zjpkNh6outRD9sSHlXEizI0NI1O5aYPqmCqD1Ys
RwnG15lPWw93BY1mtZfRODZxmN6jxHECl8JtmMznM3BXjRTBs8EEUUu+L9LXd+u9
maZXkObldNKbtvMc3x+OkPLGSPF7IXfQKU69QBVvAifC+OyZGonbzJj9qnxhoAgm
7S5R5CXSwjw03qVhOhWRbtPh+LH29PL1lwfTmzPb3Ec9nCCAQ311iWUgaJjCpthO
9S+080nBj3TU1lvOXjKK7PdtFkr4rH5xfs+NQdLidBqiPf9mPny/m6xEN7Kq6OCh
dLw22HNzgTTgPkyLh3ZdcxbTlAXdcWvUD2w0Hz9KZDTtyxQetjbLyf+7HN6+6Oo7
bVJCIYVokhX1wLlHe7Y847eubAiuUM9QkmdfWWiZ2ReFdypu/XpcpW+eGi1DYAOv
cP2z6nE53R4JyRCM36rBV6EmhCFukq2nQ5trqEWoPc8ZW8/YkngaospoiZbLPUve
0oG+hppgTG4wNUjexadL2claAnvwjbLj4ot+LujyAECgRWCAwkXlFA6Fz2GyrBUV
A/Ozlpxzhci46SRudbWO6uDKWxM+pOIWalGQGkc1xbGTzJjGC3FEhvlRcIFmDAVa
HkaQlZwBD+G2TLynlmmY/fFR4ru424dSPEinRqEH6qLcacdOwUTTcqqGa9W6DS/i
9sE1MtgMQSnfLf+0Cclbtsnbo7EU0SdWuETSOA/hoDL7gPUxc0Ly9VrsTzWKIjDt
aRGENKhMeBI1gy8y8HHwwW9ckhNos9zipJwE48QRovpD+li7i0B59YM/zCV+v4Mo
BDoQn+Qtt1d6EtzG+P5RkvRMSegq7tJssNtkyaSCojjBXV4V0nhz3R0oBnyy9ZfB
b620KFoVXKdcG0E8a9l1+8CsTHGB3FacOMwaDwUWwmVnQVTRpCIdmGQp43yA8qfv
hZqi4Xnq3QCFZIzwO5+Hy2ACo9LxfF/VZJC67pczbgo1nAVmfptuwpGb/cfgnej4
rPrvLHEHbmh4If9l4STWfFgzEKGbn779GScpvekMiVKeDSJ+oVybxs4sdl+j5YNT
owffYHQsX7e6XMKWraSmO60xwNMyaCakfZtPDnaYLudFcxc4/bcC+p6s3DF9X1Zj
tbyF7DDjSpuHf7/8TvNPkKVIlOhU615BPKWGiFbkaHsg7QUBGSluVrGbftMeFD2T
ILpCLYVlaJSsRMN0CHNscoM+GVR6VK4GxK1HRNzu1jeKwfI/n8YrrT4yXHzN08tN
hzACQnknekjNGRmVZRLE645qPEaOOWH7XxO/dppq6N0oukallLhl2CtTAsyKuZPr
1tz0xDfSYS6qAnSZ99CjiRoYLGjBazjV2NhGhcoCiTVZoLHsnNVczY6RKPWFu2il
fuDtP4adIYakoV43d7v5zCXW7bBC9u9xgvOXxpiRFakx6Rp0LApaquX+Du0y3+9/
otKLejogGipZ3AJJ3PjIgQcmflPItUSs/krNU6GPfz+ZAuO3bvAA7Z92pRWREgVn
mjK2QoOgyk3VaQZdJN182GrjZ5unCQ2/kwkcVtHXMDkQ6s4YOLHJKBpK40coqvgL
X6hMY77KDTEWE2Qr5d64jJ8X0ZDW3Jtrfypg8CCMFk8sJ2WyRkFikp5oeJ7elly6
q/KsqRa2b+b5tjaJpudQg8r8YmgOWI9TVOT5z3H7RC9B1Pp9TDhIDKu0ye3NW2QY
4/jD9UT3BBoDjVyDyFShXG0oKnSJR8pKa790QTUQemhz9xPTRDhmbN/HVBJz5L+7
zPA5Fd0wTyrxq122jR4vfZXWb0ZnKdvS0se4oD+eVNqqAHiZnHEbSRdAIqX5H0u+
QmsY1J8Si4XsZaYxxf1XuJtf05FStYe9QEIHQWttCBNQwPLXJBKOEYDh5x6cyIZZ
oImfzWbOy8vppG77pzLhDYKmZ0+ia+DB88alAHbMo6o8USr6j+qnO/qsiHIbKmoI
CkR7YWomMO4WnTHpWzVfxK3ufjjT8Y8n+gGy65XFKsm16QYedwQP+FKXBr1dRRiY
9psWgAqF6DLG0CxqhLbW671nLgEhtW0VlJWbhfvPcu8Lx0c3o+Wi2nAqsSYAd6H0
+lXl/Ez3L8bXIai3nZdxzIYkEJV2/icDq1PlNDv1IrLGi6p1dyfTwiRZ+e0ySUvV
Pz5FsFEcEizlLUD72aliwxjawtOPurTzH5hHYQ/W92Yp9Rue3W/Fp4llrXgQ9+OB
iaR+XI1GChbUn0mFSwo14Auo8NO4nObRZWYou6ztKQbG4vjAwuqvlGHlZ09A7cKj
O4f57SRnECTdm8aXn06i7MjVcCfLpNoFyr3mGz9Q2ApLF4YzdDvDVcGqsxK2OTxl
UhHPP/3RKcCfvPYpUZheCnMEDyT1HhFt6qcs2BrnlcqPbCsYTy6LRshpt4ePnCcT
pFV6Jbm3UlmowgAtyE4rlFTqaCSJweTjVpzueWlf6LbbKjcSdBaryVrOkoXxfLCP
09cmILqmKi/vSR102aZZO0XPJ1Ogf6fnh5my5MW0liY3NacSQRP9FKgHFcHQE3m1
78YNil7aaqKP+xwOy8NXUeJR1r7Cato7UUwlW1bopLt4rTIKxJuBpSC9hynw55ZB
DxDqZlO5ujMqMOTpgxen4e3q7bhz5KzbeRf0CieuX25hdutSzVydWOY+wEuGOti8
6tAc/vH0qU3rPkryEkIhbAGWaOUfBoSeya8Dx7EIIJ2NhwsuVVRd77hbIMOyzYBo
M2lCt/G+3aibUWfqV/b/gEfQDc8R1O5sch09mB2Cyv2z9/Tpgi+SOzHgb2pqW8Yp
Jj58nHSiM5hbNoWvKzykznXGbHBIk9esj7tsG79Tl6gre3YCgVpWuq7J7ZGIJ6Vq
YqENW9tOMdmdq+3ey/Zv1SqK0lmaMqmN71m3iWjPwwQmGPLw1NLLCTN+hhcCYgQE
xRgzGXm9pW46HHuVtuIGUREyodJLFZ7RM3dIHDsKF0Lwc9FQDo1YdaoR4t2N4n93
uzAGiA83+/63jQBDFYHO78dhP3AJsLn9kZAeLrZimyB5BSGGuHNDAEoSyY4w2Ooh
3yZT0JX17F/ionxEP4tzS1lZw6qUXGCyc2fVI3Zp0hjowXAWhY5G6E4tiTHlt/kp
BqwS+AX5jxVZFFgMfNbcCDCJP4MvaBNxnOuktrLpz0icce66Yhvx1FKJLEJSy+VT
HH5znIrxkZiW13RQQ9mWWTTb8SnwXupTHsc9ta8tiwZlczY1hXNX76K2P3kGh1rc
Y0QouqK1lJefSE986x6b0UUNfZpc1+moZavdMPlo3QZ3OYHYWy8VJrS1MazrGp9n
6mcAv7yjmaMDba9RnSMJC5narH0wlLcyZ6qMHoH4UVJ4qiH2oixSnKd/ElHY40Sb
suWb065S/0EK55POEKW5ZoIIlBYEBORthztUk2BkHm2w09zqPK+NqDUPXUyilC3C
8kaDfZJCQxB9CsryXHX6Xz2vr2DaU/G1LsTwx+kqFxMH7UM0/zCEomXiK3f8heMo
QzQwohRfXJpDnBtG6luKTNox4KNwwAXZSmFjZCitcpF/012zdtLkMYlIDWejTq5I
FmY45SZIwfKTTP4ik3iOUGz+Y3qCwTJfJepDV8dCGzOmD4zQkpcH3I1pRJ2XSGe7
XIrhoidbzJqF2+mRST/hge3wVZrwgU+A9e9eZJksynm0IiHSyPXUQYbHASMnTxO4
6aAcKVCyh2TxToh1HbphfAKSGJkX27F30zAXsb2ie4oxJCx19z0wqRGKO1/xITbF
JzKbS4Xxes7LI/ZMyKh/KhizQNKUgd9qf9sdG7kECRSyYsHOQOx57bbzm3VjvaiK
E1z3zGv7BblCP7hYngct4Op/r/ZUGxMTU1D5NuonEj06r9GouxnpxHySE755+y0a
s566gnm2HJWJ0JcsH1+LwVCBiCg2xS7rYD0mrSS6D6SxIxHDDMMeWjh3bbD90MRD
0yI8YpDqMywXC4po8IX0L9qXDWPhyJ8qabWZlAZ0aUNEYsB6ybQBMaQGtx2xjz1k
SQhlqRL0HYLNEynF+XZinmi9/PEa8bkjuGHJXyi3eDlKO/pqDQ5RcSRPm0/pYAGU
Yna3MjY5q1oRnp7Hf6lFgjFZ7RfyCtboF50+54MePdsdRjWCxPBAqwJkLyNuu2/T
0bXlKVLoUFJWctiP20NFfWgRXUeUBeehOLuN5eaM4js61enUptiCc27gOXSUMpua
Pd3Sa3Y7BhB3ZFWlgFdrsKNWsCRSfEhyu7ejwn9aO85kgvvwgy0BDyRWlICVF3CM
XBS3aA7Zs+jYH9WsUZHHshOpKzN3ev+h9e7YnpLa/5iEjcrsj+dBHJNdCL/jaRsp
Q0yCs4W6UYu4E6y+Ibv1HBUbeFdzxEwsv4Mdg2X6qqYLFjw/7iO3X/xpSKGtyyRa
uL0iKB9y2yr3GMQr81+G49R8GrTbFeA5uHqlbVC54wHlKRWzQEx/VERyokkeCM86
RvWdpGTqwpasQBs1kc7R+JRjPKeRNMNF7JydhCTPxblPx8C1BvDS6vWtehwuy2sb
LEjvgbq6Ru4sVlm8AwzzGziQy2k2ehNf/0NCGEaVIVKids9V4Jw195CpuNsf9Vep
j0MfoPDMByQ3Z3f4P+7R7PVzjKKALU6HmJgJmQAcThdiW4guIia1HW5hWNMliin9
seoNtKsGninY22A9hrqtZSYeTBmxPLAcl+VRVhBI8eqHZSTqX7MvHrgUbSc2J9Gy
UT5qYhcR6v2qnvXe+vydwAFuKyUKn3yhFZrtH78RrwYL0r3vszehsFMy/xFTv4JV
5ZBuG89xdBUTsccWG2og0+JRkeVSd8NvjjyzeB0RCok21jIRmTP75NkgUwJIkq3E
mmiU/+aMb/HnN4E1u9zU/pjaKkEVvy316Fbx2KVxWSA5Fr94xpD2fHXN5+dnYEHM
DQY2AHkMqV6UQ8XXPuttkK3y4IG5BNPkm1PXRORL3+SjQ1VUv573WWVZ1HkHrdkj
gyma7LPmz2lDgnh0iGyDpGScBKnCoEMTnlolHfoxn8X/ta7M35iyYNFgbWOeX/Tp
q4E9VYoLQ0i24SMDH65MgmqIcmdTPYJ5hsysnBbXTlI82+aVEkkT/2nm9AQnbYrg
uWZ7A7ciX7DnUK5POKo83XPQK6HU8uzQYOhU2ga3VVQBzOTaiLufWtl1iF+Vmani
1RiczJxVTcAC4EaZy9UEnWx8FeZJlMiiiw+mE/MjJt++NxbvGbalgM5eDYOqv7Ut
HMhYElRL8BV9xdeP+zFagmxMjQibzAKdLcE3gf2V3J5u4z6/byvPuALqicvgu25q
tTDoCv54tm5zynE0I+tuSit+apqgSZU7Df9nmxBbT0xvlotZBkPa3kxT8uVqehuW
O5U+cOI63PQbt5CrAd6VtkwsK6F6N/OEZ7bzu1TCDWAnM2SacmRtahFJw62JmOrx
hBOg0Nno55N0+Rw/FvAVmTBcyXNFMS5pAhaalZevw9/gyttnTEh1GJph7aaI83Zr
RbaRJXR/fyWpjE5iWtQ7AfUOjVrYNwKXbE0GyYjM4kWunVGbjXsscgw2iu1MQxsg
jynMX2XdQclwTuNuDfix4ncgIys7BrdIuEaP4sY1A1RPMMA9UNcqGUWNdY9J/RZz
uAgobkaG+RZMfYbRQPeC4vd2nbSE9X4yqjm8m44Cd36JWQOW9wI5Gfqr5MZwOf3H
4YCWUOdig50PlePaHTEWOKZ6I6nRQkwJDZnCNbXygH0NjMed6h5mChcx/1CV8np8
IZAzzzv4AucA55o776SJrnbPs8Rr/oSC4VrsDlPh7zNdqM5nwbBokQ6b7jVCaVRA
081z2dhOSrrfHtEdglXnTFrkRP0GnPBUye0gjh0/ya0jdKApI6C5ys7Y58AjuMQ4
T4Z3QUHKjb8Ov3o5EynZP5Hcf74gGznAcUF227LP7CvExtpVmUkF/tLEjYWu9KoR
1lyvPPpmu9Kirq0qJi5TIwN1g/WX6EYoQ8QtEUGHzmRG009htl3Dzm5SNfPfqBLS
vYA5v24YdA747pUNy0lhNfE/omE75ZW1vrTfOf7tSySO1F1DUiL8Pg1mhUtrmEbS
EW+p0NfMoGHFQszpch4X7uTBPbhVsaMESMqinkRV5s+bccgVyGAPlRdHtIwpWSr5
H3io8TaREdQOvSGoA5Cj0gvAE4hazbfsy4pqJzIOm2pzUjZAJ/PlJ5+LiyMvOHk1
7KrLTWBL1Nos4O75ZMy0wY5T5sNAZxOGKYZ5nLF/8HS6Si7qprrAoytDcShnqKJM
Jw6zpw8/zGr2RW+dTWmY5QQkBxX1ilSluleUt3p7ZtekI7ynj6VJC59+emPWbJ/l
/m3/uL0Fz9ZvEEODQuMwvRu8RQh9O5m8RNl1ANIh1KYhDJlCPxosmG1yygKXxUJf
BXOsYa8LJTOsHNPwW0Ca+jQf3cIRW+14Vd2oHC/+9Yj5hTkaF1WVs8CLpKHLz1Jq
4hx8eqko1CeFl0JuWC0LRHTGZ8kZ2j37wqKQxJm2q3oanZmNiOgTY7WLRjxcPvQx
RjnzS0wJR2s/LBOL4H5ey23aHvycA8uIWi3OEKtEqk80AMavYDNq5T3d9PXPMeaV
vAMnLHFnIN1vVwd8+hfxm5ZA9z8/LZ2yEbHhRHAxQXMG92l8gxY89dgtLT331zmj
mvbEvK7BOwRmr/22RlvgHXLFIq69gB23wIqjPz03D4Ps8cVJA6V/MrQwoc8QqyjY
TqJ+M8Na2kp8Z9obKdqc7uO+ZeZsYherEMVQI7pCUuvGKfL64Mhyqvy5UXgRA9q9
7lUozgTpRDcJJJaEOW3caWXrQ0MiIFwgS6OZArPsjvGD8Kr634rDjgmH+dE9IyZg
lHjSVUtKLAcNZfgivmU/5wDgh5FIW2NmKft8ZbUk3MwxVb/cN+BjwBexIcvrvNyU
ndEH8gbgc9KoLOoQ89qkk1RMOX/XMBENPZiYHAdxT6KpHUT9Vh8JCOlrZ7YV2Ybt
5f1FE9DMA8urhiT9ZV/XlfZ9HfCTB6lT/luRfOFCrYKpGhSw/MKIzOv61RhVkwhR
VVduttF7aD6nutYg9nG6NSJvDShrJ2P5MFMoxPTJDDE9wObi1qSj0hspMxtr+1nq
72ZmYfg9M40ea3c2RBtrCYMNnfhVZ3BK2X40fIm27J+UVUCeg2bl+B53XJbFVvpv
32lF+mwggYfoogiIvEC8yWTRGwFIq+Iz23q2PPd5lYHnVbMmBjtJyyrvR8/qAFVD
DNg0RJUnDBFrhcHdrZLSx+MbhlBKmWaoiK8cMu8/QsiK5CuqyOr9038rQWUPCCqa
vzmq+8NK/R1uIB87FfhTwtACdcAthqCZrO6P0edfR86wBYxd/jpX9Y2E+ZHp1/4r
Wyms3t8uGfQyEMY3k6iKU92nP90ywtPDZoC34MRe+3SUCv3x6+vpMY+eEsMMn7LC
F3/Ngc5szJ4abwAWUgjagL6ixQlF+lFX9g2w6cEXUbkVFbW6Zzox8vv8vTBU9tin
NmpWxN4J3qeDWTLsLmnJfgd/jFXff0O+q2SMgVZ95bzbK7YBvi60hNf9ABGMIHqf
RI3ukg9fZlWyVkO4VAXqFol2YBz4Q3oxifUmBc3+YOyXDLW3wigmiDBUKxE+CNKd
+XGQkQgE9f3sFguVuCDxInjnll1RUSblzBehNkwFnJMtJ1j1VjoOqiSzYZWTxOsu
WT299HS3jVyRP5zGRLVU2mvb4I86pfvZidSB7pmdnG3fvQ0lweRfnLh1wEm00vJC
MxUbpVNLT5375MlxIFDyjcUQ7B6wX8+3GMyx8h6z8+sRnoBIDmEcNp/rUsOQu//b
IwbhYFJOl9KHSEnmcw3PnihZO4QnXDFV8y+8V3EnKbyaYY6oWBXYyTROpSzmVObF
VWAtUHxEfyT1yPO+0UYbahQEHWyibWivqHPzjIUdnR1xhWoGkoc0ypcZFsFa0kYh
3jF/mjACV4BdRwIOtlGJWX7KEGcUHdvrud20gPb16VQbjDfU/tqy3jHalU7urkpI
X43t6YBsQnGE1zjuxy7MWImjkDg3UTTgvpOHOtJCDVyfyh4L90hUnZ0ADztzwV93
agOvRZSsmEGfHZvOV865BjRdAGrhgGR4i0+begVg4xyYyFu5voteYE2m4xuQmsvQ
ql/aPFzOxJppRjlbtndocCJbIv4Fsd9SGOjvQT8WM/SLM9b4BsVjyp3rgQYl+Ytm
GRRgQw51WlfMMOGUPRklbAJ3ZH+BP3wAn2BfJGTli2bH8NXBChYWNTKqcEsCgiJi
Hj2+gDG/gXzt4lzYwi9zsysK5nwfWF/RFoBSAdH97tM31hGn/VxSd7VrtEHYxCk0
kTNBL2ArE8eA4X2XuEHTbREhgrnfjVcEIf+W2R1+0SvxNfLKThL6hS7QVRyakufn
YFirApn3UgBmyp6Gfosaeeqopej68QymPcjDeizbT/yuPV5IuZoRU/CK6xaMbvx7
R4BmMiYuHtkee7B/0TRdMGDOPmNRrPFS0ylJkr7Tzfj7zUL7/rMn+jqlc4EARbRX
OwaxZmRQgj0sGdXRh/JbpOMiUfyah1muitjQ1NZ5PYskgaiqMkI/WmFzdwSiqVis
ix27W8oLDWDun0ByruZj17KAXDAtj075knhWd1mIOL8d0OJYdHcj02ykDT0NjtRA
P8csPqo2MX6ANnW59zEWAbSd2AkDvwVu8YgfK2YVR65Yp7N2ek4CAPl3X9WgC+bl
D5WbjsvTSucqoSVdtGEQL9Vn0AT/wNVEQv4Ecaes6yM3cJtmwD1HfKKBuRkS/HJT
F/GRMVo3jG8obvggk7wwXOvjdDrSp3A6nHxHc6BolNqp3/yAhul7tjdTpBkt7MZT
8H43L4dKSvwb57jDK9RIl3KCHHMM9ujG4Ex4W0h2Klc98z5fR6SPzg7xxUcz+iyu
pVbZfm/SEMRrS2supQjA1vZkhcB11HpF13ugfgdaDbi1D0RepvhU270glzvIrTCO
wOIDYEgt+yycY+RvU9uKCQme1oNrJz/Ge3dP584e8PLAmJenVN4leGi3WOZN3T1F
ugrkTx8Ojyw6C/oKUY8K/FjMqSCxkqTpMTMj0FgUy9060PaQdLAeXcajUumYnyhg
jCHfGku1C6AqtJYZRH5/nRYXLLL4L0H8zbFH0HvBJ7/OB5elQ2EFu798qVOyvBqL
97s4N76SuT2cNmDZizDGZvjWPBmhBgKa4bQxronuDThCxrS20dNmkR4iVsx3iDti
F/bgm0z2xX5IyML2PprzglfiOuZcU+/AvHAIWZia7UfN5MA7KsHo3oAXqotD1cAo
zyjPLOZ405cenNGektKIOFE/5M3p7OAuaiQJUulGFCe47O01fuZOnECrc1kTvHuc
KcTlllLzPcxAZJ/RAxQaHV1O8cdmvbLaT5LL82ydQfw9dGkLg+MGimcBBtbNcr1s
A1rauXnmjo646yjc37DQAm2ksxPOb+X/ujBXPJ052rk21i7o1jZLGPHx1aKF8wBs
Wp+e2k0ogb/2SYf/tNi01oprGVWDCYQf5f6qwUUxjiTHw1t4LZbm04vhryTWMVui
IMJsFD7/8Q0YLaoazwx1YD2GanTD1PLto/tL5mQoFXEhvtzywxpZrry9U4yCDTcw
UYiTrZCv+c1H5TwCPkfrUlT6qtVtP8zWMg6NiC8GjcWei0QrupQRlSf0n3V1gNxv
d+Jc+nQmqDZtOHRcLZPQPewhoLpld1XmcXSMd5t0WUaAcBPJj8zKObB2mGYAyllR
D+NT10NA1zqWij+mLr7Hokw5q8AyWRxD3zKAxBb8+2Pj5QtI7rseAhnZZ4KiIUCr
VbxrMa8CdOA1mWx6jgZ8c7X7v6mNXZGE9FwQozFxSiLa0r9ifTf3lJxrfPqh/4QR
SaZuHe1DaSPYxiMbac7AaSoP7vrSGEazAIeE9s7nHnB2T4a6VblsP6kfBEziMZsC
EqUxkC/b7baQqcf0G9dX2xWEwt7TumxB1TGX0LYeZLdQvv8NMmgdJtPbkd0dI8zU
KdhJ8yNDdSwU9TrQvoC7ks+eBx26Bk3fQ6GJzsf1YJEck2xPaQV+DYe5DjFHJqzs
EOMSBTrv3tJPdug1sqnBaVuspEBOLUv6f1d1odOSs4iorWNEwDhqP8ogitWua1V/
v1tF3y/W8v8nY2hJhue1ElsXCVvDWTm3gOoFDpnxZCVo8Kf+qtah3rN1NV7diyuc
slpOOZRSEG9e4j4ekGyNJVpr8tayPhYd7u+Mzgw6KSZ3f1GevCbJvmUTRdseGSHo
eXNvJmFWItKEuhN5lKazKBEXzxmXR+cScxKVNtrHJYtYvLyj1bd4DAkw1zM3H+On
XfaYS2xCgRhCmdylX/dPF+F91KSrvBOwArQZSoeViqnncPTklTDhBROhev6hNJNV
uHr8JQ3oNibVdF+nYFOo3DCO1VMuC1e1m72WOzdl28woK1nunTQUfBzipMcIPr+L
5e00Y9XxbxrJC7HiWoqbC3WjJ3+d+QqaanpZ4bXcfbldw/psC1dr9DCbygMz6kl6
TujW1Zk484C/FJn34zJN1VKMDKdNx3f2de7BzVLx2yHaq7LgAZn8aC2zT4IxWlxg
aCCQXSEXb6QUVeIYDC0atYTvLcLeSFvzBiPhEkv4iZSr/9Bs/dX+m/kwAVwHhnQo
wCq7iqQhBRXHiiDPFN/3FtSQUisyO0WnCCz20Cvwup2A0pdvrSlRbT/AS1ieWB0S
fyu2Mf11oG4HX+EPQxPFVFk+KROVVpQYea6/EkegCQnMWYj9cDh1xRUFPM96dd71
uuwv8eCMYyvhHpRFQ0jzpedAsBHlkmN9C2EDA3AwbX6Tl2ALTb8KhwnRsizp0gYU
Pl+WwMMmwINOxlC9E/HuKCluDE+s3Cc/P+aXKFejL0EQdJNwGv0J1ylhTAHcKl0c
4NwqVJyoS0zqpb9Yxb5oR9ComLoltX1EKFOFjOu5LHMYMlzeazvthfH4+XpsWeNd
8Ll+usEV84RNuBDsmkTDu1qf5+6XIXIjCwBo6/l4M2j4Otc3p387FotLChAuk7pp
t3MglGLP0uaOGSIeZgC+/MZoVs8ZrjDX4CIEiEPCmr3P8cxRzgwVGpZ5nauTt8jN
sgnm2qHmAAdo8sLbbyBEj76aY7y0Td8TCbzI67qVqbnJyMNLXWenB2tGGeeyUz//
okaYhXljKpdcynrHOX8Ii5PORyrKOSgKL/SS9Nm4bJPd8mmP+m0QjokBiQyfkmPe
DAMKVe6OQ79q01ho8VxiwsOI/CVaeTaW1S1vzSRosI9SHcUqkXxSiR1SDP4cq2r7
e59ZmzGrQOATlzOw5vIHJPEmmQILD5sxIt+MqzLa9HVIAB/qxDupitbgt+6kFdIl
NzZ4UR20D+o9NLMhaEbmVYB041kgkWnyUt5j6+y9lCjqcr1RUofkI3AMcIPgCJIE
XqgKlTHJJk1PWrgVGRKujnL79G0ekT7hPUqB7Y+CWXnuUwQWpLDrVjP9g3pZQTBc
bT0fm9tQSNTiTD4N0vkxOWBEKPc1XCAyqNFuSQ3p+lL37x2/tDxPWw5rMmYH1/JU
Z4JIQTi3V5q0oebULcfrzjrJZMTVM40SMtuikllzYaeTNbXsmBCB3n3p3T98E5fA
qq0t+RdZZOcUTUvh6vjiSrfM2DsP4JP81TVdlUxRNWbH2yK5AkmR/4vxkdLlEKCj
KSw5HvJjbsCo0xsWnH+Fe50g8Y0ZU9CYMI48CnXG9fOboEdeNLtUx3JWw90BON5H
assaxUXTNj54KiGPOoup2ea6OmdPI7pj/yH0Rpyxw8sJpIfAx6auaihWUd2FnOWH
497DCWJIw9v7WIA+H6Vo2jD+T8GNEqHwCE/ycuDPXLprftbNORFYRRSdbGcJEb2R
890dUsEXnCPZy0XuQ3RFCOnG7CC7Ecu+kTeZMgE5ysiT5kmxGgK/6l9OQG53Z4Lv
7IsDI8+PNvNt3NQ3sKHTi+wKShwGo+7IVxP90p54UyBiMwRCpm5m5I5RfmTld83n
/R0EFfpueRactZlEkhS1x+ElmyVKPi5nUumM24u/3SfzjrqZpAukm3dk2JQZI8r7
UFtjaGt0OhjKYrKysKh3akffVqOsveaVIRCzdUzDuaaQRx0zxqJfpB2D1kP9QPrX
xHmU6im1W1yxFa8xI0ptLnZmP0CYrg7dBE8Y+OGCku8A12ii0UtfIIRWiAkwUNk6
UUzR1RfXUiRUCFiTEsBERxBLAYYc3Hk8N7laGfr2sYPV99h7f7OK5GYRYsQVH4tt
Kp/SujYFVBTJrePGfBb8RNG0BB9CMWPEIGURJCT8uQDwedUQaKLd6i4nSuHW8v+R
eMey47ZDX47U9B4E1C5omH1SvjeggiqN17/EuHVa7Uk+DMiY0chWESZi/jPg/D2Y
9gSO6e3w1ZqymisMaTKsGxfEOwT6UXru70BEmdDG/erM6UVIznpim/EHOTCI8rju
q2eJj7RM4TJIrEOdT0pJXnm0WMbZx+KnyNOEGZOiS7OiwHLH38bh/fvp6tOkoyf0
Ccxa4nDh5pmMK65OAwvOFkinQgfAI1LpYgo3rOS6jJZRChXczgq75S5PkkprNmqS
cU7HSdjH9JZhRixt9j8UTUN0uKINx8XZchiKrRqrCoR8jyslqOl9n6Yubqs2s8F/
JgRjBX7ASpq7MhEK6bhbwWUkYDJwYVqX/FfiEZw+CK0vGqAUcAG1MKMjn8zkfpA3
mWTnV4ADtm4oGWYlsDckLvVHeHgYvij5weqMsxBlCx7wbczqnYjTYqkPw1ATb3Zo
CWHaHqQj5kjeLn91lcoy0fet7m2YNQBaU16RBX84acbDPDOIID1YNi2Wf6n5b/p5
jpl1zRW7gSh4UmsNVL3mFAkBCg3bkRuFy5f7dS2dvq2xtJ+DNEfK80msC7x00cNY
XNl/MsZeocILcyIj6+cNGW40w7kQa4dciItkCzZwaLNixMpdl43H/aGmABZepsco
FTt9O+FrZr7U4MxL3rfJaz/plGld1xNyp8lTYwha3A3ls2XDhgRgge8/55nXGe0Y
koqgB3kfaoohrigEhCoZeoJ7AI1q3XBpRin5zrlazM40RUAEDyksrIh0+DT/rBMB
+pUdfoeE9mNn+L5p1oaH3gjTyGJB2NBhEzOnXfcqxkCH4zGdkAB1IiIOFIbuUHQ5
ixuInEkr4MO7hQY82YoCahtCC4XH7h1Gpl0RYmTc3iLn8iBAwnQzn42pg4S+3Gu1
+icYMCuwGJxT9SHtizcSdreAno0HhDSlL+Dyg5pQRSxxQtwwMJVyVnt+nwJdJStO
4rncNQMngrjk0Vd3NlHSF1D/iJErstsUCiPK5wAEgP8fji64LWOoDrp+FCXGCPJj
mtiQJkj+YcEXLHvk2GV3z5f5RvG1ahteJ99w1b85iPp5SeUspdvwD7likECIo85t
4kPWen+LWH8zXfPqYJfbhO8kksNpirmTDN3FPPFNOuYbfpE/H/+rfZvM79PSaA0c
wOUbQ0JXgg0KXpLyk7VyMjSjN3zPQ4aZvRUXfFmWIQFMBCiLO3GeMua3ZeJ40CSu
IxcfO6Nmwaa6DrEJOz/RBKETDQtqueC0EJV5bl8WOcx/y45ycortIKehpcL5b6PO
e/8GZJKt+YUmuz/WGElv49lvSWkU3G+lINlBhHsTo+g2SRFg/HvYCajwfBqteT8j
pUQE4C695Jfkmup0EmAqNZJTic8dqxLmfaA3ctYIs9HkawxGDd336XqUTTCGbJhg
Nhby3PBaxf8BkHxxw13eh1ycfQY+dpPd1Zd2cAkLDZQBlLpQE5KJlJG37ImDjM2K
RrTY+bQFAeglBo2qohCtFGMHDqqlL5RTW05tHx5c0sS9/R6OyJfWP1fty6YGCVif
zJIeHd2t3TpEgMVkw7enWcs3lmZhA5At33OtOIbvx2IaXuki9myZgMlJIfCEC2sf
hqOTWKMAIdU8iiMdXOhaYKEF28MbfIQmPDMfWHVwvPetWz45GspMZDf4wonDnzef
quqmJyAvWCy5eJWX6vkBgN2qMZMz/jSadBrM7YAYzgHOUGr9z7H64bL333EXy9CU
eaksbF0DN/Ev8auSRDgoJi+xFOqMwqlBN+D2Jr6I7zq+fbOLZeWIN6+tm6ADo/fD
hc1ZtZBt8Z6arV5woJz6z3U4z/aricEGr6ag7/pTMPRvCGU+4cF2JR3vG7qn7iha
hleXAfJ3jG3IKMsx0u/iez50eDcKYnx5cvEyRu70Nyq4efiddpK9fDOHzDC4FGkt
7PHL6XZJjSzpPouG1mrF0d2OohypZ3bPRZ3oHuW+YkBWh5Qp8tnGQ59tWsSE0dfZ
Ex8QTOWalCcCqqRHXm2eli6h+loOwTutMFDZoNTfkOPcmK3OyRzWYHUMm/ceeAVN
huxdqrue8ekSMU5bnlj2bzoNZGKDpOgS1y3EcoQR9GW0TkPH8mW0eCFWSLBKq1sy
6G1RpCGW2+YiqZqA3x0+cL01u0bPJTVxz6TJ0wxBrvPIDKgT4I5z05FgtbyIxLtq
iVT0A/AkKYtIVv07Otk9wGeNdR5/UtRgiT8HqLanjuQSj3qcgjr68XaJ4odg1iqw
wysQ9GdGS0RYwlnWd26xqXBWytGS8J44AQIqL5BR4dIrkpzAwlF7ecUA/2TBL2UR
wvJ0sxjSgi78iVLbK7aWRZCJNlcd8LewUaYJ/deWcKB/ek/rJKODoIGlQmIfMzPt
Z+5HUY7jtuGE0h+uXHLBEPyzDg+Zu6VdsgNszkhrtJKqZgDxJ576Dcu8uAEmqL8G
atYAV1apHVhbo7Z1hUclU83SiZtRABqBWwlke2MhAu8MiM8h/UIUWR3yya8bALFg
Iooo729OaVdjGSy8kPo4n5/UYjPTrC29vcWp7Esju78FmpjEPIzHuLJlcWOev8gp
465342SM96r5HEogzPmWnuMwM3dzw+nozaGmqGYjwQDDDG+GJXb/cbJ2z8/itWCK
wi7yElnzqYP81ataZZTGuBmg7APJIl3ijKS1Our05Vj2/PXUUneLE37pAWkZBu9j
3wMmdbXKKhRyC5pTzqq5r+qdIeZxfJKfDueef1z2bzj/6Ab4fnSTbiMcnI5oPUoA
S2rhLH7vrvXMjl9gqebXBB24KIq7+dEUiqA3mfiGaZOYNmOVSvTq9KOCLd2aYJbj
weQd3xLlv7pLhXJyAbRQ25C8euFAZG/9/ypdhd8fSEE5pFnTP93hq8g8f2l3P44j
AY8sEKdUOCk9MYIiUY86c45Ni7Kbea+9ZxfOdcaVAusipU4Kg8r4EKxVHq/NwnOW
xRCyDgMTtD2dFerH3RnhnINjs/hR/gsXAOBepSyvYq2waejXCStkBYza84xmxOqi
evxaFzKiutcCeM1ZMVE5UldWO4Xi5KCCaf23zx792LDj8tuNMOKnoIYd3i95YyxY
2mvkfrAvcy6rOhLp3LXXj0rLgv0lJyQbWREw2VmwHcg68DJho4P/t68EcHOSDxrJ
NWTADz9e5JgIk0zfWmOWjTrtdd2jXycHWtqOfIw88h5RJzcFIxoUaFHC5g0Lv3O+
3pjrkwHZWRF2vuhgumFj9Bt5StrHiJ5wwZAAdZBizorapsqXsyIcdY4Qd6MBn9Hk
S+T36n52JvLGHIyh835A9hm4NvBPOlXoNtIBZnTOKqOkAslD857O5aOJGpQF8F/3
ROIwK+OUvN6vKRauIKa1csw2/EjvAOEvfsJfO7XsS0nlgUNWBZHimKqCNCZnjIPN
Lm9XzuFaWivQ+mOXoT/r7Ke7zMeinEfCCDjMyiPHhngZQkVfiQ+wSwvYT+adcmUe
Pu6B7AO8KOhIKO249DM9KNXZ8owvUU6VE1inbL/pWUa+BAP7yDTa3PMOt+XCLqfk
toaXeVkRfp4Fa6DFMFe6znE3xs2vGGMD4GbAV5hSkreFEpFtQn1JKv3FFuvyfJ0c
W422z5pT68WuRUl+YZjiNi+Vh3EZY64QxrAdpbFfmQXosLmy6/4X1JZBmLrXU3UA
DLito3Fj+x62BIbFefJiRe5bJ/xHrUm5QwqDNCeVeWwfrm6nq/rMZG5l6923Ham9
rNdJ3Xzm+pKHB15OtZW8GCtH6betryGJmOoutl6hlvKAIYqKdZdaM3j/MdyIsYv1
4sXnEl84fZH68ooDq5tDvPvTshi7uhue1Jr8+7R0ZEly1yUu0usi94609hWdgG1I
P+GSdS89nRAZn1GjGN22EynSCTevRVR587Pz8RSKB3hcsF4pSEPEkHBQdfFaM5zu
OZBSGLhgtrrVQuJPSFF85Z1QdRPKPh82NzUKvOfm73yjzGvXTFRwFRfNf9fq2+wU
pXXP93eNTqOo05RL/BrvFseI/Ea0oCAFFU954o/X5wEbgCxAYnZ2s4xQisNc13iO
OzEZaqTirBvICe2dKpOFHJIYjNgHUj2jrRYeaaVRJKGnIExmf+1skAadtUxydTap
l6K/ENA4SevEqDs4z3haWu3ShFYDqvIn5cHJmcDG8hyQ99uK2giokAlhkwhWd4uC
MF1cPIRFz5payZ6IXwpqVMA52/WU3btfL1gB30GCHRjXQrOwIcfn+WdUZk3wTwfN
Kn99sbDnYRv83P7SnkY0NErARpgzDftFw1BJ7PsCf9pNcOGEB0j2s+v7dO9KZ9RV
IGULwbBAlrVEeN3voVbY2yohsRF0YDknQ808I0Wu7UjMbIWGKV2F+MOorAPuphuL
ngsTmTtLgJ9OAKTh4UriIrZhaLy/CNAW7HE3Tfhyp2DhEV0xnpo65RR9UiOfezfZ
6BrOScwAmkBRAuQwhEKBmJegtCFFQjQBMgBVauF/zW89PS9D06lb/7oaAJShKbT3
rjXkFkZKCjTiyPORC9IeYwNoO1H6gvjFCYRMeSI6S/fc7yhSazEctNOUMOTnda5U
sNw0ZAGORq/AlH/4NNuWxTvdMIMNMFzqoNOc30KFJCWax5coXXSE8LWWzNJ1Di63
ASoiTMjn9ZznsOwbmIw55sZoUm9/VNu8Rp9jIggpaRLPcJBSf/8cYMhykHllYkN1
X9mgf6AT22YstoTt16eWFb3MPmUv1WL7qkB0y02jAjZpcblJBRxzdG81h3X+k2gB
Z078Fh8bi8PuE7dp7LJL3l0KV3KUWg7srNkiFICzWUxXIPQcn4nXA2qZnk8QTyCv
tLs51VCjMfpEZrUIOZk3qOtBp60q8V0tQrp+XmmNQ49Qs/82+VCSDs/oLHQquMRD
ECBArwSnlo79UWVXud0l5S4V+cWp5Suvaq5eqmG9SK52Zo0apjXyNM9vB+ndIus7
ECrSfTm1mlZ6xlmjDwQlpqCKbiZsiJ3jwcGjnzUwmSoYI3OSIdnEZRhrK6n9v1H8
u99X+jxnYcjNnlTVnUCEVxVFiHZ2Rd//xMnBDE1Fgh9uOB/OiSaOX2MajGAkJK6y
ZmfZ7UhgMf1hvcAqaoF/PBpI9CUA4AQmi6fI3sb5KKf2hslKzyYJR8UpxAYra3Bw
VTGLlzJey6E1FewgPqjvRSrqVjSltI3gYUjmIAFBqHH6rTE7NP9TIBhOaUwZhzh8
Ct3RyYCzUhmGbvIGgVG56WIstkNLa/Mhtfx/lEwitfXRDKGuYysChACf6y6blqaV
GkDMa0w6VPQdp97bMBAdSp47E9lO/QKJH67gaxxePYJ//OLjcX6iMHALpfFRJ+NX
lIoY8GVcal/88bRI8d+ujIeaHPdk1LtOKqczVcAvOSJXJ5ryxxkIBEWU1mzGOerO
l1x1qkBpHTprOqSY2VThV3ljSNMQNX45bX0EHKPZjkb96HXbZNfV1ITqdosXZ3oS
Uh8Xsg1XZmJCGsYcQtp0IO5p1XYT/iligsogDxOKtEM5M94YsFVUp/P9lbRgSHxj
LvajCs+D5dYecLGSVjrBzyrvsZt7bQWXvmvCzvV29pdv2gL4TlS+rJJxjgEl6gmb
93aWggldE4p43O5JZkvdYj5s0DM/xSLRjw0Z9h76UUL4uypJRobKehotR2FpsV1c
WJmNly0+WibEdWLXVN8ieNb/9AzLA57nQHeH7lkKeNQZpoEU3y29y9YK6DmmZ2Re
TPv85bGPvAIpCiuxK+9MnelH7vYf4ySp4tbXyhyINN7mx7LYe8NjG3hjK+XxnXU9
rqlBd4HF1p9dV/04ebAH5wn4QVdmgxDp04ULjPKWTRvMMxcS7S2yE4qUtsP0i3VA
uPLjtWH5//1GeNY2jYlLB2Ph+rbrKZgx8tket2FUJDsjMu+cSHmexVBcu/uUpzBE
U+2fptogQ0xl8nLWM2Xj7Q0N1qr/EBNHFxucdKu/vOGVR2ZI0W0devqTwiFHdp5b
A4SOYyf+w+iU8JM37ay24ycX5K5k2iqX2w+4/DbtA2a6GHf1anQattI8OOAk6ofK
XpgQpxPxIqwe9adIiNyJuSZ/BW2pcjlAmSnSdFnrMry//7F5Ry8oUHTdpoN+QvOd
Y7EspCYweDa3G6dRMFrtF6DavrHXbuvoJabFLvB+N9X0RFHl5tPIKE2r8x+5hNd+
Dr2JgRfCKGvgo2oLlZUipM5xGUD2vMfrFCzTF3buujjub933b8lUlr5tjGJ3TEri
YUV30imHoBTzRqwCKyq6DzCA/WZYPfQZhVmQBs2bRSN3tn2EG/P+5vyPWfg8/OzX
3T12tUqQ07TR32BESGH8bpTK6870MYYCDOYxG8U5LFhcZw7Az0S09ngk16VYkz/M
KR9XIugY18rck1Wc42BKGbRHgQmBojNNA5Mpoz8vBJjarWnAJpi9CN8xSwhHIWqW
ThLu4c9Cc0XKlzOtqHPyfQ7+QnkmestGmgs7GnuFoQY8eiwaSyvy8qF9NuoSqyGm
iLWICfcSCes+X5SX84qis4VLt/M84JT8AMNTE4+vC0jVdNYwAThnf9cZndhevB/y
BZGHELRDaIa6y9odsU+Q5VZ6Pg5QjzgIsyLWxF2voLi+r+R0L6jX83AS4EWIQuB1
L449V9VzM/oq5V3QC26n/cm6xxnhgqOzC4sM25Wiqqx7ICqZIJKSfg6Zv4OewaBu
EOv+/9gfNNPC6b0W4OYm5zSsU6REMhYOsJAN0JQ8zn1sYuRwCpCpFgWkyh1lw29e
Mw+F6ExA2MpzQu6SRbAX7j3N1zZgYl8WricliT1cGtDtHgBd4UQmDcU0L67BZF5P
BTD3usd+SrXAA+vKCLnUKEQRfTuz3YR3HfNF9AFkgoDP1i0IS0aLc/j28sfNNqGC
jK2qJCIblB73YNRZpt8ktq/cfdQ0ZvGWq+JlE8ATxXkvjmdSsiCwiiIxWabFWWSt
6JgRfrPmqpJffJQfHSG82+Y8WvIbQ0t4lDgv4wfXgZv75mufnx3WTxOGt3SGLG6a
+K2GT9Y4wfTjdnY+rT5pojSI2rhCk/7SIXgRHSWL6S+4MgWE41l9PseDwGNSfEBe
suiJfqnCE0G3JMI5q4vT95x+4FXi24Z5zLHz+JZK/G9gsnOqNAc/swCtksgr0zQ+
1hFqua96TM30HCw00LlCx7cHI9s6siL0sEdjKyozYPVoU35b+0fzPV/PML9b8cQz
Vu1ot7UxapiFFVK1rMkraSIn9EFfjmEOV8HgbrhvNvU5Fo/b4QlDdJ4LMTD3FG1h
z957V7HwfbERIzQ3gps81Cu/nnuFS/HChwbtbA7ryirprSX1FTr8WOe+tu19YEF3
vnwYhFMH4tO4oEOGypt4to26RsCy5aDLGU+p3C5SWT2MyPxcf9d45cDRoA7ncCEX
lwE0BBz6TOB0yLPXKdFzab8HMJgRQNm83ZcBB4zpXPnU3rxXT7FERC4udkV6T1Ow
bcFuRDPQ5wGLRn7XEgNauy3yyTr/VdsIXJQ853druLt/7/lanBsv66m5Ov3QuOWB
G7kIyYZrfCFGtaCpyvG+3KvZQS3akRdyol8MXE6I1vx4oYsNSLcS4Ki4GmnWTOat
ADPc7ukuenOpZKZZaNLX0Ibjfr32apYIaOKm+JsQ9ba331qKyD9Y84zq31bILjdD
lmQZFzXAy1H5Vd49z3RhAbd+nHyfDUoIrf/rvaycuJQrd0eeSMDxSnFHSDPUK21U
HWDl2ZJUvtvAz18K2D2httik4oP+Xfc08s1/ypNs2Xb5HM/RbSGZhhXUdZC1tkx5
Ebhvy38JK6SL1bfw4I7wULSz72Kfzg54Q9wvmCE1JVSgcJHRmsXQp5iJXwPM4QVR
oPLtzNWVFC02H+RZOCZOnNV3kGcoyAbwQinyARJkr2OM+/24ANl/UlFBjsjI3tjo
4mlx5gsNjN7UGcMocutjoWFb27zv4nvSbdzRRVp/EsiqCInO4kT5VDHQ1UbVrlOn
Bu4AY1xCI+cqVn3U/gFbc+LiGu2bJAfxoRFwiTBixaoUVVn/9ZCN9leIf0K701VL
OuvtvfqX9FMnhN16Y6O1Vh8KIRlbkE8D4WnVnzf8uNYc7JjP7nIvY+YYfgiaQA6c
MrQYrCLPCzFP0+Wy+LAd8WGssmFD74U+nYyKlvJ6UFuXcXF6Unkx2bTyTmWyA0gY
D/kVD0olQfdUd9CfD66PZyVUooKhwdhpWS09tYcOWD8+3HwhWX9Qdy8S2FblEBfi
4uyc9c2spRkEdy9yhPjcsVhYEzPT9Y26XdryvhhPS/+q58O5rMTtskniKXK9QiLL
dozWboa5W/EOGDuJTttnwBTNqslgW6GewLI1BS4r8T2cw4fZ9Bt1R+WCwn7JwPxL
kwZ+R70ysNT25+O0hJD+gm/LskPM2MuSm+GDefdm8NPmjJGx6O0NJ/8tV+BWb02J
4BvbMksT7o9Tk/g1Ydg9XZc9TMQSfydTjeJDDkpDdXwSuoD/dSEWr7R0NU+9y7AA
Krs2DYzS9SKTWUZiky6o0ku3KhBDHoXMPGPuGcdUSrNat+CqYN9wldzYi/VQqN+y
ej2qyFmXocWzRPQZD5Vqy9iDYiEm67QqKPZOyvLKluEJlAyCEfVvMIaPeKwLmqsr
t3BK2oMeME8vd7B0UOTRULGE044/flXNWFq8U1nCXpCTUsGkpAoOyAx4PD77SAhJ
Obqssifk9O7BchDwGhwPQ5OaPmWZ8INMIug/6VBZUYlG1pkM26kARHMCQmUvzocq
4PRY7Y9Pp4OyV2WCqJOApvxR1RTBszaLdOL5WYreEJD+b+9R2v0XUrLgwCaQPXte
aNqqlZhWUi1jgSSRvxds46+HnlIlOB4mm2zmtxwkSzxTiIAcuKxLnP5ZNollCmq2
uwDuGwDjzrrfkncNalUF7ni1wlQ9sWByE8e1D21W23JU+BWdw0bArcLmlNlaZxX0
1NDyWR8xE3ut+YRSS5t3Z404bRjRpMRHKayerdJLgxFDnTduxHO6UIjAbKmiU2GS
iDkRcB9r2ro8m43RimKrCwk79EcBI/UM4BouoFCblu99TP7whNc8FlJe+dWgF/ku
xKKwpH+85AbuO4vNAP6xOQNM4XpxwLIL6Fg8xc1/QY3vGfalZz/4VrdZ+2s+lGHL
z3WOhnSNRqdISvVhNCorjvcl9YZodv4ZtVQGifPkGH4j3Snx6WsA5D555c8PCmyd
0ylDzKMTRUQh2nSAA0iwxWzPHTDfTC/yVAfDUiESiDrZZ6WCpbeYkGm3fUhuiGOo
Kb1ZNVOKNMSGDzJsFUG0xm/81IEnmZ0hNowowB+hLG6wVYoelW8EPYXasOnIYsCH
Skq2md+tij2fOVGfjCQ4j5TO/YSasf3FYGKeGOYNLAIc1YHrKKatRfbpCIh2dCiZ
H3ONXt3TXE9YOKzf517bGYirr3gzk9K4CyS7J4R/ARdQ7dpmyKt13n+rLJuSUVMj
TpYWrnJY4aKWb7rBXHFYVcMtyMHQ/jqw9JSyMPLye0oT8/nP13Hgc6HaapJ3UzZe
0cqYtjRn614RRM18vTwDkcrxplb/838Rl095JS1ofjmrOhyX54j+joOU8kbyo8Te
W6GdvjX+RWl5jVRRwjDYWFym8NlME1jcLKOjz0Echcz3RyrgaQUhbGh3hkoiNXAx
Wb1Mp3y4uIBWsSsd4r4XMkx6A2JH4JBHrynQrutRrlyCiBwVN9vsTV5JI2GhgzsO
WjGBJzjoI3F5F0HNGmfpTySOOZtUwvdHxnwlgz0GxErqpOFSs2/LmXMHGnu57YJ6
uMSsZNyW5uzAgUerSdqnMdR25FECnQqH8U5rlHAF8ONGP7qpeox3OL2/AptSCLcP
MMIOjMZIHT6HXGAWmcpouEJCYKqX+Oz1xeHXnmYM8fXGyhl3hvkJ29uw3YkURaYP
6eKXiPNykCnGOZjO8te5kY8JF5U7TaEHgQ+xMRaA+XvhJeTQdjCHJkC9zXuVdnZC
1wqdqFgMkCMQBaDALwJ8Y00Sb79m5c1gCYhZPiwKfJX5jZZ0oWQNwt/57r/Rpn+n
dxWMnlP6kkc8pAfLKaKqRfwDguDu19FTil5mFW4Lat+x7E/C/uDiySPj+WAeq1Rw
wZ/M71D+FyqgURJlr8DzVJ0lmGslPnvkDSMfqWs8BQvz7dFEso9ETThZTt/pAkRM
GHyhGRKmvFaJ1pdfByWdSXm5ns4yDVrX7SORcaldru7iSiZEPmpXeIhMyFLxu+AP
Qz4OzA+KzH+oTXqlXaOtLdOhugBJF6QOHMpGu2x7JtUPtutNb06zffdrNFyfZYyC
mF10Xs/NsQ+JiXaOtdKib2bYjk8xx4/7ImRTtCQ1gpFMCQ2BD9iZy3yAK6dXS087
68BfdqgtaFhWNRtLmByBEGM4x5V7uiGJMg2pE3ApnwgvdszjIt3uGlfaSkO19gsQ
W4uJ6teg55JwV6wAN2KShCoY5VqodbClbvSdWaRXH5/3YpvqQuEVXyAcq+y4heZz
1FsI4WBknocUyqgMa21PTNt7b8TVebPfSkozUh7q15HeYY472HVxP4Ck1vjiVJ/Z
Ad6hU4dnVApAGrQzEgna5j40ocfqGErr5c/D5bVLebFSidJ7vkUb8+QvCJVhoPm1
KWIeocGzzd6unljG6ZgwilxiZ44dJ+A9F+4Zg3l94HKvcBkX38++ucOxLnex1OvZ
lqrUzRdQREpcA4m3LW/yhDqVmxXh0wvVdU8pN2RJRuaUUsOj59JRUmQ8Ib2TyuhT
0saF0LXW93iZoDjQ/jOROc6idjZdYt6yMTeimmPXJtLT3dcdGETT/Uxqia9wWGhr
Gudx2ia96vpFwl2TBoDciKlz4N14mSx+Fsp3Ru0IObIdqioFVdDjAKNUB4TL3HQh
Mnro4gDBtBz2G9iF7bGo22MOOEQjnqHNba66tmTneKNojoLM3EUiQqihPa7yHRzT
WOLeIqbv+5nwYFTF40xu0vLv2Sp3DOi4OoTDxTrm40bgwsv0BhoHrqDdAEV1NnAy
oxyKK3Sc8KpOGE01+sdnbFSXrxBvZDCk3k+9SrksLnG7ZqsbxvJLXjyXFoyRSobm
fE04g7LXrjBC2TQCD9RddSIcWiy2jEylUnkt//nLHyh5AWHIFPCC24CzKrxIILtK
2lEmYnmy6EvJPQsXEcQlI7gd4UxLpctiM6s+dtmpbguV+Ycjv8fAhmLMKpg0BX2H
WOkmsk7tIAuUHd6H5Jb7LmSUAbOrh68hrr6vLlgtdzXnYW4wjFP5eCppfRbhxk0E
yf240twxpDdYC4fYq2IfWqcpAOtDEzuzpfvTihR4sPUKrTeKSEByhXfb5RsNYJcz
J5hlrxmx5fKDep5l48JDnSvEnyOJHXDj0+98Yu1Nj1w9SeIQ4MVPHwgMSE+1WOX5
qkl8UK3/NrfDE1WsUeuqsDUo+Pr0GNmfV0vpIrdzZNqdZg6yqjfMFwS7HGMVhEOw
BfpMU5QXsw/aom1rCj7dBNl63dpxMCjBGpH8E9TcbwqvR0bAWKge4yI4R4XwlFox
hyHTM/KscPvQXkDQexJ2JT1yIT0NspswjEQ5900PGR4xP32cZjV6dqEEnUZxh6I/
4/7gys7Y/f43r2aP0NKcj8j/nm1sQ0ezE2d/2K3rWHkyhvOWzTrSPSatAx+f9Cc3
6hO3zstm/P+5ItDdxCzZQ/FMpK+InTyecgXAm5V6ZW34XRU5Ryl8cnGcpXXCq0Wy
3hthURX4saZnDhLvMR00UmvZmGt9wGY0fkJWHgUMSEG/mELGulu6CwPRd3bIX1y+
zXJoivPhFMWrYthcYfS+3mXs5CNd4BwkqHJliimfyZ6C+f9vBudMPMG/vhBAyzTM
AoVAu+sW2GR2mMZ/SGBAG+pK05Q9FsYqBKxtun13D8X1eUqfYqUSR/h9nrFhtMjj
3WR3Othrcv+7bkI21hFgn9tg+/sS9McQowA/M+oSmOWIDpmzS4uDbButbWL7NWw3
0bbWR/ZbYO1Gr+bBLOXiM9opTt/EmKgVrWy373RxCMmF5e6Ti/6rqafF9GUnaKp2
LrbCMPrSFgtYYUT5/DC1G+B0F5f0GteVT8i0m+BKC0WHUowAhtoyely9DoTCpZdS
UpLk7xIXEGr4DuoxydqeXMnN9wjlNsSmpXpdo/pbl4xgkaGmhLKzOUgmWrjnsckI
IqlEUD8T1c5ivR2vlVl+G6SIuf+04YVjx6jtPqBUV+ACekvlgIi9Mcez4B+YT5gA
2HvSVc0JX6rcn7Q/FxWMk90Ho7J20jbcL2E/2HT+JQTy7iawMHxfLGK6w2YMUZsz
OC/IMqNhpZ6QRsesa6fGjhWQocPdmisE8TS7acmJTCQUv8oS0rlYA0Fmou1XgPIm
fEm7X8QCr4Q7DpDZaYTtmVTIyOqxOuJ2L5weliNVC7M30gYBZRTsMkyf8+Hhwv7e
Mh+mdlX1rqhwCXsjT2yFX7TS6lYtJoeTqGI2jevLHNoTzNRmW5i2mLbeV4xQwYfP
eYhXjk+7pSj0pL69dlNcEl3xDNMi5e833vs5cIZD2EPkgzUrvIHswLUl4tIzjpo+
c4CHRH9lLhXPWh3llwO2FIRpXVNYRP+8bQu94qYDoHP/iwLneSSADmLIzkxrvfRd
PpefFnmTXJXxtMG0oKxVD7MKsuRzTNwdzaIdNxbjMr4zTdpHVI14UfsX89s0YuuY
fU/w/lXM95x5RqI/5o8Wb507GWQu9k3S38qLse4bQW4J52jFenTCoCUpWuR+z6/r
W/WzLthxQoPFxL8kBQxOKhk/tATDqUtZh255Ys9HCoa/l3qgFjngxngfNSmruVjY
Qq+yD1sVeJBEVbLEiKYeTVfheBOsggUZWPcONrNk/+cI86i+4/1eWmaH0lwMVrtv
sHvGenUWri8FGlN4KGITLAsvwD5gYoC0zrGk241fM1q+kys+nEhTtrfo3+N5M0My
9vGGju1HcUsv4iAZLwkk0B65p9S8xDyCVf5LS8JeNoMDopJlKx5N4zmTXKH2cs/c
oAeMeIoQ+zemPgxCj8eYmUneylWDGiN37+OtLZAABT1h5ZjT3FdZugtY1B+5MOIG
sV8RYsDYcch2LsqP2BarxT7t/FCcU6f8YyYhWo32ZlUm+nOYJlfANBXM/a+IXKxo
u8tf7Kus7CAvRSYAbHP1bF4DdSTlLIKbwV5ntC1RRsN1hsO97R3N2x6Tc4vOJ7Ru
c/Ea7qykw6IXArc2KFrxSkcQ3FM7q6qHg2vaqgcxBRMrinUB7N4WwNLT37os1OpN
WyFLBbDBiG1Z/YhPyTCAqn4gd+xB27+ZXQx6D8eNS+r7/+XgOCQfl9T55QuYKepP
7gNyuxngou5oKHgLZlZcN0B7K671zvoHCmRzJEiqp+JIM4qM1F1qI/AYeqBmK+Mm
DG6zFkWQovQjlpi+tRgqFNMOePqhTXBzHykibsV6NwOWF+BqF6x6VFHQ3jrMevRg
24/8V6W02zfuZquC6iPgaviCoAcfWv/GCjpbFOktgl1+U+9f4gZRJIq5Rx+9QxZQ
ZxFdtbnjNQPBv9HVnr7/lCv699rvZ2PUU87zEExqxon5OkbS4HTP1T9keRanBrbH
cg29x5E/9BWBuff7YOaj8nx1dOGy/i+j9QA969Uul3fLtRF05CXR5xUiOdQ23Vve
YgB+LInM93rGgtl3OVQDODEBkAbG7GKSgr8Suk9vETL6Iqc/nGXvXrKM7EmZP8/U
RNqPCZiAhJkqhMFB4vgUxUBBvNGT4luhzDWg/MzwKZGMYK1K9EHYmXwz2Di7f/GM
tZFIuQMUTOwjY4vc9uY5G325sh1Y+t6fSylgkBEhY4/5jQE0Qlzx/rQKBQbXJiTM
9mo7NCsjVOXegH94Kk8ej6xVkVJQeYnHnzua9ac2xSX/h64fF4eENG6g7O7K9yiy
xTU9cuA9K8olslzTtTJQFAj3cqCnYovLx1Lr1aFV8uqSshe62YDcG6yIT/mGKE4n
lH4h1SDfIYmeyBSPQo/C0x5Xu+iofNebK3Pc88nGbRp8iux1xyLnmrcm0thyeRZn
Sn0SWBRSFlo4lWh5ua49HIhasQ0vjN9UckZ5rWnxLeTpF74Q1GnK1pWQgbKfrmc4
qcFREONvHMc1WkJ7JhM1ISNkl2e7+xzQZSnmg384zxW0TkPhp1TSN5Nbe3LBbG31
oSqmrN1cppk0tCKE9CrzbOAcaTMkmUstQV+nUCiFK0vn9k8pVhW69gHOoRY14BhV
vH9B/eVOucOfqdJB178tiaASJ7wfTqSkXfs61t3SgkgkOltC6MhAVI7G++pzfSU5
Rx4l8b1r7+Y6IS+9zOy71pTpUZpsnxC30zlaxp85xb6HKXZ3nyjLNtvfmpf2FjXl
7tq0EkwdVOyBl7fGjUB/x/CUi8lpEW7IZVmEKvo7/uPzmtf+AhM7CqaiEvPoUZ/1
E6H6H60GOuJqENf8fahWo3U58yDN7zYQ8jldum375HBa1KNEcSuvLhA57vAlRkaW
7zliU3rAzdumLydSYuOOfqPMZKkXMhVAM8FQh43fiOuO9iyH2F061WKCeuNXoSCO
8zfEftwTcKQehNDdPDVA14FYzzxmJ3JnCh7Vas3jxWTeLAAK9MYBVKsKclCR+bVU
kjtnyd9JxPaD+Qll4UynsGxWfX+ey5h6l0egVakSrB1HYe9/9/ma+xUpzZXW+aQg
pjPCjbo2UWMQSanBCX2tmDb4lv/MO45LoNam6dwUdhCqOok6rX6YRq5L7/b+EuvK
OC0mkq+pJG3MMSxGiv716IoU/dkFDCM0lM4a15K4YO0B/nTpi3xsxbgWZoQKSlRr
6wp2Adg9zA3WUofAdjcvAJMr5WdjUGuI3eUrzd0iqOhVy3LR2vEvN/Eeha85Khg1
nlgdYK+hqq51C+RQfLFMkBqB2++sQBZLcKErC9XY7rXBDGdK+krjfuewWVSqPccO
qWX1EK3Kzt+HNT4NxsqSZTmbolL632CTVdNcfEp/wV9m02xo4IIftaVnm1KTlfs1
YlN6olfo7+2XBeWRl87/+umj73BP8YKYW7r35lNwPafS0MBjcpZTh7K9NxlkZJl3
0VyGRd0+naVcpUiZXvACkpF8pZAL/iN1l6l+skH6sn2iny9W0lYlre+TIyUVHp9H
jfiq3vYFOKDpkWqMv7QS2gX0C8CXyPM4GA33CSpC+B8MZwccXKQUbDZ42yUhrGW6
eAF9AVVNkQLPzJl6x03AeKvINvFJyj/KLb3OzjZCg4GUu4H8/gVKw6SRstSeiWrz
FODfjWjDd4CR1fnbnPbuMj215dldd78uLRdXNEHiL7fIZ5tWfRPExUWBDVk2UlTG
u6cKfFjW79XPzR9j/acRsbR1OkkvNG4kRING9Rx6IPuUZ6sPWN9iQU3By8/bbt2M
qaO5nqmh1N435IRJEEoQmm1X5uI2eu0tTjiBVR4i+ru7LtcC3rhRU8jHvD1a/YiE
AHusYI8/NoqrRvWavKH3MHPvas+z9sgEpyq+f0HcOhUElqU+PY/bwwv1hWjY2Tfb
HgzJvmnyCGkAxl+u8KwUhPWURaJ2TrxwsmZvh3FLEosf4T+avEFZ3B/e7jKlOgkK
4IF54mPFH2zQVJp5hgNml4nzTR9aly6fo6d7Y42jauVT83ounUqAchcJ+ikmAMXb
eZctIRIb9PTtiRMcVBjQEHvBAkfgYIpIAX8cb8wyMKbwbZlpErJBhbB32lQXjX+r
19l0GGvQjg3LU10Y0o2ahuozGnP/YBGy0Y9DAP1a5uYq8Kvnyx5b61Yo2O6q8azV
ROY1vOO52ud6aZjOl5tQeML1coupKUIbrNkWV4+7vcx5Ghplb5abMoaDfJlQ2HwW
2DvX0GmWPaLX+Jgo137/zxb/gZdczgx53UgsfF3oeQ4CEVmVTf4uFzIUd3Q90PtX
8Z3PCbwHozq2aut18khAWROTw/ROuRb6Ak8viJpEPDCqebanzvO+RILxdxSBWi5+
2dBc6gQr4mQ+CR6rxp2FYwX3avO8QhVpvPZWgBxoM0vIVtouf4LBikg3MAovgyoA
UWuUX9sJhDACdmDKM9ZEkCyWJ3WqAaHAusZXFZB/m6XRQhqH/SUYePvpr2mhRZXS
0FLldWj9fZWX4gF+UB4gH+avNMtXdE++iZl7WkQVev4V5zalpUHvXvejnbCeEW+b
e8yYorIUaYjn+uexHB3pt+mfJJXcN+m7kvC7ulDt8EFXw5eoSBEHJ+meAmppQdms
f9RNbsNziDGgEMUGYZQlK043wAOjDTmSwUcC6HLfrIuQaECKUwMegRRElWk3s0Y+
xxvnAUmyEXgspTSyLiiSZgR/8AlnBXmKShqbfBU2hKUC9dfdEWP6sTiNCX6PSPrh
3qiZsX2B6oVsUFa+c8aOqsMSW/OlmlSXCBO63G8Nu17wKSrR3ATV0Ersk77EMYaI
ZFEtnh/+ELOsR0WxPXWjomHQ3WjgFjWf6B/mnl7VACpfvImj7KFR3lRxBVO9cm++
dF8ZOo+QHmUjIFpZkVktaHoUhungp5xMuw8A+rEnaxuEVtJacXvXhVTsFkB9rryA
EGHrPHT+DswmJOcl/De8ohdchbiBlzI59iSmF/UGnBpVptTHpMwNaaw3DOQ/aO0y
y1G6GN1sZpe0YujLMMnMdGOif/Na4KDJN3FRZJ100bHHK4N/ZLwltI/YFfcRCibO
YNUnmy0izgRzXbei8lvqCaR4HSuPFTlgN+rpWqwcH7khWpw+nWi7wToBDTka9afB
91cr0KMehlPIu1FOl0G4sNM9zidGXOdcjTC9jR4RLwUm6Ic4eT4v7Ta2eLRTaRw6
HdFAUBJ4wVVobXQ2lZ94iJKkil65eQjUsj0o0CsPuOA+AtZhPIlEqoWRfjeulF+r
nWqAwt+rNzoDjXFekr/LfB9sM6vtkq5CCv9uz/Dk4oyJKWYqhIbXcIYd/rXMMYy/
Psfyyh/oJwpjjxV3zj+9fWy9Z5JYmK+yKKWOkIo2/ec54xH9/tMpv/4KoVP6GVqx
w10wIeZ+ypNmSn9FaoxigcFpPqJQAiDZxxIjc2dVFQbZ0XQjtmaY3YdJnLRd1ogT
/tWOqgL2hRHQjRA0LPEFyo08kV1M9q2CyrgzASh5xt5sS1ssrtD20sNJJ/xncxfY
0/5hVPoAxjhJOZG8Cgf506p5uToXD2hyVI/ejmYtuOF6pLUjPS3nfJ984JKEjDvd
lZYIilzW3xgkXbfTxsEQ/Ugo8k/s6JY8uCloAT6oRkS02+vGoCsUpo238bJM3w9R
4nmiM/l5j94acdZ1mq8MArt4ydDHEyZosqyUXM9a9wz/u36Yc/ERTWN/htvAUv7f
11rn3U2+BaSRRXQeywkSvBk5t/37S2BPBs/4q+bCf9G52qSzh8jA7DY0gBtoCf2z
AsjdJgupeok4ngmeEcgZS1k+simo9NPlNrHEzOBssbXbcTopXWqX/lHTwHWFm9Bt
93cd1SaHrmOuPw6at9OHm+iZCSvC96UnwcoJFa4TsNAHH69YaO2+gYWz2cZGPWlm
8BdtS0D+rmW7/8XDWxvNz+VmJZ9dAO04haoAXtc2hq9otMpDjhF3a31civvCDhHt
IaZ5DGj1jCc4B+RBohnG+Bad5Yzr4lV6X0AJhP7OBZXRiYeJTi1wYbFzOI5g2XFj
7cwasc0ckbrRem6GhVz858Sf8gQ5w4Xk5DCzYamOR3kuJnfKDdrBQLdh/w9LlEeh
SdRwYx+MrSQ1pqRVJzsF/IQaC0pzmEnv36Z7UqfRzgKphSfHNKidGZxMxtPgPHr3
IgQjBQ05pfe5RYmqcK+LvcUGHG4vBBpHfwgg9MOIH21ZgXmxMSICcciwveW0+UD8
iCamnFxjYkkd5Wp1HCvI9oC+p0QS/HAVtsY0laFIVsAQRk+X/ECKe43XyJAD0V2T
5Xi4EXHaF2Ev0HTiSZFgMva6Fjk7LKueevjsvHEi+gWHXpXM209RwvtlM7qghDQ+
I72AM3jcGMjaAHLtjrNyx1nVIFtibTh6z3pGn5SbVS9BeqL5UULHk8kZohp4DGVN
aKYjbvPSzDQ/hfrWwsKiwBJ/viODzLhM3LZMXVX1x2sOd3oCdBBlgxUc2xhHYcjM
YCRL5qKcXURVUxfDHCxcpEMrJf7ZrIt4n0ahHsDHhYFmpLeYYaASnYos2IkHQeaL
HvRTaAU199UF7I9pRHlnfebB5v91viACFkDaSxZo4DfRFlLwbPLc3bsxINx6rOkj
puYAsgjUl3yNQDqezXJtUby93Dn4FJpsbIzzesGcIeYvyK3R6h+95X/3e3FACoft
8SjHPLvRM2DeKnGmWS03Cu0biAFKz7NIUam+6WbzhA/2reep8kSDPyw2xPe0DVSq
ga/QRAqj9eCVht6QEE+TZzWIkDmsatc73XfBDeScEIVqWinNmVlAvWbC6PAp0MRt
kdwu3KPf3RRJ7FkxjDzk+xBLxSvwoi3TthM80M0D0gR9vhTgeSHQNWfZCn6HGX5a
ptjiICXMfQu8YMy8HjZRvgMURPCPFPJHlKjk0+N6juZ7FzBpgHGo1YiPXSz7AXvG
9cueNHp0UyzAux2bvNyxrIAZXYe9FNRoBLfuMJbaCCWgj7rjPwgf2aQZlYwdngWG
haCqn2zV3Ux29Vjs9YxddtjuHUDllc4MnraRzWk9k4zaxZ39mEkVzoJPZ8Rnn7GI
dGLTkW6oObH9gTBQtOFXmuLn87omJA7zakGtoglsBANS2abvICPOOcjotmpXIQaw
4O28VAjHDp86O4TXaUu7bN6UZM9TayMTWJD7HCZGzsET0zSnEVPdD5+C5lSbyCCC
dRC+mLxmuK6+z4/rnMgUQSBObmeseuPC3AU6vABpYlEn/mFNTewv7MytbkhA10qd
XbWNZQtRJ598Ii591rCVgdGCb/mk6tDqaWjR3bNWBZd2agUChtv0zD2rU5+oOEVO
PV5s2rt6UF0Zr3l6BsZuRLWD7Ju6sxP/5lSILVZ/lOz/Lg8+qNPMdoCoSt1N+Lp4
AsYjQ9J1FFv861NwbNLl4Q9Y5AO1DY8Iy3lBQsAE+t5X8okVjNcWAkzWuyQd7y0i
BdEtEeEMTtewBTKJ8SAnC5LUFomTpXkwHNA1WflQqtMO+h/YdF+bz6/iW6pFadLW
Xa5mjrhDQiX+cELmXEnX1i07KGpa2l+YtJ8H6WlYshgXGVlZadoToYOFDku6SZcp
bRPvh7ed5fmzepGPbFojzn8ZpbaAByh5PtyNq6t8lFnPY8AYWglQbDz4hTGi18ew
oXj886De2X1d5eGd5bQIZwjPTsPxmXEknQR+YOU8wljSCXN3pubTSZj7a9exvMzj
RIM5Xu0TcXdFAiZyTxsw5kKdhezjyBUiZQm2HaZcZd6D10uk6RCnl5D+LV6/v9KZ
JIEKo7jzVX++2ML0m8XYuuE4JBFD0Id7xACvkfrDEP1CRTKRxkgL/N8ZjYk0HpM9
HV2ljaWDz0kX3K6sXI9e7jZPZjnkwDi0ko/6BH0oeL3BUAg2EtGY/bH8YqMmUYCq
yzEkrCTsqssnucEAUOTk1YVF3Z0j/brNrJ9usUqDux+lru3btLE5NF9vT5ZI811n
r/lTk/nWR/ztpKWyAieJZ7KWaymOTKf8vP+B6au4cJ5ax10bzfPcVq4XgtpTgvFH
tScyn51znuJG5Ve1+LCIszhvjzGxw1C80MydsX2DTYoPJEXytmboZWgKA6cUz2rC
782x5J/x0nwO9nxm50ShGJZQX5MQ+Nk687f+UStn9r5nPJJIuVQGUThuqIK2a3N4
U4dvrKl5fe/vY14i8UQOm3B317QZDkziMizVtS18ZUvchpAfT3nReTvW1SMsG9hf
h5myG7agjvkPkf46aVPwTOl0T3dzyOkk74rOiljrtJ8wSke1KjZG6U/oGZ6qwwoU
Hw2GQXQAM2Ksh/dxNyxyyBVFRyE5EJcifETO5PjjYqQGmE2U5kbUcH0eYMlpzc5T
OXC088HlKZlhGVGam0qsZoMQgRrCrPtU1y5WjE+/0eWZJH97euGoxs73uPNilD+V
rQqMRFaFTpyW6Iw0+qHjszEPLGYXNo0aVMTDiED438D0g73LU5LKcPCM4oeRbUht
khGxAQY+RNJAz5Vzq77ywL3U+RAHxEYcK0MJAXl61LtMbCJsah/vAevtcCMilehJ
QuuKU/I65kLX/ApXUEa1w45HXnMiEaumss6q0e+ByX5hVKK49WM+sgc0gl5rz7zA
kBT2o2pGjawokGECc/SL+EZ9Umw2Mh9KSI2XTG7MeOfKlv6r7iJp+++UuJflu6ti
qTgiNAFn3HYvQZ7b9yNZnoqeW6iFPnvyuGaGfFAusDWZDQedTdYukxuaIEb2kdtd
vJ60hLxP5T9NY1Du8A/amv0N3rPLneshHk7GXR87K7Ht4oi9yrKHibu3s8I8WQTF
FxNWm2QyYLddO71v/yq7oXkOG2qpeoPztUukARyP1Pz5I9RwOEzJXHlE9+irHZab
OHdpjMpXrjBJvCcpQd0MiO8TDw2ZqmjLn9iS2eon44Mv3t7JLZYCn3pLjSqNgqOa
HHe4DxqpaIrxyeVm5nIG9+skxjMZjGraFh1jTdwvHXs46eKA+/5WyxWl7cQfD6fC
5/bxGKIzWarjP8lfxRd0JY4bfeLPx67onDas84cSnwa0hVgFd9XclUbbcGMiF2Xp
tmTXle28r7D830MIKSEkHb/8VlQnKIYRQpkk0rTqWwPvDUseM/Vyixz1Z/x6NjYm
iuDOt0yJQZR9PMkS0PHNtpVsV3b0ZUCwKVi18Ke67jPVDzHW7blfYcDwwJpl0Tkh
ooSC69Db5f1sf/rgOYv4zWeiCUcExb/oQ6EB9JxeMkwgqtqjPYXkwng/mVZ5fpHi
l6c+SoH+51i401K0f+VYePIE44yYEw+X3CSzuB3qtDuIYkWoNEvaHLGwqIHJ7JOJ
zAKFhTzwG8V9xtL2lhEgJvIIB/tUXDGwrOqu5sveT2z+eQuSK7vY2fv3UgcqAZLm
nOjjhuc0otnEwpkGm/rl9ktTUywA2pPv8hLwmdV/bbKtJUTuyu4emaUZFC9jp3Ds
QnwvBoia+FQ1GJKLCIotQkMsJCBg8UUD2ZgiDaEjDKjjJTFNA8tGcy16vXMZ62mJ
ad1pBygOvqNYrhCYGnqVTB1j86M46301KwYfITb8c6yt5jNsNtEjzO0eBu16WwDI
uhBPb1Dk1Tk1zgpkibJ6dSh8388k6GYltqvj3kOi1dqWOHCDio/MbJJRN8D6vx3I
rxkVDSfW8rgNUOkrq2PefvgFh6Krfs8o6OC/NWYFreAL2eJeur9Hc8gBKjP3JErs
2AcAjrm9PqynygR6yeQuJoePAB7BooXe+3SolV8rK8PlAgYHjArOe1cnvm7dMzF1
yhnzPCtQ5hc1bdX+gXC3USRJsz85Tp/AiYTiZD4mT2DtlukS87L+jbHPIvrYfEGA
ax2DVnJn98LEPZLcEuEpXoPCddshRbl3vNV7r0VB6ZCDINxwR3A0L6eeJJoS5xVN
UkG8FJ5i6NgVUJZcKSfqb8L6myAI6k+SPz3CL8oH14Hk2FkFVSjR5x5VevUZowpd
i3AHV1z+AFq5El6yT1NvmU164uhaXB/kFfag5DqaJOLiaO04m/TvGvVdH0qH3Psp
WAJJq0AW6tOut3J0p16yhCVPBoEBA2DNJbf6hFPjoPGIKIvQrnHFqwVs50iLV1ny
fLIiWRm0hMoIIHzaITi+YAUskRb9VXHaB5F1WH7nf1NpRQZ00A/EpdbNE/Vyq2cQ
5tYafKYGN1X4Blyb7ChhQDnUeGmyYbJNh/TXJ2CXGNIJ4NKi5Z/VrF9JBap1jBy7
+UEtrtfQXM57RnKmUDDGicXX/ss0kiGP9EviWd4l20TUvivzoEXXDIP6PTGOAXrG
n8LfLeaKruCD9QkqooIj3pn3BwH8xqjoX0HCmLSSFiXew2/8xDIQV4xy1uarTskJ
QkWuX0NWFNcyL+Dg/qBnEynqLiWuZvjvv2jX9MMwi+3qUSOX/UiICXLWaJd5Zj5F
8D4k1znz3EGEb+G1xp7ew+HY16gxbVK+Rckc9XajchvBRg+GweTtPmZ+2lZ3wyeu
7gdx/FEtUL0z2jize1jYq1KEufve4qK4RONJEwdxlwXGLNRVPXaiGodopG4h6a+k
ei6Ye1oVVAWNkpEuAC2A3ChcTE+1YHAlR/KyI1z9CqSPwsdQHYlNg5MYi+APtBDs
EgEmhyxQySTC4OXo5c/CVxgGUVEt95pWL2Q0Ba0Sqen3aonOUIscMyVi98acuVTG
QEcvj7JjNXd/Sfp91mH8zrkBQ20U/qHoUUcNKy667e6yXh4Luuyhs6r5RvvM7B1f
9iO8wAHbDbJ9Bw7n6Dc40H/pXZYFrSsV9CxHEmWrWQm0K9Wbu+fHSzyTHHwifJ4z
4+VMlXchQrjFwt1IjHzCbzN8xRW+FZu3KJ6BCqyPwUSsj8LbkraPtchauwBcisP+
qTpWF2o1Jc9+OycTlw8/OQaXMjGcDVoBjlcI0F6xpVPToZW2JE/AD5Gha4lAhde9
uSH19cSyGAG7zfqByH7J/l3bRq7qHxhl7hpNuzoiuaJ5R4jYg+CDKWnXIDd86+dn
gslJ5vUM2pZF8RF2MwdBO5bRxBkbD2uT+Ugk3ow76z6dGlulFa5pyLc7rQInt4JZ
0ZD1qkrii7wtv/yInq9UEWOtTPo7sfh0t0eUiGB0SZKvrwu1skkvSHMsMzSv1IBm
gVhXoDMawGXX38CnMxL+7/Mdqx9KibynMEMzmzezIDKzJhfMWk6unu+MgG6aMJ+E
a81gZ4gLc17Hg+Coi+v11qdLP4cSX9csCaCxxhTOc2SGhiianPlCoIITtMwRvkO7
WaLwyai5WrhAnDQ3QOIxCE61rJHld4mqz3qYmjZJ/LrfXv9VbJEx1LL7Qpdezk67
wrhkQPqIwTe8VHPlBszfuZNJmU1n6BkXQoVqo+J1e9p0+EwzURycRb7KlnomKxpH
jaxXyq/FQxmv9dlbtwh7rufHxqUgBR0cdMCQRinKsoZxGVagFamwUZa/sKXCeHrw
m2jQ9vnMXv7UZmmFe4SeBviVwUQiiUK3Q9Rk/OPDkzPQyTkl4/U6BkONaUGnoyYG
3/QgRhuWiZOxi+RhN+5hx0EGJG2fh30ep1z+qD8ilyd5DmN6JJQ4T2bZF/ME1Ltc
l4YIK+E8uW++DDi1iv7YebyAJ4Mq0APq4fEQYiy5eAS7gQ4gS6UWJodP6fQrbpKQ
CtOVd31FVynjPgY/05ioF3w0iWs+LYUDWU+uQD4AtI0kyGb+bV82+UbG9fNu0A5M
iU/47IqbT0R4TCiL6JcLFBrDLOLAGgxzZdGMkVqvujQSRcUsRBm1pBqtrqdWuRGv
nNHLxCGO5iLpJV0x4FZ0t38Va1HuTWjhf5qnsQofSEp76k1bfVdE5yq3BZG2JXqt
aogCqPPgldlso+N8f0x2ysW0maO3Ef1i3pVlbKxblHlvIkHiQjNVZiIMM+T0pn84
OmAMa64eio9pXgzoflbN2Xy35bnZomVRFWcH9HGpdcP5e2t632pwxoDIM7ayVuQq
RgYOE4eOgDxc+2R9SqXSDydfsi0f5xth/b8vP+3YVhGjt4U4g70V+3JciWVFUyH5
UgEp4xftJKWi7WhoD1juY+TFKE3RNwqVcBxE7pwwGiwwAToeHXoAakqQqzEiTs9f
ubonuS0UC3Pt+R2E704eDhaOrvns6us3tTKL6Dlqnc/mpbuNrfecJ0a8cp481BWn
3li0sAR10xwgQ508WtoWws3EJuIteyQT2jYxSBuW0LH3CSblsB8J48qS0vI1Rkgi
276uTjywo5ds8SkCWveHiqZZtieVg3wfSQvj+ChY3BJ6lvrcwTIx7TVKsBAQ+asu
S618zDkiAcxFU/8lPWps0kJYoyINKArvm3Srx1niJmfeGWXLqyOSEHcwzlfZTisR
p/kYgsC7dJmBRJ8u6+2Wp5sDqZh36JtQFW/npRrXFs/ee9oP2D211dwfWr7jX8aG
PDwyu+JEwrNSvABylPp2wwGVH9mLga736lmoXSxlETwBbZg7dGxtmnK9r6V3qf45
w9FkYSeHV7UtmM3tG4Os0MHg8/hkZsAyl3o6kzvZgA0+yRO1cYsNAbaZSW7Y7/Ug
aUV1Pqo+PJkEeudtF/FHXcHGOPWUN15F8OrLnVOEWgQ7mYYVh2U3y5IQEaMT5K9j
Sk7+v6l7skQtGRgoAq2KsaDyPaA8+01DKDZEFM8IR55OoDW7inmRyFQSVZA7qQ4N
yr2Aa+I0Q7acXm7GaEFf7ACBZd8u4OUyfN10iNCn/I4n8FS8947AWGgIrlL5YtRg
cClN0xmWNruopkgaHnS/wiH71Ow5YLoyLmmJIxnCE77MPjU1YNKUZI7a4fiRkPdu
DT05Kv/fOC4TTRJuDgrBAgQJBWOZpvFaHPzHX4c+uO8MgsxG/5nArVOxObLaDBvY
0acPgeuIftA4WQa0f1mf4wRYT4L/bx7yPyAaGL14563xEr5ExwKmSA80W3rJvRhB
1bqYwFJSUAJj3pl7R7+kT0TPsRoNwl2MQg/nyd0QvmH+321WXyscalTB3cfC5SuP
keqD6ra09TMNV+V7/Y8fOlzQfYQYc1KfVkuQOUT4W6AkTWeMXnESYfuuFrPcizfU
Fk4DoOSZ8Bjw1tp+58roBi2FtgR2fAARLeQ3pwMr4FiLjEQiRVD7cQlQvP8dX4Iz
pvmWueZWOONIYQ7KehoNL+HeHn8T1czWuBC48hNXqTTLgq7ah8/bemjwtx4/D8RZ
BPXCU/3Csl5zJRrIiFHTcBlwkC1inWlgjCueZyC0ENEAM5SHxCNaUD5b1eNlDeaX
mIweXiJUbSNubI84qxGXDbxiwhnAR093ivjCNbAssq4AZbp2J9vmhnSa/RQHbi+c
355ovrXcNcsFQGQNiwqDH/h1oAftjiDVMPVNQWg3xqgJMGXXeIKbYSSoN7Okb4FC
UbA3TwEA5MaV2nVZn4oWEOSfaY6zqZLzXFYd1qi4AgNIPJEPyA48UxElgRjC1w1/
xLe3nqBXkS5losmJ9R/fC2FoIsJuBBHESHAGmrvoPseLckE6RCgtha1dme+46QIm
e2MH062BKZBBJKMBiFuJZadMhWGLNUDAhtA0cuP4kRomx4ILekYDCdL8XMbHDyY3
tK345OCJvU2HBwvrVQERPBuEr3sPj0LCzVeqscVR0/s+7wr+F8s5/2gRKno6Haki
0cuDSGxAkXmegqpRBsVMEI1b8hkWBhtuigN13Cz3j5ymFgvVNNYBh5TgzGm7cKZ4
rkb/gEE4LTusQRRBJHFghi2i0UoCDSijHP+Blt9rOJxsomsDS4ByiztWvfoCQSub
/qP/az6wnG9tcMw1yfQNjemFpQlAJv1yCBBuRXi5VoeRiSc7+dPi52i3TWVjCySr
LfVk+6d4UXZ26ctR9mn4o6X6i8D5TfqGwdNAcQX/I6p3YtWRh0zKgHjUVLpADAfP
oCW7JIMmwc8kelsF0vwQBM9OI6CRh1WFsoEz8UNf/c17hWbM7Ir52Z2f6IKTIR8Y
bQuZAKZAq6akXc2YEhBui4yx582oVIc8yMu33g6U8lQ20luvbu02Er+QdHfJOgBg
aIgRrRp1wVZoqEm6FQ9ymLCD0g8pYzYQTWmx6m5bPjjFe53XnmqImwVjelKxQpzt
rbctQCARCJY7Qwy8Q03e3KOnPvkgTIlqPKbh/QCVNk+gI3pTAAfGlCQsVFqweHtj
FiPU0H9dqM2fhEq1X9hEf1bRymqOAScS4nq3oM/33j5aw6+wOIVvW4buwqOIH6BX
sAcE0v7NpLN10UE/zwZvZfznT7Hv/JYDJHrq3+F71L0YtrDoRc2ZcWfW4OwPlaUK
LIZ2s9SspSjr4BqKINRJaEIig2kvRpGb2k0r0/LzM4NI3P2PdO/sHTmQP4uyn/xS
9NuKkqo8ay91NUst6FcOL05pnoGue8ZWzGndYBf9fYPtUh/xHtDirvvTo6dT89Ud
unuABDqlHA/3r1zUvcvb2eAx9LtnRhLu9+aV85cYmCV0LBetBR/bGZ2VKY8upom2
DkFTbbwyMHxDu5v038W5hw0JeFUhYppBdX/oB59D/3N0ZUBEkNRGnOVtzksLBKcS
7hrIV4QpJey9/CoB14c+3jOn60+ab2hXQLkPP/HASssxyNyg7a4d1WQYPbrljN54
EwMtzC6ayIW1+jYKh7mA4oZPo5BgK8IkEILrhuIqwrexcjQ1vcbbcKgWbFNem4sF
e6rYRfGlTLF/0aelQQGSsfVeeQryquNPRY65cFl4PLH2IACIXFMLV3ikbea8ee+J
Dd+B1+am84E9Q4WoCf5Wy1s4Dlka4Jht8vIRiGvs1UlEstSB95BUcqoOGReTiwRg
L1YdIwkDI+X+Bw8ogz/10RidYXv+4tkqkRL2dXr6n0cTWqJw+3jQuk1B63onx7TK
7MfT9Sv+TcKXNsh8eIk2sGuDxeULzBsvMY4lK9Vxq5nEL3pbdujZS3tQ2oNGV0X+
8dSGdfwXNTrQch2eh3i6sNF5l9Ul/gLtUUyj03m0cOI/UbSHX9XlnRmydXQyMf8E
eMKYTY8Lq8cZGfwPzBWb4iKgxYyMiw3zFQdZRVZQ3+r1Tg9rnskLeJhZP9ZFjGZ/
+Fs1Bf5KyTJJpIgctQb+Xu1uNgTnhVhXChM0U3Z3ohG+8JUAm6UtxSIEVUBVMaCX
8QmvlBVcYZni7JfkoSRZfz/sI8aLh6d2FlvpfVGqZKkt/3xtJgvAcsWXYl0iCBN6
4UJlT/54g05KEXXNZNy+Q0LCnfE2oKGbXnJikhQ1prmV9W4YvXtLmgb0Y5hOmr7T
2yfjoaqPZG2wxYmK9wDRFBn7WgAkPCbQgqOGXsqBqXLsNLZSWLAgQPVnhZk/aXL7
YFN3vEYt65Cd7gRiJV8RFoHndUs1QKUwxZnnVFMtxPiv0A4Aonkpskhi8eXXVZ8u
lXKyDVCT8ZRNxf7kj3OjGL6m9NfGt0CRDkc3lgSQf91MBel7Q8vqt1XS7P5ZSNw8
dqUm9yqqMbXKh0gehF6iCuQi6LMw7GAFeIUo86PI9eRkUl69lWUEmoJaZqvFXceF
RA4c6Khzz090kENzRTP9/dMcxfKoDrytUaB+dy6axtraTb519KiySBRGmkLytxhm
lXjWwrzsKbVwtXK2ccDOWH/8Wq2vDqgRcefQEMpm1J8z31JerZejtpK1U3VKRvCX
FAlh8u3Wgrzgy+24tQ+4Rw4ZRkHHdVGr5p5jSJ70ZAxY2oT+bnLNqEy5+m8T93Yb
SpOglf7vehOXVRyNUdxdGTxATu/jwEaiTFfxa2SItmPaFvVr9czOor44RVANlMxS
0iGsB0p6eYO0BlE5i+EcTLYKukxHH4tsPIpDMMRIrU3RkjmWfzpbvkEtTA1ejz9f
+/PoV3R1N19KgmLJBOyrn8Jp8/+ie/cikLOigyxnG5uuo70lSksOGkTcl/c1r0UG
hCtNik92WaCen51nNse0Qc1Pxkp1AaJOoaiwuu3fpoYtA+IGXWFBIYc6Ed759nWb
Eq2EWe8TYfuYMRF0/BjgfY9Yg7tahfNuBLweaXDEYaO2TmxMfiXHFdhQ7JDQVFiX
7ZpDftqng0jRhfQzt9AmhYjAMeWVECS7GrhE8hVUWXqNADXfF+DHGgZ1ddE+snjo
FdUUqOsZL9/kY4En3jYVWx1Wlbs5/+Ep146nDyGtjauAKOkp/cZ78A9e+Ai2isLA
HGP5nncBFO1wBIh5KT7upB1k6n+n36EIF/CxehudW7uSsMGaLJHTErP29asLJof6
lcimwRtPqv8mzwwh/Wky+AAeyUUqT7ntarGiAUhgx2eEcdpmlfZP8vKG1FLGonnX
CarP85lLi2mXEU/WPiJyIIiVs37tmoEDF8Tw01je4sbKM/BFnhDH2XDKDcJdC+HU
bhY2O89lIGW6PAjbOvmaFLOYDA81oZyMZhdikR+eMlPGfH3eNsxKiwazuetV4xpv
aIvigyi3yXPmNrC93s9FHnNiYrhPegzfhIdjN/pxrLQ2eieDcq/AK8N4o8gkt50s
BcqzPyEBQsTkjJopbh0hxXVKlz1vfkIsB8VwcUChAHBeVHD+lpszZ4TAJNOJ/sHB
iGxWZdZVN8c0umxayrho70NBrUJF5AimFo7ah9PKB1PJdoCcKA+q9Rhy6xFT9G13
39C9YBKVJn8+LBWm8kxrIyIzRxH2HopdmmipzlF1lq1GGSi6MfUmaLE3p/n+4ieH
sV9TKOn+DLxwrzlFMfJ/qr8ad+d1y2cdoZxr+2RTqgovejHpeDsp/yHYEEb+ApA7
SzZd5IsJTHD+fAoWVeTN4qGQ8yS/Kui+p5BH57BZK1TzW/8jAE0ixx7J+smrOqrs
b6U9g5dTjyVKgG+pvgPYdp+mYsz7nYNhRMfWVm3c+xwXAmhdueR/fn2bEPeIC4eW
dr7tB5fNGjYwBjMEz6UyLbufK93tHY5l+4EzoXHFZwJu5W46jeOCBIJGO1ptqehg
gvc9QvPXith32+OIwseIzM6/YpgwetCqhi1CM2+RDlNfwCaeHeGPNSz/JiewrgED
PMxr3Wx3VNG0vOg+LOgnNZTuBGFs4SxAulV5oCESJoF9UmH1Ht8q3eOOwZhBY3zn
MRyV2nMNLJHDQFszFh25zktU1EvqxWoaaECWhWkHCQwZyH/kpKWN0DdZj0BUYkfP
VYpsIOuFrfyUKKYjQPtarP3mO+q5osqpZFRiGnn4+0CfXeJjy98nb2VId6apcXAx
I7T8gJfVmZ9TCJQHrGcK0a6TUdL/+wUmDq3Q9/eVrk7DRJLMK9UTcB7nBgnNOrl2
tC6nmz8+xVPxB+Q4oaGXjO1t8FCoE0A8Icv3sKG8296cj21GSrxhjPRf79erK69Q
WtrnlluOm9lM3SKRMckjTmdXce2wv2Fon+NPab+OxVVEYw25PtVMwNlG3izm6jJx
ahWhnej3mCQiWMUeuWaMQIMTyuy1IEd3rMNZQZPzM6m0jf2ChPQk7ExIY7zpacLN
weTkW9lxMzC65Sm459wL6IB3LCiP0sVhYgt7WnLmJovMU2k28cczIdoLvt1v5OIY
KunxUoGXIcbpXgxJfrCBsDgBeGqVhWtRxBQxVvEJJ7+z02XqUPrRhmMQRJjPmiWN
7g1LJhiUClOw5Vl5DRiNzOvZOwUlgvpDTKEmXtk8FGKEdq5u4C3vXA52jagkM/jG
ZvvjbubUZ1HZXR96CUsQM2+nluNl34WEjLpCCMxEZQ56r5fNkU5gLlO6n32bT6hL
pRZ7vF5nv0rhPVn1saAI3usCXK2yEl9AVk7vkY4cAEQNTiAi506MUPhQGr4AmSRY
oTgxTqlW8C03977eTqBZVV6kcGHx+TnJNM/6ExidmftWnIcMwahVGRlIj8+VAE1V
TpqbuOFVCDRPklr66eSavOfYZ0xJIqSWNgil7ZdpQosm6+1QPD1rZtIJrH95KimI
iqU2zxRkKcUrmVTOcw4EMNSj9U8kJ68F6BXQ92EeWMb8FaV1IaPIG7B8ERu0teVb
7vQKPrMbZsSU9RIUdk8jojDo0td6lAmtSAxtQHmEIPC/0JnrbEZWWunX5kG42yJo
eqNP/GwKSxHRNHJU7wW3SNeq7j22aYLXxDoDrwSnbX5tM5Xx1TGCaDfpaRbTIJJj
Ht8QuqT/wCBsPN4TvBPtwPHyYbPDZrUsT8UNOx325f3Sfz8EZyS1v30SJaFrBtIY
UGdth2EruuPCegx2uSY5aZB9cMwTQSCUNTFJ8PZ9on23s73ohQoUvdIJa/DoRQm0
bRFdoHcNxxIb+gN2oWv0OtIJtuq+mrSqkzelNAvb5fqXumOksuPkznHaew+sCvqb
JExtXvjeyIcHCW5c2HtI6+srzqTw/iPZW4yGs5dXL5w3FRgkrL8P/2DKGd8E4QSX
iJT7DDO6vPVsLZ4UkVWtY+BPtG9DTtClwCTB2SjHu9q7wttBXQkg8PMHoNabeHlB
864cn+wobjdYRTYEEU8mqywlebK8BxBIPdeWp81vhPgNWRg+Qt/ikBAH5d9/GFxV
4T9Kq+UxpNYnMTXyNzrkKCzVy1F8NQdwJhlhro6kNubJqA0yYKt7giFXrKWP1PZy
EpNpollLwzB5dskWteg68cQo70D5eDhjfztz0yucorYBK1vZydM52j+Oc/b9eFn0
CYwODix+a8OR0GFwAShX3DYYdx7EGymrCvurvwQDLFq8nHjQ7yPje8MtaBaf9jj8
F5vu/kzKfjWw5Ga6mr5q5NvNsa4tgNWGHkhZklBLbIYG/mkXlc/Lm2/1foWbEk2D
LwckUlO6b1gwFS3WlSRHumkVdN6Rg3/Vlq/oKM6akCJetZMIER2rY3vTgpz/WJp3
tCfd37EEgDh7Q8oTgCz8AsQFYJxae0kjTL1qWpWRCoopwyd/3Qa4cz5o2ipiq8Nz
N9t8MspfMr55LZ9FrSjD0X2mGN5tWLXPMiu6QdfI6FIjfNNpmICBXyTCfYclw9Wo
Cgn68xbhTaI07JYK6hf6MNJCIivAnZ3gGKnR8O8v779AS7jYGxeY9CpLvi+Gu72i
VWWSa0gEq26Q89QRSBfEpAq3GFToVJGoriICyuGGblVtBF+Ql2cy2rKMCO1cm8Di
gyQ2ANITnWXUkdg9FU6MfOyav05McKP1nOLkP7iKqHheRpPjMe2OqJTD3oGdMODH
D3zbPzg3ccoZHi/jjFC8G0dnZ96zBY9Sw2f3ygdH+4W6axA+cqNQi3OHCQ3r++26
8AzmaG1PbENtRl5cg9VUX79UCpm6Ongd366j1tLU3fcAudC0TE0ODb9A9PQ0+2nM
Mai8S8XXbrJtSZC3T+sBt7ROJzziIlyWm1uM4vz3tZbZqIn1MMoKEx33b1qAovBc
esGa+55LVxLMo/rgLAR3+wA1A/R6Odf65FPng7YfS61B918Y/WqtPs3E8k+f7z3n
GwcVbLhV+kcfghDBAF0KhjhWtxbcjbhc/weBX6h2upH9xVL1RroXliMa8BBjWt1d
VGDisghQKs7iu2jjRhmdtcAjgKfnS/bJy9ypcWzfsAw4gIEvQj06ed5VuwZTTuIb
AdV3YypSg3rOkqvX4BNqUnpPulFF88IqHtRBJGi5HgE9Lt5rxCa+YdDds8eiT2Ld
8Cf3hy3bvLYW8srkBhtxPNF/78TKRIVTwvrRh9UsP1w/H8cczlQGquh5Du6hkpxN
RWTFWuNdLz9UpjRtxT4Hf5B4shNxBH6n6BPgswxNmBzn59D4V/XmBwUyfBRZF4J/
HNqeu05NyWsGieIuVzKqIzvuWK+E51+rTBckD1bHzgaBYI7iLeZDG1bORuCaUPXS
PxjBilpI/jYhkBBW6DZzJ7U+xkk9PL1jmOfqxFeJuWMspf14MKN8uErjbyel4QEA
CxMcRJsYNN6kRXkfeVQuQFSwivXe7TtjznURc4BwC/8bsleclz3xaXJQdxBSMLju
/FcFYGHwWPcutG1FmCCs9RiPh7/nyMxRAXfP2f6hzDZ9Kxd1ozOdIdJay4oyfwjL
FXhvd5m5Gkv431ofFHU9g6g6fanW7V71+YlSbmLETcOrrzfecDBvrHUfwnsNdzsP
gqpgfljYOFZDDuvn1IdJLd+yrDs2oNo0+6HQACGS+B3enPrhGQX5JHluBss6CUSI
HroxChzhW5XKHtStAnTFh0FJ57/etEc5cro4yqN9h+9oMLD4x06jQUttn3y7Yd3A
4mtCjfAcBUzgVfI3vSTrKzaJtx0LN786TvkDyFpfA/69jmtuwSUwI5ZwOKylTD/v
rJvYNAzUXURaPHHJGvik+ZFomOjQBjJDDTAbYJuXPcG0ELWJKMCAp+ocWfC6hINs
uzknNCmXfMtqw+4NYY/0COdGOoOlGBf5Dr5wFaS0l1zxkaeRJm3SQL5ERvlDUDhQ
DzkDxdPKE9RnoXJ6AC+OmgbAPI13FL5iylz+rl74ysKVrfvwtXPM2QI1InGd+kky
cFt31SyLf4E15fahsQT7RgrRmIyh0jxJhYzHTZ2iF3xJLXp2iNRHrp1oflIHZg4C
RsH0BYRRt/j8dR2txonSj6cQ52Pecr8APUFnFOAsgQTGnv2mRMMdH2xxuhMP8q9M
S33pOh7x1orR38ayFsopNzAjdYUa7X9U8KFHEd7ZlIkfJGKJRwXx+VZQAjOm7zH7
Plh/fmByOOvTElcX5BMTATF/8vaj8faxq/KNS8EoPX5TUoZzYfftKLu4cG6d2Ehf
i8u6ApMn8/qJlos/LGz/uK0CAit/phgu7eNhhT7aYAN78NxXw2EDAo4tSc87jyX+
Ybo/+GmGcCeYg+NWKGF9g3wIA6AiN1Y6kmZpNGgADPJd+c1rHJYMivC5zvZXKp5L
F79v0tdBQSJVmCnlKP3c+O5l/cirDkxQdJQmrzm+haEl20gsL70pr5Bh/nuDK3KE
lO52tM6laQljOhHhPiObWhpDLK7ZPVEQQLknk56odFWk2nf1pKuvkQusQOd/hEQk
zWwbeKE9XxG1SmTDCeFH4RbNvbZl3p3O7cHbN1Jt2JSVKV//stP/919iStBjE6xu
PprWAO3AXDi9dXKnLkaQ55VOJ6u8lT5ICGcLsC1MWmjp0ThO0Z5cLrBjwnK7LOek
JGKNwBowYqPS35ZIgI4l4dXRM6h8b0H+LOgCEZjDBE6+96dRdHYbpnC87gcD367S
PLB5mxNeAHiF9ROFPBlqNq3gipT2go+qAQqHFsHNxh/cRu5xRw4Xhm6+Gx18zAS+
mpeldxq3FqEvbNkL3r/QlVo0zcsMU6VFyih0Gbvtzu2h/6FJ95QICFAx9FKmgsuB
CAXS1C021N3GTcsLWmxzpEw0P+Ro29n7b8MKxIyUXdm8jJS0lQdgg99rw3VtxFrW
fmVbtSMRVSrfbxCpMvWL1UJLbyHTBAHZ4aKHfLdUgVHANOaxFFiD+3yp2lVBwRJ8
DJv+xG05CytBsaUqui7HHnhnrYrgrgwpOHp1ujdQgeNq75Yq6bs3twJeGJhJON2p
k+LOYFX5vUZJ37B843poBSyF0OTvrKRGq0V44rq3kqNvFXzLLKSKaZQYeb+0i2MD
mMztmOXpR5m7ADTYpp8M1TRcnb+AZdY3uGHVr8Dv6S1ePC4dQDspcuhXMANbBxF+
QmTiwdQj3i0Z8leM4LkIGJTj+CEFgiI8gheCz4vzty7P3Ih/yWJ+AQprJTxlEtAy
gTpToIu+iTljLyeUDTLoI/e4lGNI/oA+ojvVrzx87P7Ys5WrkRFkf98Y4L2Xx13L
vvUj6OG/wlgsEk5C67I2Dr3DDuy8NGymm14jNQ1dKIIwaqPcS/w+q4texwQ2QN9u
5K+oKhQX419A7chF7vUH9Se4vC7WCllUuFcWK6ZpdoPHc3HY13AfRONWV+l4i96V
M7p6jmF4PDD7X2JS6KUyoufpActExznQDRXTIbs4D3feJT5OupGEJIcyVf9V0TnH
8zXCHgBgeLZZ+x9Wv5GiSgsNE3qtc6U2RBtkrCO+UWL7MivJxjADT3my0MwVg/ps
P8wYeDvuOdZNZVNoIRfg9cOAhe9XABgH13U8ZKn5HdSgeezsKXjLY1A5e8gafR3z
gENzaWQ53fg+3sBacIBHU8rGt43ej1SeSWbELECgn6qBQlOR/uPzve4/bCoeU/2N
4JOpF88VT1S1DZ0tG/qiqhpzipaGbCWRiyxUrhUAhD+KG11DgqFWYVMlULNmUlTk
IiJnUUpgRC71d0W6QnSRr+e4jXL9dK1JFRXTfGYvCuH3YBd12NbqJ4DVFtZfHPsm
QMi6E7mtDfDcplnjYfDq6y3u5hdT71lvDOeeSsbr1iXezwd/i/2QeKWTHn+HdonB
IxLINROeaSEb03NjHrOwN3oQrUYL2gOK3MScBps4KCbhH6ZqEvjRz0K8m29IW5Ae
VuRtHNayFVYL20jiwazs8m1avD8XT6FeMcOB/IcA0F3p6r2d2Pk54e2pnXblxb/E
murnc6+PdDUiACHs1HYIy1q/1yE89gad79MAzSQF3cPHdt753b/86/kp3x+N2NPp
0RvcCpLUW1IxuvEq/CxHvx0Lk3N1Nb6K8mvBjiqqkoEPKJp6U01NyyFDu8VA71Vu
vlS2Vlj1yyNYqzOZxRY2DNlf7AC0fHLBqMmKNN1NBIUe2zGHhGDXzVm+FkRJBjd3
ltbJdwzz+Zug6mrDDdFQWCiMGs/13WITWUArhHU/VWEBoZVBdV4Su413NL2MT8D5
w8L7nyvz+IfUKEn6XX4ZHomnw00Z4g+sGYPttoIlGNV/azFci5D4uCH+QV2OSyn4
TK9skQJXkxdcsXh9F0YNrpktb3r0swym3VceFBUoEbaKrk5One+c7d3tk2RIJ+JX
guuqHCOQgxarsevZFqARaSoV47S14Feidwemijj23LILPiMZbik84OARG9LOlAt1
oyr6mZ0k1OyP12S/jti8TxzOllIZcLMMQE46VlpzNLHsghxej9TiuWfbCyjWU1ql
1eAs7lmj4xzXTY8La+/DY19PuhWMmVZ/0IVzYBNmx+W4tB0C1i6eAHz/3DSvo+lz
HePFdJbxwRSNeyeetAaAHDzMVvOHw2tt04aMiCSSdf9SIQFNAUZDjSgMc5+sAY+V
OLXAO2X9MIsQVKF2dWZTTbGGvruq+tua3lFO78jOdYUH0VuD1Se2iCE2uairKkHl
kYMxPi4nLhtFYjG2cw9aM/YxnfJ6pH8Z/cCxLk3hIB4AD1daZ9RNhhV/JX94k4My
ylV9c/Lnq5PAsy2wrUP7ShIagEMQgtg1vDOcVXTrH7on5yLmr+/PSdfZHF6AiUHg
CsTrQqptMdsDqSQgXiWACVCpxbVkHdtOqUFj9gEhRm/Bv860BwMnqHNPZHSmBozF
kCKF2B6JwBO9+E+Cof/WAERNjjZv+Dd810iumx3YHubZJdqG2N2hNnJYl7ipAKlx
f4cbGQKrKQwghgJcdNPizU3jqOSsqvh1/IETN5HgtJA+Uj5A0X20wD9MuR70UYJR
cHn5ksxjmVTVxDZKoloWcI5Z2ljVZFDrtE8sCKZ3uRuU3LbHNbSWUf34hRZAeXfj
eer5tFXnAmACi6uw13fLQWMTdG+ENedg1Y5x5MNJ4PSEU1G3XmWCxA+I69kco6Rz
WoPnS0aD96eDWE9bMQU6/Dr8jAXRbaeMgONkFC0S8XEdwlM9A/vuCW1SSJ1DTcB8
fh0pZa4NJEYVnohLz2xpcyJlz4hUm8A88YbHuOhPlzvG5zv30ziaSLDxwBgwRAwP
ld6DTltpuFe5frn5OlBDVIZptxBEytgUIyqRn+DqYM1wpNyb/vem714nOd/cDtt8
7DEtbmIEM1c9f4DMyGJ82A2J7Ueq4pv6l8xYzCU7HceFIXxUrTlTQLPi35iB5wik
XzPKn3VQykJjpD+5sb/mw8jxmZuPdUt8JqL0szh4I+A+zS0h1Y0wP5Ae14YQcLZj
IS2bhFRzk0ov6+tKO6xMCaNbhBldtMkq50fSifBfRN9vFaxwzWNN3NEHbsuw3ip6
vM+WZEtgFo85MVgFYhuaz4VD0HhWSA5X6GpDUhfB1UJVnXtZTer5P3TEa1BJCkrE
CmJIsk44OXA5s8F6MSyf9q2yJ0GVAhla7EdJ7Mtcx6buFe3TE1865Xgl2CcgOka4
GygS71TRlGcemuakbtf+PhB+6jx8bEqg4r6t+B6BD5tk6BhGKBpSz6cHWf4RbMQP
ERwUfOk8XV8qUJovKW8VuwmVcH7cz0+e191I7cb31V5qxwgmRgFuYv6sc5hxCwoH
CPru6r2FmVBjKbxCAaks77jzWeoT8GL1ECUMhNgDh+dOCbqodw65PG4tsPRCVGbr
sc2I5WQRmcQy+AqcYUai7BDMLU529RK3jr0raJxcKRAqmZOdj3iONe2PTYfAdmgF
wPUmpB0n2+ktRNeVQ2wQ33Df6U5yAgcw02xUxRPuVgfGUgbf4zcdvCyxVpO4ll2Q
weTZSpzDyiiWPE/bAIZt3fPcAdsstpUZNRKkiIskAPniAlgvNzADCyta0Wom2kLC
yg7QfTlhv6ONIQYMi5PERtLir7QxacuuAptZikgwvhka8E8dVAmBdSGiyEpEaX08
Rwm4YhZJSj31TQFbu8CQD3n9/5wBBjm5bw+nxiUDfIjcxqs9baymvkjKVPV1Qep1
T8eTJeC3u7fxRWr+jprqXRlqcdGABSk1xv3yPA2TsT9A8aSSl6tzLVJckEm2ydA4
vGx74dexA2c0DoBULnUzYIJOaytuHKrI7Uw09fS/FsXXc6S5sMt7/TfVoa8u9Ktk
C7sCIzaQMH6APpPXFSrPMyxF/xEaFS8LcOzgqVrRl6AlCx5UZKEPkQiCsHpqGLSz
Z3nIrspz2UA918a8vQNiMW1UwYdQL7WygIulf+OBe2UVTE9EdkO1lPDU8ZrL8fXl
QubNG2LeVSthDFOEjwJ5uioiD4Iaezqkj5XEI4+s0DVEImAKR5aOw4OvKRjwQ7yD
yFNvJLA2zJUqhK7JdNC2NElHb4lFfYyEbbk9vwAohj93rP9aV7Bh4FOK6HLXq6zl
yWtiLPYJTuKo5cqIJnD7Fzt9CcK0+9KbFNVcLrl6aA+084+LaowU2vCpe7qoQVXS
y1qS9S0gV8VdJsqRxq+RfVuZ1iflgDCwk5QBmKRLJxsJl7zwP8twIjOKMuVLnQAY
1NkCQG4m2rIoRW2CC3qPLWW3+NbGdAcswG7x+jNVBV1v++XWsRIgTAXtlEUBkM8r
IHdK1HZ96b4+H6I25tdXPlL9B07UrlGMALpH+zoKdxJ0nM4LucAHLzgnHREMRu+d
/BuNq0mOpnk6VhntuPQC4hSk3wHzBaLUmoFya1ZgCZO8W+Gl/3QkKmK1Fw671gBe
WnydRA1CG4IIPcQ5jjDr/ZAuIVoG8ZCTfaPkGNJSy3k3ztcKl6Z+JqWDj8BmV0mw
Ze9Z77HMtydUpr1Kq7pH83bZIhnV6IQluiolgz5K3P4Sa89FV2L2LZFdY1OTQmHF
pdQJEBF8kyxKjZtbWOb8RnWNHTMZWulhM92oasOkyu/y6lXmwGhCJesC9uY9bHaP
CR484M9CUnPyrY4/NWeAE7OT3iQQIWT+zN5p3iKKMUMY103Xid7QJXLd4IbrYcn8
wL2++zzzPsl7WlmmSZPJjaGEyXhpwlznlSZnk/szRUOSfjOhvKDvtTarU5Q5EsHz
8h8B/15C+uW99vAAy8XksZ44izTSaBhChdOyBcVBeKJc0d7h86QiC1535RlO3Lcy
n6kBPOAfFHzI6LhaNE6aYDxRBsx13tm4mRuS7DYG/JZpYW9G1cBRyMlhEH/x4SR5
IHWpUuJmCdLmLYRF+wyhN06lobSt382N3DzX7nOp/phQivEy19ZZQgdSzaOx6Kiq
gdpwrIxsSpfORXYUZjtzfTHLVGccOsFICceR50C3K9cb/CLFu8vMPzpaeTlPzAzP
S4WEypZKUc6cf6QnXqgppMYCAoFWQXjJIbq4Mu91lvi34qU1fK7A6an2Lv34Mtpk
DkRCa3J9HFQRefLmu16mwBlR+J9COepU36LvYcOVIJyk2ZNi4U7A26ZQ5pbOb3Ta
tmrI+egU+RLaJ+q4jS115gXaI3RPv0ZrQWxzVhZh2Kk9EpBZumVm8EQaG0W2gxxW
KkB44vUcFo8ByQb90kDKe5oWYV+i6lbrYd17wcVGGJSAC5XqcTUZzRgyMonTrMxy
r2BiceLXaMxGe9pNYcLD7bQaCeUiJk5XukjJ2uWCw+Q5Q1jWHi//73inJyepkvDd
MRpreJHUn0U9stYkzx5dnx9mfuyatnGIS+8qwf78k0LdS2WZEHc4VEUlFYczBmlr
IpTxL41pKhB0+JVzcBvU4JW/rXsXAJRBSogq4CNQ72cXvcH/MdGO5TJ+qJapzuOx
/uSbIsYbZx03AkXghZa4irEsCREe/XIgEXDRnMEGAsPuuhLpkHO2IsYS1ac8soVB
zza9v6o8nEhFXZJTwuapOUtePfQD2QJFLBpBITdXFfXftQhxsa8HD1wqG+fIH7je
Oftx15cxh7qdyckvDurDCC/p2RMPI2CO1YJdrBsM+89Z9NAQn1M8ndvGq/C4TW27
apDO7odpPTR65O61NQkp9rLjdMxEQR+ZTbwiLtPZl3Mx82/2caY9lkXa/rAokshB
XIoj3bX7ldG2Xqxdyl6qbARmRlHHxdyjJFK9UhQ1Fvk+R6tWCuuQE9fu2eRExSK7
9ATlpkt8kE/h39zqmPq8GIoR9OBY9j6cqIhWxKO3XIlzTQxIPB9XnLl604bDwi+T
/Dcyb2nqhI4o0xKmhaRdUlZlqMlAe24j7hA7SKjklY19k3OFaJAVgwgFXyGc/7OA
WVjy5dfxhX4zn7MdP3CCKffYcEc8Z60jwLUt0qWeqmGt55OSW2jZhZiQr3mnbaqb
C3C193VURmgYtkUZhFTEzf+dFuzFzLgQ3EsFw9yI2OFnwMyph0XXWv+pIm8dc8EE
Rpvy3DUJERDpDmyW7KC6dwT5lsp3FQ4n2Xsbwsa6mkQKuC7jQxS8VDOPKBDPAqlF
kMxYnpFnIuehBXjpUUvmK9lL5zlvpcNYFluteMMJYSm0k0Ta/YgPPRRW9QCxNLs0
RCZQVfNyGQ/WL9fgBDEeBcfw6Ilq4iaye6dieHPlRrsfVlss13r6FHbdq3h5XnG4
4j+i0rxFg68/lVhvFHkeeBSr9jiU+ULXlKnItkG2/ouBKOBHFe937Gi+08V1lYM7
ce/b5mEjcoJG5RC7t7oOp5Ubrr11cIUMyM1o4x3FMHFLdu92BfvXhupi+cvC4vxL
tXzi542zbLrZXEwETaEA1gn2UQmey0jW5C4E+HpDCBBpWWuhGd9GQtixpB5CQb8y
28/lnnfDmI9RfIdRs8XbUJLGDDmdKHQarCzE37f+nOGFNpt5NQRaPEz0WpZMuKTf
2BRcIMgIaq6U6+cFequzlQbj3MeXwy0MpNavFxZnBRwewf7hDf4+6W6YDQqGFSzH
i7RnWI6e3Eaaofe34XrelicneFxD6uUNLDxsNRz7dEvLX2AP1LutGF2fHpZYmsFH
eClTo0MEoViOe3bqmC4sihYi6M/Na9O6WuDASPEgDD1uNRe4dau0YErA0MzJg+Nq
WlvYRUHo0pcmNA1102KS+uE9V3/9Amxs4Snwn/Rn35dJEUeovkIYODiFXo0FVnIG
bCslulJyvN0tZfJZCLYmjRiIuUPSRnGZqnzwuYWiL4egCWRRG+p2WOKnjgeOkHdQ
V4zwYet5ieM2fhonVJjsEHkUeOLz7zFrnxYy4Y9Wr3KXuCbY43QU+6khZewoJiN7
0ku2WEHC69KPZ8STHq1mFEHUu8HfGwS6BpTytjML0ivT3abSCU+w03ZasgFFgpyp
jm3jfpP8dxKj0F7FGcN1zrQea0MzMFZwCeb/Hz9D1aO0gLzJQDpCwd+4IA0tEG3z
VMnGedvkGQFi7mC3uwmQSdVehwO9uc//iu1C85mc/ymhsCGRutpLbl6Cd8xrnWBR
5ieY1jbIN4gBLOMUmigkElac6qKbetbGkGyTAw68wnqK0VPPFcvN4aGCmm+YGtah
hmpk4uxFHuELNydiRmb7WEKpMrdXL+Ro/rGk8Vy9J0PHlLGWOOueaMagpKC+NxT6
HkiXzv40pbO7r3o7ZmalfUttE35ODy+Z1zKk9MXEB6jddxCcpBgl1ZNllcdN9bM4
BJYt8PAJVASl8+tfOMD25lJ7KhuLUDw+Xl06XUcae7GTNL+Y1Vw1sPEzZRsYurA8
P6sAKKoKzwzPVeN6sakFG3kZewWyWpG4sirj2g6pQBYl5/dZATaSLlqH+k1Ee3QK
ZVMy39egIfRDIlxa+4NvDCVAesjKpV6Rjv9H4y1m6IbSiXv186OpzHffLpiUoGTv
aPLA+v/Fupl3Gx4oUZNmrApZ6dWjv0JyFV3t5UvDzF9NcBRcKRFx/ljyTeoxSVbh
fdQccug/DrXXRYRZO7TUpbPGV7JHlOXhwnKLEBj2EVOdzYV9nBD5TLFWnaXBeR8u
+H26mEP/hRs0xkoPytayKxO/8IYLXndHMJR7SXhwSmR/9I9E7NKQmvxwToBrZSr3
GNxdCYSI3bLc3O6SJSyO5v5tfuZsRl/otAKfw4P6P6uTgYdnW4iaDQnjIAuQzwwQ
ka0k5guk8pEuBJpZfnABBlBTS7uYP2bi7X37WzEEx1kR7DcqhxzdZmlVrH1I2R9B
F06oNkB8AxzdHS42hmfycbrpBmbdgR08cSbRd/VCuGBHGNdWazGe1Z6yzHm+G5y3
OOct/cGKh9mmZlUA6rQbLlsyU/8u82u06joj7nHRLPm+LEy+5dq0Bpx/no547IwQ
LPhskFmKlzo+LWqBbvxLKmeAitxRoO8BWkKd+Yjc153ph3Bsy9lTPX91OgjjaUUm
FPRoxefY0c4bQmFoumQ+JEzo6rzM7YiXz1B+AeMYQMXuQWPZXVI4gyCriNzslkS5
ohCskVSZud4Cyp2lCT/vkluCFjuqS35EryZXjz2iTCKCBSYjC2mhmOOROS8xvAlH
t5sz+rr7MqH4MfSizRrN+uOcow32LO2fk4kvV1GQc+TP6fwEqUQ4W3PJbl5EOVVJ
MCNkaGvcDT1wdt/h3y8V1tbqjVFR61RPhFG1LLsp4o5rzPwL5MozQYP7qluG4/4j
LdqqXREYBzBytEYJ9HpzPDAvkXQD7CHbvKSAbRkdgGINfDIT6PuZsUAZcl57LHIJ
Sz/hyynnVIVMYLUNHtUOo/Sr6l08FVGneFvTLrEQFiepaEIPd5k0s9IEkoA/pUU+
O7C+gVuoTzBJIu2ihlJVPi3LtPCcJfvi4tytX6MK55wR8tvIt4DY4YQQLZnpVsAW
VHUsFwkO12K8LKf70tC4//sCWm/3X6D73hYwvM/aThleMv07A/GQSU0jnkxN/gU/
c0TuDzHRHPUBL2JY2XZrGBYMziqhfZuZTfQsuYF4ar+6g6iNjSWTk3Xs60+Ag9PM
GX3M043DoXN4GlIOou5c0vo8qz/pRRpHgc8iM+koIiCCk8ke+5wP/To3oE7HsRt7
qJCcGaz02kDkM1zVzMWzX0A8jBJF+08+9Yrh1V3Y+N1rZgGeuYG+5OWFcijJBAIc
RgY8/YuWudS3XKNBI72xgHzhgtMujv/db6IQIiH3DxvidzIZkJ53He2eARnqn3ob
4TOvZwpPuMgUjsrp/FcEXX4JiJVOkrkd5Baf6WxDOsK9X7k7YkIug3rhjdZf6/ra
FhdNfaE8Tlk/geyaxIXDl0HiVSAQbIkC4/8tUzyjxEBMOYt6WKwcl5AsdQMY1GjR
m+6h7LnfkIkHhTb8M9L3msHmEgyW54fc0OUdu3bZ6XF1tJ7WGs7VZ5hB9aX+Vu/T
/a3ZY7lrj4ACmPYtBhN8XDb3q/Pd0l/TyMoZdj7O5J9A31qFiIzehkOmwWgD+g+7
ZfBi5535GyHGoUA7s1gk0IJ2aaEc9rgVZEj6wl5ZzogBCVlil2lTXmsTjVIzgRCK
E24fQR3FS0s822WuI7QqlI3K4uOlN+8ZBEp/W7mqgeHNY23SVRfP6rmGkaRYS8oG
ghBqMUDX6RypS2NmQXl06fyb9qvQ5SImuyIx6A8gPwl9GPFD/FNwgoEwOepyITaY
KN2ZKM5O91I7UeKsTqmhGGSW9XJI4fy3jhF4wBa9zdLx1nZhu29EfnI6hCE5cjOX
Hi8RismzpblqAuLnB7UY/ZwChfvEjg/22as8wM5ZDnfnPHqehy52ruUKI3ue7YQ9
zoFBLrSKl14zEeeij+BI5LnmOClw1mkHBo9aFQ5LzcPqhLCGMeaRIxy2hAtC6Qe0
HINxX0u/vtRc6DPk4GSKLEdFwBNrH86+x3yCPjFRxB9O4G9XN0h6iY0MdT8VKvaV
nAcMt+5t0DmLf2WIQmozxBFcnJ/6rgulBCjeoItl1KvvLyLTQGzR+Ge9R7/JQuGi
bUxCwcFSYQvzMJVRA0F9S1q81NAermhm8zRaMo1BWFlBTiiPVs1Q69NylzPg+EbP
bw88phZXHx++cMbsvqwVe6cL6PP7Z7Bu1z8bi0Y34p4NfWsblH0DKWQoB3Ll3i8Z
OgjR3niWGoRXgJunDdF6uBDUMETZyiZmV5RX1tKJIXwOAIVTFCd10/2rbTnizFCU
8A0sRJ1nguto1/gGbQF2BTTiYOBXdM4gooUJVdVnYFxQFUtCBmI+xe4u/kVVdEZa
NQJMjEUnySA/JdFNGVFN7uzZyGhbQe3cqfAtS7NQfVhS9YjRvhxd8k0aFyGVzzRm
LroFQAWIJ3YxF1ayF0b4uxewmjh5oPBQVWt028+TUp0lZEcoXsnsiyCbRS3g2Y48
imNv40GDrmEJ1vdFO59LwssytNyP2dTUIZfIu1mLOIrKcoLfiTUc8BEfSzgppZCO
rBV/lleCEwth9BVsaS6DQo3wvY5fuFF6wKC9YhLJJyIEJWdmmfGka1W5wd7SjT3L
Ve2dj/5ii9OKpdrsP4CGdJk9WquHGcwDFXyOyGUPMhd7rhIC38QYo7AFUILhdEql
dD8+9jqr3zCH5n5XdxVPZQva/f1g5n9S/vvUTHz2XDd0cYhxZWqjcgZe+FjHv/3B
u218JXXM3zyBdSv3RJV/kXA0WS4rm8XFce1jmVwf62b3W4S1EOd19FcSoVJ1wWiS
pO/6I0/XR+HQZrAcRY/k9nw63pgUAQ6Rb+6aF0GnheI/jE30hzEC4aWF52JtAnyK
kIejN7KLUGJc+pbU1KcH6iQggp4sqEK3ZcLWQPSjDGZ+50sd+F+jLwrWww9M+m+x
CWjPgBllkosI1VqGPHvRUF973wrs+7ZxXcMMVP+vCQijpT9TXpEl3lJmyfz8R/9h
uLpqt8QZlb5frHN6r6WkMk/GFRxuq4qmx+ml46XvhfhGftUuzSbrqYi2tM3lLR8W
sM1AQHEApOhZf8hKUI8sUgNijM51Ynd9ozImJ3Ymr1LQP5mk5GseutwcPVSIc9Xn
NslNxNbXTMBRfxfjJZQtqR3Y0B2I22yEsUnQVAwINagEiBEkYsH4bkRiqu1RVMpO
Av2Dq9FgCCipwvPR07b12193E5BKbCvWYDPBEIRwj1RYOCkzYVPmYVkd5JSmxiTZ
4gzXiQfdUsbBWJcG5amA8n4Gch1G1fJXYHJBDOZt6bGRlOFpvxWUh51nsvB3UZPD
5FSOOQMIcUKuGaXMlgh2BtkNNnzO2mI0FY1sw9m2/cvUAp8cO9yqSO86LWkInm7z
w3UhdemfKYzfcesXjWOH2ydfbgtlLkKv478g1jzXz4ieMrx4hZbUQA66tUoIw7Q7
98k6eCz2CC3esPTQtJiwSYzI9qbwjsV3aRvVvxCeDwHJrHhn4b5xnEdQmV1fLFzX
JxWvgNQEmXAVOtC3iNigIbB6JikFglSyEmQYjLMp6il8/4W6zgewCqL8kEj+45mb
4Y367hGC1KlteNRJVKISNyB7IWIvChrwHicJs54k0p3Ph/sI8ITwDUqKejaQq/Hy
OA83pcejNfe0nc+n7inyY+pLo0vwkzIJmwJI9LmxtErd9rWW90eh9eMJy0NRs0DK
RP3brtN6afMcLJeUiYhxWh9AyLV63EHUYqDm+wpnzLEAOOux8VF1M6Ab+X6jJKa4
HuDHeOmIIhhKrlEnBHaJgnVYFJ5RVHRsMGER5cVZ8upFc9mfzULiWz3crvVi1wpp
eucm4FIiH+JePxZqjYft+fOR7JMk3q3xhDlFXKM7m/+sgIhwFVS6TaG/PigOcCUM
VK6hwfs72VF60KaNHKLsVYJmam8xq6QfhNHvJ3Y7RRg4whLBA8XcgiWS6l+bEPuK
ReLBsTEeshxXA1+j5xXeHcHs5Wxqmq2ZFK7s4648IB7HwriSmGvtUdlxE1JxQ/OS
ddE1wmjnip3czihDqcsjq/bId29fWqwP/QzPjgSJWmD4TcvSknN4GtKEJ2UJEajr
cLnnxgfbvyISRorv1ow2kSCHEs1DXpklln/Y3Tebt/AQVKmDua25CjV7H5zj7AAF
lAYC5DIBlYQpQB1WBXFkSyc6/2PXcoXxpWXMioFm4B7VokdYkfYdX+lYUr87oew+
sjeYaDyoA2Q3kOsmkTH/RyAmbg7bJ2xhuDvY6KyGkAQVAIR4J+noF/Nw4W0b4zRL
/ykHsqXjdmoVOXoX288HT496vvjTS+qzhQdIAvK/kiC75VORAvaHBXUXsAvCGYjL
W8vRuLQUZpR7dPbqGqrco0vLDQYZRwhWAiQmSAWcECw13FtIwGYkcMErYqMVecto
frddgsg/ehzmiRF4jvCaVRbGkbTgIFgpwPuLDsgtHB76tUgR+WWjuwO5+V0JPIaR
U8quREzcU+kz1DWKvjAZI19q1/h2ly3LmMaDNwqIcGR6DivNGBqyNSze/xPSz9mI
xlTqURgi5QoHECgx+KNFzWC3q07fhCOjOuzAqyhNXUPPBIBMozQe22Ge7IpSwxxI
99zhvZn3oBCXOkmGKRpz16eaI+upAeoDOsOn8UM4h02+CWWPTOMBnkkRmZhk2X1U
mW1L4gkp9xx6qtjfoZ+V1xMHY23HKOvf2h3oANBqrFGfeoCYZLheI2tz2aFzEH+p
HojKvk5bFuC8xxudI8vmf4NIWAiDPgcKAT3JXSRyh3S6Y4ROVfCmPgKP49SYHdK9
mgbaU3zSIbUZ/+/3RjZpmffo3ig9E7A9raXYN3FbaBNMnYhCwCz9QU9dIhagjH7o
8+sm3zJTJhaxqGunatlFS6TqzoyBpgmGLs00R8Kl0RjlI/YBqNbzV7V3iS2KxtoH
PCP+wKzbfvkAOtcrGq3z74FC9NkdSi/JISiNkqs4VePBoXrnOh/XE6af+UyYsaxy
SsA2q1z0owPUNZQk8hIy8l2HO2XukaUYKbLo4sBT1FZemDqDzc2V6Zf30UEdK06e
iuR3q0IRWCFAmo/AMrl94XyP4cnJFT7aYmdG3SWOnXtIAm04bUZgpHi/jcLL8F4n
B9q5qmKxfxW9scMOndGq2UEcJSjrxCSaD+GYi6yUqBbrxRK6sG2UMRBCQyrWgUOd
Q9J27ynn4Dd4+oyxaFCx3BHFzCyUyfxquoF3nSsyHuaVdpk05VIiH+37iYBx4Zz+
gSQUqbMSOma5IAskK0gvuy6RZklUDjuII82MCgXnLsJUbZye0jFv9ZrcrSfvS4BL
9oxoflShjqSdcyPDqKuPjibYciGOnJbvyMCqkZYpf2LtXbIgT5SqcgW9k6ejO4q9
sZEQCD467c9I535PtIjdrutd7+Z7Xzl2Rc7fwH2HLBJX1KqoGWjL3UJHGJ9fNyPA
9WkdlXQNpvcxU49SF2wPsTgFhPZrdiQ6oVttfdjgcoPmE3LFFVDI/jk/cb2FwO4E
k2Sit37ixqJVPSNMQJm/VoyGK0BHVTpx7NMFO/4ADfCODPGyTKucbRFSdo2G8dMB
cs0qwLzywOqax7HR72Qu7itJqTENys3hnb+BgCz3WxWCKbbltqOH26p/gTTEQiDW
fWQylCkfxWnrra3IsA/RzIBdbd46ZrJiWq/KUHoBXrq+R64eBDU7vVZOJ9D+/va7
PuGOE5pa721sR94tGTbOC9rI5fZSc0Dj5IufBnM8mmPDlu7fHEmIGT6mN+W8rVFi
RzgYkhK5eT01NyS9ofCuAL2wqQo7xJP5ydpd/nF3Rr41xQZPa0SOGzgclAAvZnMB
lehH27u2e2ZSdL0Pz17bDHpToDYjGDZgENmQiYsI57CLKqxzxDzk3Ep2k0IsOKNA
jwqDfSU4cIqa+VXLM0zAZqNaP8yw47w8bfgsHI94vE1qSuxEwnOMFzBe24TZiehQ
WTAAzMkKO3lfk8b/74O/sAxsGg6uRw2uCxZQxhB6aTw0VV2cK+pHMT5tpNpvcUFV
v3FB1tDxycMEp6dC9+ExKlWZGMhap1RuCgoCrN00ujzT/PcUfW2ys3WKPlOC+9c/
PJ0IcXS2iTPFM4bLL+cl56rJ8EvQ4yuPN6Y8TdvkDOZvvJArRguIrVPAdNOY9sCN
f75X2exLQVAcFXkiK1HBToNRVCfWtzMa/mXZiCossa98GoFLyqWglWE728poddkT
0byEWaGPq/XY3C1yxku35Ui0f6Fxc4Xd5NgJzfDS6ORPpbKBUPxLhm4NSWJ/Kw2f
JWxsBJ8q5eSkNN++7P5S5Hzo/ceKWwGBZKeWDY7EUqt+LrgttmHPrXROKc62YPId
ldwO8MT604alSBdQrvqwBgx7r/66hjXT1Rs0jttzsSvOkQFku3XkapPQ1hnt1dvU
WrXyE1z+N2MQYtXZMh/m7GjiymbyF2plllV2WpfNVfHXK5ERgBaghlDpuMvCUuyy
zfE10RuhretJ8h6wOBqLmEzSeJ9kqgHXouJ850gUG8Tzoufv7+KqDAQaw9aShBxb
afznZ9ar+PcKS9+9V6aG3ainbAXnigOztfMaMKODPXWRWpTGpqbA2uJOh5cD1B8p
09Y/qnBLySfS/vauHhO6nhLrEUi07/Z8v8YCis0fplViJHYAx2oMSVkxIFH0PCo4
soyScYdxEN4LM20XaD5lQXkuROsXUWLdZTkf2k0VTeT7bcPzDlc3cvlMmnu3KiHt
jQAJ8KZjhaCD7YmTNMNjq/VcjIcPgzkumZ/W+tuaG62UVOAqEXOsX+Ohpu9gAcjH
en5nMrYBA/J7VzLw+uOcbc8va+Yd06YCCgeCf0mMcxw0+z29BrJ8bR0l9H17kbvZ
wJ1e2ILF08V/CS+9Cy0sHSMFYSaBWCYN86J8Zqoit1lmltEJFjdN0Tb1w2pP7PUS
WxW8eSjmGQJJiJV2Q7nUp6DBxfjd9x5pKLhfft4XhNfXwTKOlojcYqeD7k3DsGCK
Nng+jt2zZZmCbZVPOKT47bIaAsRBrUYxfRvxUs2iugwWpMC4y/VJCHUaF26Rdrl1
tLq10ZCwF5EMG4zM8EguAKAoZIA/jz18qaAuF9I+Khg7BZTrL9iJ1l2vIBqhpuhw
UcbLskSaIretn0p7mqXLWYAKxJI9uF9Nfy6W28TB3ZYnKjeSPWiwGggFwDF24jpb
rYbdmmd8s4Ed/ba3btJGkVbfBxlJuwweEqGLRQ7z++3Q8tyu3VUMlscPVNUM7emQ
bIUFfD90cFVEIQiXid7UfsM1v2BJ7gSqE3F8RgZ6mDWkCgCqzn1kk+SmctORjlRW
hnX5/TgfPlbQma+6VbaIlRCkwD5hHenP7h3sryn+6Dr3cQlHwlJulwo00LRmS9KU
83tc1gsW5r5TdbYoUuoo3pjMwrSL7ZWnKUlMlltyS+6/h4rcbVPbtwgwim43RvGP
sa1ScAmp4Qn6v+vVBzIGmeUHjNcBSqVonVkMwlEmW4Zu4hOO538hS1uReICKtoN7
hSUtwqQbFcYqHMukxyx44HEYW9FBI4AifeEaDJoQMvOx8qWO94A4fhZ41FIHs1IC
2f7Zq78HXCIzixR6y0G2zHf3HQHhMcx2LrTLSnvsgr3lVTSInWhzCj7aJ0IXNPah
PJ1VkM5D3jB8atI3zMIiBgynnysy94lfkQ9KHL0nS8coE5tMkbeQ2i2zCHr/G+g4
6bg9YGwE2GMetsmxAjUwA5CR6sQs10GgRrT1IH+fl+2sUXNO54CFyeX3zImbm+tc
gTvlW6JyBNoR1qiMVIPFWfL8x4YEZeCiTC6JZccCK5SJf8BBMgDcJ1ErV+qxgO+R
9b1yEbXvbweH3p3abH5WdWWz1MCQl9kKyX9NBYEaDdVQ/B2Pv8Vu68FrI4Xg6UZB
NaIl9fILCn+5WufLSkvQFm/mIIeNljIleGELXhWRgv4xcgczkl/GRFTCD5M6RABl
XKTlff5+WudZya/EvZziPqas4c4wLszJlVXT5aCz/ooejtpGmqsJj8wQYb4wgH57
l4kgW8GGCwz+73fycTYwuyFewB3xPvGqXa/j2waimdHN6a7cMcK3QdjtCPuHlSUL
s592Ihhxeo9N4Oct5NTK0p7LkfpbhiJjKwEFs9nbo3phbB/Rabi4bW4sOPV1/WXm
6bHp5lFJ8khOwFYhPvBE4KPwllokHvGvlkRKlYgXWa4aIq9Ja62vEoVy6aHwu8Z9
3dpPKekjarV2lDjUDmeQpGu2918mr+Kgku/MydnECfzGjEy9aaf0vbMIFU6mhbSv
UNjZqYd4CwCW3rbnBCTCPYtpACAHJWgs/IylKdTAWv7uLgjF99scKYBj7CZ94FvE
uES5IGm+5LoEFTFnyehBxa6/+JA3m0u9j19W8jXeu3CNdF1mQ2t0K+iGmTZ99Hf5
VT0G3GoAiIII4XwrWFP8qbbXDWQXbhiR+2Vj8sklNDy8JAuMRVvGvBmbHqNbYqe/
t9c2TRKrP1rslG1WUNxjIHkLCpPgXeWDBehbzi1mHBQlVoyK6YLMz5LCIDiAOA+T
p6P8jbZdvmm+hwtXj6jtZzZjxnMcZS9YcoU93O92XEzDaFybBEC5pjv5nrou27xp
ZYkBGJTvc61s+xixAOuMsXNsf511GPUti7p2Q19Ntoay1S7DS7Ixmgv1/BzHep//
a1NrJO15QOEOjioiAYT+1uCwWuDPgu1TfZpZew0YCnGEtMVWWCoFraXwLeWK+s4K
mkhq8Vnpf+3/irPzbqSeOoy13+ctriTXzJLs4tohXAE3f8K1g/JPvEL7/uZq4Ax7
wfeF513B0ZImqWY7X/8dkRovtydBdxqE6jWS2mA2x5ai2xqZywg2ihtCxnBK9hhl
1tysY0qO8Bk61D4YihzHR2NMkNwoRENr8dDrpCTZPguw5gYwWg8r3f7AB8T2nBbA
vfxhX+6RuW8vJayYcXkmhhBj70w2fGXGf1FX8WjmrVuiLjdvowPpXMSlg7etgDbn
+mElPQRt/jPJ4pMXaFIg397JUpKYLWqXM/qAMFW+e0QOYzZUC7vZdElXh+XSgDjf
s+jUTAO9Tovu3oWveSfObqd9nNyKi59vo9AldT13Cv+RpgUDGXsm4A13qQFjp5TX
UXkQ2hzRgToXOWlxgyyA1iI80isCW3MP3R5C1+Vkvw2AcYxd82eAp+BfkF0lBzmZ
kW0bZTwnOVg4CYJmZPdsM9zxVR2/EKn6zSiDrJGKXJxgcMBF2zO4z0l+v0ziqH+5
xAJCduqR5j5tz6rgZAoJ0m+vI5gwWRevQOU1DgDDQhk4BBEbxVHxD9G5ctu8Snz2
VgiPQQR38/6QRYOsQrs4OP5XhK1BfKVqVx+fu1LoaxvBGXvMb8OSv65EvyQp1RYA
QPOxUZkc7OGI+R3/TUGEp6oCjhZ1UlyTuwhkrNzskaRThOCLm+Ibr4o2Qbito/WU
NIAnO+Rz5lFQ1aKh5Qh5rSEL4MetXr78jyVeIXDZOe4y5qmNBuuOerdE4cbqtDXw
k3kwghhTVjoV3GFk07y4Y2bcdPjWgVDXsfh4ZZ+kH9ZcwLyWvIUHt7zVaqiiTIl6
9L3wr8g1LI6taFdod4Cnlyxxc3qwouRHu2LEu8ZYv3D2TZn6HP+Y9Qst4/V1ZpWZ
QiXCgPmeunceRR7vuSZc0uQqKD5Tm4kmY9kHL8D5MTGwDUJJ7P6hsoTY14fodAyz
/KIOXIsNusDbOsW6oTxOlH0x33eZ3egadX/2WvCSSKaSaMV50A3k6WBk7CpSv8XR
DUKxOAMu72km8/Ijwswc5I/S3peOIatHU3vC9yXs5/0vpJPcZzpzkAeJEmEHrIzY
/iEgycJMulpApX25CyBYwkZRiZ2RmnPlyMZng41+lwXqcOhBYlqq0hOSuQ3KMn1w
RF4g2iP1HE7Mwl0XzVPdXAKuWRyXIeZKCmef5wWWXC65O6aWdojQ0NpaioiJTaC4
N4VZ0pBd0yUZlZKv+07puJq2wlpoeY712q4gRVhlc2QhPpXLO3vYW2ScPD+Yikzh
uKfgrw1hjJPiU34Zh+IbGYdBy6Q4x/L7Bt+5BV4Bz/x9qHzPSFDQRJHKawzJ8e3E
U5lhq6YNF8BFNdInC8sZvADYotndrrHQEHJai2JIQ8FdAFiY6uL/xwrG3IXfAXKp
FTkIEUIasT2HD6DKjsjMVNkfsefz4rxlvv6bagw8fjcw/flX/zgkLr3WYZIMpSCn
K5pLH1RuJ3HUMgI8sniUkMJ4k8MqvDetbvxfq4bMMNn8xDUhpFKBldJ9pFfjYyON
RPg4jfvgK4LMGjxAcL3XN0iYGTl7Gv+29Av9Hp4h74gzm83GoLDSBtVJdq8CEMDd
ahX00vJHI8wp8QRvs2JElDEtaOiE4dWMN8tnFfgVjJHxUrRmcpoB6XgTvD7uBgS2
IZrZgT4CGC1rOPJ74gaiy/fCRD4S4MCmDGE8Hez0mnrg58zwjUfp5rUCnBMPL6QL
n44xqb2A3HtzQxlyf6Cg2oPQ2sE0vGG2DWd5qCF8RAQ5Z0LM9LglcKcv58KRZ9Iy
0OnFxDhnpTe6QLY8FQCpQ2DqGKwjcrAihS1ICqMX6AfSOcOU3T5NofP6Otf6WQYp
vcdJNtKXeK1f6GYHjC6HpsHxBmokcTrhfoNHkwvZvukz8sf/0jIYM6VNdhFCZRWT
+w+te1OcrMFnXMP8pWHPuwCsOLKu/MzSSJ94dDeMfDkTOlhqzkyX3P1K0kCBrL5Z
zV95MlZV35p5ELyLPuLjditdUWTfrsAcxBS9oZfCoPcYpWkk1iW1wdvBbgCrsfZK
nNKiBqa0s47JUkrN5NGO3Dc2EEYPrIfC9O0sNV4IGBOcpzsJ9LrWBCv9LWBEMspl
ujNeen3Wxyt7fGqf5UUf/F8nRPtwz9ubzRx3hXXR91eGgzOTkivKx81+TQSEnP6+
rwQ/Ua1rBVYCujYrgE6+NFlFwZREKId9WIULbjzn0i0PJjHm/4Tucua57NBxrnFw
3v8IyGvxUtMzRPHu5xXdkJQAwU3vij+WhU1DhXWTDQmk/wmvqbp1YvwbrJjlSgc9
GI7pOavjUd4wBoXQUuzn933P0Fcfp/YdrkKX86vc53rQD7J6qFBcPnar6NNoAjEz
kXFFPTapPmsZnflXtkkKZjTY8+7q3C2zLNp/nVr3EZhcSDxh7ZIT9Q1kTgp/ofLd
CAuJY9LsQnDDcVNLAJ0lI34s864I80Id0+q0Dpc7U0mPQe7scBPgZhwWaCchOPMu
KrKPRt1nnhywYeXjKCKd06xRCFIRbCE8jEQkR+sOD2dLkB1gyX8xcDupLpcfo4M0
L/8ll0R9Vi0c5YOG/yurQa7N6NsOuXowdrrW551THafN2jkNXuByDpcTnQhYc4dH
OcioC9A9yUXhzP0W264Tw3dD858qqKagvBCaLHZa0UEW1oZMDUyOvZaI7/zAFoH9
qwUVRTXQh2ZVvbbHx1CSyK9R7g20WI3QZYjchJJn7p9T8t9VXJElPj5KiXk+wOdR
islRE09hzw/uqIqmcqsIVT9eH/cJBlmO/r6vUKsJYbVgMX+GpuvyuRMRZEuwvbhj
qDrXFF2g4YrNkBeeplwbGB3cxXewI/BckZsgRGp15q58vnmMJ5UHDGvgZ94G0O+E
HJ9TP9ZjeomBWCjyzFs/PPMBJuWJNZkeXIjbYX73wOMR6Qd2IYlbXTwH5V+Sext3
VCW5ZLHRiRyVYNkAucid07M7qDN8SqRGe3XRjBZ+mLKJ401LwODXamQg2dgf7JG0
doO8cIjvmSWhRz70fyFAUVhjJLP6LQ5qidIE9aG+5r3lExQHKX54KVxI0wVcJEUn
8Ytia302nHV08D0kKxA43lIGSGAsIBebrxXcWchrZpjA7w4XmyAJ6EIDLYrP3yFa
ZJH+E4p35Ghc6WTBXUfmHW66kzMpoaELuKV0U/KZlOp5KFNL4w8spOnOIxzb5LsG
w7mgemBkrir6z3PEExACF9kT3pFz5PleG/lyLj8RsxZ2FjSpHXub+QD14GcIW9PM
DlhPdi0fnUJA/ckGb1rH/e56qrqIeeDYwgFd3qoD7YFmuPwl24nDuA40RNhvlIhP
kGfahBQ6Rb9St3LH9kgG0wrP1G59+LR8q96IF3WwIHNIVUaKMQhOUaMP5f1Az+H8
2iHwaiU9ugqBraRpUQvYQqIVI+FMcBmS2jlHBkHXKjqy0JUYT2n409TuUk7RtCsa
3mG69cZHnhaybUJbxCPvyFMGLyVbQW2pVQvgseEKZqyS4GMtoKeXsp1l8pzq8+hi
TZNfhTxbBox+NWHXHqzyxLKYrhvJDC4+eLr7itGIdg7a/42MFrA4MEmGYIGsAMKI
h/Lk4vl+d1LOIFPnMkKFTc4Dvi4bj7SWG+/CcRZnI4xrCJSlC6aCCuPCdtoBvPJ6
Ti9knSXbtQfbv7T/DduayJ/pSaGwHs4pBSgEVzLbXpwUGxhzocN8dHNJ229ljBJg
jYMf6/rQcSGUkEHTFeE5aqM8glbH26nqYxAryFnHX5s38lZ/CF2fa1nDmLK3lkEf
iNQv9CQ2wmvvJ9kKBUD4Dcg8YK/2xpTT8UyxyItt7tbllpGZ3WGDhGSXcK+GlQFA
+2+alb7MBp1E+I5kJof8tXsgXZmDk9irao9hR/vswIhP7HGaaRwZHfhAfm9u60h8
vuMjvF/YgutX4ut4kPSe5JLCB+PA8bc51PBargK4VHQipMlEs1RJCTjM5cb6Gk33
D6FtBPXKdtPjT6KYBAulHMJub3kWeIfX9RUemyLe8eOCFFiYRyjdODZm8RkeqNvK
dx+alhwGYNpcXVzdC3nIFKtctiXL3a9AArt1j+2By1vP7UuL7CyF8kY8H193RI9e
+t4ydzvlt8TzH0hgcC9t1xvqHY0UuaqILrGzASo3nRTSojiUoSzfZySO9lxvkltf
oGT+8a9LeK6Ww4aLNC6/J/SmcoJw6NdhJq9cMx7f1g2TOKIuJfzuXf3vxPfzVHxU
dFBQHO8cXo2MRYRBYFM89F06Nlcqum+bUImdj8XRKgluH0eiIogVEnIuGJh0ize7
3Gj6vj5OdGBF5QuonPzCHUHeZ3ehvYBFiNIy7JeBl702wqUIb8XpdovvnGf6yh0S
4wWsnpIHdrE/OzhpA0tm8rCVN6oN1o55soHmLggpkw5azo4h6Hk/QB65cfWP0vvy
jKJa+UyY69tNOE6nY+iTqqCOgoTBJv05BvJQQXB6b2ma4fZccOCpMk4O4VqtgoZF
EqFNhGLKgXv1NZjvgdOKMZQ9UZhjiDIQQRMU6YXVlrocB61xzvQ76XSglI4S4kPl
IP3rRGFL9p2Ek8+zkmWmfnWW4d9CZeDggMq2nYPxR/DOhaujoMD4LzW2OwtvFFUT
BhuILYOubWKA/MhgDLYp7k7+rXSXB5q/z3rP1jsQNxNHUe9Wy0BnY/WUDxOsoAxH
AVoS70odEmFnhJWCjGFf9OgucEEQmhNKa6gv63J2yToi32EqcCF9ssSPPSZqsfDq
HQdLJ+geUDr7WJQQc3IK9B0mxGVYiELB9xdzc+yJCignc+W/C2NDt3wptEe0BduP
wtliJbVYEejFe3obfuU2Uaw9RvCvwb9vCNLaCC5UC0s7X0FgDQIiEXT2XOIBFd37
lIyQb2lhv6s7EZGe2pa+Tgfu0km91gHcOx+G3w/pu5H0+t5DPYoERNGrk9nAS2co
yMSoppuo3TN72Mgd3L7TCMorClxEISjwlYeMKjqcbEyYsIX4gjl0voZZzUAnx7bj
rdvvnhIoMRoACk4w4w2sY5ZDatiusa+pO4k0wOWjr8NgtDB/LynlXz4sSK+AQDCU
a0olsl5t2GxRfVx3YrqAg8c4w6HKbm8h0nyouCN9ESbxkKkYDiHCYzyNvcZCXwCw
TcDdvvPlkoH6RsIMHWPLFxac1sezkCDUUViCEmyhgKhd4nKksFkVH8rgTc9Y0sYj
AU4XhcABecKCYm53Owc3fLScNXbTZNosW8P3bPB9vEmMxIUtTEbV144/Ogv1yJp9
G8/Ov/MeZotJBAulnjDqyiQteVGlWxB4CENnnSJEQcbWk8aMivUnyqKM9DmJRt7P
eKsC4ukAETMWcaao9EzBLs2zJPZLw4g88M2/vZ3HfjtHOySYZ7RcBY67F7+QKpe5
x91B4dIQAbG0L5Rf1S4CJgxZSwluI2CeHJOgMTKqTgttHhEenZ/z3w/87cpl6Lz+
l4eKP38iCXwM6DahISZSo+o1FXwxYkrSuCBb/Kmb4TiGIRjPNtHAqQ2CgSgB+C5c
y7uvkRn+iKQHdXWXMXmnb+/u5I+FP0rCzVui6wS2jaHjshtNFvW/yP0ME7cc6c/r
cxFCjP+6QbvwAbmY1pJ6BB9Fg/EAnZINprTmueH0bHKc90XlSkF/omef1c+hDYLd
ALRPvaV4NHPg639a+rTzRs+Qi2K0lmKhl89KJeEmt+EtV3vaOk6ouZscrbTv/O+m
7F07NJj3/dvxWeh4y4H7cE2OSst3zLrt9N2VmQEQb7f2COrTRBqZinAly7EWGXsM
OiCocjjssMDsvz4A+gEw5psObR274+8yJSZaYfZI/uiM+Oz3RQaKXmiCy7pP6L+i
gRQ9q06xLln2ByHEVfRSlcDCbO2XtbVN4gtANVzyHWZHIJ9cWe7J6KcD6QQs2BnO
CMIgnzjVc7iHegykB/OIApwG8t4oyhK0ECYI1hM9laQ8z7YQmNbihoXaL4bZjrKw
eSyFexv86VSmR47FbtG0A99cLpPbsTgdmSEiVUbTdBvSz9BAVUGYlSu5nzM9QASe
+hNiJS/+HJqoufE7pVoFAZHTS3r4oJ2YVfujygICh80cFyGibEjPDSzvVcU8MCqC
RfypcqsGFTsSsoIEXO6AF50hwlYQKVS/yE0pjfufBqaXlyqQxbrb2PJVtZS2dTz1
yXZqrygFoZlJ+OUet6YNIWvilEMFVMlm8AgJwVQ127+cszMCwXwihgW0kuVBaMcd
2hpKjupyO1Ha8nL3FizhuglLA7egPYnY5xL1O3pjDDBrpAzFt5oVzEN+oRGJ5UmN
I0pkLvFWsRxJoqy2zhKGLwkTojhYvqcQlfAQ44jsK+6UfJW4b1HsE74Z4Rck3dFe
W4h6pJ3rFhnYq48E+p8HprKL76XLQ7fh4N3FduQ+cjl+4Lg07WjMC87+rgebjhym
mCIZWTFHzN0LqVX/zjIl56STYoJY3KamccFAz7YJ1g5GbgA3/B9NFZurUO7jg/mF
pp7EgO6KT582AgnBqGuEfm3ichcUs0m4OW1FPKWVaq6gaxOVWtM/OxwHlM/Lwpfh
40fyZ3ejYwK0CLhEl839MFj6Qws6tiYXLg+t2L6nXcx8ieP3fTRDYRckpwIMFMPs
b+v/IqftDM8y0ItSx5QNnIRqQSmn+Qnmbr9s/gSFVYkBOUgnsg36mkvOy8zwkFfQ
TmZPo44kHMBC/ln/J9UutVWuJtWLmkjZ3QgkixtTehgtCN3htm/nkyObWl2Pnk46
SH5PSElJDVnD2uf/J6jb9wYJeMV9EdN46yoVZCSfS2NRGKXe/oTmLzZ+st1ujRBu
1WsZ8YARMuu8luFLx8emSquOH70WMeL++Gr5hDLe/khKcCVHNejRxG1TChdvpXH9
Ghf7W3Nv3OAI5W4YX0lnTvLXXKU170oEIKkRv0L6Ltcgr1QZFxrhcwkAMkUVNjzK
6CpzCN1WCoSHWrbW56i63zT6OKb3/gUujsvEK+lTWm1deIRo0rWtiTYyw1YBWg2k
ogyTAe7DgURIXz14PKQzwQ==
`protect END_PROTECTED
