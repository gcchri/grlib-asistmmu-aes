`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YjPpRt7PayqUmK7y1vwKhqDyx43+Dfe1PxnLbITscA8XETkT+xeJmBvFI/XhQJcn
0zU5j6El/IHuMsBulg6Cr1yg813lDAtc96WLD1DkqUgob+bT0GIy4CGbg1GLFb2t
PxQksF9+qRyFCoESweGqeYCm9tPbaNrcp80+I3l9882/D8qq1x08je82aGtsz8UL
Ot2e6Sv6YnYcFtzKdzZECL9CgxqvhK9me5ZJo450xsau9kFZpwTNY9z7wIXmaMh8
3U36MLXdQBq632wUzndrrJI/5KqvT7plRQPjw7wcfgXPhyDHqs40tJp8JnzE3dad
oL384nvav0Fam2Gqkg0PmCleeoixSrJXI/vuObd7SKCrPjpFxk94pwzbSu3iLMVx
Vl/XEhnODGMewII3NhY4WpjjEVnhMLG+mnlbO2w7QuBCKGQKzBGGmX/TpGg6S/Us
v1mDAijdGJF2xkLqBcne2Fg9cJze2ZHuzLE6RiQvRFfUicLwBgEX5IWcya5ICxwJ
hdsDy4TZiW7k1zT4qHwRhFfFeQIuU67h5CJ5zgKyT1zX4d8ADLCl+2eCCueodHrl
FcfCDYcMdGpaXiNDr5kSWwJ2X7mxdU5w9sRif01Kfv4h1qbUNDzJz20VJ4hZ/5r6
l9zGLoyvSQ2MZFnDu4Ab59LouuflJchQt+xozQ5Yh905ajgKik5umkZk3UUQ/EB0
/5HMgs8mCP3G2nboRUAcBOHpXfw9va0YeA6kaw9e4OBYvNlm91IhN0HiU1M8JZx7
hF+RdMat7QK5oyZVhi99NXe/phhZ71+wBMi1esQUYoHR3nFCi9ceUqh58QwCDDJc
jMa6O3rciJald2bKC46+TbW9wM+HZ2MgJx9dsXl1iAQ=
`protect END_PROTECTED
