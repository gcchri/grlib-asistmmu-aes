`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZdKNhODamfNkalRWNT+nAGMN02T26Picn1RxUp3alOEaE+MFBs3iPqBJYxH7Y7Fy
iqnydU6KrcgB8ef3/Ry1ej/EN2yHdJqaB3Bda5Um6e9ARlTg4EbK1e6KX17NDzhh
A1uu7Qoi9ta8atQtPsEhUVkAZTWgANAmT1r05+NcgKi8ITw/ApH2VmpbcTTqmfWJ
pgMqHTtDgkdnwiHkqtqyxGkGrBJkqlBtVzijFz5my0dfe4RvUViSKc/ZM3L9Vsr9
AW6AdJ8OyZBN3+6//VZ1P8KMKolHWamtyl10//n2s1BpaW6vQ3/1tpGET7NQiF+U
R6rBbYaffzlu1oE2R7/FnpvEsxx5LdcYZaxObOtFbGP9kBOOmJ+n2v/s1/dcbXYW
9fwRJ6Rn7imPrvXbNdL8DmB/xpJ5b6iJES7FWuQNfWnuyC4g5vFNFcmHvbpWMO3g
WUgK4tM8nXTOaFymzAGtsH5tFrIf7hGBPDVN7PhPldCRb+F+AZzpnY5bgjKcXuM1
WiHIv51kPZBiLYeqfslj8WVkU13CkGzootZTD/W0rI8Rdxl8TkDSvrhvio2V+s26
y6q71VpFRlRo6Je1CQI5OjFLkmkLG9syo44CDs95Rr/jct8FNM6S61Caqc1I5gFU
0w3oqVMTH6/9dTVOqJTrE8Dwvt/gG2mR7y+HoYj6jt7b7nN0jpB6bHPSkFNDj3Gg
k40yQXB/MaecoJ7QKtzKDesmVjGu0phOrq9oHr8qdtFRFdQwvN9IhPkvzAJBN3FG
k1yZnhuuLp0xH40Xfov9PMCebF7xjSwoylwkwOXVDHfxHWXT3v6Ez9F/KTyNJCcI
DsOky5GOaGOptvsZ6tbDkbRjntDnHpVZAukk9qTNYmuIzabL7PvZyPr09jRm2rl5
`protect END_PROTECTED
