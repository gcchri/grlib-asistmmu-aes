`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oLwAeo6N4z+sR3O977KHTxnv6kruKW/qTnxaTrH+0JqwsVtev7Qfv5uhs3up0Jau
ST41fy0WZAQj6p4M2LAdN92R7nIjOzgUU7qaS08kCRJ0D7u33VLHPyG0YCdE0HHg
1nxb+wAkAvpZW+hvTWZUA4x7mpVf91twRiBsBWQ+RNSdnm7Uwsd9oIQFWF2uwGPe
NwGQks8pjuMBg8ZV4GEnOmFIFaQcGqq/gyDV7wu1ELNoKY/VQHOt2+YaN079hDcj
UJGsxykn3TexnVCIvgGLO++CM9NZn5GjqB9/3aHuEQBrjNIUjH5ASDQLsXE6iFM3
Si0C2us033Ucd2GLSWZ3olXJ1GEfXxRSy3pSTereMqvvZ7Y4bBxjLXaf52ihdI8V
EMeLiMD+HXdDXR0xVdOewg2pGNYS4UVh1txxCbDDNZoUjaS+2Uj6QZICvT2s8n07
vDBJdz2iMyL9mGcJtlM6iDTpPebawV2T0D7CViJNVJRRK16v4yJx7IKC/1OpeAP1
`protect END_PROTECTED
