`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BC9n9RVNkruHSei8wsxO1HNBR8jplaqUJy91xGPc6gKq9jcelRMcm0T6Lz4JDtK/
ThZ9IqQsxKgdi6a/1078zLVO+3qiQLXycCThmgXpfpRh9upCgaYTLNFZqANO/ra1
Sc5k6+F5NnMs+tBmgT0pIpIh5sPy6zTzKvXi675zNs3tbJEvrt7uEeZcRwo72riG
X4JewwQ3uPj9GBgw2TC8T676xY8DaCgfKtRUPOG1lSX/v18AHFQJmijQ+DasDK7q
bcGH2lGr/ymiysHuKARP5w==
`protect END_PROTECTED
