`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RvZGXEtimeJmsRpeU0HE+vz4kZcjYzYpMCO+ndzoqLD/o1vqD+WLPsD2UQGfPcxI
9V3dwPaFjuH/k9FwA/EvgN3N4XwPXQvBodQ3+9ACR078tVut7i/gC9yDmEfKfvkM
KUF0Z2Y3SN/k9u+3jnHGHmirzO1T6p+W6ivzs5SzRQC+di95ULXw0vpu/M6djHqt
iJF56cmzIkl9PKi+z7bUCmzP+QoCW9URME+bmXYGv3DdLPW4NoSOMLOYm5AIhffF
GU2uMHA8/BGjtIJcAwlOcKATt/oZDV2OAKcwSzW/p6vFU6CxU8mtJRr49MO/yRXU
KhZ4y3jDB/6dA5HabrK+GUjJQ6uMrwYIHXmqS5KnuVgYgkUb9N4pZNbacWl6R4kt
jHqNL3VhUSwlaDw+58bN9KGlSTNWg6HjdFmNBowODVsEa2PeiW6AoQAWyNqJorC9
V6+aQfl3cTUV5P40rJcLDUfRLFAZEpMQdrKpRXTDBEi3fV1QZxdNmx8t088ip8S9
AAtKlSlrbKXj1H77Uq4Cd+ezPFhBMVMTtUuGLiKn3ssbqdNM9zGZZJrQPkPQTpCA
oYSeBO4HMiXtO61v7/ZXU+EbGtIgMJoDZZE2PgMWwjSeV6/RbThrv2kJRxLE7GQl
yw8yEyXdy8dSxDGd++oye8KPfKTxAH4qqs9SDYQkH9JUBMH/+5qhIWLqe0PXt6di
CY12kvaVBwoPAL/xBqc/sBuAQNmZkkC+PvrW9oltZI2kiAz1gngmFLcho4hDd4fJ
FmNi9Dl+wfJqgGyjeV0wwvgs9VB8LWpSZd897qQ94YB5Wgm5/TlBxSujrfmUvyEX
EqR4+LVYpD1eKvCI/6ZQb8C5nn2e5y5e/WCwn6ZLRjtwoYzWebE0xc95+TMaoYBr
d+rDxIEq+jWyTsHuJu7hwNacjJGGy+vFXs9DJrDmjn51RrDfQFUiGBLgE4uxr1WI
XJZT6nkOafLCOTJXr+Mpnqga8kSq/KbP7UCP1OpJTtXJFmidRycgYNUUMc4sLZso
iolS3lnj+3q197d/3jwPx/rpSEoh5GYjXrvaSv5Gc5k9PdH8OMEA+cLQiEjYfUNq
29SUbaqO+jG5NdxgcPZ6Ff/hrHLBu4iq+hS2vsxaeW0ZMhgbJUCColI2LT/l6EUS
Fb//1ir6cEwTMg8m4g9xYQuRJPH2cFcU/72+zcACG1NmtC4pfoHlJluxhw8OMcO7
7rqLALzXazi1hT3epMn51zPB6MKK+GbzFYJMvIT/JVhc+IorEA/zrQOEQ7UXSF9w
CI+CYc/rvMrcrk4z+gphkFRQbOPjaxM+2Kpb/2s1kpFN9IpD3gcrBhqV4n9/r60G
CFMajA7XnujPjA/HNRpYxo4+fdjGtzlPU+IyUqyZb5u00G+2QOg2IdNYsvZ/SqPJ
j6R2Ihp1yUv7eZspVG+LRiWPHDhCTDPulgJztL3w41w6cBHP5YKHWvE/Y+ANZ5V7
JK3YYAxZ1V+KnQgM9zMLgqgvxYNzq4trY7diNgZ4OR+/8YhDI1IOubvtpxdj+giK
XsCYP8Pb9Z9Eub7kgpdJJ/+OIB688GBxR8UZweYUOmdKowIAkLlQgsY4DPpYkyUQ
FWiEJG7oIfiVkIuR4Jh4EUMi+CammiSEoHmlM//ibiCjccYTy/yMomBh16x/Q1Gw
YBMH0t432BGq07buQcO3anzAaVP3E+dQeEN7Ix0DfONVZiO7SZsHVJTIqtEUYmLc
i1LXLsk+VcTqBbAIckkSVk5Vzbc8EFa2PIFkupoy5CjyPYLYcrLjc/DUJ5lnlBmF
ns1tnLiwKbO7Sp3p/RYUeXNGLPCtBOC/LGKO3jGqqjFZCdsQ9Gq+NLN/wqYTCnOR
/ER4PvNwGe8zPiXYtKOnofi9XKA5NX7dMK1M+gEojx+E47smefGv2MfwF8zsshKj
7K5IV6yfMHvgrAxWyDWKWehkuBU+9UwhCNDiRIGnDZa+KJk1+1qCmoBcEr5P7D+0
1VPbPmEJYRZju0KN+PaCsfPK/PELAjcT4oHyrmqpvuSEKACo31oV7PsAcDqsUobV
Pgn0PfUrHXOdOBjOJmOgCNslf7SPeIfrsw49+FGJFEiDLnVoKu3TipcrIdI7i2dA
Dkci21yoSTAT3OHCjGxxoBWHcgRKdcU99LhBoiWUKBKkkZHhsKKG9tYSE9XgcKNH
8DxeZjWxkIvOOFVUgfHiTB2XEH0X69OrksKgdBISISq5UTecTXPh+6P4gE/LMVaW
KXj9F9h22uHSNpQcoqsjFas9hSzj50wUmHpoP1VAU+Xpr+iPx4HScrOMtOioBaS7
1EmfNlmrVq+ub4FtZ5/XyqqV0/KQo0IEUjquxy+bZXM/8Wf1QKdgoVnU8yn71Q4G
15phHiAWXacd/0zzeVWuZxp/YYRcbqYTbmgax0hR0/iDTkbDZpmoELPQdJRuicG3
O9cZFOojSh18lu8TXbgPdw/kKPe8w/8rAJruy8AjePoIAV+rlgVIhZdtq4PgcleB
rInEY4I+Do2BEIaSqNdKTzoSFtAUq547IkWA37B5DIh+oDyYAFCd1W9Dq5oga5dY
14VZImopXcdRh9Fk26NvPhCQZQL/Lla87cP92dyJmc5XJ+pHCkCk+AOmrN06S3vv
t7vh2GkRvzGxPafTYdaAgWS4VDkAarIzoKaib5Y3rxK50JCcdtxLerCv5mzt+Ozv
Mv6gaJx8XooesRXy/vprp17deQnBoMRQwXBaARo4CJTwvK6FzKfdI2dJNuRkrkYW
YLcFHynAle8ew8unFgx42cFUha/E991enWE8YyQ24RcxsDADJ0BKhVOQWddlmOyl
UpZU8YGovb3xtpg6T1iSjQ==
`protect END_PROTECTED
