`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q8MMJ9M79M7wIbUgxLr0mFYjc/OWv0LE9V1tLry9GpjAMuh3SZn1HEduF5MLxFse
8aGM8RE7n8l9kxWVnQWi1RceOPpGTtk8BfZM30ybq5vExpCibVYrC0h/zc7feQkw
iR2B9k/grLNizARBreWKuVu/osKGdALN1JjdxO0QTlVKQ5z1+F/QnXai1tH61z3T
U5SjuAAYkMwg9Ts4f+HZOr1zwR30cmCdX4s5ht/h4VTN70x3GUNpl+98E1cMBx24
ooiRmQO++oZEvXupZrbmOICeMS55TKWdSsuu11WlGJowTD3biysg9ul83ZIOLbfm
RjhP3AnnTrpSAgN6rlPioDtvzLB6EXMO5tuKtIc9QGWIcY2hRF6gQRn2ELvHiR8T
C5hBOHRhWkkCSY2tpyELkXFB5AZytTaXo+OG+IdMjcseR40L89a+N2ON/T/4a8yC
/j8VJQd0IbSdF+NUKaRabJT5E8R5Iwr0E50R6YlDuwqlPa5RQWBvsNHa94eyFqL/
XRjVldowcud+vAr76ovdyUJhPjk+BhVmQdna0ZZr8+PrsclzzvlITum/5SAOAKM5
3sFRfk40KHe0UXKhbonQRE5q0ECOBF8Ezq+YINilq0AwX40kxySsx2bLdvE4QHE2
L5KL1mUjzi2s25IsDREedAd19hSYj+dzCWGqM55y4y9tcOnsufA9UB5/GOtao0we
Rgq3ODYFNI6JMCTOW88Y0ywK9C25Brd7jrkAe1VvwyYqDPqz1KXcQFffsYR0uuv2
NWIDph96RBOhWzk+QxPO7Xno2vdeSL40BluoS7V5MGSFPoT7Kctm/jqXLxUZ0HL8
gEwZyRzH4sDnDZ+1+qNUi87N9aEaLf7wiDphPwwqMQCgTFOj9uRMY5qT19j1mV8A
2GIhnYLpsj/WViuvppdSTfa6iip6UOScYB2t646yawN1v6EjGv426u0PPq1qeTDB
13qmFkWKItW9fbHENQXbk6X43dqf6b4CGtyXtdQwAieWqaFQGaeMU66F9qRDCT//
RaA4THfj3I1litvhAUoUNj/mIcxLFfjrRJiWyvd7/R4LWostl6uj4BufMYzS4Eez
s6aiv3OwznWN19hyDLpOBVLIy3qQNGlxqCxnVFIMrsV9fVcthvQCvK6BjsWBnXSg
I6wHLbmy0Sp5aE8kUfmP0lnDnn23LyIA3VAoWzWn2gIWvZ9OLrt7EAyMuJtOoJmf
C+CPHKQ3ldM65ujgMW9Fq40JBCYnR9WoPypoi9TPV9syOuaE8V2XKuIvaCdPDSXe
JF1yd9zwAjdI2NVE56lIEFVvBNfSGhOBWB7cK71+3NhnpPMrqG3p+9/3m4enizhe
t8R3wlTZHizozr4P0Vr4ffzD7pl5czTjxetsl1pxW7f32RkB8j4JH6V/UHJITXj5
aWbmGaFM625Uw6MqFS1KJhw+Z5SHYW8OBfEhbJ/fGilPnMwrVKWuBN/f3H6PtNyr
gC1VfobUbcmXlw52wEIQ0wVoOVhDOaUXwMb/Qed+Kgc9J9ANphyC0Oxcnc9SGkLn
sTkGTkCLlQ4mRH5u8npFMp00bnQiGlGUdJXTch4fzXHYIZZnPNM9CGQOBb206z10
Dqc4I5/8j0iDosadoSO5kZCQ+FaWrN3dR0RLW03ypBp9wgD9paevAT2bnb/vFAz7
1rSpcqAuMAmMdUevCUFPQYU72ysNonOEFkBCBgqVU+wq9s4iG0VDY9rV0Xv/dX4Z
yv/5CYBcXurYUg13mf3M1USV05YkE4QAMwRVj1uOd/ntVV5L91pRzpHFzOHNcPTL
LuKcY/avrcZYBZ13ZwGAlgtN25gNbtIK4o5toI8xEuASkVfLYRTPDqfx67Zs4u8D
oMCJo3KbZt9noCNLFqA2BpL1pVdfoQuFzxgRiqOnJ3WUBf170X4LwFwtbTnAahfr
O8NUhy5UteNUTZsJcRm/xA5Q8U17OHczYPiS7UVxEuaRMf0uqOBHUc5WLDx/pGah
SeyAGuMeFJF3Glepu7N0YEQHag3n05g+2VTAYMxcyXbGnkXeDyVKDDxIsfvoU1gL
sC2+EC9SmuHmCrLBmPvsB9s5yvMJ3fQpPtjfKKWrUZMwVSk1SJVbmqKIIXez5+5s
YJr1XkjvhsUDbvaEi+tthCv3IbL4cSsWSFVzZoT26TfdO00bta/4tkEE+zpbVmVM
hAsjdH+CqctNeFtqPfHvaDRvUvSeKW1Ldvf+YpQzD/9yIzQEpuqv1gqwQL81kp6D
LbjarVmhswC/ICos/u/h09q7LDM607iM+9R6vstuaS+nOaFhqmVTFYFZ0q6luLVu
yBp9VFqVjfoySzaSqiDIyE6FcvnE689sdmTni7gcd+YToVP3VnUC9Y1/pqZPsd2d
TtYlPfRpndyghGStgZM+fIYZVArzQfShseyozDDJWVHJTMoldMfvlxBGFJCTQIKI
hfydUsa6bHXL3Ckq90bL0EgrTFz0TKHEhbw3aqG7Su3KzR1nNcvuw/ehFV0Ywwe8
5KP1DsqbgeDGEMtImfV6BhBdM2EktgukmahI+s0QPQuqL8BCa/VC18o6aj/kfi6h
9v3gYEbe89lWwwEPPVLG+OO38cUNRQxcDSgQeQq8oWD7gjqiwkwcxlr611kC0Wht
R087Crn8QAd14qzuxkdE3EPlna3xfZuZ8g7/VaPxaC+sB0AMiZd9L9Q9c6925A98
XuXc4jTgKS5UAzTsUc00+1ufrU9R/cC5GDB5z7gPGDxdj3XgcY+lNb3x4O+fXJKx
iRWBQ8VHW/47HnXJynRC9APRU2wUCqcvJh1VZubrgo8Dp04ZBNLmdOvSB1bVAtcP
xOUFyhCinZtjBh1AcDv3IUl5uh/GzclR+o2ST+PsITM=
`protect END_PROTECTED
