`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ahCSXXlbZHw7uAnkQAnJ1rNhDemwaLmlQ3DshLhoPj5SwTUDtC3Y8GloHkeV7qFg
PGX+Lb4Z57eALVAHFM2lCFDUJd8+aZn4+FjQUcCYnCSYqNLeBR6d7j+OD8bQeshB
3zRt4KCAEqjacKOBovI7YD0k3eoBUW8/EiF5f3RlZfl3GPLu9JwysLowCFXGL90+
etg86EyKztceHUeACq/wmzD/1CVjEXVr3NrKfm9nv+SnRqBlF1B8FDROZSZJU+d+
3VrxFCur5JMhEXZqOBKj93dwWQTeT3X/ogdDDcBXqhf5kVAqxPwnIcRTih7mpbIl
LbvVBBFMMSqs5hM6FMad6MAfN6UipA+CWv/rSIgxEr/FX6CcocLD3NOaZrJBwo6Z
UON3RyI9XiY0ioj9Gg96kuBbV1wIp/UEJ7XFIQpuUKaaqbDHbkCPq6harY3Zf2fA
QCZPdTwA6xHXibcVZPtmMN2FPAYpxHKgm+fUY2maHGpbbS4ifYwPLE0PgeQj4ge4
36Gw+/3K/0CLuwVFOe7TZzPTAOOwOG1BRLisAZ31kwqWFgu5YauSG4qP2ZYXF6Uh
kXPhLmopBnFVkYpExx/vNVNZc/GClIRTutRzMxHnjkJ7voj0Muai/T+wQxrdu3lm
cvax1yFG9RN6PY3y6fG7E6OhpjCDe6+sV0YDfbBZuYy8DAiwoxeBwWY3G5Gegtf9
dXqcjykN0iMv6OEdN/rocHYjqaU4+mnse9fN6VEgiiv0e0UtubKUSoZMXACFa3Zk
J9dfasUJueTYVkzetwPUlC+vqOaTEnb+0+OcsS4oQRz0S/KlJ49vkhg42HrSz1Gy
pKlzlVaf5hIeXREoOZfE93amI9WLB1YXbUkpSYvDn3ADgw3QNCcJIub57caB/6gi
ccrY1Le7DvPoftjnqteI6tDDhFYxsm1I0s3/pw/G4RRYhOB2wNBpCLVzkb0kmmMl
3asrHtCeNYp7nPiNfIdeIYuJ2sBF1JMOpslX94gbdyGHpgXIWkhvsZlAmtFu/fXR
k6R/X/wINvtuO+mw97eyQgG3F3Ebmgvw0saDrLvgao+0yB9Dwslg6idhCTJ7hbzu
VZPl+H689gXQhGXfqWSfwd0xdyJ+Jdrh0nTd0LCmSrQ6LuffD4DDTszVkQuDBit8
gjn22THpvRnZaLw21nri3hXmwhCOwAa+SQmW5/yd0lUQTI0ZJyUKq4iJA8lRii63
iHkruMwaQubRXSOqqjbYlrFExXJqod8G1Si6FClZ+9HbmErQQiSURaKS+fXCvqJc
vpPQDEdBMU466Bzzap++shRGoOTRr+Cm38VFHhv9g7B0XLCMxYwk0GZKUihw51UI
AVXfrL0DXD4oTIQPB8o8157q8wi7LN4U4PhqnC2sBSXBbCSjKl+uX3hylpG11ZoY
50koJTFpjOAO8uzKdasjgQSSrIFtSHYf5xVZQmvLkTm2c39Y+iS+HxQR24Ubu0KL
NPdMc/Aji0SNVIXRcgBGlVI4bBgM+VnE+I9LMeADxtexb7jHYFpPdAjJoLrnbWfG
Jcl4BXM+vIsEhyOOl7gHfQyVdOvaG+AdFCq2mRGXgStGgiFsDzR1kPUdXq+QEDe4
Qxq1nfAf2oLCm++P5jflh7vmKv3nx5yRrLDjPIaiWhgSeorhg9+Ov7GGxY6hCFwo
qDR4f0dpPsdQoHwE2f4x/kAnFR5JsDn90+jHJugiqQzbW1jytoWKpyZORRZEog9O
6PqtJvb4Irwm9bI7fR80KFfmtLsVmKl6ezJQoSoXAH2V0AJYlOEL2jkpD0GB+Euc
H716o7L+5aFpiCpfx9gPlr092pWePLVHWKhc+Io1xbkVOAVMXd1ollLE7/bcY7/5
6C1mSZ2v/4pxIbfah4OsxHSHxEaDSeOjiIWN5ufGULCkWgqyAMA/svdfnzxf60Gn
MqpKjNzSmTA/o01+X4ZTaZpxKLnsnEyB5ucKiWHDr8SpQ5kPqGbo/9M81rOipMR0
NqLCG2X13B11MGP0kxGy9A7Wfj+w6TxppC0IX5S6BLy3o94sQ7r17qh7b6whPLvU
MuXvhRoDskHDw+WfOpzBPUZtLfRAkPfnGfSBYa4GHOKIC5KHuNH7sgLYGXRt+kUr
oicLkV8Obco5U4LqyPFVzaGqT+vR3m97g5XqbnUDmHa9YO5jOMeo2vP/CvChMgYY
j95V8hUrFQOjnKfkrOmOdoBEfkAYxhfra22dm+OquTJTDEHG8diRoqaV2az6J1lr
DSiA8z/Xuf0UsRqtD/cGqU4dYHZE7+JH4rSJwcRd8LbUOYkuUGfKxJtCuuZpmabO
uuVHVDq8xvIEkeNWoZHTtdP9FxanpVsZQCqQSH8A7PqnLBtggqYSYF/HrFfgbIQt
1MXqRK++Dn29Z7jh1FDcWAXKq9sJ79Z3lURo8Uz+7jgR2Qu3aEUitx0rvmTQkZ72
bOKJVBInSxWXV/Gkc7mL8TsmW8XIg0kqqQ98sRQvDYnALGq0XAxjpti9f66H2eyL
OEKqLAfM+bkHU1dDSQSNIOJDpTls+WzHCvsV/Ti1g6ppZB5k5/3y6wIvHtDnysDm
gcUp2MvdtNJg+wvscgOK7hzjSQ28rQeirCAwf5KcHLHVATyDis0cvF1y8US56enD
r3eImuccKcVB12s5uyw6UfyelqYeyTlPB78tGnzoDEBygoFVGIhJp8215fAuYC2b
caXdXKIMvbgzivBj3EnGF3+ufS7sy2RPb2akopsYkCnrp5+vZV2Gpgu97ODLabUx
hPukuqNqWf+Q9IOKZTUozTNQ+6jMKzb9z0EcuVcsNz6vDGdtwq+3FAzZezrrTnoY
xBYNlVDgryBgUWHLjyKVj1ijDfz9RkEeZnCnksDIwuUhJT1yB7jnVAjNxkvIGuSI
oQ7zYNffAHqrUS+LIeH1vcueXtrOOF7y0hdrxGLmGB5i35cek3mJBdcOeIzbGE5W
srYKoW6jBNXam5Aq6qIpOmnAzDSCcVKF9au3Qu24ENFDcqRo/Efjzjx1GECWFl/n
EubJbqEDCmOed6wlVGaIZJU20TkenDHK7x8liYitbUyISVOIpx9VJLQHblUyRzQe
N7+xODKuBS/uJr//Vq1LbAoOKVqQJwVCzWWWtPern8QGzvYA82lip3QVPDh5ZWRP
t/ZBA/ChfJIvmhp6tliRMkZrLFdNZMgnYt206WPF3lsmVvmEgLEWWcHQ5lrP19uS
Q6aN2iI+75IUNkjEL205yLqict1OuHuI7Xdd79XlTPgnGeUBYttYoMzbR75n8Em5
3y33eACFedvbyPVHziWWWSX4s9mL+l5hMPIhnkbzYGwDF5qR/gZ05cbkWSBTVUAX
yB7f8xmcgm5WdwtisuOCHJGL4fQf1KLtc3OuwBOLK3XO38zXBJR/UHIubR9SsmY1
uxWfy0IXen4zrpr62Tn+nKma3ALrx3k1OT0EAA5iTZVsKL5TJcgil9qJ59JfK/yM
+EMo+rQs1e2DYC9KPvXs5KZqNXnnd7k6cx2VgA0ncQ307EdVchTNJkyN+QIuoDY5
ZQVlYqny0BqDxQpjQstzFvaQbuL1A2r5QJrz6/ryietf3mH6LgqgSRi5IkOGEWcV
+G0vJEZF1TXUp3nEL7RxqZsK8u1UKiME7lhYwmzeHl/RZzNsG29prqX9zdN5mpqR
S2g2LxpVYxoPBGp2iqTbMyk+70eZ5pyMKHy8dst3RMf9TWdLT1BPHjSNmboq/TQ5
D4Ly4wd4bj0YVKjhWmyXGryV9A5ZlzTcZ07yUTN1gcYYo9syW8tViosdlnXnHRC9
9M/aTo5F26vtlKOJmOZoE9lJP5fbp8ZjCuPLKJsTb6M4VWVfSIInwz/Mj8yhcc/x
KR+kHNtMvCvIrMKyF8YHVei1w3Z5t31z2ta6zfpCXCVVlNdpDSbJKwTBZ1xZuG6F
GqW4TI+3+x12LorAuQ6SR9/U/vLqg4+1EMZPuvCg3GequS01A4wW4ObuiEDyk4i4
XeP1e+C5vTcJd8zQYmmJk0kxHDAYTy8e9kdpqkCouItvO1W7yajILTWVeir5lKaE
KfZH/ywSXsTJnFzsDajhIpq+b2OeSQWyI9fl0tBv5xjZt7XP5VUGQ0ik7iNU9THb
X2pE8oc2Bzkx0uW83rFwQHPCkYReMez91q/NnhevW7umSbnApqlqf6gpzQZwVCQk
KUFwDbnfmHvrwBT2BQj9VfKsoRqMNVC0eCTT0kI9/p4GsnOGnlfkGGeBHZxw6gwb
WXg1LE2C7Crhhsyq6JpRUnzoaS0cjMxKNVtMtZFDy5pqlxB3uAQYwCLTQ1sEcwmz
405VxpaOT10WDCOvbDW9yXDlKXUwQFL4Ize/27W60b/EQo74aLysWkVzeL8W0EV6
6kVY8jVSq7a93kmom+mtANsLSamnPUdgj05DUiy28rDOQKD7pdjeN9etTZj6FBPE
GSlWK/jacjaDHry+kPlBWB+FFib3C13s7wSPQVLCJJ1OuABtn5XblfK9li1HI3x/
FGArXkYloV9s9zH9OXFmPAT6ZYGMrOEEeuFCRbfZRLCUGjsmaqgSln24s9l/6I0l
haGaq8ClRxfsUjoeV/9uW/hvUQhTrPWW4vnIy5yi/U5liMIl4k2I8iTSfqxx6dxc
9Ob/qaE34oK47QU/UruCYkr2iXSM9Jcy38wV3AINlWmo8yzlcy2kC8yZ25ouqdSZ
e8ddcFP6G0F8pLsGn/emNBvRTzriK2oVqzzE1zfyZZkg50SpWCh5ZqwOnHhHnAmV
DVsRlyuJ4Grjw+WLrfNdj48NXmV4JrusBUdYLxbRuVTL2O0OeRMOzrYLwU+D2BRf
DdnTqAlUj6uQBx3FSzbyql738ewkBopp5m+YLsGKpo+h/FexO4z1pzKKIRPbc7iR
rrK3f4qEM387u2n7PGOLdge+1AD29gG/lo2/7nmZCIJD07tH3jTUO1SpOlrVQaty
NJuBw1MTLE0GhJ5DzXgiC10nDmXuuc6fvnXjJdUzCOIF1o1vOEZfTicpiha5bVpr
b0J5PrNnqJaZsR/KJUqM1jMr9SnDJjql86Lufaz0IcnJ/t9FKhRGCcWdTBSJ2pp4
lwLc9nhK+uyeJiwWrvH0JkJgOpiaGSRBOEwJQehsdKW7hqi5g2xPo1hQqOM4G80K
tZQXgfn7oLq+Xzw8sJYDz4oaMo9ld48RUVgRWAJYQFY6EbWiHzqPx3MoQkKSVm81
OPosptZYoEUN31bDGuQ5NGMZnQM8XMoBbQn/BYpy/GflSPmpouqlK/CLDRDjY/aE
V38OxtCfiCJCM3kFiBcgon7oh427H6RQyCJPMr/dI1pZf4OS7PPP87HSAR0fmsYk
/+CBckZ964qIiA/yTqw28+78xY/1rasdNbdLJS7PQFm8n26RNAWxjygW6OGVumgZ
YNdNZurM00aDazWM2z17gh9SP6+eGzyhHRvSYrmnyxEGNC9wj62PC6Kg4Bb9Z4tr
PvfbjgYx+AMEPfI0zCPdwjL7iEeG+4aTkEgIQbweEPPNwMcGGPiqvtrOhowSlp/o
yLqb/oSwkav8Mmmab+fvqR4zdnaW3sapQCJeDkAFWKlvg6wv+QjipZQmc0ji8i7X
+Uqr/6u6u4yGN8rNwEAC2lmmG2STOP/IF1+tAGKTdr1CN6I98gyyJclGOyV9FbZ/
0VG8Az66/17do0qert1+NyM6BHzP2KLR4ulKuxoVeRrTdEGZSXPuBX+RXpQ+usZ3
nDKeurSsRAHnbJ7ugbpAliqfoV9G6iJkKN4bcHYnwF6oMQZhann/WjTfoae3hsbD
6k9oMQBJaq6Y+okI22pncjKJckEdsZnrxyz7Zn8Z888dbSVG+K4T02KznqoWvrLn
q5Ex/Ntc1lHW2vPluVtyC/SdcMN+XR9TQGdnoy11LjKzoDvvI0wBdJJ/3IFhTSrt
kDfOam6QDzYeky2N5dZ3/CdUc8rcWiP64wxgOwgMS4duB0fF3jkCkTFTvxSlsPAA
FgLtI/077Y/W5ALIQCV5/+DLM+G4injpEi9SUb7etpnbiqhXlgCzPCKYT+5r1lKH
pdftObbinIcbFCgdmfPtJcELcXSn06c9pHglSUj2C9lhgkIMPaJ+bww8xhmqta18
HbbuIJJFCprpVNV+eHID20vj7wQ4hB9fbByLRTilyQ1AyKLKVOlgnyjoykbZw7z3
Rd2jRZzC0mfUwImB+WnCbBsrfcwDo3EBF3DuIk48o63muzT+byltm7ZwfPIhsZug
1umcowpNGLPE0tHun2K24UOaU5dbiTfHY5d8HlskYt7ZySONMc2AuB2wrcVHBlx4
necychKEMPGAczNsBksbKc9jbVBuAWX2YLI0u2eGU2S9Fw6SX4Eva3ApFeaWbepw
+SmEdxRnrMolHG2zkv2zOt63v3I3En7j9SoZ3d3acceCIS4eXjPZJu2AqrqJJKdr
a0BBm3pIZhroKE3TZgwfP5C78xriRfIhSQ+aieUS0aK2qkGz9Ua4vo+0CpGjb04E
wTH4rIUG5mUpcJblx159mhSaPBuLlEhxQ3ZXX07seZd0sG/sa9z4gptxreA0HR2i
5nE6YYP5070f0sjg+gJUKXj+4LEQ/Qbp2rca1NNz1qCXOpRLSQD/kr3PTy7wnvHe
hBQJYELVbIdKjID5hStMONBl1IEhG6GVQN+zO1AZpjZuHwvcR0wohNNwuvmNIWrp
B5zRYN9m+snOmLxlIHfeWLjBmS9Z527TIa69QJwYkF/E0fEOBWJ0Vmqa/E0vr04P
gN9/jM7huOhU9Tfj7kirbPrezRwZDYfyr7ouhnSko5iFa8MvSgcZ4m6fr4NQdUNq
n1UtwUzUHjJRKcLCVeLBCOeCMtfOUEiuE+BlAytldAzAzsYw66W7ZtMT/slqH0Cl
jVCic+NyUEaBd34TOWmNbSaClTLpHPuR6A2y58lx3YR9/4/vkS1FFGriH+TgohA2
Mn6MvcQcRfp7qbhy57ok4fZnrJmDJZdw1d7q+w7egtRkXSKz2Nh8OWv6v6HjkAiP
hwGIjTGvHNrxTrd1bhvOyYqxqljC7buMaz3GyrLRP/gx6hCkLXAreOKQDKIqSzkm
pJluVkAXQl8EprIx8jSPygShMETvnmsoOztfE94nHcjKyb1hbvh5TzuRLIJSY3xv
iXrz6tKBQDnJist1HXJNGvGIVm06G6dZ/jHX0xduDi1x0lkKu9N+NLVx0eXl9Jis
l//Em5qkxiLMUw/pOqvV+n6om2S8cYWh+g5zivpyX4vxklYlao/mG/YH3YnVebVl
BscW8KzctCb5Z1nyEY+FHhlm7GlspjuNwjXjS1Dx4Bm738mgvc/LvgJX+u78JtaX
U2ltrh9eeGd8d1rt0utI2gXL5tV93MxxXtadOEYPM712LChrLgSQtV2N0MY4Vln8
aKGnNQoBsywosZqpNZjbCfb37nsYvtvr4aM6UMk4P2myVTFJtGNmB65pvkIN+KLS
oEVOvhB4cSz5MWzrwkX1Yw7e7MoZkzDUQtDii+ROnARcF2/tn243B67AxFZ4Bd5p
EziCOGDJdpcIeAl8KvWgiYVBoJHqS5mylCQ0DCdyYwqluEL4OZEjNaE1WYwhExSZ
jl/27WRvSb2Y+ZJHI9kjcIGbVN98SLnuV65H68sxOAn9ciHHqXZk0EuC76V80HHT
MJvJkiK1/EQY3Irtm+9L/jBiGehsTrtAEzPbdwSIev2G81HJBGFpi7EuIDL8tXNT
se9b7T03Y5jPbx2YQi8BXb9+2Th0udKK+8Q8RMqVFKrDXTtw30mVAIqtDDCtI5PS
2coWlZy8PNdfV4ycwj/YLVRiHx24ADiQixLBEWkOLqkttagLoX8N3RMGpeR6/DWK
xLRfeuQ25dxWpuKsoAaqFm0ZsuGxJ/2gurAjWYtsQszMtwbSOpsokWOpmDPthePF
EfsNJqw0fioyzME0KDh0P7GRXbd4SZiY3ap5tMOZKYgEQPZUhSI6XS5YUUF7ffni
cBClLsk+NacCZp1nSDlgbAjv64MVwyA5wGcJbbfpUHebNOHeWr71J0PdYfnU/rdY
67Qq6Tmyk4jnjXHDQcZogz4a0he8lAoKaKqCS7dIFpVsbvesPm+DFwZlrGRDb/3B
oG3YGOtlpOII1hC3zeDaOuMwHupH4h0FH6FEcrXlMDSa2OKKjkBAD/WYhroK1kdL
TrJ+Jf8v2sUDTHTAgwLUuDZXBiLowgMYV9KTkO9BziBDStvIMf8b/Mdwz/ofSRkG
EVYsqmuUV34uXP51WXjPb4eq3Z/2LdfICqEQgfQXuDlwL2OTH2hgOuEjdpxfHVjE
FiZo9ucCp0nBbnmsBefmAUFakMB3Nd2xdkL9CmfGzO/T4wkX3Ge6ElOEoI9S3Em0
7AyHWTWLHFxv3wgZoC46vpjoX89GWARmUu6d7zuRYlKVxu0ZVpuNGdDWGib1zoVi
lIfqWQY1K01px6M9vSSXZWtM5vARVU2iQ1AN6Th7O4HLXFgfq9n0bCOoyVcPkiRC
zmfxQW8JEx5MVPb08oSAiKrMqAhRt8svL7Rn2o9mjps=
`protect END_PROTECTED
