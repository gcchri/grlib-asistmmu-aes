`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wX+DKeko2RVE64KAUlzVXLEYjY55QE6xJwFUpGoHz39Gu4GZ2CzsMIUxGTZpz23E
onoxnIi5HKu3E+XIzj1Dfu1z9Ux4SQo443Rp999Bk/IhstCDHKGNjDcbjXz/txml
8B6J58Ksm3EL7E3hCPNBF3wDnlQ2AsoETnJxcu/PKbcZWpguwuVz9lKgeCPxsmut
HghTFlKlSvahjcCfGVxh7ey5BK2Dqqi00IuHDNidurNED/KTkDJPgnek2Vz8amEE
xo/EPaMCRlLcOZnV6gQPF3zNvCHbOaw96rI7+Oo82Z5HYa9CANeJJ3m5j/CwtSV+
Zswxpp0i5lnaUAaq5EPKItDInmUMiCnKxFPM0seGYa1/RUYuIFwzoULRyqVSAd9f
qSXL1xnx42nSUcH3S54+KA==
`protect END_PROTECTED
