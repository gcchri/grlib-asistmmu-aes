`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ke1H9l0FR/CYJHGIvYc1uu4lpsMNL986vV3f6VP2GqAahvBV9gOjEULrf7iVUnaN
0XuzPywTQOx1RwZ4GbypY74BTPVVsghnNGaaGozS+7oUviuzLPlFyl/0DYgOzxHq
FRlrhIJqDgMIJV4aQoEeLxv1wo9CKucJDO8Hff52Qjft2BtSnjdZqNDzi/2OlgSu
ZcVHtMclXSMaDKktbKVDiqubspAKvR6APeWJw88rizw5wUOMEv+/9pJHuvK/3ehb
+Nyagqw3O7H1qZhM9WQhsa2ea3Qd9H9diLt/hkRI7HQfWZsfyDMfvpq4YW2BCeGa
lNXgLmrHJA2zNHulJ3r6k4FhLCbVvaTEvHa3x58bbsslkFaHadWdu66Ny/HuGYe8
cRNv3JBsvhLN9VxX8Hg9SIwbdYkFYKgztDjNxXUuQd3EOQCd5QsEv/6RS7cb8a9Q
rc6jewUNVGEDhO67VVmpsCklnEDKYydNwZKDm5RfNPV3R3bHbgX6W0yObyJDf/1F
DWRHgExqGfbt9N76zWcgtmGEbGIzrAFxjbyEOn8nlBqi+Wl2tX3hrT6mDOt+ML40
KABWerC2012a4RKzT+W0XkW+nhFb2okbmMEeJjJshUaOOpiB8oUHqVHZPk1RS+zI
sxe2C80O23IPmyGkVnx0wNxplc6UmR4TbV+ypF3d30SRSooXwaiPnfdv/E01h41l
wKgVvCMvkZO0oeubDx18Q4UGxwTxGAOzD1XHEI82GEyPTXdM3hKaYHUVoItNNQYV
3kQFS5uFpzRLBQvg8e8VdB1x/0UlqfHHgeTfXy2D79uHoAhz9JgXfn6AsMPJYvJr
0L+e8R4VVJF49aJjSEPGjc72XxiIoxnCj+fxXEO0375toy7Op4N35ttmzyIiqKQd
+6Vb7Ph53AcOsTCeSRKzfVoFEP2VA2hWW+WCSYZub+Tkpps7m5+0QEHlJ9uwKpeE
fiThaGZQXGymelIWWrGnkzvddV8CU0iTX+BaV4wAZpT+3iA5/YM/bg7SFlcJdUbZ
stvNTZaZ5USKyi8YhSl75filW1WvVME5eZ1ae3/179ZWQ4CBYqySRAcqqwgGOxm8
eH2uxkfoKiq2MidQX1syns+h8ppd7WF2rPfZCxUmEmMROw+GWUmDnMJZw8/MUTaM
L/Qt7kKnMhfwZeHypm9vLDDYe051QKiwrL/afd27QekjH5wOpIYix3XuBqP5Ulqx
nnnUfTfn/uy/YCsC6xeurAJc5XHou0apKeqnHOJiuVWtoPSf1Wq1IECwOd+TVQOW
QaYRQNsShEM48wxtZxDbF/UD34W0Fuk1wa9at1GmrO9t7SNC8hDxDqwQasCgYHQN
7OnGOKnmeJ+IGMWYDd5eQt29s3T3ik+OzkzCEL1u1JXSSd2ybm0s7es7fLXVB2AX
7iOJ5zaEdwsUlbHpEF6R4+FwfjE57lWF+kmmwNkZZpAY/mH++zDNtiUXISct5p5C
2arcQhY0oC4TW7ByglfdtjyHO6wUAHRassco9ChG0zs/GbV3ruudx2MuINEhpLVy
KC5lEfmArsOpFLMibEhreja6eIOh8zKC0hTmgrgVn8eDlomJSghJD2lEVa/4EmSb
S4WLHvPOBBPGpmiueSxdzhTvY5YH+aNIUmA5WBvIdMtjYdG/gj4jzNBRw6LN47QC
JyhZ8WmS1f6r5dOuM5qwR/IgjWWzk9s9XzaWRH3d2embYpm2BfUTO20Kan18+XRb
zrPgmAI0rG7oh9FSt+A+Wl2s5NKMYtpT5o/G82jgQCsY1w41LMUm5ktiLYRvXhCd
fwcv2HeJ8kNmlVIkgVwv/+RXPd+awuTUv90KLhrBxlMxgRLyrrk25Ed0Uiuyp8UH
bBnTaRC6xTpMBQ5zjuCI7Vqitmib2xaY5HSpXfFtqqsQQ80i4pV/VuNT65EhRtXo
edWdk6Z5mPPnT5XxXWNNzCecTJiFJLl8yl/E2ZE0pPpXKtJ22MGZ9C1m/ky03r/O
5TSpTkefLCwl9mRlodFIYbKKRK1TtgqxavDV9e8BaT+oPG9uSXeM4RSirvbpAquO
kRb2Zl9+MqFT+24N+u45yAZeQ17Slm3k6KOY3JofRxPgrpWVkz8LQU1SyLwoLC4Q
RtWFAGilN1lE3424yBpvwBv3GalY/5IGdmJdyYdP7uBLTuimbZgrkYmQtQ/W6YYk
i6uq4WB1+yg71mXCeXvoCwak8K4Lp1ZlaoAdSOUDIs0PugINmc5Ks58jzUNHNL09
0RugNvQeG5WOWE23JfsOhoCLxltmZ976YmoIMMF2WxyqjhzMbBTo8R5pbOg5kSrP
cm2j2QNLr7scGCBj36DgiCxP6VxiLxs+k8TztkUoZ04HaR5QYPn4c2rm42l4I569
q4dcd2XFJH6GnJVFTMlxkzwY0hayGGcCDFqmzAoMFUbcuDk3ZO0YfYRYiglEoH8N
Rx9jUP0rgNvy+QbLX9gDk6xFeFBzudBv0MAa8oa6kN5xM+Q7FQ8cnBTrZAXpUIBb
A9IYO1sNoQEd1GDxDTLBQeM+3JqUh9dwOGQ5uxIavLBAzk43hiHBzKQTUkZJ19pJ
CiKiwQi/99VVWqeFrAfavx0SStrR2JmygVKsIqgCJN2r3lLavfxUVlF7h2jxumEk
jHGjT5TthxtVaYhbMgqxmLz0CqmXhUSLtu6XxSaFyYMnNOtrTO73FclnSDUdxa4Z
G2Z/YiI1WnyRlQYcWBlVhv2H4Fc4QyysOr9H3BKNyYsCtDthHALWFHqEzRbIISvV
FjkekqNAiFmvwx811ZTXajGU3SgAb1mI8kaEQ9kqy3ZeSFdNx3RoABc4b0e9ddTa
012v6jyNlbxoQbY9lxKp5nox7swRvmGfdhmR3lXT2S0qM/ahmdQ98V5XMrqdSHuW
GmvV3xIfWyh8TJpkysTP8eiwj4DWdpzx0ghYMPOiI9CxKIQBF8tOb/zW7iUilh06
tm0cnHRIsQmfab33e0U0NIrj0ucyLKls8UY1ivxr2bSDCAU62B7ZIdH3DYUFnULb
qTQkjHz+5nfdb3ti0tpfR/iUiEXeKFHSC0EfbdUWePIbsQI12FC87QLU/fO+8bob
ymYBGefH2HwUSK1rAABOSK8ATtqR05xcaNrehtjhHtShDb9KgSCvefGPcW7W0vKB
tdCGA73NZqZWhyDaumMaDw==
`protect END_PROTECTED
