`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CGfn5Q81rwWvtQ88Vrd7WutyKzreaS72OOw8Yn7YJYBpbaKf9tMXcZzYq8sfzuQG
vES3lHgakc8LbjZoz1K43p8XrNnu+56Woi2JlrilLUyVuwYqq+/pNlgWrnhc+OfR
TyoE3A3878a3RP68ikuSiDRpTDkrEKMgqE5OFU+SwbkGhnPUZqJoOETx73JBTeZi
Cb6hYZfJsX3l1mfJIeQctY756XmG2A7FLOB86Jwu7SAQIkYIyrfMey0Ewt2/c78N
Azuba/i7Gtq+A7ONm9/LbE8izercNYq8D9reIo0uZMk=
`protect END_PROTECTED
