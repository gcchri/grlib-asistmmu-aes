`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
spCvyw124C8TlNQjzvsv6OTU0zD08Q2kY9MdXpV14SpyRMSvIudhhxaUoAAerOe+
zy7S8XQqL2PYxSHjaJfemDy4DdBEd3yaBf6EnOMXpBaqTUbzHyKaN58GQyqwqDoy
EsoHrW90JvCmjcRSl7wIR5Cm4PL/SRWlxIqUUSz3N0xceN5tw+IVXx5EEt8tMPXm
plSH4R/AqBoNYzRJO9l2gwraOgrwPJJi9MMkdu/hlaz53eG0TkOjAZL6EE8k29o7
qWESQq80AH95KI+58Cr+gg2kqSI5pzt8b5wZoHD0uLjwzS6gVOxQnaTsJK7poZHZ
SjHzoq8mdVwDrqyx1n80+nm912qCXW4W7xJ9MM8jcVnPuDF83PXnV+nSnIvY1QHq
IUW61wIFsQiTaAo3VKhbbY7mOYMZWaWAtGU4w2jjZsPkmdKHjKz45/INEg48lM+E
`protect END_PROTECTED
