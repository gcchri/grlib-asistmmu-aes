`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2rZxCahdgq3R+IRXukJNQTeezS6NIUlEWelccOHf6Yoio5WejISSTYNTvG51COT6
pI6L4JF8uXaeRrfQhJpPc8Sgxs7WTMAV92GS+bnFOya6dHjfdriaANdYjTHtijqM
qzYdRIIGWSiBLtxr2kOAhFbxrmSJTA1Mo3euDZ3Trphw1jW6Xp9swudF1GeLsEwG
2nzj+b6nsw//NtzmgVB2oFs45X4DWldQ8oYIwhMIYr4FqAkWH/QbryrUBsDyz6SM
FxRnL11H0Y2Ksyxrid3y4EYn8pVAGcoOERftsUYzmiNnOqeHZAmOTPoYSCuITAuf
4nPyt1Nk/NVJE1nl1ciBtyA5iHcvtjI728msClaxql6890kwFW046IQyquxl5oFF
`protect END_PROTECTED
