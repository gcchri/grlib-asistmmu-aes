`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9zjp5yjawfm7ojHfTYJyuCswTW5aQMTHwgquSvJbwtVDcOEz8ok3yztpejzlMUL3
xYIfiCrxTb0P7VL0ZNKgaPPdZ8Wjx1y325atVLY9h5Qxf7imi+kXnebOv52O8PuD
U6FGnrXbl2WkYV62EPEE4kH5Wpj7AMaG5bHE63m24an5ccwhk9c3HaNncD7BUdZC
OyiZyYE9+B5URtWMstvBBuY/kVYBXzYU9tbbuadMGtcnlL+E55EI0HoSf9PO9EMZ
396tUKP66qXbS/F3NSR/oQ==
`protect END_PROTECTED
