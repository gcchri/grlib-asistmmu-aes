`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YRX3bZ/FG/RlGSw2mNjdV3mOT6E801EnTVqUhc9YGA4u3B9Rp+Sx8cJpkfT+mpW+
qQvYg3j9kLfQk/TtJKgp/JIpUdmGNMQ6Q6p4BGh4AILR3DR5FNRGDFfqr/CFILPl
p8QyGDY5jd/zy73wDG69jv1tkQjcdIA6R3gcmUKgAdc3LgWjNFCJU/afR5t2AiCP
tIQS6oGjcI5yyuit82ED+OpkluwdLb4Lmc1ZH8DjGv4Ssd6k/A+qL0guiaPeA6Ap
dOqwTVyMUq8V5zXG/Ho1NxL3YVfH6v5eBg5tR+4xyrWEQot0GxcdMOSgCFiZoBxA
hX9muFHBRXAgfZMxSu7wiA==
`protect END_PROTECTED
