`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cyVdRpadfBNzeHS1L9pCmMz8D7KaA6WqdbcYWhYO9AJCBA1Twcmk3Vs5denH4ni+
7lEkZJyuRGL2diMZ9bOBsTy1wFDqwlh7iepbPFQ1/yc3ARjpSHqizYWtvnYKAVFs
xrbUAa8WmGQ+uciyyRQwRB9jvGImV5k/5ynYBS+nHDjm9cWP3GngLvviN+qRkl0m
5fQ9ZrbGnELisIAzRNoLGEa9KxumAv5cry4Q7G5JnLiuFVSqYR3GQkuvyYKxzTPl
WPTNo7noo5OubT00/bAcvpCRBn0c5a67PQ0HRgEVimfs7Z8YOZXHZByXIA2izifP
1uzIFcq7K20K3wRXzApY5hTxz+8m9s1XQQsx38zFrbizFVpxoeoAI4fNO5APpLYT
DxNPmpbLRXgqHDXrbJqc2ipAX7mcsikslwP8/Xq/sTbRQeI09f5tNkqTAp+vjBG3
/UTDdDzhAK/cvbTtT7adC2CJZ38kyugpzSqvIh8ladO9ujKm0WLXMjBr+6LpmW9q
m4YY/f1/DbnNb+oSWON/I3/Quhn9U2xE7IGTn7t+7/v3fNBAyYrNecVcuv8XdcjX
BkoSn2QlS6Y4alSNnOwOZuxqun6IB8GrpQkliZbbAUnQE4fQkhiot4C58pxypUuv
K08OQZnpncwVmrwqlngeYYjIKjgA/oLLfJej7hYD+nmcwkbxFHqmJWpoY/CA7hVK
zZG0xZ6S3DEn4iSe7fJwpQ==
`protect END_PROTECTED
