`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uv5geCds085UajNyD3774TDZGtWIbDI4mKvK40NyQP+/a2pLxL2/c2pT/8Lwvk2H
8CKTQB1gsWoDPBz0NPLO5gBMIgevvCPawo7XR3HiEjuKScwalbYi57C9a51ravDD
bgLX2Wn9mvZPKVOowK+qAuefhA4Aqzog16kPJywG63+2z4O09HP1Mdf/0mwSKMid
wUfJKYmNzx0UZJDDHNtb3se0CNfDZ+yTVX75ccbKIXxfiammqoblMQFwq+KqlZeI
3UH6/oCVUO4hz4AwclkT6dSrfQTASXI0a0qEYEeRmOXaFQQaSMEJsHP4AXffZXJh
PwvAWZ0EYapahv5Djtfj7eo51+w2UjhZ83T132Hl9qT2fw4ECLTQEodSi7xFL56k
HYQOF6eYmsa0OZ98aqsqjrO/bquV5gShQr9CLZFBZ+TM4JK357BEjDcbRI+1DHAx
AKq0ZOznKBdBUrCigy0p1kqhHPKt8u53l+fkg43Os4I=
`protect END_PROTECTED
