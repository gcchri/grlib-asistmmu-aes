`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O7HA/P+ptIVNH88MEHsytQJOCMV9AHfMl0TRb9gi9BM9fEWYObDsMUkJO08LrayX
8K95D8+5Te1BS1/swZMMRi0plM8aDghVciuPkTTsiucN7toO36kX5qyPu2DT+vbI
bKRvCbieu0GcLdm7xs+GoiD5MpxiDpLh6mDGcxcgeEHZGdYkQq1Gvmy22fL0wz3Y
XINud0TGJCk0OjML/4586mfd5avsnbuq5BgZ+hAgxtizEHVEM1tLLu1IWdljSlR6
Oa8Hb8cmoVXFuTVVoyPQYM/FtCv14fLjQ/Y1qDzYkFqyUYtkAWtsv6gvISSAQP5N
6VldKjcFNISfbQWYgmvRzw5i4lp28MUMGEyTxw/CRHrogaEQlH0G3tPkkiT/Vdsb
GgE8X+C7YvEGXJ/hPAuAPnQAUQeZkzBeY7ceTgjtS8HO5CLdRBTUJguJ8DWabQV+
st5zbLI+JSFu1gHjY84su6GZqKEPM06tO8fJE5ucugwT6ZUucjC04OmsmKTQ61gb
aQeMpS3lIhRT05/bTYKXRN3URtiptP7xUGUUIGoF4i+9f3aJU1hKlDj8VwPeNzPV
NOZIitJdyHM8iFB1x2XJXnz96CXfMRQcng2XQaFn51Q=
`protect END_PROTECTED
