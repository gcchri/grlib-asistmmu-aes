`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O6QdQ/B242nBcqPlMxPAO6mXCWAPenvEnBG7+poX5ysvECc18AdtVF5WyI1Lf/ZZ
0BuAJRNK0ulToM2y0pztQeuwWnxITS+I4hz2yfUE+aHtUQ2KdWapO1WbzMa8ETpd
okcBF5wR6/LfzQvs4uGH7sDlPikcLo4u9Fb2DVMcuzzfu79LH/PjJ2kX5Pg5ie04
pWyIGvOkZs7eGeP6OKFOC9hpxJerJGs4Ghw7u9GY0txtDP+xVC3wMl5tydLzMPjH
mSQF/bj5uwpePVOqW5sLrpuSr7XMMbgDZN+DGfyQQXLZiheKG9O/Aqo0Yqr6gRmH
OClA9yVlkRIRoCurWxdNYYNvMF9dycimPHcd+83G9NH/L0enEMLvXgBGmEmK+UdN
uwMpzDhhX8LiIFeT9BJQJzz/srZhxOlvRPcA9pdHzyrvT62fgze3vAR3I4N68yE5
3KKSc5QPuYIhIYxHVnjGcNvgBVEd8E2J+dp6YtvTa9jkRAzWxIWWKgkntL0YsBKu
`protect END_PROTECTED
