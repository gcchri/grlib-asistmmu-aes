`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CHkSLEB+rKrqFxCNHaLP0PcItmMjsVai/fxd4C0T7q2lfJeyuIDV4I4vfz5DOoY9
PH6Au4q1wTb5Z2vSU4mhWaguYdRfZMBcK/OphJ1KAkInJbupN64uoLctkvWdztUN
7pKNid2+aIUc1DsRFT+u87LEXqVgzg/ZKomGf9zL03pETbsdDLQ4UXppO4uXSOYo
CVu2LqtJdXo7MSnJELJkY3t7/0y+rtnGfY7UkAY1EDNClE9XVy+Kxiv3eGXb0eW2
3xY0QUTFA5/vVLKLb902QxsSeBw6JxY7HcjWXGNaCxOP1q0W2QIvmB/Wu6hVn7v2
Jji39D9TbgNtemr55+xO+ZM7ZKz2P1nlibFl/iPKLXIaNNwhjWsW8l9uq4fnZne8
Z/42ceHmEPdP2dHWNywYVAZI3U+K2nYl1AW0vtDwBYO6atLmZOuhnoHR/sdJTD0V
vKWAOEIDwOHVQYNlBTIBllp6ZCvdcu+qJuzd0ZRPDyvFwPaHDknZcKFTlEiv5IWB
`protect END_PROTECTED
