`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JfNoCstlUmhosRE3JZ6aVdFisyH81lvogSfJUczfA5gp3CG10jEz7USQfFnlYRyU
juutdBkr7J3rbwBlr2og3yoGt2Q/fNFQzGWGeIs/6EEU3YIxGgxdj6ieb6NA6Nu2
xBJdYoOBBTr14MHEosKNEB7qZZSmDWpbwwsqBx5ZLvR31UlG8JCeUDW0LPGWOwkk
9HJHDUnPdp7uai/+hEf6D5E9KDPGSjIrw6njvfrovz+FOhLXh0zP8hDqbIx3RpGw
+uBReXXUyadv/IzTAeh5ebhRML8FK9xjlx9q0oAaJr3pe95DtBECPMaK5KTBYPmJ
4pel52apan4fJeHkaxSVl5/M9cmY2ttsadAdODWFSSO4hEAajAPDBmfMt+Q+4pVj
50/8nGNHGJo/eZksaV86i3mzuzuVlFsrFQP88lwRzt840LMm6AFicOAFG5mHP57h
FyEGTp0Xdyqv9zaTnHN1Xy1tj/zda2cBUviuQ7OhTThCma1hyhHlLZRpYTNqabGS
QNrgW2y7Jr9qgvZgKN5vUfvlV33IGkNrzi/M1Jn+nryHbDaTdXcUvY10P/6qcnGs
bxnXFvl5R0/rgVwgo+vhn1AaQh0Is+xCgyP5epTkNt2VgGpA3cEsByOm5AvwtJQy
O8of1MuGYT2Qk/N8/y7+HR4WV+IPnzkegUEZ81x4RP36vHFwol+37Z/m12C5K63R
AnnEITQV3P7Al2TNI5JtomRtINEa2WBAFZitOgPxZcEODaSuP2oitiPb00Phk4wt
qdc03zbPDebB9ywjK5fUpoB1U8Sg1RDKSCaIxPejQWq/gdsYS8p46NiTKY+bxbd/
nZOj3lm0FSZfIaKGA2HStUDoejirpAFv7QAdpMyR/H9dwpJCchWqvOh667Eq1Dn6
oQJ7ahDRHg/sEYX/aR8uFGup2J0lFbbKGqASQSHgfWY=
`protect END_PROTECTED
