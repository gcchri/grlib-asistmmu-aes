`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TeiFxNIAqXAYFKmDU/nXIYDmB6Mc2SRo8Uc6eQbu98i6RmtK7aWXEO5mhsNgSJUO
LsXhvXubimjqYJoRrILP0ecppq0yo6FKtnfS2TQf52JL3xOvDSLLaDzwHYil3ey4
Vt0fz6POz/tT8RytuRSks/9nRmrhNqdLIGhoEuCvBXfSTY79X/uUd/qg5POGwkAa
pplpWKjp956+0p4LqgAaSqtgT52OfkHbFflTmCmYbB5rBvzOSyogLHo+ZI9EYqgd
9TyOrltcvqwhBWiFq2sdCXDtQZqN7I3tC1zFq5fs0M+ihBJtR/wd5ZDsQWDsMahB
HrKY/I27XXoBYZx2UAvEIZEoYr9Za/h6u1Zjw0JjrE9r3CyL6MhOZywnOEqKLg8h
GtUDUxJvEUvhG5uk1iYDdcmufWF7EGOgsO+zS3nH0GhFi6Zviz+FQl3ykFatDSHe
UKOu/JsCsqtVWF3/5WTge9JsaZ588gv7f1nbyynlv8dhDJ6N18Z8x+kSwS3/HLY2
NJBNqeIxhgCQWnQrJ3mUKQohK5KeAtHbZZl3+GVFH9tWty2muapyQzfo4b/5OoRD
`protect END_PROTECTED
