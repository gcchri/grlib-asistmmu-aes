`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4r3kgScHcUjlJmf7UtzL1TqoODMtEI4BNlL9MIXE7f58ny/xzTnTeNJ7HTcreFbz
QBMtcjxaV/gufvnePkOCqO/zK0SzCkUfPQ4TpLNwASYaCahjtupg7TRB4DEEm4LI
HPD37f84XekLARPbNq6Cqs8irRoxWdc4TY3gMFS3AoepGzMpFxHPcc3e3qe8eqxq
7s5NtMiS05MMc7/lkARevYEpI44SZmRU1njZVhiULQKvqy5rypEtl6BheI7VYMdw
gnuYlsE2rYQ6fc2UoVl/57ZGOTLIosSvcxNxNdVTz6PxEmxKHLrEG4ueduKMi2L9
f9yV67kr4C1g+Y6pWVXiWrH6VZrOzL4OdKtiOQoaMeAEEdgWeBPK/0IZNC6ds7X6
`protect END_PROTECTED
