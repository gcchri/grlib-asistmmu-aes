`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P8gbl4HpzgrhkP8LyoW7iFEfzngwN2j+giejwTSQNxifBF1XllD5IJOaCIDfw71c
ymdQUajJWDZxuVlL1tifoqPdf0VzOF6/O9I2ivvYUiH+jYlVq64uG650EGTYSABi
exh6E4TM+b+XiGTRo3mcuz3WxNtojt+XpZKWnvaFYax+N3gzSL3PYZmiyDdMl5M+
Fm0qTjPs1dzIVi3OQLXQ5pbhfzT9AyrXnEJc4A0e8cKJ3FoUk+XHPUvi4jsNsaBB
Jssik9WWArgbKLWNEkrZXIv2fiDf+/Ct9nVRG4J94JTKyJtDb+Zm+cJY1pSogeFk
oTJRqsgiVlbtD/3EjIpkSt+8ly3FZLnnLgduYnhfYXbg5CzZbtF7NaC2hxNd25BD
`protect END_PROTECTED
