`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
biKGV1VoEZVFAisFuOReRgDBCTSqDmxwXdsq/QU/6bJwU2JFOZAZHxZouojIwc63
+ybbRZxCKE+bmw1Ne+UTwIYrHPGIzHxlPm/EPPS743Tz7eopSsXH4u+OxLzfS+YW
KD7l/jBvHZW1Wi39M490Xwb2S4H3j/oItmjN5Mcs114acKCRyt5CY3muyD0Hkoev
s7DR/tbSM63rXsbcMip8T9no5dHaMGtFi3mxRGBqbQkfCbM4fZDWgvOU3Na7oFHG
AaT1/Ui8pqr05y9NDmZ7zw==
`protect END_PROTECTED
