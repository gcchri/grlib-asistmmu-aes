`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bmdyi1aColFculveKJfHoV8CLjVUU1vLLp7//LZtRye5g+HuVxyED2atGouBq0lC
nB7s/CeDEatWydp6cM/ye3N45luMUqApe5eKqFovZXP2iDfCgmcbNhrUpRrYUHmc
rY5p26TFAAXLmbOlynquJTY6Tn/xKGRybaBoF7JumvANUlawiu+LgPWW+lVR9fKs
rP8ThT7VEF6od0Jhm6j6Ui4pJppSRt2Mw+asqCUemSx9rqHaLL/QaFVUszG9Ezr3
rdQFMxD3z34frgRR+QCCDgO0M6lihgX6ZFfGFFZ+TN3z4McqFYndNc8VjHCc6saE
`protect END_PROTECTED
