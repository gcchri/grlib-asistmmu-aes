`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aUKXcVU7Wk/XIsKhUOf9uONVT6kDE3zrV5NL+iY1EdXkTtHvpMVmZ9mxEjf+uYaK
DV+JoegDb/QgoxS4R7F4m4QO6JjcRhEi/hf6fV56/UWLnpWl1NuJrt1KaKAdT0zX
rKQ9Wg68QNqi9Zr1L9/oTtFF83EqMDzTFMd5UtgbMNNDUu+y0Fbg3+BxLn03tFDf
mVtXkGeAIsIhdD4CSXfKCm4itLU57vlhG+ahpCdCili4YoDET3r80LbINnvsziBc
+rtOllY2Gb6nu4X6ovS0+VwZlxe30u2WPZ66ib0LkJum8uqpkCjLI/lwvqxrNfkS
frhMr8pQL4C1GjQM5kXmmB2LVzyUQuLekycGGDjkLS89KZYxkkzDVcaDeW9GRCgK
rd0yN0c/+zKG9aaz12dbGg6UUdDLcGlbq37wR2dbMf62ZXM4DlcAoohFhsSsOCDh
JJpCoM6qd5KxEPD0uonvJFyMkKuDmxRRQWeLsKooJAqOCCQzCuFBZT+lI9fvxh61
i4QMxTIiNk8u1oUhKecRLvTjsrXaFMrDmcx461OezFYnpsbdp1zml011PvLCXdcR
FD8Q8RecAl/w2seTAAD3MIRU3eWD2Lo3EEPPZvRLUIZ+PhJR48EtjWSqalPjGpFV
0j9dsf6OS/bOokeLrQQNdXak5BDxnlLknO/nIJRTo1nd5PWRPXxth+2zM5gb4ywN
IW/jVD21fEz0XEYfMj3xYs8Sjm1TiBgSsznvW+7opOXo71IOQbvwiTTZCLU6Y9Hr
vWO322291L6DvD2CiDmRP72ItsIEyMgRLly7+QIYGOJqwmOosbwRPl6iGgOZJKOU
89Q4WU2hXgnrjufQ5Dmzcb8nL4sP6aeE4+nnz2Qk0+JCCJV/n31MGeY0BABqBgcF
VJ9TWz2FJFh+bGKREHxoGf2tlYE4UCcI4qUF78BUPnFRdx/NqxovNQxXn/LRb4Ir
oeLIlgMKfAWwSoBAZkXnd+Yb/NBwxMWpxobWnYRag+U4XgXdSNrT7Wld9Tp3OeBh
fRdOTzfodnoVbmmPuum0cROJ3gigRPUhKgYPCDlymeMhLQXHN17LckipEvX3Pxov
M6TZc4ELBM44OCAlojFuFZuUk2Bs09xL+tOgfOq7JryNuPYUDShnVol5a9x/x842
PLCwKRSA/8BUo6JzNANAH8Mfc1Ygu+/S7X27h3las9zAVL++E02vfgx5/yC0bW2w
UXaoSpDh/zfDLHT0XKzjNJ81Uyo7DfWgQk7VTJJwwU0pXKmzlRRgYpqN1CvonzHh
MODEXmIw/vAQHzvsZLoRTHfBRSX6sSrZ4aGjGIgAr4AfxQEzU37+2x714rOmhTYP
OpUX/XIVNpyYkUQIneboUGQfqrLtJRhxy3kxpQ6jhPRv5zRW6jrRsSa9NEfwkKwR
xwJikbXXpExlaIfIXFRTburUjuz3QnS3p826XtDW6iWNzGg01q+Y4smq5kvnmdcl
mEi9LftyTVAAJQ0/MN91d3wt3lS1iEaBo4JrWcWHyDHTg5fLOjWYM21AH9V5Q/i3
Q/abmelpJc6n/dBDvoAziAm2U/neRpDaT8TGhTRXpARsM4iuLSDGJmPIMKo2Yr4S
4INrpnioe15T91+h71fdiq5azEM/vnQIlTED5Um2GYEHcKCV7vk6TWjvtkx9K5uH
FlYRyFTEIemswYnrJzL1c49KnHDwmfu7Z5VShzKmag40LbkzrjSnEGFyxBYLzFfe
oFXGO6+goVMIN0wrcZCh1hxVYDcYGSGnhIlH21B8cVHK4vD1hN3vqr7jMywj/bTW
aoT8Vx8H3ejcyPDvPN7Vq7k8ext1yAdDU9uQDAtm9CRbGHOi5PjCQcwlqqL91kQ3
OyGg1TeQyzETQ0SQjq6cvQJVfA6QMf9WIpltxw92OCwiDnLKjh5xlBzByzUg/ezE
YYgJckKhZOoWIvxxh7n/He5uzk5cm13YUpFTrtGL1/28pAd8aDmHxTMO1xeBKbmo
4JdWCUtYhDCUsWhxO7LZgUpC62CoyWh1SdOT62xBfhUjF7SJugPkCQJ/o3olHBjI
bz+hH5htm4jM/nwkD4eVnElo+5xU12lwsWdRknEQVih6RDmQu5Yt2IKWJ8l5bsj0
GqTe789DEr2eLf4DAO8m43voZkcTayEwdqmjeTSJGytBliEO+kuaWIvn5a7QBOZN
LNDo5T01OXU2+HYhE0QkwWh0zZcwmYZD5dR55RDmJWBn5Z8Lq7jJhRJeYWDM11LN
r8IZOBn78HKl9u5SKs4rD7ycJtwA+URrP/yihhEWe+xxq/6auU11qQJ8ljfAcrrL
NQL+BknMnop7xUbu9ANzPACdGFcSHVkFythzxYJAF9Whhk/xytSSEpQX/+QO1Bpj
YrNbG0iw06rWE2x5Zdf7xgwVk4KpTDVdH/k2M8T8sTICjwKdAioWsH7n8xeLGUBu
/CnwZ2dtqgWqRKbX1++lbzz6cynDJdYeQSlk67fFpsHw/+F5mbsPEk5Vjd1nmjfh
aIcXs4W+gmPcili6VsbTLrfy5s6MqEblsNGDUXdCxpIjpLQD/0c9duUQuaHw0JnH
Ygx5cQuYyou2Ppw4+7IFfl+hmdi8zeFtc15Iy8Qi4BABem7oUNIWOHVv6aDR6evb
0+q2kdU5EdddksOM5RKd/zs5pQNhnzt5ASDh6Z3c+sErWPQig4lc7OPR/xeQ8/PQ
nUQeOoi+0N0wmfwBrq8wbl9aXmU+mbiQZnzDoPAaeN/oDCZAXDw7rSJ4LVqygQWn
CI2Hkgi/lvdcrbK63+yXQ4EvEDIFFaVSwspUmV/0b+KL6Ck0qtYG1Kt+OyCJQH5o
4O1Yo6J85Jxof3VVZNyXecIqO78KG9x7Z+1lQI9JbfwF0tNhj1SMkBOslHKY4muW
lE5SNyJKhwmZNdnrRBnkfivTnxwxfYT6wDdYwDrWHfWVjoUp9fUXgxlMk8DmTLJm
FrR2R+lTQvvriia+QmS4i22Pa9dWbXoDwdscgrIbKGYaVmnJokctst23xZprkrf8
HzWVaSZk6p+G42qQEt8oUPZbBkdIn5g7230uk1lszIdhLzHSwCIzt2HkJahTGkow
P+VABOl4cq95lSvLI7hUGgEPutPwH+8/JGTQtPizB82wv6KOxFL6mHflKXquSYxa
P7BW+MXbzrpm6+3o98cx60jhcFWK/yHRqifeV+i6BLfTo+hSnewlvoVHO5QEu0pi
Mx3JH2+Il5bU7IQsbIgxxwMTfpBjHqGbcawpCzjnUUbO/m+SMxxiyF7Yd2f9CSS/
rUBJ0OS8LVRCHTrM/DUeaV4EACo9xqcYwN1X7zHMVuaqZBXCJ2Roa6fzPasfvxtn
tNRUT/vrXuXdjq7NCkKaWOEq8c/Toz1H8eUCfECtx9cAHBm1GEozFiol5DrD0Rs/
HBPDvy55+r3kk/9JA3OPZUB76lfNGevNIKrHomP9R3rzI5gRilQvmNkhYLzluvAk
LismD/+kynk2aIgX3rMmn4QJb8JVkKtVMqxX8+xe1dSBMgrepCcQKeoPQP5J9Ahj
Ur9qjiaJobji98/t5TnC8H4tX1fDHv/B8kmLK2T7LhZpLoYZ6d8ywd9BCMF4MRGM
QMAfyzS2FuJyH+STiKxfzwt3LZ2cuQF57YvtVozWBSQSQEOT5rYxyMEhQ5pMs8dF
2ZC075gLGcgea2qA0KLFcezwdnLPAGXpMxUTFrZBmQvYIXvxnLDpqwBFAmZx2HWG
Y/LzCB9gpnHq2mU7TGPpTllrw76qDxDS3cQOoYNiq+3OrnKOyagGvYrVpwRx6Xzu
YYVflM0sPSEraRL6Fs7eUP89bufBiNnUZ3Ohhxopc6ML5IztDGYWo0uRQqmbUgQ4
gGRTm2glPZPdh47wkIlsHrTDsI4w/QzKqIdl4Bv4Qw9mjJT9swg0NLD2SJMHBPZ/
a9mnVaMhckd/hNoH8BxLb3wOK0KmlGIO2EBPRt9CfeMH4ggaaBwA90tnBouK8LU3
wzlYhQw9AhSBklmFVRTQw5OMQrX/ggZeJC6Lsueoq+H2Ozhe5lcTTskHOfyY6ZrC
b9D0c03DwfYYDmaEK9pfN6k1U6DM+z5Tj/5aMiKiS+D04AQvc3tVZY//2YSCPrxd
mnKTCPKeu5dwf+p6nah1oDR3JYfepr/V+kzcQ2SgacQDNd0oPv+O5tAUnKAKzE6b
bsHoXMithwQhNdAnPCyDyQtQxYwrc2UqeKyKt6ssxk4s4NBy0+33hIjyiNH2e6zZ
UlJtfbDCvkNvPEQ+3ZMGT0NnO4VjMU9wYUEZxDnODnkc+A5HlwXKH5+GnKXx0Hod
bwWyIUS0DwDrz97oO9OJZJd37+3bjBuR5tjPgDfQJ/0YY1/PIdYctVNWvpVuaQZr
csOCTx3jaRfRve7ADbPGsMeFdMD/8pDx/sjy3Po6u6vCY1A5pt/SMMVTAg0PKgVZ
Tpq+dcs6r+MDSBqm7FazXL2YOMpFYSpd+OBaXSYMWH2pXKT0BHGahBlrnXXMGZbm
Axjs7yzYxRPd9flLA/72cNhxCgRaRSlce7J2oqXYhtQ+3l9/T1q1srkWvoLIxWtS
haW20VX6lNS8UFeKoTqidYEe9nXhTRBouhsSjJ6MwHafRhHUgW5lTqKOUlphCxmV
ckD3uFImO3D87PWd+1a9dv9bxW65pFUnik7RTjlka4ALLN7MncV8OB6YEIxHTsTL
MjU6QLkJHKzWCLecrtGvGWnKsrFgkMBEXyo1MtIO+y32cYwYx91+8+7fNLADud9I
pyTNChx/itD2KIOTHGFSdWU0/3oplVD2KRqHCBQB5OoYYkziKhttgJdmHBJJp2MK
NciUSprjrhL+b7A5nQLzD0fZzuT8iv2NrI8A0mjcOCgrIiWjiDVu7o6PykyQJFke
mgaAbBSBeA5RJTg4DTJRHbMTYlx4Q6PLwsV78Ff208Am68mAw800YfYqfGHqDdDF
GTk9plgyqWvcx1tCNpeP2oSedW/fhysBUL+bTC4tUb6KWbGislcH+Ig+n2UMiG9w
DlHWOcH03KHZPv2IMJxlya9hgFEnWkuva9YciePxPlhM8VZkbGlS2viEjhJSOqAC
o5TYYXe1WksAQbZV1pkGcbsz1K/A6eMdp9R9oduk1xSAXx1a6ukHy71WJzPEdvuV
EQQuMeUPwyqSa5H0cyQrW5hje/meWRLYJwhUswLeQMfVtQ4/6GUWYAlbUFHdhhPa
/L2A19XUK5I6bp7gZbicCErpncVIvQEtRxUmQYwFdVUlbDhfDxUX1ZP5mKHEqrEW
TctmE3sM/iR5JL+loJsPJl6Z+5sZBNnpPiOWmAgFYcmjzk8UeWR5dAayckfiavu8
6idl7n4pCKjBiQi1GFWquWk01V7u7gtLNKHDq63z/HiCFVkg9qEGo++dv7baaneA
VXXqB1SKwJpJRjoNjsmjtwE/Qu8XfGwJvpgyzVUK1ZQkr9Y0WvLAJD2Jl0qXp5aT
nuOgQ8neydVT6KC7P9Jg6wvxJzPM7EaAYKR52eGwt0JVfDVvYaptYOhbNU9pwQ8E
VPl6MYJAUOaZXDyuwINoRtvt70hxGcXNkcuPnUy8GL+JURBNvN1lZB1aLDqSb0Ug
AQ2v/fPaTvx3y8kPE9lRbCaAA6Uk+C1qCDyQ2C/ZtY4dT53P/eEQ25dSHya8RacQ
x1QhUbixcCxOMOWfHqBzJUN/wH/5YwQiZsZoK+BJmS8vfVB1JtuHbc42Vq7vOgk4
1Qrli6a9gBADQIeAMJVXu0k7r4wjV+NF1rmZMoHs906BEB1y2qlWBKhH8/dXCUbz
m/L6/LzKnfytxDCRJfM5DhDiwS7RYF5PiVYkK7x0ov7p00ujfZuO0xH0dIByQQq0
5gzH3nkQpsAmA8SzfsZ0lBZN1ZvkTgSgbzTGbdc54HZ2SLWIT7cGhducFU9Rkrkn
kZP66tcHsQJJZDovtTzDrjEWME4Frn0fL0CHTK2RNrxhzr0/MlErlsfr9/veLZpx
+stmVUT64teiL8THOv+x/F82ol6IbSf8VPCEjfjvf8vP7qc2StlObA3tvzjGWNgb
RCyC2VX96zVzzeLUiTany+TKMJzRcZ5YMF1wKVIjc9A3YCirNQIqE9AQf9SlODiF
WHEpEBhj/gT0oQnek6S0e+xB8ZlXw92KN7VrD+tFnf8F09amrUTWTKhTEnrn+KQc
UAbMZXO633+urCfdYTlvaVHJ23yx5j/PZhAf1pN12UXaCFgao+uHTn2ZqNEuF4GJ
eoz1sCG/fm/2smDdYlF3JQ8v4qhnf2mEIa1W3Vz2f6UdSLWNrAbtTwyUfWN/LOTe
AGJ1rHPXIUFHX0NcYbS+GNlOnsS65i/tFusYHkLCqFocF/gSeCoQOW4rl8nxVKWY
4XJkg07Ay8yyZQFJgLz4Md2IsTLZ4aJURw6RtryNtMCjOf/tWVtY6V99nTYJSOdT
f3Bq3QnymeYl8oYx4BoJqW5EoWpZEUW9nQx/8AkfbzeBlKozLDx9pBWOinrOe22P
sb8LdHYF3fvLoZRAPiXE2ZHOEjLcs903ie8MwJVlG66KirUVgJwHxfTs+PRg6HaB
i8KTEVLYUf3rz1XdIoEcwQi/SUPgYuCQ8Ydko/XlOAfaNUTdxJlrmWcGqC23yDt/
ztXCM1JI2wo8zpE6o6zu8RvxYoIZHGr7I2xwf7P3ygxdIy0Qi/IQ9iyBcAc8dk2W
3ZZ9zTsVYI/kIsZPnrglCtwxF6pjDt+c/DrnNWRYhQudv1gwKA4Vhb9DzX/vvdz+
4FNDPsH43nQuG/+TZDlMNQYMWGP1Wbfs1BV5efmcsnuykA+xcChdJWVlJk0i5D6d
bEwyJoxd7l/Al2V+e31rFR4J6DFS74EtdNhrKcU4dXuJQ7IfXQ9q/kqm7TuJu+Y3
/GTAxf6DEPqd9QyCTbGwfOMKmwQHVtVrfwpOJmP8ta4gl73z7nbLabDWMZyp5/k3
1x5+uq8OpbKAzdzLO+cqYYMq6BLZ3t1kbMhx1oHaD934zd/AKhBoDwGtTZNbgibG
HQhcSnL9MJKrJAwamtSmtUzexxBOTQXQS6ICGIn1OyV9ZPdS8hhmw+sJP2USe6Qp
s8YjfruoA5cKG8yQBQL+rVfzSRSowrPTmij+cdXqvCnN/7F2ebzJ2LOBGEwU7rks
/4ossE4JUHjlERJrktF4eUJGXfC0oUxZKc5fyut8wqsfe1q23GSY1UqQynUPTMhV
+tybEScqGyC8XLMRmYkZ+t/YmEDEnpbECU8/bJEPchWPn4VIw35NW9Yhe7FKUBTp
qEO2WaoM1qlMb8O6WuqTFg3ccSpjLTPSq7DHn2QMfHlKalSAz8B2yjySpxlxZFdw
CFcFw2SJDtuuSeSKzLqff+i4tabZlKijBICz98e9uApBwAot2sfuHZs32huFmvNI
AZgBGMJJUetN+V2kaz+LSXJsI5XrPiWEaKvk1wdx9rwe82vRjn7Ko22heSrvTCro
uS0GDABtT8gMUSnR4twbyjm37MsmU6/e1zFVcpzfy4KUxbqL9+1MhHgsC1Kgnf3d
13XcC5ces7kp5zNwtYg6+Pa9Aj92HVE2SxzqQs0V+SIeLJ++RKDvjty2Zu+T4yK8
hJ16Zo3B9BeJSFadCsmSaR+QNsygcNZHD+KdLPrtqj730C32801DglGfV2/3y99b
Ct+Oykctp6kRcpMvzPEQbDwFfZfsTT7WkoPkDw0Er3/fMptnymmFEsLYpgErlsFn
zBf6GuaUYZXXimyDjAW6gxSXRobcZgHK2li7H1FjeHe3ECQb9n9wAtSYAun/omQa
CJSssiu4cwwUltVn3KL1ViplgHVIElCBYGYCcEJ2GaTm3eQWWxcLLrh7oYZx6Mjy
y41/oF+rI9UgKJ2F3e/AtD4hjz6zLe9VxUP0mfQxD4MA9L/vt2ZWT0z52sGwFZyH
MZu8T6Y8yePhKKhFCrcJNE5Bke78iB3F/32fE6f2YgR4dKeys1x2hQqe1mj4kUBo
paLHV4x644IBu7GALzNIGbKwkHbZ6qJLQJaG3w3CHVS4kgLkc1z7lWcuSQUOmDst
nByWu7/MVUVczLzd7TmkeNFw2txY7V1KgL/jki6AU0wigDCP3tzW7Jku9hEIexQq
OhoaPQJGkTy7BhRwtQNNR058bbPVmPs/+sXEe0bOqzB4C2dooQZL9nCdeuy1yEkQ
rtuCcss13RA/9CeTXhTk8jrU+dRFCRm3DF8elld4UclAuiDG1xhWT2ipedBI0+Pa
iIHMjni7hDjXi8QUZS1VFOqArWhlHDTryiTRRzfCxt6Dspg8PNOQ7zLEjq82Byz0
WSGEVLUofuDfSqySc8G8tEpDMbosssulxt4VTM1lHY6+chCdY8xxSZkflQdQZ3IN
Wjxao38Gi2GUxztnN0o7sdmfRN82V7hs0bq5QTaJnp/H6L0TgkO7t+GZQaKABU60
Gk14VZBCB9m2GbGZhA+EBLOkjS0R+4FITS2lh0IjY8TfRewmTbJTOsESfoJc+qjr
oq6Rg6j1DUQnuW87wAtHnKSA2oZfbL5vMiLSyy33855bMusfk/xEBv/djq5ETe8l
onl8gywAd8xl1bA045KS8UiA8sh5/EIcCEHmE4ttVWKe1d7n0d0KfQl/uacxbhv8
efzdHMtjJbp/Qh7J/JS8rNK4KL4IjR9KD1ysn+uKcUMdRH/AIZR/NeoC7OiK3I8m
Q+z40mjFQ+AbqpRTE6cI8GaR1J/+R6uWJEpJQpKFXju6Tkap63hG41QotqjtZ3j6
NfK6ZUjaNH038wDW9MVeThNuAqqVaUB/HWMbma/15AIqJ3wqLxovIErVJj11G4N0
BX9XwxnoRXkwUBqQZ51t5dkASzkijhGltYoNb7+OfQn5F3zA6bexvVtgEyj2Zdz7
5LwvKOeOfmOTzIj7+NXKgMXQoXxRoNGf1+2n9UzVoE2gA7JuMw5pDZSkiEe8QL+F
Qpfi17KixfSnBM5ZbYwtacL7hInqJwu0tGKmC5OHT9YE+8fyRtxihwVw0Wo061M6
fv/KaSSt30efzYDHsyjjbxd9BS4bUR6SfGB4iV+dnEqaiSWpLPy6/Dqdca5U5lpd
8wO1FZmpY5/WyxNHrS+b99l5Dl1qjimVKR+iidK7NhoOkKxIOHm/CFxujF9HP/F7
+9sPo4UezwbaIi9HP1AtSm4SZEQsfkFHd8nc5tpAnz2Sk6eAC1bnE+J7ld2U9vru
jO1jgGcfgdbK9dbtVVyFQRz2KqASXnMjy5nw7dTzHIEiqyCMarOUGT8A4+lT18GU
IEQc4EfnB+HkiH5YvPD6tlrOgH+oZYzOV0ZFfbwsXxfZmWgrYL5oP9ihJ3wXW7i2
z4dx84A5dMEfYXGeRVAnevPJcN4LAaFd5mtzFSl8/JZgL1kd+AnDqavD+AR3NvSy
wmDeHvlmhv1nC8/UAEr0ruD/aaOa43ZJNBlOXaJq7YDd2ajEQKwHrcL5t2KqVslq
MCP1ch2XNt6UwU7ykbWtZKtVoWEGZX/bCFa2XX+JR/4btDKdpegZ12Z4hk4jpm8+
75R3OfTS6h7QawJqHPYEz8CMl35rRZkx5Axswb27Oh8bo7WUEp8ZqtX0QPyngJ4B
4TNPjHajWv0cV3fmG1QQ5v0bS1F85gzN1l5x6VWG3S4/yp3yc6QQHUgYrWI35tvP
mfR0O7DYJJLanOOs/dQt9EMtseyX+0/RK6uViQCbk+nKxfb19XjfYA2hkCeHuYGs
4bQwfqg/hWyv9WNUP0VochnNZSvPH8MR2JSqZvO7VeZUhQVHHVH9NkYS5VPHfq9t
P/Vhd+DCdCppxBu4kgPMbnk1DV6HXwAbUBXVTox/O1yFxJZsnAJLImaJTMBdLvZ9
6Eonyh6VjiPXjAONgT0J3aJ6cU247Me3lRs/e2FMpNb6Dy99vz+S+LtsF6Rln/90
dh//QuB1HFYikAXO/nrthdz56tKZRLG3DTijTr+GEp/yhCWjtRCzMqryDHdKZDgW
2IkeoIpF9vxjN9RoLIGtL2fSRcDhG1fwSEOAz3BM4XGTkaGn1uhSE7zNQ6KAb9Fm
yrY8kJea4TyS11t2s2giTr8HLeUt1JEDAIdvHoGu24TUq+/eXml7wOHL87RWW7UL
9pvdX5mAKIqNGNYErGiJlv4PhG3+nN0Kx5cibsCAD6fLC3y7tpjHFQVKbg7U6IjK
scecA4Qf9DpMddoqHpWyH4pvrg9F8eBOz8pSbtF3Mf2aiTGy6RV1XzWV7+QI/4bY
ffutWoQaiMGvJ6pNxubDLu784CmbOIbyAs5ToPMmq0SApoxQkvA+SdJ0p/qfd4fI
xdMbZRprueQn/S/1r3/2aGyllXjrLFrIazoyGiyDWeZLd9/vNeWzShZaCW8T+QhP
sRiDmd2WF4Aq9xLDcyQ7hv/PpFgH26QqisIDox9MCZqVKWIYDkC/zD+uKmfGy4aP
oObPiPo1QkmtBV8U60mWLBaRlnnBKJ9JIbW405Q8nnTTOIF6NF8L4I38G8M49V2X
8QscgXBtKWeP6KckNqw3XPmGVHT0gJaW50l8wocZjD7wU4g5HFAwgc6jwqA3Wkrx
VF//Wquk3S8f/sD2fOe1+b2R5q9QgJEAbAu/qR2xbxcMFdvj93zIQGKuUcaPBv6p
Gg8L9gVa0TiEpIQjv4b6hK1rgjoZ6HEW/WnUk/Ra7tAxFQjDJ5sjwJ+VAXGKfebm
3XQr99ue0IeScQvIKYZs861JTGub0Zahc5A+5ZoOVCLmh/QQTBqdXEyQ9aposiC+
YrII04659nzqRcOcpisrSpjlWgMmyH0EB7Oifxeua+o55etEAzloCxuBVjV0bsLB
HgoDRZuQ3+gvT3YYhPLCjTv0xpxtHJwYhaHHPAPZ4dG4b3feMEHBITqzDa1wR6BD
9tpnna/ZaNN0vRtR4JUG84ITZlDQ3CdIbELBFiyt0Aus6zFb/+zcD73v8QsPAu/2
+d2C13PTPAW0DgmP6I1aE3lslSL6FF7pvshtzOHeP5Ax8gx8jYFcfaw1qTQUGN/d
qE7QUgFQxvCmvegpFn4CBzKYLT5GwLciTy8hj+Og7SPwYO6spnlLYMj0wEmOutjZ
R7qb69vLIrIuspKM/OqqVBBsdWyNmPyzZw2Gdhiqkmuv+vhL33Vs8evvgRW2F5V+
QLr4RcSWB1MRMwllxgkEtvniqR6wsXc/IPMYbBbk4V5kpjVtNekYktNfuYFYcUAZ
JM338GK1LZHDwwxzZWcxdQCVp+6ZmZc9DYyt4DEzdrEfHpK++iKIRKltJHL4ACcp
rQDCIWQ1gDyX8Pq+6OtCpBcMxFqFWCjBTd2DVTOoTH79ja0/sqAchXaUSHoXLQgh
QGwfZnduHFlHTW1FTP80YXjx2o9GyNLn6+2VtnOAbHXaK9CNoZgSYSE/EztxjJZm
TctLTzZrmmtdK/cBPNAfrb+uaEWCHr5BG3m2+IRNgVvShRtuKe4V+vjA1MSjUg8p
t1q/zSR0qAQwFqBJ1kbbn6eCiCBFqgaeEEM1F+peBZ/0fJC+P4NZ8rKCvAmU3tJ7
5RJvKYv29J7LnretjpHYwdemRiIqon+k0S8oLUqpWZpdN1mW8az7NRWO/iwnOC2S
P6u9PcZKWn9yvROy4zn2/ovgjtQlqC4cnZm7JGtjSe6HNvbXN73ygZ5ZOhmu0OXk
iZKX9HavhhksJhk7BYNeOp1StHG5dSPz4d6czdXs+rNqWWKoZiNiSr/AagfSwjoq
2I56G3fvdpR1AJBgECUIpEFJuB0aVlFVJ7D6HT8brXJrpik5bfGFG5ixvHrqG1A1
527gpww9nS1FgVDmr46JKMiUmrmtm701Ba10hOlhy2ieVQTpj9h+9vVAgLrIrg1u
z06kkNdXxhxeAlCYX0SuVqT6ef5SK5tPfMXj6v3EWQKTV990F6Z4T3mdqrUzsF9v
/F5VHGK7SX/PqqGrUU1FRGX0jKn49kaC4dqUtKF+3yN+PlizNG8GYX/OpWqnedt0
XALaeeajMGeY8C3pL3zAGKXBFGYIRxwDxHmCro3p/jXoaxr9U1E2AtFcDri1HwT0
0Iyxnc+M/d6vcEYsMD48WsYb4gWywy9ng25PWlQJDWeVwiC/bRhTgyYRXswflCN/
214M0jj3otIu3CC3zyx/cUK7u8wFUggpTWgZHsovZwjx85P7IbJxLYOOzY1XA8Nt
vTcsnEU0T6ZVLcYWjwB9AzoYrpqQqdXo1Dgl2P/VUwCJX3lr6vMOsxCF2Sc66HsA
ytCrxkTCTjje398IiMoEXGj6CcV6zuO0aIpWBAAHVQR4RJQ2D1bgJ7aBq4rPBTg+
p9NrkTHqOF14V3ngGOKmJ16uFB4uDcam64SRY57NSz5g344ycd7tgR/xlU3vYD+M
36qexU22q8LNiTH2LnLJ7khE/8ktmBxaT5keLXTiHj9yKIhSdUg/4c4WJGNdByFe
SDa5bzg/Wpjh4/ql5iwk8CMBgj7tmQtMwGXJQbSPFp4YOFPGLu3N9m2PIk4J1MTy
5vXCu94jiTuUyjuZzKIL1tVGexRvsLNDWbRC9Sv+3Z4ouoUG23Q0cUOpG3kzsoj1
u147V9OCSX+89ZgZ9pcgez0P6dv6f/38iA2JCjrvni49Xnt3HT28wDrIiqshhqvQ
UWnhcFMvhn2SK8bAmDcRxY48+FVNU126J36no8wktfEUg8O9gx4BWrjmLPg9ZCm9
TTRiSuNWISIKAJcZ7rmmnvTcCmCzIdXZc2ipb9zIJ9NPu4sHRBSk/WOa5bOaTe2r
44Cnq/xdniMUwnQzkXPiKDXCh5obkbYt2WLbupM7Yj3DIgM+jNRu17vJQsSWMmwh
HpJD8CTySItATsahPv+FvKL1nKSAEmylvGRGyuDEuge0tD81MVmyj/2ODMN/alUC
zFu2iTooKdc5nBSTszqFPvKRHQAYKZSgGq9HcMg4t0c2hTdlcBH2likiNcC058LA
yM20Kbjib52eZXyQkMzejl/hTehAlDODuoDo3qH2ebTOxX3i/yBHBdOoZTrKHQYa
kwVSdWbuG8vflJcnD+DEavv97PuyQCrOPZ4p7HXaM9EBUKnH1SzxT1JvZ+GHwE7Y
7SsWcmLoMTsAEUQLBMZaQf/GRWkvKoYvo4ssd5yXj0MlnpMhNSXsyLmi8cOrGJ/J
EHSydB7vUmyBlK20AjO8PN5IYi4y9vMN4cgNuAqk+3aflI+qs4t5uVMYehm81SiK
q0FEcHXDk4QL64gN46X30zoyWjeI7RA/ixJQURQuc2wP/W+mpxqvo911tK2moltE
lkf1hvHK9RCpuCFB0B9gDrYPJ5hrH2Z1MAfK7t7dmCILtGwwnElYBhb2SyvjLI+A
72OmoKFKQ9P/RS0X1KWbByZ/m0KHt2xb9KXYkblneneKPs6vx+cIGgMz/2Tmy7Jt
d7w2TdjtXbV1CPmDR9ZDSWHz0X1wejX0ns1RgyaAiRF75+9OvNifM1UIZQZYU5u8
e3E8ROWlZcxH39II5t/35EkhfDbDSWxnndvYtgPsYAPVcj5mOoIpX7AgxqJmF1qQ
5e9na6ffj3ibz/bYOhdd4WNrNytionmj0PZwtTD3E+qqhmoobcEX3t4Vxce59N6C
pQFkMjV7FMoWrrTI4si++M6tljtVf9zNUjp4rn9SHlw0L3Lv5jv9TzXgUVUlP+I4
arBex3wJfMLI8FWw6U4PN4uWrqqh+CAou2kSCFJa6DudZQqU3DcwGVA8XxJ0+YMO
1n72g+kWhr2r+dtfTT8JDMyPHiinA67nz1Fxkn4L7DliSDYlv7DSPufejrVkz3dQ
E13ha7SEqeerpXdZDim0bETYLb5n3OoWWon0y4JXqq7CxV3/UdcgUFUIxzMTgr51
EERNk4zNPhSxb2Y8q4XJrOEXGkOA7wCcpMR9ng9DIMeFHl4v6tuaQ5smGknXQYQ/
Ec8pSezxwKvhgiefqygUqblIZjJoUmJufzA6Ot9emQ/IquheHDDID3JZyTNuIgq0
6NWLu9HAjrdVbjHJurwxAaCNLadgmVXWzjzORZFQsnZtPf9ontjSEHJ+H8ZYchXZ
zZGe/13eLIjsdaWCOuxubR4e2Cjg6bvfkV+dRu1YdGTtW2T47R/OXAOZVqynVBPL
n9nCRUN0RGQHV/XbeTz3KjS7LEpTTcUF1qAFWfIL4Cqd6ADGaxGl+XDTkP+W5NfU
UW+l1AiJ63SzbqvMY1HuAPxzcrtuBqDywIC1qj6abzGy23n331ot4VMn5hZMw0md
/H89gOr2STie53obra/iDG95pTiiTmdSFRQZzcpG8oD5gCtY5cQScPqAnIlr11/0
wIJpoBxqJtPLR1V837KtYFkjfsPeJWYjTgvmqiWoykVrxprRdkcKtFDJeMLke8Li
MpOsifpTByYUxzpVL9egZ9hiqdb9hnPZV61CeDf5u/HOhxpT9Siml3Bvuc/wUBZ+
E6WdLJDxDWhPPuW8thA+109kAz08zEt58alRkNEcdItJClQcwd/9hNY6+tki2ven
xKIJQnGAd1OwWwAXiQt29U3Tp/irTxK7FnVgo99t/OxmUFmoEhVv5ptZXk7cRu9G
FHoiZWD2FkZLQyzZoUAOUTCS9qb2D1tZOMRwX8mT0pLJygzrqzFXjl20f/7e7pD6
LBAUyXgYmgR4OZR/rhNqGnN/Ekg3Xb+NSAk5+U/bISlY/euflY7n1pQHLSZ6Yofb
4l7nLkWm3SMALIbw0NQXbF9SJF2IAoURE0NyuwNs+R5Tigm/sxHHgBI+ufQv9jJm
tK4wnSKKFSB9n3w9kED09A==
`protect END_PROTECTED
