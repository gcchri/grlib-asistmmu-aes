`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ypTwxS/qwehayYmrBvUaq9M0AOwTjJiC4TYad1ygCyXAgWU8Yd0kj1ipIp24riMi
tm56h/xiHycbetHA6o1jgLyPFg4XVISeg2vc8aSVqaLqj4hYODjo226F9ztolLCy
auB3cF5uKYBZp7ZFMlxZq/fUU8YW2vh9GWO4tTGen7VLUkmfzvw65FAgfl1JlgC3
LIDcYdbbQswE+PncFk5AA1UEdNwu7FlI6u/Q5AmGwUt6Q0aY99+lC/m4DBF0XJz1
XPQGD6+3PJFzN8HiHC3t8glXt00kJJWTWDI1rnl2R4de0I1wWYp3Q7OjQ/303Ims
z+7oHffTAo+qKPJ5e32DsRWZJUObON4E334LOSmnpyc=
`protect END_PROTECTED
