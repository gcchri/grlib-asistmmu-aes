`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ViALYrZRGGabFfxqn6WehXcRp3xessvsP/IIBsRE2yC9nAdaJWNhlMCUer8CKlG+
7O0UiNBSpcoqDVppOOyiK7lJPMWi1VdZyQUILkvcxL8fhXYfPxQthwKsUxWpKYqu
mTwQB1fROE5MLXvv7j7tGwZ5XD6659l2UVSofGoE3ZD4LolQIcJXg2x80VxOum+N
EGrNppdN6jk3wbWFs8dm89e0HFxa0EQCpeCTym9/Ysgen+WmFR3GQfh6o7yRmtBk
A/dSrKuT437bxj9V4XZP+L+OHy8dDBNfZ4PejBLYJ/Xqqt6yqsnKddtQ6fEQ02M/
FjC018imfEU9JeYFo+v/3gmaIbYQx2ay12lLf8Olr1qxVdn5CkgUriNy1bLOGOX/
08HDvdCAuAWtDck5exGy2AEMWm0wTlKKny1ZrLNVUu/rVwUZEzfE/1kMqu0AaAfS
jCiPpivKtkPqFeAOOgE7roP/6cuSaa/v+QL+qwxVdmwMaWdgjzN4YJT7RWJZ4I/P
6x6StXJtvDWie0dpGuDO/f39PkR+93Zzb4k8C/U2cwrzsAPevrnYyPz3yo0YT5Z+
oud/LqmNK7k3PTZUP9x3EtvNCYjwIRcvExMjvR7WJn0=
`protect END_PROTECTED
