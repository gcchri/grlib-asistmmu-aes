`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q9zPzkFXs/MKUVKngCzRuH3r6kA0WYSVrzG2cDBGWCZ0YdfW4m2h8awJcvs6RBnU
aBrwIhAV+l31A6dj6Vfu5BUQ4x8X+ZLztND4mwjfzvXJ9kkaBXNlevEoqtqtXHrt
nNEEGzjCSlRst1YEGETAsw1SHuQhv+8P8Yo5Z7l6zRsButWcmaH//7CL7GWgQ6/i
YZVDS+bjIjzrNmRiGiSfigLGrIrSs5DtYSs76ysOHeg9hi/hQD21zGdd/Y9c4NLO
zk7Xnb8ySTmvyjo+qw+P3ZxnlMIdxjlOoYFkDrX5XoR4c/tEybs01195MXjR0Qzb
0lPcnkKnNtggh2Dw4AzrFJJDVBaQlK2PHtU6UwY/qvwFUF7mXila0oBDudAqUfpW
ptqRC70ozbRFQa9LXUa7qsHEDrAProgvXblDuH1aeUDXF6K0pj6dNGvjqvWg0KyO
UoHBfSKVClHmVVudHd15HkC3sJE4ae9fgiBmgcvtDV5J2Fz7Uc87EH51CmLCMwz2
lBBrT8rcu+B8FGhKnJWBr1ollf+hIR0SZWdisvzhgAdCPn9QItgBXhD2IDYuhM5Z
9nxiomE10Ld1ZL5rTUD3ui/0xzbiw0q5mMe9YQUu7//nL+nQqcHvHDy+cU3o3LNt
3FpwqCeJD1RryHvrOj0o55Is55k/moL7jI/33nfI/67iUnQ3uhEwYt05NOpOgNDb
SVVqYqbBJEqLUN3paHJ8JJSQy/suEqESLW/Y6dSWdkG7UktHR9iXaRSyLUKUfza6
27XzMZ/GFSBgIsVpEoiGyqTk98mS/Q0sX9PxbPuyIt27+RCEAUcn2PbukK7nrcWa
+02xPxQMc+lqkD94SsIm9Isf/GGGJNYDA7o6KqyjNS3nxt75TfBtAuqk8kBMp1Rw
p9lJl876AJeIHlDIxoIyc7cWS2TvQ2Pxto4NEMKKLpyh70JXGd0XT79XqYpM5zqP
1HoB4W/MZ4riF9l2A1c7Cetihy8TZ5pWRgpnkOCZUlKZjGGRaa7IW4T27z7ZHt8s
WtSsYefHU3ep/x1a+50T9i8EbGV8oUdNPI+rP85GUmQBxvnVYkFKDUSUhWsLb0M7
HtknpCnGS4iCQDp1wf8gnvI6kV+0aJN2xtmNnq54Vq1QEGiKbsTLsVTVXBWwSgWC
Zlpfjrc2LCR35/SbiISvlyL0bkv7UO1xoPv8YtL+EYUt/wS39a2gZLjJI8elfAZQ
GPChtZlh+6f+VnCpA5KsvQ==
`protect END_PROTECTED
