`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UyJgX5KUAMVZWBU/HVJhzehzwKgX0Z+Wql7nBlfylhWIgxF9Ta5oJUIRu8NdGv/u
VZeIes7XxJLvz1hJr82VGcB6NTMBTWkl78SxPAyriRXthiNzG30JZOnSauRL2Bq5
5cTu7Pp/U2k4rnSJvyiv7G4XM8ugl9DAaXmY6wjp7NldXlBFz9E55tGvu5OxWrCo
Ls3jPYG94NDs5NFVeC9hEEJYxior+E/5LGZ1rjF0F6/oOqnjAPOsCHu/fUnpAujr
kgntfPCzMqT+aS8MDCK7lIBzVAakS3tU243z8HAvNtTL/2kGAqIoaIomjQcHfREX
cLiEJYf9A7GvckgmwTKtuQudO/kpaT7Xd81ow7P32sCy2C1vOUD+t65QFqdQkL40
alMECJm1saGZAizShETzHFdJ4AGeQ+C7MCXXmaPSXhkuhDBNEmcIWXlAaGb2DJzO
O6Gtfm5yzJ1paK2X9LsFJukz4kWgqjaIitpIWNO1cr1/xDMvZz9xNlnOyTxDhN+k
wA2K3rAAn8264Cb75Ebi6Z2eubl+WK3YSoFQq7TbFxfRKiWTzTPi6SBWQr0eW6ot
9t1sT9I1BzD61KYm65EyRGhi0vSjZ3Vk6L9yKzFzrVJCVVy9mbzcgF+WtiO6w0tt
iQVCpSkknekL6Xg8R0nwwLqCSIwwTC8blaqOjY12ChKMY9IeO8h4rjrBygRvZfNl
tlz1/yf3TXXE1ASIQ2UO7nR8T71TCfyGUx4HQ9AaIzN8KBVJ6pOLN61vAW6yijoX
+UyZxn+6PvUXenOyLAmJanXAZamKflMYTzsrK9pfnD5N6/tbO7pn7am/osvongio
I3ey/y8bCfmld3W0YcXdF3yrSNqm0mHyXEpVlrZ/tPKI5UZU8uf9PhAv0s51I42P
2hvWru1Vr7d5wuiCwxi//w==
`protect END_PROTECTED
