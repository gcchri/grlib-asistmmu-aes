`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/aWHXfIELHhMwi2lXDB+2R5Xedk77mhECi4CvBzabzrZRH6MRCv2i5+nSazN0mhc
+IyJciSthRMZHvqHJjL3orAghRX8b78HhOKWQdveSQMd5k3FuSvm12/Mbi9ACsu8
AiS+nObeAlkw30VqYtNoPizcYgfSM1iKDa66BWRIm6KADhq/fpN0FLeAV90pRJ1c
N7Y9jOKe62h2gMWPvdEDQhIvGvg895VBBbYWn4tMUAzYW2N5ZP9INW6tZ6GiMqSR
r7tlr68I0DaifVsWrFEPa902MTtlCovqsSgD1tpIpaqng2h5aGY6U4+MWiIpWB6W
6d3tDc3i7PmeEgSUpOVuXD5m98CgJyD3JvWs9H3t3bvnCZkUzZk4tP5NV59hcoJ4
5JZI6nsabp51jy161j2B3A==
`protect END_PROTECTED
