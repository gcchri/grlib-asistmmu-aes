`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pPNIKLk05xqFhKLGQA0IhQvkUX86z2QL/lkbUeucTzzIYozPf7xxBdzrmhmPPriD
mcKwBXNuG8ea7+5lTIzNCwbBh0TJTsKA93qrjaEK4BRTdkKjKWV6Aqpn5BuvRw4u
V93USonpEVIJWZXAyf2C3NZWlRWxENfKcp8kPTk1QWaUMDLNMdlAWK85eSBOodvs
oF5QLq+6oOjGlfUkORwrBiUrlXYbQiYGcq69XKY/AKTrnfPmgvjQ6LK/daNiovsl
pJrnqYFXL/xegP1hNMXEkyipVEww7JlhvJ4vjFLevQZlPMnAeZCT9AlrqNy6MduA
FfcOoDj4TifIVmFGGE1Qej+kCY0Vuo9Sq9S0WKlw7MFBImuXJTb7ZKHlUVj8qNU1
cTKjYkNl1MyVbwSZMzeRgKqtQac5EsYWXZLOTBY1bRp5p1mgov6+N5I6w/BFStBQ
5akxl5UpUH+r0/Ek/OH/GRwbFgJVoAc7eYjiVRVvrisZUZ+jSYvsut29mZqIoash
`protect END_PROTECTED
