`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xNzN1uDIQXrP6qJ8hNJcz2l6REAsXkc0vsMg8dDkS5KTa46/5jZM9hyEgeiLrDEv
QJbhT51Sdqzbk/ie20gaNW/1wE9kOx9GI14wqqtDc1kr/IOzEtKZBwLocwq6iR1W
ZLVoE3nkyd2IiMLu134fJet8uPnh/Hr/+eKLpAU8gQb8yxq/IMmdNyGpa+WcRmcA
7uvifkBVovAS+S/gpIuaxpIlwbxEB/LMksXFgy+UneDF2vM3Xf/8J/QJNKCWcdcy
A5wRLAaIGTVN433QglstF+01oQh+2DCwQ0D6Tk+sFDbn0T+6ryVngt3Bcubu9I4m
a5v3nRvZeVTqeGRRFFzSAbFxULKhmjo21PbQovdUjcZDyC1IlhUuNsPBIZx5tJLi
CksQ18eWTOJR569S8Uk39IcrdHqKkvT8i0EHZzR5z9BLh/XRWo2FiNInhS2l3Qn2
lvy51bkpqKCX2LjNDX0LcjybGiby3x8ZNsjmHvFDLPooLhqZE8OcdNrYnQlDRBuc
wsv+vJ+s5768tP/CYKkVC68qu+b/9j5ezH4Z1GVhXhQHt/APS7XoEm6smNrfPA/s
G/098EB/X0eNgzNxu7txHN4Wr+LIM/dNrVEoMSOZvvXgMWq3YxlZr/y2OXSKrN8t
VkfAl/zgEMKuFTCmLm5ymvA+MDx6XzWFcDRvFjjbFHRt1ShbQYhfnof5vuQafa7l
LNJ3Z55oYq/n7wuxt/yZA/nNoIdonnWv90KtAJN6We0Tiv1FJuZHl++R3eMJtUTI
mi+cx0s/vOOE3fiWeC9PzfndilZZnhxU3unG6iSJngkpwqsVebn6uF5DzdSZoxf8
hhAb/wE15nYb+MUW3BLpbIy3yq3DaU2V83ZVmaNr96tzMNIsN19igt5yPOZlkseV
U2/53cuOkqJK+qXytlNjT7gQIx4DtIXZ/WJoz2g2ebXWbr7gKeGL8SLt/K5na6/Z
rjsj4xQAjK+vpsud1ermAqVENKvdzX6Wj86KstP1Ntc1aEDMYluuBsjvNQry8kcB
+Y1F74rSqLXZoZ3CpH3yw2kO4DIdXfjRox8TQo++P20ip99yMfgZJN1KHc7cQY79
VebgTI3aDeaMaBFJFJvgbVOK4+4LCMfgBtQhnGMyBspXgeerEFD865po8YMOnusT
2repIk0g4SRzCHYur10TLew63g5xlBV46sisXaR9QFn4K3Mk0PUkbTJdJ16ljPj+
FZIYYueYB98+RVp/j87vNwHVr6GA/CQE8nYeQOwi2tjlv9MJku86TF7EFa/KY6hd
NL6QeqpuL0uYt8/xTTmufEwzAJ2+2t1DPxCDQpelt8kfgPQb+1z/lYS/ntFQ1KOY
bH+VUAP8NQCuML3NN9qoadrdGttVMbVs9Lcz/JXXvuIlDtZcoPPZK3akhKSxkA3I
YLjzYOb8bw3WEyglPHehB3UUYJlJa8/0xSrUfAwUVwCLw0r3sQD/FqA2dFbU3cp0
5AT3Oqzq+PcrVhoT5KMo7Mxi57pwIVqZbAti9Ck5q/JbJ6nKPF8R1FXJvxUmNodH
NN6TPwBHUNyijnvL+40daQ9yPaa7eUu83uexF7pE+KW+32PlX8rNv3t6ymhIU0dd
sHzNKuiI37GJ1mpQ97HV+HfyNUDlTGsth7cwY0Vdcp5vTZPVJbpqvNOE1zbUmUXK
g97zznfhvELlIt9S/fvvd3rlhVRrBfSMnWEKNSJaq1OHsWcbyLAhsek8lVYZqF1k
+MCCiPUc0urdtRcOi78lsEiZ4lSmpbIedhHuQ692jjk+M/prDoDV3Fb/LdUmPgJv
o7diyjEVCQtY2TLESmO6fSjdumIzER9c4p8SnRCcI9ZcryjEOsg7fA4WxR+/tV7I
MJ1N4zo99i8WYYqt60Yxo59fwI1CkLcMwcv7Mc9ksKSL+Dirl7jKCbt/Lrh3jtr8
VS/fpCWJi0OWYq6i0O1UcSTbWMfKaAJBTBshL+0rQ1Iy29oawUUQq8CGrptu0rEY
Yr2Isol8X86rhfXttRT4J46Brts5qOCaozdo+oEjgVYl79YS8ScvTkjk7rLX+EjQ
QHdbLJq2zNsKEh5f630/0R/p6gv2+bfryT6sIYq3Bqs34IFPOrrTT8A+CuTt6i3U
pq7hE9bptRJYpBR3erC0vREvRCR2g5UGNiUJ7CuRLXV1wZsXvdLaVipuxvsGjrxw
yCwq8976/k9hYEHWbAleCB9hVygUWIpZNnon5VymqYZ7tkb8ZlRB3eL1G/8Exjoc
ODWemUgCoj4R33Orkk4jM2trV2WiTzIqbD/YgLMoIV2U39fROH4l996mWB3bj541
6FELiuC5vspP/jBBnJWHhedNnDzycuc1WFwdLG0CCRAMLQ10NVq/lcQP3RYzxtmb
N5u7W6MOd/bI0AamZznPZ4Nd47KcCRQ7nWjNUMe+Bmh9IyNoB5EUcWhfblyy2jjf
6UgYuCsB+6p/bNO2GGBbD/G3ZsRYa4It4fi9pMUR7Qp6uB9O1JT8nu7YBmqnLPMx
LtjY79rLvlW2jZZMoYq6vqkWds9oCGEUbKIdqT+P9t5SQzEgeqW7t6WHoj26uDQD
oU00BWNJb17MPlTpznUq6mp4LEQDAAuxwznEqfJOQJs=
`protect END_PROTECTED
