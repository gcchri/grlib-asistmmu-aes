`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QP4k5i4qryg7CTYv96BfAPc1r5Jfc/BPPLjptnas14kbEu7qhnmw01IMt6yqQlap
Zq08eVa/mIwotnnOlS7Rc47DDjv4mJNH4tzLAgtV4X2RYD7bIWlvFI2jgxuYXqVQ
mCSf0eD99IU2zeZOoQwm8UJSbItKFI3x5DU26djczpc6zh1CaWASH3D8VTE/zVs/
RwD+JWopcktHDR8OfHBjJm/ws5p3UrbxKoXO9NQu2AAtXohJYVUcD8yusraLmRr8
oBVWWX9Lamqvc4ZgHJbnvsSfM5IRxBnpkHOV5ebtHcxuA7XJCSoxcsNkBIQA+EmR
p9QApA4OM7vbEV5mgOYJ7THYT86u4oktKF/Y0wg9FQz/q9X9RoaDu2DoekIB/5Vj
b67GVIQWSrSL1VPkEoPviAbU28gl0PUAcc33XKWfDhY=
`protect END_PROTECTED
