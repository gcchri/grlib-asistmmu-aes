`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HawaH3JcmgrjB7l7ZtqtrkCVmEnKuGxoRYz81x1wzR+8g7nICwOSio9Vb+haFkZC
tV0+89GjSQ3OLEBi6oj6ZqC+PQt4cgA0GN12Xx1x/P0MH6YuDGCvS+GEiWj6lUlo
4HP5a1E21jFHhTMJu1ww2XfzWDokExg4a40Fm7hOzronRIvsvd/1G74vb/4NWBv9
X76+kBaphxcnSBqY8/4i5O04GsxgSlUhPGHUiyogP16ctXJmxxJIJKYs3KpLHgSI
ZaNPaxUuLQEARMXH3I7FuTTD3P7H/XvVex1Se8P+QXwaAOCZjff6qkOeSSKJbm6/
CEHk2UCbtMfsVWpHvHomM1fKvK/SmKpRm15DorC4Sg6/yEl2YSzHf0vqLjcilkGB
o3CnTCRRqDSq6qyJLzo6YekxMwWFoNiJd4V/qIEQtY4u52geKdo0igKp4XFCcFzn
nbi4GqFVgm48TVQhZJJ/GwvYvy+Q96OCG848EiElbCB2c+VdacB1ujSIzsCAGAU2
G6PITkpRQg0NisVvHtSDWFbFhdoPgqAroPI1T6Bh69FvDVmFSopjiY/CGtYZPrlQ
H/k4BSS3inUKd3/r3EPqHrV8qpL4MFTnJdQgCoX/d25k1jqQ1jSeQGeB6LfzsOEq
GAXJBrXasa1xnj9/vMiCgg+EaKXi/jKP8ljF8lg2iceUoyxk39HkzAwzyKHAhpo5
Z6Z+kN6SF4JzZV5bAqlJlfALdKQtC0YBGAI4RVlNpSnaujEPnI+tzfb/86fueA1t
/NOr6F01luldycS54nLCdt+crOBTtZ5ta6LBwaJc2i8=
`protect END_PROTECTED
