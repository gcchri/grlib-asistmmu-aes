`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U3g+AJX1VZriMLZyT7ZGZsYDNtdm8FA37sUxfu8/ZblIDPP/vFyPDTI4Z1oeE1Tg
Tf1RG54dwr9zOJHalb42XSTDKF7jabV2uvZTEM/mWg1ZHt3IaAFb5lkcxBsh6hS9
iUk/Rafzf9toQfc9XihEsftdYHhEuHfXbjRB065+Ep8rC8HIjLrhp8lb8K8z4x7K
hgJVcxeP7jxNu5vqABJWNS9fiKvLTJOzpbzngwHHFZWx3v0uxxLH4EeQOS1T6Acb
QPsIsosfxFXZl2pDecQSKX+d2/wvwS5u3p1VWOj+dQ85zyzDN3GrOLhvh75+y5iz
p0vBFpNm9zEBiNh3Ipt0nYxj8+FMNlF/tGG2WOsXSJwPp9/4WVdQqG7RsCorRIKx
wPJF8P1Xa3esXrMQE+olW0wHZjZcUAzuscJozN73hdN/1hwbmfz/zvTlxIXTcp+T
ucJZAEqtT7cI0PMWK8qExMwD01rdfqIFiOYVEUCuzzkn+R1GnLxvQ//Iwe2PKIq7
Fwz0/EKlKAdz7Uyn2GYQDbYJwYY7yelWS3D3b6H8T2PbGH6hKuY8jkWQQ360pRFn
6yrGh8KAEOAYJ2fLoQ5dbw/Dfte1gDCtq3FRQN5Gg5bcCjecAOALlj7f0/L+PZdg
VrXx3Bwmrs6BGSrX81vobO2hm2CHvqXH3ovwNDrapS57b0s0/Z9K3+1d/1TWmgzI
53VbMVahgtts2UJyEoX2nj+NhRuNUXvGc4oA1kfne3fxMK0BmSvOJm6y1EqG6pnd
zBZRZFgfHgQXpTV/VrLhPzLSlL5xprRg4xx56B+9bYY/rcaNktbK5LxUeLWnYN/5
3jYGwWUAEV658FiUdPuWxi4kDQaZdtDNYVwhifHFal/t0m6XEQ/POpQqf5mCMOXQ
VNnnqroLh9MUpRQALyEHo3PgUNNito34dqbASF5C673zIJKxEUyD9LvqD4W2Bdt6
Ed993dYzoxWX5hIkPeevRVKb6tYp+jUJ6yBEEXFAUiC8Avy+ecjQV/bNAAfe3aS4
6whoZURnrUV9Kfr1m7BmubS7iPXR2f0HQVAHUv3KNAWKbXZILf5gYvxFdOaSu4zw
phkijPTzLEjUviscYPpvkmRMd0zMjbVkEIG3U1KyHWNznbTNmPOluoDHLQHuPnmB
PZsuWANzd06OALuae/5GTjRBRGDOM2MHQRCxtTT1dTszlK578hWKIDUpItk4IOK3
o0L17lF9oVheG2ZdI8Kdp0rUKUEYk9JmwGT+NvGT1vIZ/vpHW4XcArEimPlYGU29
ewOCF7X0Bo+8Gv0XbwM2cKJozXCWxiRv+6VJRs8OESSfmSoOfUn1BtU/YcWOCcrG
mo96gsDa4W+jLZwewPZzdkXiBFzKzpEGlVDlB+NFF9MbHCtrwqXt5JKDNKYYob7s
mvk73/eXF6HL79ubv1NVTPb3rnRVwxwgKWuLUXZhpDNVRVW3y0je+Rghb+fIu0mw
oBGvmd1dGDf9UNrfY5e3coivb3OyRxSNK0vuc3827OLaotWltxAEXTPzMYOrOCEY
QuKAvpRLdBfObNscVIcORH1NuScNJPr2xFwUUHRc6aMmnrSm5u4FEVn/j8hKclrV
3TZ2sKCnZD2cns0+2A6qDmTz9NJLGqdRcIu+gcpRcsA5KiOngqQ2OHxIZ8BW8RF2
1fKuBJDTS6Qd2XXr0kyvivEgJWaBfMBzLVCVYspv4FCqsf9F2PRV0c7haFMhHRs4
1PifTztNBJ4oeBulUmaiarnaK18K33VItzJVSl3Bj9v6ej2U78beVk37k7PmkuJU
Iear3BDtW4fm4ai3voSsM7odhpqUGBgvOSfZKA+mN6cNYMbBsF6AOA9AmiJD819z
YPtEwo3idPN13wAvrtZWXbvxKFeSKGwTeXNkBT/e8QcQSZcAxP6UvpQXapBTJL19
4SwCVPAU1+U3NMhi2gVdZeQ05EVoi1agYsc+W4folwUFw74Kv3PuL6ckisXaKAbk
7CTBmqgqSlVBY88VOXaTqdsu/QVl3IQRQJ1OOR2BzTl5Te3Ty6Acp+skFwqJhF+T
5gLQgKT0reekcC5U3VfsiT6LY07v2+Wuc+ZMSdbli2PRnUSl6djvPExRSPD/aC2x
FXLrtPb0ryqJludkwNeoFsqLR6qZSOgLeISewEXzRgiiFOEwe1GLQb6uH0Xjf4Bc
hcf1y2WXR3GAEGt62oTGfV/nlJjsCexcpe6pi6j2FgmnA3pol20O57dU7k0ZYoqw
OTfY8cJsvXjt2SRjpzl69gDR34nu4ijASYuIpwl+h4FPyL45qT9B0jnB1BEzyftB
IsI8IwZ5BypsE0iz5HwNc7pB4v1/tun/Y5NsXQ2UKuDrJx7B1d8ktDbhyhUSzsb/
5DMUEZ1oYTwAl2AkFiD9IObzOJQkpfhWhRBGaIdMdwZjzj4mVEQa0xp0jreyIzlt
VuSZ5Wd9Vaf5tByjT82DWXDZd2P1Q5odjwutVpP0hWGWwgUQoaeZiLQ+wUVQAy7V
9s/1ivsQpwJ62k6Jx0OHanjwYTarYt1PiZkjLwGPcjaONy+hUFHM035fOdWizXSf
QA+dXJHns2ZgkI+9mUiweDBBWns0k7oRXFEkJ8fBDbxcnpUOXmYSOQDLILpHf0ji
LrSXtSgmjtGvNDFbgLq5rst0yVjvCtXwnLXkQRZiDYRQW1bjszkuz2dNK3WJV7BG
x2Brsbbxe9sE7fQ7kmihh1sNHmF/1n9SnWJFzOHCBeS/YFSWFZamH9W52ow4OMfN
u/MK0IahRU+hnI+na4IuQdbxTzkcpuZrk+nkvLhChhHEOP6ltusCADCO/fyE0l6C
GNCebde0+9f7cmyuS0Vq29eWidwUddAfMM1u72L8rXicEB43BNvqHovxmk7inP/M
mXbLJYc0STFK0mNKr1dZ8qZ3f3J9PhFCeayfYPpKO79mFnrvzdkJl0/pOODfWAJi
5s3Fl2H6N3frYup2P2+NLTwWkYTnjTyh0NKwJCaDNgTwwqrYeAgMgxKzcKfXhnol
Xhv2+yNwKGJpnukza9sXDufQgbI19K5XHTP5/pWo6NiZcE+jkmm+4gc+0lHE/aG8
MwmylOsH+Dn8jCKJsjbEZ/nscXEts/Y9NvzJza2p1iaCW3nwBkGQNIGRscJjaTiJ
9/OW/vgu9Sg67rv8EtV9Wh9SgYgdtqnbGxsVtQHTBpObQEHECY8bDgVIXzbiGb6k
S6DSu1eomwegYfANSyf7A9xnhhIvxrOGnFu53lAolt4=
`protect END_PROTECTED
