`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QURjWwedfdClfqK2Lb1CS30lq7O+q2Mubskdl+4jSUoGm5Y3JPcE/ksOZMblHoG4
3CyA566NuR7SgLJW5mVsay7s4EkQiSCbqAuUU6+ToHtA11fCAeFAGmWLTk4MSlcu
ssu36uRIOHPHfcoREDL+0PhEjqoZChuFywu9Vagh2ZsW4exEehxF8Cx1ud/jyJoc
sD080QrO3D0bgXpCBVBfztxeg2jW6cyPmhYcRVsG8vnlWE5E+NqF+VYPTu7IczsM
5wzSy67l7JKNwfUrqH7t7RKwJQWbbsjhTA8l1OmfBfeazPfcFyr1uHPwEm3vDXrW
to/GutLBVlGchZ/bdg42DwFwkd/vBWRETzRvAtuWwIPqtdPaeUX/egiPQlJ5hF9X
TsOLtdIVbxwCCf0C9ubmZqDoU20GTAGgxXr+ooYycCoDvnk1BDmTn8gAK/QnH4gJ
u+Yb48Hrh9wFTaXfj6zuJ+RgQTvKoHjHLMXbqbE1m2EiIcAhCVv0em+bJnZA3Nco
F1rzuDc+nUK/NOBMbWoTMMvWITfMTsPJOZkTRpgYcXq201e4LCAhfjZR7RMoamyh
bqKzLoAs1U2+uJakUNJ5NAIrPIeZ7er5COyRNjF3hXSZTObg+1XCcjfpv5+wpIoE
q81ZiVDOPsPgOBXSsBZzmfwJreCZuYLVscGKtfPK3Iq625WS3wPVT1B8AYiGNajH
soyjfi8KVcoLYGTSlvWKYG4bHvuTsDZ0A7dFwnTREqtIfNmRUZ5QClj/xwl604yw
hfwfSW7J00nz6uwzfq3QJJN45S1Tiiv+GFZgkcxl/OYdBZZDafgbq8nFa1mQqCmb
8IbpYmmgmJZsIgWrQ/Egqr1s5Ke9KsSAI0y9lMDbzwIt45TVAko9VHteX1nUV96h
5UkWeQGPSoSd26amwB1v7v3SM8NQiMpRj5QhJIe3lT+WW6wkdTuhAm0nl1KW5v7u
iF7kWjJqubcFUVAvCTSk2TPHGh/nCJ4vNHRwrzZW4FsGFq0cMqPQ94imjLHNcoWK
Pqxfk6ejiMeCOhjBEYjUvV41JRxWb/cnj5IarcZr/LmIK2p37DVUflnBFNnEK4uE
X1RWe1Ds7CrfItA+TDyQ+xHubioLC+eXw+pjkxtvUXAggpgu8P0h9L9j2m34lCDx
M7BezWLo8x9fuOpxIsbpOvoQzeSrhXcjsmv6PKdiw5J4UU4WfF8AhMy8+23j2Nnz
0fjAK0CpT3a7M3tP8mffi6HRgI2KuvcFYIEC5cwY7z5g+NUW8fMnVbEOIJe9lNXR
knAAD8DRmIJVkYMhBug5aNIoojfjnaWQcIsWDm9IcjtJJdwrUQB7fTvB6+iA62DO
tSm++Pd30s2Kgoz0pWJlPO5qBSIRXjy0beZEYVeNkK1XF07iema28zBwJomNECsz
Y6W/BqWuWNt/52o07efUHRuP2CrhgApVN0KQRjt6qeDZTGgTI7KNkfC3CCE3p5Tg
Igp6FWqpXqGyNmJeC7xmKDiFL5TtMlETi1MDySo9d+J3mO1HYFtn7JYBa7ug1hvj
KaosSRAb6pz+eK1Cf3H2SFBitko6C/nQ6WS9l9oHQ7tDUGjEC7MV0y8RXcvoN3TA
aX8oDajY2kPZQEf0cGmCW0ZyTsa/H6DKCww0GoAASG1X8hfQrLxOzORC6D95MNyA
Cr6ICyCb7At9AiGyHBxdyuTlLigPFrtCZ7MeHxiQIVdbk3b8pVvkQA/mHY7BIHwr
5dcZV1xKoexOlK1W+H1gEgDyoYDcOC6W3zXPbAh68Dm/fQLfUcB6Q45KlrMA38hn
fQ+WSF6uQmNjMncGB+8kErQziM28aDf+NWq4URt6o/yonXpUO2HSSvkaegov0p8M
JlMmdwsRDojkPV7KPz/L8rDBQcnc2LRR14rU7e/zZOwixfpEElExdxMUqxu4EWh6
XQaeTIlJiYvlpNOay+D8KiU4wcLYeoFGUbZxXTErN1EL5YJhBhujJZWt62bEHTfn
iOrTXbpkbhPUghb/YZC36ANKwQxu5gM81bVlkZZLdF20brsEW44OYoiiWSDQxd9d
2k7J0w2r+t7cHbAyf87A1tDw6odOqC1x/4Nu7XSs6tFJjrGBFzF4PweCSmH1TMxZ
ihhU5Uu9Nlq5BU7WyAEgTjQusHo+nNuxdQZvF6izPsY=
`protect END_PROTECTED
