`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hdVbWihYF+UoPHC9tmpIRjDZvEy3fuuGNYoMrsX71KuEqBfzrWtFRA9BcQkCXzLI
WkbnSGwQQ4AvS/nYt3dxJAfDQE1Klxf3RzwYd7yyOs51M4MiluF/n3HRBHaDgYj8
Jy3e0ErXc6IgD8S33ZlVffI0Mjv4ZJWfjBxnFTbTbrzEJif1bBzu8uYGplBCa+1+
+I/UCBJAMhYGnyRRGxEWF3IgshOJSY8DnhGuNWH3Zhg9jJDBVAN3PvT/09QDpucL
SoklajVke6PAqq6vzdk5smeVwQ8vTAnz4lrEzDdFEegkHBu9+nyelI5GIoRSwDXp
NVMgZ1G6A/BTNTmknDLuVnXDl2q3Bg9dP00OxM7zseEGPoh4qqAhxAKEOlkhbfKg
UH5NsstfGa8wcTSvJt4uF6Wf6fSFbRwI5Cicm044o3c=
`protect END_PROTECTED
