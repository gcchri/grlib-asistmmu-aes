`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tZssxdiCsjtu4eYNtG1rhrBVOIkheyfPfYoPmuRFHGSpY/W44ej7TiZjGJ2pOe2o
CULDpdLjbSsZH0/t2Kwan9n2ng89l/ckqus0laZsNptTDb4Xs5amz8cGUo/cyZ/M
TWHEolBGLNAxOTIMdfNPUWvESqenhvXA7UtPTLCknJbsxOjTrB8EASHo5e8mCWOO
ZOGlKcILRZ6svhbn3Of8FhbF+CSBvDV++9vEqa/lBsAXHHCe/Gzbr/UtuoVyWCFY
KfgTIrTHmuCM9S9u5J+fhAdsvZjq4tD9FyBXyp0u1kH9I6gUJCYjUnP+2cJeulvW
/i3hMXUGOz5ljgL0ejRLqimyhjEtL6NWJaThqqwzHW3TGU+VJ+ewSrsZ9j3P0Nk3
njlYquRCoH7VMuuHomfYP5bLKh1l9Vz6KbczGSxYge1r/Cbt6V0LIfmLcM6JiPnK
AYJEBoNWHwoiZyWr/1Xy/X0cLdAMELrCXUO1r5E1XavYd5u+VfgxjRdZrJQKB0cn
`protect END_PROTECTED
