`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6PM8AnEn05LGIfZbEmgX8ADuyAtrcNrOCzyUcZ9P33VfWwUx7OjmT45wQcpL/OU/
DKXNLft1dPB9M+o5ae5UOYvcygSNmGUnx71Z19+E0S1iqqHw3moe1X7ION0p7kj+
vjQIpYvO2DJRbl1Jqh9yEboqzLkqLotMqaighU5oToKPQHBWClglM2syZfZnbDZc
zZkDobYJc5nkdrkgPFJjpiERrI4mmzqEokb/zleGG2JDOGX0Ih3Ko0hPyVrPmi5T
1BfyPzswaJGkK8dv6UHgPE7s60by8NtRZ/MKTmOltnBhnanGW8E6QljrHDfWE57Q
4GHWI3BobDzs3mKnV3JPncdOeErQzPipaV0QY8eJK6JFa9OINCisgFB/syWSB+Za
v3Guw8ZH4ZvvNUChNb6u2htOwtrjtAJlj3Pv6MDscfbt5/Qitk+x00GUuBqfskA7
vjQmqIgQnNcmuxvhtSN6hP0maRtTa67ksxi4Oazooq7IQyURcL0oCOJ7HRNIYe/i
YIcfZUd1M9fTcnFyzBZwLOKQxIcbVE34GoIGeHV2D4WNYTVsSlX87YRFlJg+8fmD
s7JLtDRjUZ6i3qDgu+jEzdx6KlJojzlijHMzReDpvOWoZFGeFnt/Fi4E5jbahVFc
aDgU/u9kFPH7TNoxwYTnRe0v/SGAFifQUjMk6qkwp30R7AxuPBrj7ylN1sPdJfq1
Og5fOCGHqSYJkBxcuY+ziBr7yZT2W7a6n0B9/UCcdMY2u5AJGUSBqD2Ny50Vf3od
hhvqhta3FfFOJDKUjVPAC8CftPmiUR1KUuOLLhHAzUB1CS8NJ62Ct3XkL8OshNQk
+fYIpFo5lC9auOm6saZ7gl+UAOolCGaP00Go09bCs7vh3WS5F9WWqqPskM5nWlUn
sCX6HaTuTdX0KqrApE5xRLYXqldpEzvzJld0x/JThPs=
`protect END_PROTECTED
