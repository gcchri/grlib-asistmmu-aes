`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cUnAXs5xjD2gmawo0Hn2VBpy7SzrcjX+y/nsgtG9ERtVMoH2lNq0KTm1Z6NYY88Z
H1Lt4W7CuMAYO7LuHlMElJ43oqdsHmigsmgN2Tm3sRbaoIjwKBil6sviCmZhJ5VO
gPBnp/9ZLLJSAAn1W1MabVtKCMENZ9MmWqQDSKC0wuBrWue5CBNx0/3nqEcvBe+V
ICpYjvSWErhJt2JMcwwmbrluMyrKz6jpP8uQIphA360=
`protect END_PROTECTED
