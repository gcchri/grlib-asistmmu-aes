`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ef0Cn42+p5xXnmTDicCVr98vikom0WQLtcgvkuh/8ze7XoYqCGkFg3PXufbetWHz
th2YqKoVVqO53N8uQadt/BBBpxT/nWfN1M6fn8IAIad2uQLepg03KSxNqpa272rL
bds7rC0ToVUo+j5RS+xUBwo8K2c5xJ/mmjKMpd6KkT7uZs9IxQSy+j+PjKQiZllu
xhxn/uzR3X3G916Lj/2opVVNN5FJYfc63xhU71raaI1V75qyWe1xM9XqnrC+pswI
AwgZDtp/I/3qMPMDXuNYwAh0nZ1OuaFLUwvPPoeOQ43BTrSyCZS3fnFxjB9A8Pj3
PKboRNC2EcTOoj6+iBiTlvo/gntL+9HT0UFKOm7NXXOQEUJZzRNHrd9ytc/maKsO
tzw/xf34NujARlpRSdg6BBUpEy//1s79k9BfRRSrqTwkL5zMTJlr+Ih4K139JII6
cSGpdEupaDYfv9dkABYmvHYPufMYDTakRkH2gV0AwtZDP+I4qnR/gcplT+bDJ190
nPgxLreiDpeMEQA/3QBWMRHbuV6AQfDAuhTDVe+xGxSZOgzvQwyT3biwIuekQFdw
zXaJYmZ8PEjC4JvNpJAePJkVUOcXRj56CYCIjxUwK0OrnT8GUvrjDQjsfZKRS8Jh
gJfkCH2NGvPjIMFqUY5eqYqOXWdHJr0zbRo7EPLOD8E8LytMCGXfDOFYIZcLQzRq
WJZtku64OnhotZ36bjwO6ODMNjKUV/mQIXDOi7LZYLci0fbzuXY67EEXHzJgHZFn
YrWrZJUsIOTl9zQI9ORh//14kJll5/07iCv2D5eZyvVqWv+KFBBKVnZ+sXUimLQ7
96NsLlpIuJxlTInr3x7D6IMKCS5KPbX7DiH2f/LZbFRf2dSZn7W7f1CGsS9uKrcT
KtVzfQJkyPsR02fm/CD2xLfEDHKLNDo7NvdW2Ba49dZEnMPiGA8y+nhiA4GMacH2
2j3x6uIXM1oJRX2//SheW5T0REWJAP7eXh1EojIYkNTTh6k6wKwzeFM877bV6DqE
9IgZzpY6VjWSbhG8sHu8kSoN1FR8vZv9wBAPwabuYWv8C+tQrhZniKWJR7TEcLvL
gKbS7EbQIGySmQxmcK3Qv+/wEbrXA5rVWxsufG+PpRP+rnTRyvdWa/Vp4FLtNAQu
u4lZZu1glZhNL4A42nIdw/nfzof0cZG3fwa8Yv+sCMN0NO2/n47J6oOhm3QwIkEH
k6kMHyOrGLkrEI7/B3ic3R2yXXa4iFEJ72s8IJlZ49/SUVKQiRUiexf0ISRNSO0W
iDgWDwgk45b9nld5gNS4d7q8IXGgxnP9uoDZoQCaRGx/X8vDXSoIRPBy3l7501YX
tiJ6Ifmya0+5lXD04jsMr01HlaxE//Eb8hTH3o8Pu8krvqujKP3SkP87Xvr6bo2p
m/z/cNeNFiyu+Y+MKxLVBLOZ13FrhOdWyHhjWj0eOx7Ell8ROyk9mmXgdddMl83I
CURWU9DgXQaa001/KLR9G+sZNi0y9xf2Lp2U6bglufcxCISvoXNnkBEgcJVGYmEV
8neyV0FGZ51hOldd/D/meC9lwB9ZcS6VEKlsJtRFEgwa5vutIUyXRKAo6Z9q0SFL
59dLcZgdG4ROed4Z2w3N+dkew9CHp4qQd6JYDmQCeQTd/ZdkB8RxtPSeZWyH4PxF
+thUe0rMprYsCOZLbPqjSU4cu6CorLUoSxzjNH1WIUJN+KjWmadbLplZIDlOt5n8
KQEb+BTFnDr1DoimQ0LIsxSdHsIHzGTwxWT0sAgLhmGANWNlkhXrRSmqtYo+Lhuv
lFEEjnhfIOsgAucQBYDPxkB0MDlgaAkubu/bmQInqwhlfbX4Y1VtBqzI+vl2rNEq
Z2OpTC59pnifhgyl11K4upx2NUpxE7M1E3IpTOpTicM8gRHfPpYPZCag6aSZLmlA
d46AAytKRSFnJ4npVfmaZb+iEKa/Ht6LEulL0bGah/rUMtAKn1mtHWmpfqCmQTgS
hmCzFcXzilXaWmcdHQSA6WyxWvT49D0zwomXURa2wn2fveH+dgS5TEmQ0eZgsPq2
msJHrSgnNrrlX8AEki8kdQnaphXMTGMaet1WxK/lzkeZ7k6m6TMo/M0mF4qK30Ta
+4rLyeY46ajuk/foqEHCUD15cu0aERm5OVBi+hnTKQ3GhyTFWU1frhUJy2KkDVx1
KF/S8NW4MPgt/OauqNKEl5F1hI3FwUGcqIKsli6WKnPVJeAXpfImspiHetseUGW9
nJTTQ470wwekCvNk40WeFhnnH+vDWB59iFFGt+MbJCyhtNoQZQ05Yke9ZNZBn846
WC83+YBo+JQbGGAskXqOiFjuwNkNtXWEHCDyhDrgHDvpPs4AqsWquTuM/4BiSGJb
CM40xLxIZxFYBbXYyp7QfHHFORgFLgm6p5wyEZqPSYIY3/aB7p3jb+T/xy3uEZJ4
0AtXzAUI+vUjDuUF2uyzNEg6T/I+Ov7A/+4onUgU4a7KurIXrvyGy03A7X0csnjp
o2KiTIDjtm5aX6QYaUwhDmU8LQLzXNYONM5MQZfUPUNEVCqxYWdlMVW79cwI/F2T
K/wlNgxm8HDP+OGqkzD2tPUJ90v53s7NoL9BPLpEDo3gRlnONwNx+jIKG3t7MUIQ
3oy7iEu9Q1Apc7oVo5uHCUiqW49qDnjSA19DBChhOHC83TGv8bT3nhCCqrhN+v/+
1JIuwHebVWr1Izav7Q9jrNX23TEBYlE2Bz+m3WxwqTHEZBJlmRgE6oJEbaZW8eIu
D/YL0E48ZQxNxrETN+DmkS63qV+cNmDffQx0x/6xnFfwKc2lU1dPyIloW8AV1y4Q
sBLE3zbKiE5EDnQBxcI240aYcL9SZTMoBudslZEo5uBdzDC+TOJytjrhTIz21D4N
ssOFOs2PVMl8YZ2I07oe69uCQD8Jbokc9mw5y+cnEJ47ivj0CSJeDhobaSW1qbkc
3jrPey2yq9SR12+HfrKS0bvd9gCxyhPnCsvGFHuIJeQHPl+p0YO0A/dJipjgJ9h6
+0eZ97qhpbBD9rk727jNkgz8o5xum7rkV/SohMeMCI65/U+63tZD6OHblYIgwLRu
wX7uXyftnIZr8CkpzpNhc0tQoGu9Ubm9Pb+oBSmYAjbtFr550SbAKavQ5EEX/jLy
tUqSRuOsudkkcUDYkfSHcMq0OsobsOPnmHi1FgLKre4Yb38aRnpRWOzlgkEcqH92
u9+1PDI7n0rzAUIv5GjjjdUOEL15IYS+CDbMUO3tamNaqd5gRXUaLiX+V2ah7z69
aBEHpG3wvZUarKXc6rsuocmViS3OicrLwnyxzRoWerR4/hrN0j+7EenoaKgmpUFm
mHvp7Af6dGPizqxOty/bYXnbjInYTl3Vr58NVgOGlLb3end+p8LwWdmJ175zLETq
Zug5LWVotBSD6OGQaRcdzvZGtLLQiUXZ3y5eRE5f/5slRu7sf+OveVD7rBD5DZke
vrBFCQSWqoU4tKfITSP0JOLieqbbhSAkWpWWPZv76uIiSQu0pM7DK0stCaygVW5/
TQakppGrzWTfh464yi0pFXNoRW4WflK3a42gnKc2wX2/BJeTCfW/pmuIzefMXQVr
fsZQvRa5qK6N8NAEDPChncWyFKKJxTveEzV+495UJoAwUC6kzIZzut5JLJsOKJXi
JUE4FTklldGf0QWtV2HNArE+gybls1nU3O4j5JaLcmUqSVyOpO4tuCCsNPuV8rrw
Ae+G4wQ5ctFrtcvjBoTLc8iolv0zpdmm0uzYxd4IUwOvJ8bm0xfqnDrGUfNeplSs
4lJfpFsrRsSAE45bOV43a5/KwY+vTMZidMawEyDjK3htPLRMEZ7bHk3pjIRGt/Do
0o3DhFenBa1GkMklNkl4WLB/8lFPyXnqyqI+85HAuk88o5GPQyDAS1oLMCP2pZ6N
BgzThA64RkiZye7rpFd1yDA0rrwbZixOyFNWHkCAeYYLIRQMe7b9Iqv0iegShk+n
y0d8CHSEmSkBxgPFwCxULLCw7SoNy4QVFbBU/e9Vf2h2rM/Q5YzFECg0gIptgOAq
7CsOMvzW7BwBQlq2K2QuAShCKdsPruGsLxR02O3z8hoIp6Z1tKtsvhxtvwrA/M7j
H6CnrPzlJOXp3z/HJyBohv/eaJpZjHNmImKOIegVvO9RmHrih4MpgVZODcRTTps8
eyLLo+tvqP6IW/KQm96fWt++4d/jFW5EKNpaA+aCgUDVlEI51fkGOol/QwKL1lFW
ksOFWGmwDHtzMC0cSY+DqHXHuCdLiaL95QnKdyTxuVPRa2sTOCEAii4NM0w+4gDb
fwig874Hc5F/sztfdkw+udmMe7BX7oy7Ap2rwXOI8/wGTy6Bftn26UGosjL9Bv6o
23CGB8rUkvKflgISyby+C2sCzUceduvo8v0YL1Mtl/cV2rd7J9Uh1Bd05dLvz0ts
/1NLMRWH7/cSvVm4B21TREh9EW6fmUykgoMOsAo2knPI1NTDJKcyFomDbxLEXQM1
nh4efhQAeuad4WFCCFltEMsx/Cjknd62eFTDN0G3jDBNIlfmnyVF0t5zInQH72G4
gcocZ92SC8RhyU5BcrTP/9apGibpGqtg2L4HPwF0EGMRLmxHJNv0k69DOy19DFwH
kUAKOpOId7IGNkwRqUceq4olWAJWTjApKQ3ccweVQaspY0HK9SU7Wscq6LVD2yp1
KuNEn6i5N27tcLnnVu5Z42zI96FvzEURuu8IZSP/oMksnismViAyc+0Ynh5WwSA3
eJ+M8IxEV/zYuSYjvkeKasou80luizhl+8XIklNElGsIS0d/EGW4xQvkAhAXi6Jq
bSxcZs2kaURrzxe4lImh5py8J6aEmfrt26LomP9FOVqDTha47xqbkt6ow5mW5Jb5
Y0yN7pH+5RbjKPbZX/eDRWnudmtb+VDzT+ngokLAWbb+IgnB4/4c34m/AS6avo0R
ufkwnTo+Jdd1zlV5AnyG6wTcKk+3K1XoZMYsm/zi0SOa9dFiuYZAp5mhuN3Cp3pr
GqzjDRiHrp1ZbFozogDZmE3l+x7n1P9kb1FrG4xK1cMp/WvxvuXyMxpEvXFUtism
rdtWf+EworUQDhGshLHRMVunhnnNJ1t5lDmhcXck+0qXKeIUWfveBlnwekRdkRaZ
obL9ZrrnrBNxmx7i3NDlNcnIIu0JIttQ2nqGGWFuDgNQqkDwbi74+YorgD7nuAlK
s/Br0A0NhpZQmxdTdukyFBr6BbbYoENCxQYv0xdkgEvCkvZI4K6exrnqbyC5tx66
qmCyfsZo2MaBgJIvh5PSvRy0nB3Xu3eOvRVUHP2uPfSp3YTIm65Cx8n8GdX5F48e
wTXzfDZDCy0agUeQkLCcRirayIejaX6FW+IMkDDKW7SW0vbM92irGkvyp3yzqOVI
IX5yByEDpom6Rz+c23cQwsyt/410En3OHmSIgocvgdR5B0Pr467Vue5uHdIVsW21
VxyQcIDNmFitg1Ll0Cs71GvLNk0pTkdIy7bUEyQTCseiAxjHC2VcmoEVaHci+P0g
tLNACqOpC9gbzZdLnim+sYAf7q1q6zup3nx9ALHEvxLyz0EEUBaBiCTAkG7NnkAA
AGujdN2hNi6m2jSn9jsXLwQMSIOer8e8X/vo292tp/lWLQs1n7mFtpnrMH4ilfJl
ze04jnUZezG02MhwGCzLpwH20Ib/C7ADbUDBe9jcwa0dpDpch6Zp/+04IwNdihle
nUicq8bPplECWHViuCpoVrLeNr/Sdl7B2riYjL+r/2NHxonJ3DSg8VxOMOL1J61g
xuqmDujDu0GaSb9DTmVUopXsY8fm/x/ONwDH9CPAvkWdZlsGuExeSIRAB17VEOGu
11Xac4ZRYvQDrRpL/6WDEFY3LjYDUMjmin0k+/yRx4Faz/GvANOefgpUnC7rDKzM
2ixh3e08G/1JQKtp7DqH+5hwE+CEYIT2t6k+nO7dghIoNgNpc+MnoJAZzLjSD2rl
KjmcAgtoFdxu/PRi2qCPmxdojTUKmF6fC4id8rGbtrfi4VFGNLE8tTJnmkn39YNM
eXgQrM6bZOG9mVgr4jd8sF/qXzAZdOYrYTO7XfXEP8gupcAWJCsosuXOBi8sRn0m
C8HuHcEGaynOZCip500Vi8LptCpq64PBPAf1YpKfY0OfkH4ptLw4ZLug/Y8Oc45K
pU6T5wRA9BrtEhiBY/Zxt710CNNB3T9xAPiyRX7yYnReDHOsDM3kzJTqWfn5tBSd
BZ/ABZwf7wfYCOPnpx8DTsUc6Tayx9z9/VTJjS6P0fZdSBI2KkBBKG4XebhhcLlB
QYqTiYBwBeAtjKab4WXSFRuvUFeVE6XVpY56H9BUiy2uz6U9opm/7BLrueSU5DJZ
FyeYl2hItJFFN6GxmLOu8y1FDGwiKw6z1oEZfkD32UI=
`protect END_PROTECTED
