`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CwczsEhSl8IEP6Rq4Jej58eechICCE5chTsm2mdClvuuy7y3ls6bF2yPWYhASMHR
MSv8mPUC1mAwSrNrXeFlnGgDiwQxMkKpHxJFwlQLXD6LqpzkprLRa+ZypUkEAH0V
xiAYoT1xsDZ/bS6yVdZmOGUIp3N2Lr6Cz3xUFPLr3wvSy9W3l+kcuNNw1y8hkgeX
52VXBvgOamWiZn9uRAiIHGMsaqPOjD0qkzh9OBFxxV7Lo396hN/MeJVyW1uZ7Drc
+72q1fdXlkwrq1sdSOQqsgVcl1ZDVVbhtNPlWdqaHGMuWA6iOVVc4wk9qGgyWTDe
xekK5p0pkw8H1jioTZIUQ0RapM7Ud1SQ3FBf3/n75m0ZHwKpBUVvqeKO+Nzzxxq9
RhfhoP8UFbZXF3tcvUEldUiq+BT/FGEYdeBxUa+hcLGrnzr2d2g4OdMQ3jWsRsF2
+vVkw54KVuNkflLxczf8J9NqavwUizHvL8koAa23UBxa1KO3AXVkOTVfl2xCNDSm
PrANl0CnqWj9wmRafdviT9+N9RYaNK77rBZvEkJymDVwVzAEaE45RVYPgQj9n78A
TMuCHY6n479p3a9VVn3MgKjpJYIScr3OlfUcsnB5fqroWeG1DYHsq+WDNU4hHpQ4
8UdnktOBn7MU8Hf8McD/oMRDNgrwR7zJVbfxF1ET1B2R3NipCR744CjfSaicOlMu
Q515Ilx1lvIICCO8puxKKg==
`protect END_PROTECTED
