`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NsBkvvs1hH5N7EVrpto5kqJTv3pUlDwrALxYnaf3QiCtARGkKVMifqez67yvJn7y
zI7dviWJI+QbLCxnkesmYnRuxQyvGqcmJYC0nVRALWP3DCzwUxKuQShHpIKvURK/
u672LYQfDM4LZsV8teQmi/06jxS1V14w/rfxteuywvJvSvWa5mH85TH+iUPu8YuU
mcoa+BDyTmehf1jjsem4M//gZT4vreEU4zpxvhQlcdY2RKQ0zUGcmFIYsqkBnKrU
jsAPCmr4Gfj4713kSCdWPRBq3wNmWecRiwKIPuiBzho8+I+VRMhT+ZJmi0bn5TJk
8xgTLfOx/nt+aI91PwM15OdPr78d7ohJlJINI4x3wTSrT4D1i5FDuwIgT4+mUgJl
2e4+EIKfzJb4owA+2vbalJk1mJ3+0a4k8ffvUU8sbJs=
`protect END_PROTECTED
