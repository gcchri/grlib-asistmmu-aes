`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9BM/zwKQjviriHwzY2aE+vJYpMQ0r0KsL6tfe6fYghvOcdJtbeabBuZnuVN0Ui2
gcmEdC4Ollu0baucFvWVYQWB9u4BnswqHmo6vfRzy40h7WYhU/4XceOGuCvYf+zV
nkYQpgqKxUmblkgj0mh4/RcscXI98DWereir8gStotaVjd2UwOhPGkqKQGXPfbIu
2kp8PbXeJoWk67A85IgWcb+3Ks+3bmmzTOfLlK5LxpDHdZQjlA1grn1E4NPGy2tm
2nQ3BEV2IFdUfjAV9gxWlLKo+sQS/KpwB+/NfGnhs5m0VGR5uf4NHZf9og38zJzR
H3nq9vqFYWOHsX4y030xKC6qKw7jf1nGVn5lXzZrucFYCgo6EvW8z3hAuIh5iUbd
pEx67yjJ3xC43zGHliib/p3Wu1Sehn5/RKkkTrg2nbNQbY/8Z+vM0MHe5htdZDY4
L1PCwl7iEC5cHwZ863AxK/uhkol+SlB0oVCe9KIimrrvBuWEHK+s5tGba733+nkR
Ss6mfEptJzIpF2qNFZZXusaQhbcFFUjWKpOuxQ0Iaym1hdQpOPHVPiPIG3E9DDBy
UEfl+aWPJMZp1tEgRSjkD2EUG4MEiS6ZV8kU/l/hqYAZr5Q1C953thWQ5r/xNOD0
2jSGzqKmkoHWS7CVBSk/bfzkEL9+UGCTe02yyb8oWCZ6rlFotlbJlkM7yZe698XX
yAVSUWNrzDd49sweji+q1f8TQdXSROv0DA1gJlFEZLcMVsYLLFhYRHCPuM3RtX3N
e5McDdwwflWztJ3vrdWrtIyvnorqVUFBBcT8JDzc7Kh0KqtTq3rdmA1p4jsqEFeW
PFkTOXJBSLlpJhEuZPoRY/CAmjKg0vIkTLvCb5CoDGS5va3qdFe/JM/FiAnxcMLl
`protect END_PROTECTED
