`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rRzO3/SedGDNB6Ke9vZrt0BwCKzzgwdb2sY/ASb3o2UzPHwTne09Kyq4Ge7zW7mv
l47TBwSNdhLCPtybjW8RkeSPiudRj5XqjdrC62YciBRDWOLls6LHnsVQt8m3alHV
/o2BfTh5cYZq1SKVEW3z9V9WCigNwdX+JxcZY08icPZdjrMZJnmAjmuDlnWlnTdP
1jM8kgB/MoZoZcZtt2z1xn0DmRMYfMs2wxyjIaa3AYIqUVVSgKe8HrGltA4Tm1Qn
IDCOl+GTw78QyE5CNMy3kfxJ7CYQw1Y26slMWWOm3lbqD316Ez+zvSviPC/u2vWS
tyMUJ1MO5HpSt1koBslGS7bCpxo9vdlEHfukqIEayzpeyuyR9xVXWYZEx08U2CoN
YbRhN8zySpPUsL76u+eb/tpb8WtPhf9/NBw5QqOhqXCAqFBdvjc8BVr/jTgtcPgG
FUqmCSesGmlCQgamwlghgRNmbjjz+j1XhJDPZPAJ+Hx79hQ4Yjsbv1XW+wRJBlXv
vHdBHa7v5UJe5tWc7J8F8DcH7x6osxfodUyHqC9eMHonb75yXXlaoWa2SSY4c4G8
513c42L1AdZTvj2EQQW+fS9a3VvhSg0EafGxim5IswZ/Qntcc31JnQVP1BPJKlpp
sRMS3cTHcBcTNlGw14an3Q==
`protect END_PROTECTED
