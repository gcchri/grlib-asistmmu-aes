`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rjUs1d5aLDKihcP83fF6j/Pu73lKgDqDqdsi3FAqgSkgBMxdh8A0ZZEQfs9Qg0d8
vcwOSR1hl+mctbYwhjoulUh9tT+CFRdd83/S+0QM+ofh3tMCh8prIDsn5LdSg6Na
0gVRUbVAfardOsK8MFAx3H8iXxsuH7bqobQ1TgXfd3XCN3eqBF6vQ8AJQlyzIHHS
nXfwSTywU2gLc5NNfoUuVAlU3zJbIH3aooGvBMyQYoLrq1FNb+YFYdKBfJSIx90m
IQ/OYK1a6uJ4EnZJ2Sctv3dq2DAowvOUDVqnL5qwc0YpI9mSU4TZFmva4Iw2Nx7K
U4z06nzkvtmus/AjRV9gOgZQd43wgyyEQpGTBw2S03Kzp8gIASYaEk4SReQxYgf8
BPH0nouEHPfil/E6Dg/sSy8n4sZhnBdRXbQtUrdmMNX33FbwXVZxw8N0B5+ujfXR
b/dQiuHy8FC/zPjU3Vmg4vgKnCr5nKdenktlpFSLV/9V1NRo901HLGsavEBa7vvF
6QPf95Jpz1u3XRe6uSchBAY8r6/rddIB+1nrhsaXL8sQVAUPFAWCjlsF4joMDKtr
6GFPB0C1drnC/4/tQmh0IPnbdBuRq81J4FNEr7wPMRWrVQPHOnPIf7QNOeSMa75y
VbrQ6RHAWKCYIK3KYdjWsOQ06J1ZqUV8ypUoBTwSFsssKy1rpPLZMUeWcyMQijHE
k+Zcm6cqPQ56VzsUyA778Q==
`protect END_PROTECTED
