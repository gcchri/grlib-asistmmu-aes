`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sWICKhXGA4VwlVkBz4jhi3IILezkKpKvf1tHLEG+xsFl2QwyZm0BkvhFvlayxK9G
cv/KuN0g8izpK/fKUnipESA0EGb+Qs8HT3CGR6rnOFHpw1LhLQL/Z0Ss8aqOKWPE
50KGb9mjnjCKGTpAxT+eFnJZWd58h9zKmf8hjJINSalJk1SKk5fLBFk/aeZFHsnN
lz+UJNbhZHgbptdYZEo8/uDnU0CYuCOI0eJYjh2ZC2ZdcDfpT9yDm5O39t5sGfBj
y/Jet88aIVw943564zNFtbVLvIVCwR4v3ho8U6Goes/1eYEGF1sPsNGXZgim+HFg
qgjelRpfGQmxdlCQJkpVQPuoQffTgsnezor0C8Dd/DCFL51kGsBMn2pml2+qfCSz
GyeWQW3HixZtr4HK2GF3uD8yQxXdfWDBmBNbGmdIPkj5hIejF9ExiGqxU03jzsWi
9zoEf6T0nERWL3J926WqwNvsC0xl0415lipA7cGfxFCyjoxogGQhu/H074TrS1iZ
/YwQH+7yAbGzNPOO5v2D53tzUM76os80nic5a0/kabsHkDIBgXT+qw3qsy+vCZqm
fwEtWMyw8vn5MEmNWMjSKYNsORpaFTrLU1HqCC+/fs854UcMruvVbs1F8gS9kF2v
MRnHQTVx+5nxcAIqB4+reXlvVax1dzcAb+HZApjP8ocbpnv2H1q0XMOFs9kfsVOH
pl3bznCQPhi1iqITGXTcefCVDG4hWy2asHTI1EMFsuGbbn6OEpSTXrEYSJtrUgQZ
bkXO6OiK2OB772rHrNjNDvIeJdQDzLVxABXNORVenv6hKs6161C4UK0qCWiinF9Y
o2tdhXdlAwN0fRvPitM9/ywwRL9ZkOvXQzFkmk9ZQsR+DpTDn6WeXm2Xc9mKO9Pq
zaXqZywr3Cl3Y2K1O8mQ6UIczSCfLeWGxJLYDLDKMoIYB69RoRd5ceREYOVXIyJb
Crxd6trJ1vEbZSWgTn5zKjbKlFLAosiUlYaNKQnOUnLuXhdEMBL9DzBjgXTJ0CuS
3h5KHWMvMGGkZEbw0dNrDcGfcYxXMgOW3Cp2BCmSJReW67R/4Zh9YluN8T11oseF
irjjsajdMXg9KSv3loVdBq7sV66tu2aJGcyt/+m/o8v29MBdNXl0s0GNjDdOq8Dz
j97PCcDHQlvTk6iGNDCUzSfMFhnkIlAOx5huzDSl18S3DHXt6E4TL2mn/o9zjEY6
B5mcgI5/caAZ/GSq6mJI9VM1nitWVBbR5FPR0MumkbMe9Pqt2v1lqr+SrKcsmQG6
BU41Lt8WIFUrHqjUz5pwUIGuhNdjcqnvjqnF4O5KUepbm6xEdt+xYy+lcZYGIZyr
CVoI9+DoZX6ukx6le2VjPCOzRSwKT1CXDZjQX8elgKGdNTNTXbryA3YnbvDib2VV
CZhnm9Vj1NqDJOB8J+EjCx0Pnwz/+D1rF6/VmZMBPYC30G2gj39W0Ti03B78cVsn
D+6VcVCbk/BjfyTPLueZP+RgLu9D7KMWBGUV/giAMVU7XfZggTJvBvS3j44yZWUH
Ny7PJk51CHsQfetUw/H8hrwUBuzGLCy2GDinOfuo6wT//yqhjn7SaqEE5rsHZ/Nv
NwRqLrpzLtfeL3Js70QHQqBvkmxXBvkVHe0MvwpDG3sguwd0fVfzjejNaDjnR6E0
INJf03o6v+rSrAoOJ2ILqlzr1lD+Bvf5goD5UdGiIxZz31OhpGPy3BHakLAmUa5n
aTPDdKYl6U2F+HXsh6n79bAaTF8R3nrgYYHJGC2SiMLuq7ds9fzbhIKnnGsv/kEL
QNSQhSWkw0bIIBgxaQK3/92RSnNuhMkY40h4Iyb7yEKfc50gfDKj0o2HAdw+pa35
XUW3rTFvGbPiIh9ofsG3/9YYgikphEXqJzO7WsZt7pivGg1s4H9fcs0uOOkpbExB
M3hjwNjRe3jWI51UFyUo9H3IjNoo0XXv9528CIf2Vh5qcEAsJEOvDEg49JytFgEn
5lRSilbTPEPib/zuz0gh2f+pZHxPVRq/Wg47u2movRWspPulmyVlyTCBWe02pGRZ
8UGvLVW5EV29UYayuQDKd6A0rBAkGt7NCNh2YN8MmTgGwLduiyVuGgYHt/7xjl+e
mmfr/CLl0dPuAfOnkYs+OvaSZsey9oV0Fbt7spP2BrHLXZXMgfSr6HMKn2eyhOpd
6/+K575sX4Ht8owK0p9rICkD+BTp11MyHM4a7UFko3xjasIGJNotAIGpFOqfLdzH
HF9BvvlblPlXFayTtNDrU4Ulo/pvw5T6tjeCkpQh+93skFFicjJF23TkMhy4Y0s9
`protect END_PROTECTED
