`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LeQbqQxjEBGuKWPsI+ghygODlYYhrA1+hOaeMnKSk2u3E+SG/Y+O+N3pfkCP0Z8Z
jdXY78B9IZaJz/gwWZsy8XYCx+sx++Jz4vfYDe6WVsMjSz+duYmXn9dwrob0AQv9
E8aqeBTFeSgxSjR3a51WFbj7NyfG7FRVpeXb3/xQhACJVPy9jN2HgK0jMuh0kETT
Bdk83popZrPlUOONDwJgOEtyNuRXDG/GwPo+RrrJA34ii9OzkkxDZQI/VgXLtmKZ
BKk+8KvCncCqcW9Bcd5www==
`protect END_PROTECTED
