`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4syZ2u2uE4K/1fRNg+YXYphzWLnfUaj2J1ZUYqVReEfAGQkMb1oZOXZwlawMru4O
gqjh3uzoVbx15/hktId8+rj1fX1QSiHnBBoqTm1B4ncyOYgMJZkjVJVMpcwRX0E5
bgdUSVZQsbbSvkn5tYPP4kA/ocBwq6Gv7y48TGTdPWNIoxhXHzmTwH4Jc99kn1ZW
fTFk5owBaRHkq88s0fkOUrWevYn+Pahxb4V1reDfzcy/LjiS9S5Coa4HWEybCtbK
XMVNMkU7tS+4xyK+Q7McbpuJq00yNwkXDAFlP6ulrko33J5LvwpA0IDslqqOr9m6
2rRVhoycm7TrR45VZ6he5aJ7U3GQZnU48xuOldODzlo2HKs93dgc6HSgi0Yd/QX4
R8kiT5KpKvDr5+W726xyzcWLcSFEelzxhjEfSywTleA=
`protect END_PROTECTED
