`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ha6J9CbmHS2I0o4GbpSpzDbVTb3EEaFHiG+9NPgapL8bMSY6vJJxI1ngY6lUcocx
guGMhu+QfeAkKV7Qh5PpHgGFV8H21UFJlG4Cj4ut/3XH2pFmvHbrJxhwBu5PNF+V
P35UOn8xtpsr6H50VBSLYeTOrM7C04+vW88FFscHbP7nd8zdK+NVC5Pd/7dBPIt7
12KAymS4fpajbJng82d0g3qvt/YqjuXCWl0u8tAUWudrkZ9XvrMYjSku1HEPp6YB
tSgcvAUDLa9dJHqBQ48WfUfcHQQ2nWa/z1nLPrIVXsRpSZn22HB0nbGqLg62ra2O
`protect END_PROTECTED
