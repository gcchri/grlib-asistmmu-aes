`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IEJJyrMScsrIpGkOjSSom3GovGrM/amzolJyvHNZu/ZVrmIVonHJTRqVgksFiZYX
a6RSSx8rlRvjzmzW7Su/w9Hkn4SeXhZIG1ICl1L4uwBhNZszheCRVuy9vBcETGjG
SjdvsVLB+eahEGHyrwK34YLIKyAccD1TCV6qN2VUmalM/rOVjhk48HlMXp7c8Pzt
YO5ITFBFvBanWSr+fhZQW3KO/F5jHiHftd7n+T9wwcT+0RR6xGn4EXfJs2wqdLm3
z/9JLhf4YGf+oOLRdCKTQtvKh1evGxn/qrwN61mJ5R+w/s5zt0mDb5CPoFmToVvM
ULbX7v4d89qcd4naMAXA0eaDOvxB/Nys2nhnawEyiReVhEmzGj3pgho9D5GPpnSU
ZfCYCNuF4vh9RTd3jeNn4MdIY1CDoue4x1D4lROr3sNS+i05NgStBo7a8mkLyWSW
uJhd59leNv7GIEwV4cKPPxePSZTDsPCbKr7gPJC3ZeIPC94c86eMX59NEN4jEjNH
jHtN5iPabsE1qx6smmsHsIknjqMFfVUMHBp3B/r8WfzJ/Au+1ughV8dRIIMnbv+V
G4iLNCtER6cZXSyCHYsKvtZaAEoS9CA4HC5x8YXG4x/BzO6/lbiQLtyhq8ti7u71
SEerY2NHATo7evXPR8bOsXizpsjk17z/E//1h0le6aHDXmrY00JFW/jVlYb9DTiv
eqzpwsKH5HARz6iadbuCxkFNbo8IJb2OFPqvsv6DVi1bLEQRHnCVNGNF+TYgxzDH
P+elSD7flvpNjNG4FDcfNgdFlKJvjnzTKtFG1Y8tqYn/lHzqHxvuHtx1wpRaVN8b
fv7QCPkAVWmmyANFQ82yrQBAmeJ3iHhCc65jaj4Y6lHaXuykjfjITCC3tEvM7X/x
HIwI8QjJPPa5ffyEaDMuS5ba+z7NDQNHJuXKpW5I2BDafv+NmV4QTzQcpeSMPlaL
GtvGcSOn+Kx65tPnZHq0UvgRcaK93mIlzWR5oV2ypxa9cje/B3A4/8REAzX2samu
hF8UpzjwOQA3kVKctnW+c2cUJJHIHbwZI7P8nikNstha6jTHx3K0uuSDf+oeEel6
vWuubiXYwU+GAdtu1kWp4Q==
`protect END_PROTECTED
