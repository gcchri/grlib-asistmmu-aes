`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8qOSod3rRRvmIgeM+1vUhZ68lrEdnwWdOhWMim5GRCJewETqZlFoZxu0YAx+8paZ
d7OZ+TNoYKXxORneAMBbuSnE8cwvXApx0GobekerocJaOQWyZAkH/RrLs+kF/nXM
rDcKDIbF/CWkcFOfVkz5qW3R+fo+2QJDZea8EJNwXwsjU3aLCQdQ2DtZqScMPE7Q
YkzgFy0eKFhvDgx+TTgO1pw4cr6l288l8JNC8RxW+OLZPY5k2HcPN7TJ/hGqeFRW
CLjZSnr1gzYenuIe4X5XIQ==
`protect END_PROTECTED
