`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
am1qwhRyFbcg0ZQ5p3LEB78WVl4O1Lh6N0cFrpkrmleN2IhcB7rg5UzdYlqedEbT
zp1m7AKH3HlQGZN6EaomdB7uzYUFEchv7WhcuycGjLleTHlhvY8jZssHl/XzBJBs
IdX8TN9CAJ87Vl6P6W0lc64nWRwxVVAIge1QWDJ9z6g1aW2D6LjJvcNEdxHWBY3f
4aDWrkOFIKFBTqCibpSfqe3dhLVpFbrRE5S69IQkELkyCFvUoyljkb/ZgZvPR5vp
fOpIZnW+l2DMhPcZZH4TgU6vsS2sNwjp/KgfjjAgz9d6m3eKXJe95ONio3LJr5rx
Z+vH2t4yOYVpbI+UpWHOKROK8+1p5uFUbolYCfEkT/W8s9N+JnuWnL3TovdYatQb
oQAiE6kwq8RTYjvrbROkI+lZsQvpN0634b+oCsTSvVwyYsYntVRDTLZfbVAPwFZO
VHlBSXj4Qsv1gGUnKEkJPr514EVs0C7svaB3JMoQF6S/gmD4hg2mGloc6TbvxkI+
JS8ZZXR8kC9/zZZKP2EBTXjZ4d4zSTZc6EGfP68/b+Z5VvW6FRjCJePA7vYNi2qg
zKJJdOBLFI7j7Adw7J2Yu1prCTLL9qVOR1021vdGMXv7f/wjJpJLqxc/RLc9nc3y
2EnbXP74fnz+kP6+FxqB0xP+qT4HqUaJ58N9kuhLqyTWHlBP/RdZ7x1wXmCXu/kx
oNyTr7kQXUrhbOJPI45Wk9p0yl5boBRzhjVIOxKyiuaA0/Isg9ZLmc/8eA85eY3r
a/p9q4PJRiPWm2fQ/fCZTUCCZCywQyMJRs6N2u0wP82CaKscUsvw4yPUIYrPz+M8
rvh+Ga62hjlYBv+vS8+Wo8hHfAGfDlff8t5bMcdPGZkqJoMEUl74EpbRCLmKySJG
R1TJ+W/XpNqNHHkyN/gkA5zHruRzbUkD6YWtIk2sdK7Ndgx1unTxXrvrkq96ret/
wAhbGvRiuGhRR9LgfgfSn5h6Hsa1cusduoJ5gZZod4DoPMS/ccTBz9WydNywBDbB
yLZGvTomyS3eppXQwFclcFE4dwYODzSuCIDZuecPJDjybBNr/7BIxY9SY5WvIJWp
u/F5YtJ1L++mabZ6p3J1mDXvhPncm/WzYFLYALlbvACXEwv8y8XhbOKop++dobkl
gU11AuAy7u87u+gIV61rH52xI0gAo0BcUo3BRQSDocsx8z2sVtyeTIIVajpMYLDK
MlLP/xLLMzlWYB2mM+YYRyjLiYbOFar1rtrRqP/jBqsGVY7BrFLy7P2ribxawBft
`protect END_PROTECTED
