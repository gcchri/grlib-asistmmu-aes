`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NBC1Y9WnwIAZknn/9PhcUKxgVJdV/EuZr1xzZixL+nOE+4XEDC06+KnhPfqt3cPz
GwXWc8gQaNBI41UtYicR8ovBwvdaE1Goe9S47LZIzKBAAgkjAZmLjbQ4fapdZKVf
Mob7J1vFs2DzSbXQrvJnf25DHM59SdXCrUFDisBTLFeZE+EW5DM62VOMN9Joa8iL
MKsyrbF1z0TVM0c21HhSgnWx36Esf5dyHSn03Wy8H0WdQfZYZ8xu7LsF5kCWEWIA
QUJXwSvM1K+vNXP7w25F5lluCEgn/0Yo37i8NMPjdT5AvTdDe8HtHQiYITqaPsXn
+8gaLdOIwJYPRvzuNngbDLrcTc7J7Lp9tsVEpMq+FcBGBGn7PsQrKyBGv9c7qksf
vQrIqhHRJEkZQAZQ3Swayjy+RhmfHp1y9SVHcC1iBGQ=
`protect END_PROTECTED
