`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2I1pdzcOquMHZh6Fn5sjcpQrNRKtsok+WOvCeTP1a0BIT9Lxxt7MI93tGjYJAuz4
wUeHx/0BKfsjQo2vLP5XIRYkl7OmLd3ICMOtRbL+jEQ3XTKhgOclziOUxbfCWJ3h
98Onq0HEGjqINDbjzKLl0H5S4X7RSEemXnTvxzkV7v8pBZgbL8OFsXZSGhtyx69W
yqLRVFhkAvgg5VDPk0zz/aSjB5EOJ2UCQbo67SKe9GLdUIpBQJWS8T++fSoXq4xT
z1JAtWwbiJC33xXP5GSLA8dPNmxyKGLgLf/2wqyNDpW1bfKDAqPbp3D5mMtWJ4g/
mT7llcabdKrlnVQxN/Tr4U7Gfgyl5G1mf5GoyjQuJm88cZiTAJNN9hnYEZtJW+Kb
GaLoX1xd6n4iXfGcBtLKyJmBvMAPjl0RNh6HEHh/u0FjdJ5FWYubezJFg9PokHQ5
MDT0ye5/A5bjgoC7VgGI0YI4/tyIXFt1W2ha/PJjQmoKoX8vMoC6Ch7uYkdYiCWT
Nllye0yku6p7G2FKc7qNouUqGpsR6E2/dc5Ppw0ZFD8e0SzYpPsR9W6mxzOPu1t2
mK4yNFj5mNRWtiVmoiXINEdOeknob/DLusAP+2lHTqA2xJbzu18mlBYs4w7aS0C/
8zjANbGU7bOByXPFYqMETrPWIS44+lNBqOQCIrgz9DcdM+Rh024aO9XVJicehtat
/kNra6T2RTWCAHtvdia/TsK8mgbIgsJjRAMQDsPhHCFJ1YcmW6ZerZfEXsVh+SZr
UNT9+cWxk2Mrd/1ATkJP3hjjqG0ODnDnzfrKog3xEwZdNtuRvDfw2MRRZlIPg3aW
91O2iuWT3Du5xpxkFsc8Kmpn95JeRAztAe+51f5lk7PTCPjFyYlKS3NuJc48oNa/
z7CmHnXpLPoe4XBTyYpnS0zP5lyxosBzupJNpXdGM/4mm4o20bqDI8CTb3Sf03NJ
VtTwn0Mh6oweUOchNo61AIys0oDmUHJcEioZDPX/U9iTKxBamapZPNc1p9ZM+FVU
Uv0Y4aPdjXneqGofV3/v3yUXKgTcwLeHVdpurtGmHPR3YsNfhChX8WEZwTU9gnx/
w6mbJNbUkgSYUrmngk6KLjely9eFcdxJR5zpY6ZwPKXqva9yn3f3SFicNWWWapWT
ehFClu+Qw4zHqlKVBN+ggLOIwiZ/rZx6OvMBbVix25FCCxIpwvNwrOeVFXHz1bb5
iRH3KOyVG0CpuRqCfdDvYggdM6cYHOKyaW2o8M8it74khsyUBvox/zcnRT9Zw6D1
lZJk6kXZnpjEkpsNjAw11TTA/HqDbAJjFauwl0mmgDsLWtOHy6RVV744gldsnV2r
NLq/DQx+uD397xgkOFv6L7KtsprWH/Oi1sv8uDR1wdta96oxlsXWOlJ8haB8wI1e
Hu9/kWLn3wUW1PsqhAFUxf7XtyWd3NTOKtlrVOYVlwWmf6G1sH+0pUtaa0mPyGe+
eiQMraaMG60veqhP9BYVcu2h1sbbClkPw+W2sC4H+uJOFrnbiwEFSQPndP/W3Tsd
48mXobAjNAfuuJ6ztH1PAKkXfXqsF/u/wrYkqgOM2Y+gwo58F0fXmvPp27Q5T19j
6RBQvwkjMDFhb7vh+P79hUcYz1r398H3M7J/FQy5Ab4mzHJBByEC1l4RFryxy4Og
/iIESTOq31hhG0C3h8RkMCeg+du8hvsrks/gHGVVFPqlvK1z3QFxU1UnKvsZTpE8
KCAVlfvmlBfkEs7H1glBQ00lNUCiv2BF0WUtS30n+8FaEYBdMd8eYP0m7XLa/v7e
bnFo5yQnNm+by3V4ROcx3d3peAQ9btfIl7SrfrF5lh8mRYgmm46TIew/tpwNFPZy
ZWyxjdfmOL+dx9yz48DdmRT+wMatTk5KAeMISrcwacEY2gFRClq/SfLf2fjswYAG
l+dGfO4XXMtQKx3hh98HZNE9vuZASZVSuCuxTinE/3aeNShE2jV7anhp0Y9WOO68
5Grm63WUiRe6D1705F9cxEW55/YPdqx/q5pAnnkoYhmaA7ldOJZLWDUX/QoZtaYf
2wvAeJgANJG6sIUKdPwj0Af1XoVMCnxDwFCoGHnLAuzeK3FBw2tYwJsc3Glpge3w
r8dmgtuKaNgfkkGgevNCalygjTGae3hZJx8w0sQ6fDiymQJXvf9kW9DUQiEo8yYT
vdxCAUxC5E7qwqvSn/vLmmCco/xNbYZlpQknRJvoWEHasP1pWGeYR4Rar0gVhcuS
B8GSihs6x8048FiobgkqBMktji2gthSfespIG5BUJpqoE7LH7dRyrkxKSmtVCcBE
Hh4g1KOo7eWZUmpCqxfcnQDrvWf0DUMKX4/LPI5MhsNntv6fPuTWpN7A7huAOUgC
EIvVxhfKcp6jhDQJSwAGnfrvYpgTaF47UZd9imdTm9LqicbSlLRUZuOhuNvnWxTB
4I6oavfzJT46q8UyXQRfmFF1ySIDMZ81JTH/+BzTDDcELxwF0Jr8sJEh6PFiNW44
ek+dOmWKXwd3zSAMV8muiSY3UsxW3YpGCB0udOq2HD6XYDLe/lVN38TqcnJKul23
Mp4tsEAGVklPMqFCENP3t4n2oVlSGcygAm2KZLjDctZ6tEW5l0p73tHqO+xgcMQR
J4Vj2n+PzhzOMKjflb67kVSyiAUhqaFVnDyY3FMcx65QBl92Cx49FSl1sFBj2SNM
2rAxbkCvUhT/YpfrPxcd4mMXEDDfA73VOFDa4+27MwGGUtkuaW/KsVKd/Kzw8284
4/ezaRSH5ERhztGEHFJWMZHOjQe47Z9EyYboQIjqqz1Zr5I2Wud/xKvN/bOD30WZ
CByOpW4mg2NeO/I6pBmw1e34GweOOolfRQCPGlDqFNj/z6/rQY3mdjNU6AYybygK
i8RU/F99WsPcbTxFCJSdOO8+HCpv16VQv4fR/iAXwLE/5HxOg6FM9j1nKJ2ZQtnc
/qrYGkRsDRaG4i9a25dnWf+D/vUeuOHfzb2q2YYLfYzp+A0bVqpaREqEzTC4HN8K
6BbTOkvgEvzB+q7n2f4rxvzpPW2htRMo2rELczi5MztIjz+CVtT2T4nVOGPsXaiL
hGw+aAjoguxcFD7Wdorz9XtM0umvDlGIlLmkRiTJMGzT7jnSsOF0FSJU6pSy9XHJ
sHA6/WboPkTjbqvxgp/MCGjqCX1MlIlRGmceqFSUoxOMoqq3W7leAHBblJ8g13KF
fi7H7SlkE/BsuLjRyPhIRXdr36uUTv5o3PxCsXRfYp2o5EYmSrHqGzphzs3Imvlq
ZqV/GPBQmfk1u6mQuLsDOHMf4Wn5sixoUOsbrzou2SREIoGiewxAeliYrPXU2bGl
UabiSBxtPrkZolmvTjMNjpPu5ihLFTJe6tMOpvwtpbVWHGPfqlXL/MyQgCb/xX9+
3MMGsKQiPhLHMo6Yv6pc4/VSQDkNSU4AOpEwE9Mr0EtKbknMmpJ9DAyxmmIByLB0
WhNzN48jLAIQc659sGQxmm3cFKgrb4ns+coFBS8cW885Eguq8dXX6TtInO2hHBqG
jRmNTBXgYx4jQP+R3DCJ+uTYTTSbWjSJfA8EZDTL8PkhHquixQmn88M3aqbvj7Gr
xGvv+2s0PPf3nKcUY9e+6QCOOdZTz+K+pBydsLGSGbdr7dIomsFs6/YTDnnZlA0G
`protect END_PROTECTED
