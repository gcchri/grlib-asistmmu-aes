`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kPyvc8KUw7RL4zDTPVX5CEZyq5bKHTwInbCKz13LnyPLfw7L3DDbQteEPIguuW/O
kENn1JWMnefnUQGjfIMnvq2n2hpbEG8Ggx5CqQjrDXD+oWlNU/P4QzK7131RSB9g
5qFGuSz0ztqRpYdBcz+5X+XPM2KMyJc0V5s7+WKYt0P9H7g5BuD3GMTrnq7A/yEX
KgApB6/kbw41aYCKBcsu4wCSBV6M60XjaDtvYCBWbVFvhiWvOT9Rwy2ZTvHy310w
oQRArJoXuK/I1Cf2HTG3NkTremJtILcJ2G/ovguoLFcR/j4KJqz8Y2BStmtr1xJs
LLiXZQRV3KZDT2d2xJ5FPUJGY77dyEcJeQomaSUKnKWFRYA22I0YEN8LyBKj2g+i
IFR+C5hN77vn8kDl+3v+MnR1bBdWquVjQhf3Fsxz2pVzNGBD1uHVvXj4VW/suylQ
u3Ucj8OTtK3n85j791k9zS2fCO4RxxJ6fFBhp15KxI9qgYdk4l/Rh6GRkdtJV+R0
Z4WzhZY1xDp2ir+ITiCMPw3hGMw1W0sTqsz0x70XB4lkoK9woTdNXp5MbaPtlsVL
lza6ce2g1SKO79wykmwA4CRjA2kkeT5NU/gGGRGQ7wWWtyP6UTvuqhdyUWwkD1th
2vfFTADwzo5ZVsv46GbNMSWPvIw/Ai6k/BmyRdEiwuf5TdWYRuK5vJ9Mt5a4WhjT
jncIVlD/gRUZW1eh9BheLOJ1724lUHA4wzTw7fr3449lJsPbAQRuNE0RHnBRxoZI
OXHGZnnbrEnxEzDthEHnCjYlfCJCxN18mjd0cdG37/kRar2B11td+5hCICjDLxC+
+/ONuPyFZQVryd4E2zhn8D7WFqhps0eNpBUS/zeUbcOnsJnD27IC8EviN4VpBpQc
wLaE3TX2kVZaSWjutS0lB2rUE6Uvyk17yrArygqCTHRm9riVkRd6w7UiLvZgD2Zq
X/JHyH2vApWm9mu9bRbNDRVJb9urRn34gr/y+Nry5llqQlUh0jgK9oV2pqUvmLIs
MiIgFQ3DUrWDDgR4uIA5hfCAW2oV6DQLlKr2gG1Td2CZGDtXS8Qg2KVGhmF8FaDw
PdnFNICamJFSHpoEJSLd5PqeP374TmeZH0izJlAAzEXP5Qer+9LkYqRL6GXxp79R
ONk9IRcMJgujWxJs5EjZ+rXCZ9k3njpQsBAUl8bFlFoDG04GUFsT957PmT7x3jDt
xdujTVybDOCp6XVYNEUHu6AUF+dd0n1pYuteJsRXnJG2jaw/sYqroMejMhxSsE1H
hjFvp3Y8T25H0v2JWs59woGEPmSqUl/HTGup8rc8loA1ftDNPmZSwZJS4KDqmxLK
j1DBgRGDY4vwDtXO/23eUBqnoX4p0CDudowFPMXG2gGSYmzvnDyuSVj6ZvoLhy1H
P+uKvW89QXtXWhThGAx1sQPfdhOHB1uaDO/PsscpDm2DiRp7atwMByWi7ZF3g3r5
dETPVmeklCndqKDTclw1tUfO0p01NA56z/ut05MZbwcPxAo2e+zxQimU88JmPzH4
fbjpeeir/IqzMRuU/vGkBdto0lMrl/g49AZQvehipc0fittpdS+HDWEM+bP1e6ln
+xQci3uBsK2p4hZZgFXI5nqxHjDwutv5pLDMc7S4hDN8s71rGiLaQ8wrbA+dFne3
6sZGbe1I7umlFKfCfZsITREX9BHsmVxr3+njBBbG1RQMFTa9w3VSboIsHXOXT9et
QHYlFVf1ErLuR+lrvHL9MEhkgBw997brGXX0kVl9ThXrXPf1b97n6tXxSinO0JnH
TbJ0fHzH5SgeeNh/x0zNdjs5hFjKBFP7LDGPJ25wzxMW69Anrr4e9aK0N4JgwMu3
1zqvVHONVNdhtCEhpghunzMa/xMrODzi0ZZDgtHKO6WbGMs2rCgiUqwgznGnK6z1
9EJ3LI+b7NfN9Oti/z7yPDXxfY5zoDp9yZ6fFXU5glYTaIRr6o8G3mmTSAutlh5X
HTzkRkuF7FFzoLRq6c+RlELgs2izdW++AY8V5q28Iqb0frFQGhrHIbp4qP1Phts3
MnVfYEX8yyEiBNi9ckAXIP/3r8pp7EYHVNd33rxyXcf3dnoe5wwt6WwUpezW9SW2
JFu2sDYD7iKOdhRGXi2HYMmfH+eylEuMg+go7Ep83+ZxF6suVozepsd3cjTXGhdX
xRgoU6UjxUIJIx2zRzow3YlVX+BqSINSYnc8HyrKAAP5M2TCaV9lIO8pjoaX8jn6
5OS4YLJ13D++Zej8MfkDCmbNhUWwBfY9hzyrZix4+e7XbzaAwhRZdmJdpy51Sue6
nH86HZ0Bz5wSRb30Jz2X0PSraMxOULYwCp45A4PEfR0ZoeQonp4ql4tdEJ6WbvT2
fNvjPJdF/jtIzChGKWc/AxLBRJgDVVg37alPyqFVNXkbFCEyHUPt/czbAZdrNqsU
aZhQ+kSoxe25BijQQqyoSvP3/pbW9GCzquyStSlyAVFgugQSxfSY/0JsHUU5a7+N
N/h0EHdf5znfFpmZf3IljH79/i063TXW5s3+BQAmNTrUqywcgN6B0Rw8eNPJa5x8
Al3lMy5aNryKOX1SwsJk0a9Cm9Nl1bWPprn9GtVAnKE1LfzjakhBe5MnqB5Co+l1
DKOzlLztBKr1hZdukBwc9fJ9YExSNYryWua3A91GPy5YE6NLUfKPvD21B9ocJk2v
ZqvoVSl1Tn1aqrENlrs/M/d7YjmBNygJWmtRxf8xi2Pi1JGpLMpZT6OfyjY5Zj/B
dt++QW4oMiWNY3h7vUX4DGeYos4BeRl9sItR6NNMr2p6ksZ7ZCy0dxeTpeujO/eh
ahcrBB3rGtdJESaJ7TnJ5rtqHL3DxFRE+AxTys15/+zd1JsYJO2mmbZRFTyCQmyx
UrppBcQy3cYlrdwOc92olMmTzQyxEiPUkfjOhja+Vp9Bhbaqd6nqoloaiq5fEv1d
sQiB0WBgcVqUNCH15illO9nNGt8+zPVdDgrQ3UAONbt5cQDtj0HIhMhKxviO1+fy
hkVOUkZrZCQ8AImjlS8C0RzakmMbZYW925dIUw+mDVgY7ezl/aqSklJlCzgSsxVQ
gdufXfcGmBv3zdIzS6+JA+f/CE5ceBa2nV0w9qzpTzsQGZWnfU/gk/Y5C4x8W0pD
dpd5XlSPJAu7SEllkexr4Z7MZnISbNzNxGjwONQzzlso/gUYQmGGo5+C29YD44ug
c4hwXQzfrEP3Xu/mu3ScT3uRgsIa+6hLyz4ftbi5upnDJE5H2obf8PCID5NzCG57
BufAL1BwNnxb28szTOKIQ8JgexH4cWKdTfej/kjNDd1oBvfwteg0AKGQBnlyumMm
liJMEk5NLn4x2JMt1a2NeA/lzhTDRuaLj9f2XsZQvpx9d+Y4QGjKtwSE14cNmo+k
HfEuypARKcXFgGxvkxmY2Z7IA9glp29yO+dUYJGu2xVWTSoCZz7MB4HwRHabmBjs
RvXN5wq6oCKninfwp/9f+XBJkJ+5qyMrSDmqO760J2IckSfNA7WPl93AwKyQwP7F
WfFYPfRnIPyPN/AP8BrdtonLLHex9kARfo0/Gl0ub6Zbjphl8LWOoygDJOKspnC0
WmI63xrPl8YFQz6iGzDKH2kTp4OROcSXecJ3bHb4H+07Rt6c+BfdUx7YixbSKQ+r
8xFWkS3H5KGXipiWCs9PT1LCwWzsNOU19VhvYRQAWCJ4dg4bfxsjFMJItz+cNBqD
FpibX6NkAZDlU3P6jBIqLLPe84nQRyIKKHB9kUO/C+HaHjivI/mB6bxai6riCP15
mYnV9n4SovCXEgAXGdTNLlaCwi9+5GWz+1kFMv21aYPlI84QdbPH5uOmAuXj2wrE
mN5Defpd4wgeyCOYo0+u5VMF1oWPQk6o67I+2dmgyyBAi1uW/4gZtR+GtVrKHiWo
/HbXggyWpQyQdIKPJHKWnfTBTJd3h94537iEsNcx67vTR6XnIC8u1uaxLChUJGWi
wYjnJ0r+V0lecJWy3SJgbGkxUfMxFTRmDlBjlxQkfFUPPzytoqZez4XS8CgOQ/cD
ZkKJ+dcWT7PTSJZ2YMGgNPzROZGTo3NDFoTEdSjXlcBOf2cNDImjicOAKSuS/G6o
XWyIU1QYBkK164D/wKxRVBUIbVAgbKcA2J7Lkq2dqS+z18o+/p6yDmBNJ6qFvUvB
UqXVW30tg/nxHNCHDo7G0QHEPGKfF9Pr2FQ5yj/jY1eIrsmRfzbKCjcGTBSDHNyS
weiYIp9648JJthUZPBS2VU0bciFuvQGFJqjzsK9zascttySG6tzeYQ3WswZxkDf/
wLf1dvlmQjwcgpYQpZVUHE/Dbt99pVxFE4PZbDQKQUHlJ5QD+yIB6ftBIAD9qN0i
17kJabGLIBxl2K+n4XWj0kcDoxuNutzdQtXAEDXBwnVscFTOqdQVupV7Mze3+BNt
Ds7RvJNgXJpgwYLhwk81Zt2qdPpzjbH6HTNQJF6CVDtHKlUWB092v47AnNtg/bR+
4P2o49KDZDv4TRUl/OCo/XLE1JOnTx2OWE+IKpUH+WOyOa1TwF+TDScLUX5pUoFk
KUHaJbpFncC6TgJSWzMpFy+HaAwoW+t8p7M6L5nxgBphvdD9TKnkm7A9mFEUspNq
mZ8mKCRBBcd0MjUB55CLgXOwNrCnGTPoPSLxjnWsRP/wvVQqvQhAqS+Vjf5Jg88h
AMdCtlLRleWCeXwcopo1fZ+ciyCMyOeYNP2eQEaUFgYySALLhJnRyfWKY5LHFPdh
C9oC+DL1JwsOSH4sjmD+koexjIj93TmAfx6ibhMpDDezpIoa/LJuemtC6yLWrmMm
gwUM3RSdBh8/HK1faz5L5QitYhA1hDfo5EVAZ38km1a8rkJjCMkkY4u1/RnqVJ1f
4LWQoNblFH02ML+tSHOFHckbq6WuazKlOvg/li2b9sDaystMWc2SJHiGpjqdqjq7
cnPUa9SSF7Akw4eUBsvxb4hMTsF1tgAV11ncu+MlVxcKaQJrWJUST7t3waGeiftN
7Wx3BAaoEnu6pyOm+ASJTsawye6AXXp9tYrYD0i2CKLh12EGMKo+sFZ4tUjuXKTz
hXNFqBFbRNmIMwRCuFtS0qJ+59Mwozy8/nAHCrMR2ueHy4lN0dG+nvVQORhGucQN
Yv14oJ0IVXDwV6pnd5jBjS7lx1UTrTBcAjNHlhQx0/7vPI9yFU1P8teYNjGw8+L0
mTS1KAl79wP//+qFr8BK6vEbei++dFew38HxZ3RlJM/hNLnJdF//sTT0rQwPLuM7
Id/z571mohoDMkiNVT0KXe6NTQnHmopv794rjbULwVra2z9KxDScQJ7OuRFzWtKP
YSf5oBSGobbClk/Hpnl1Rd5Jdv+Rhb79KgKUyhKN2P1qNuvOyescYSmFPorP5EYV
huYYWEFKu7NJDReQInG2lHVw1RNpbOiNLz5YXbuvcowzCH8qjE9fNgATGtMO/72T
owu7lvyDx6LL3fdrV2I4TCwdSx8omXD8Yyd+qOoYfGEirNIQH4eH1lfNKiFuCNZU
omTWBL+yr/7Qpb1BF5y188Htkr7v+LfTkYpNjbc1lYn/R04AjSW+vSoeUsDtvA/Y
WfGp1Z3YDDdyGVXTvSyrsl28qfYY+AIdcSlKi8rKiRx8DUXcn3cCsNVxsg3jK9zY
Q3RxLvrARZQ+SN9ARHhpQYyQCWNVDLHRmg/LVSKLRRrU2VWCHvqjcu0paAkEv3p2
4HyrdkeirVYp3iMr6gUjjGpju1qriFU1O6M8jro0hUINz+a7m9sZDn1jiiAT11ra
aKZuZ5QBFqJ0IaoATcFh3exSf19Wv55LQzIeoS2/EuCZoBCk0PmK5DKB1S9YAE4n
xwV//DolsuefUzXQgBhpIQ8cscFaLNQ+SZogzt9qFgm2ZTyarsxgtItbDHPp6stI
4JS2+ClAs0Imf0GkFW+Bvz5N4/8fjqNFyBuhIJZErrmbcJfWiy8fTRlUt0BuoYXC
INU4YNyLHsqshjYz1oc9014k6GBqNVPLea/mn3ixVGhxrI3LBP7KLkmEsjQJlR0P
bQZAqIJ63FAUsKBmo5jofUWAWbN60Fvw3A1lYnYmwfHDQ1bo/xF80zHnJrPtd8sw
YjRYkgPvpm5EwyYwDd4Ghrsl8v2Giy5IhkzMXeE+sJMO83KmRvLqeB3IrBkot5Ob
HIHz+0Wmvfs/4BgiOIdkvPVYEZ8t2t/Wg9vUymMflNJo9k0P6EsN7EvTdPtU/kiA
gh5xo4mCKAXE4RsZeCCppojtWsL9exQWnIoeLLheW10Dgs3ZveoHDxAtBJUZj4gg
FQEtyn8X/TxghfPLJC2tnt8TKV0fbrr/XKig7dAzNfI=
`protect END_PROTECTED
