`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8J5y1zsHAWmCk07ITopgAWSyTX91ZZINwxXN527Q4jvQjjHxFqX9gl/Air9Ny/C4
lJhVsxEWOX6FyHMC/6gxXuXnPDuDch5tRmGyiHQ1NoLGmvMFCh0SWqaFOfGVMtIO
RLShO5q6KZ3PScoH8mYfNQ+FeZalOiQyEHUW+1btL/fueV4nQlpx2NoGzmWA/wt0
ECz/S2u0AOOOJkfwnn3+SUn9B4SpZIZCGI2BZes8vnCX5aWyawrxgBAFuHcEPsw2
BMjdZB9/mmXfcHqL67VakcUOb1v0K77Aw6zy1+2niYZEfu68qA4cqpQ/2hGe5Uai
SdRwBrjYVwNRd7fP0+4cRFv9mzniVN2d0kFxK7zpUvXTOQTmxIEnTSbF7JoK5+Bw
`protect END_PROTECTED
