`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
it2/nkgxFQ8V+Dl5JBoCwQjKlKeZ+AhxprSQik4L0WoHT6jgGAN0z6sK9Ewj/gS6
H0pHSFolCohuzNof9i18R73DahQvLAmg40yrNhp9PYNuX1D4YcfvtCzxzJRsSdo+
yMYSoXYXFrNaAcsT6F3Xa7jA2i6w4ymqAyByJUx6hbm+wAgyVxsbtiIhk8rVF/ST
ISszhpEJIg60l4bD3UBXolL5UxoWRxgoMA/ZPhmd3HKIIOVcTYkDXmPRUFQGqfe0
aoEwyfvgG9hGvUqblqjmb+w58jqDHoWJRy5XFwsdOp9//VdUn+mePGEvXCzo3Gmw
ItW2rCICzwJP9+5yveU0dZkB2sFUJQOcOfLbqY3HRmYCwHTevr3xh6TRI6YXp31b
URT4YuGRS+uKabbL3HpELGOw1956GfVee0MLXeDETui7+RLYXttXyJzWto29QvjW
XiohRPJB3bBXmNzVPoRzxnaYOknI5ZZG7/mgVIyD4aW2pIC+nKHKAswQ0aQ6WGMm
JbNCApBQvC+yCLPQHxuhlD9FK/DIeWvofQmRYjJ4UvCLFdZo244npMw5GDJ+hfiJ
2DOOkmgylvSLUm+79bqWAe7+k5iOpcdAeErFPEo/mDjx+wjZpdlac4JBaqn9S6jO
4228ShK9pVdnjfGkkrEoUXETgc1bND4PC4UKqsEXqKI=
`protect END_PROTECTED
