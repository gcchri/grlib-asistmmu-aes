`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ghliFY5Kjst8+NW3NzqrioFVAJqoBPD3C0EXDRf5GSTEuYcS5Jh72TNZR/Vsqkav
rYGxHpdprZjfCXs2G9+QhbjJh+FH/L4YycD+JRtvmzx199XmosjQbCtGXEd62eSd
9L6sosxrP2Cgn2tTDmVn2grORxRHuF0cOg8WFHRSDkD4yy4Wj6BArzu44Hxr32Oy
HMZFZex6VysncBHwsWgvZlQ0XL/O582VVYh5iSBAgbGX8dw4tXNmCXpU6oW2aUfi
9qc4I1D7dkDm1sh4NSGWJ6hUMa1h1Yjr54ULM5kfQPtpqINZwYcFsy60kp2rvRg8
O2K3YAsT6lX5m7UB75KERxPHKuG2poyDBLXjImg4Z8am8UYJNkyue8K9w1cWe4wj
ZWI3DOevBZiZ8zIDKJhqtg==
`protect END_PROTECTED
