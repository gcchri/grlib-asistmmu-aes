`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ydFOwU2D1dYMV65AonGFuHe7JKbU24q7c8c1ahnckkjjKkInFMcMA6aIodRbpYPI
UoSJf5XgJWJFdMbhMZ6JiAtO/RyKkYdERj/z/mSGdCIzBsE/33h7u+RbVdwBEUAm
N1goImPNdnfUMV5ryIh4RhPPEU9igZ4bWop6HnJBkpX50dA7TlIXsT+bUq1V2Srb
xGag83t+TKB1hGJWkvel8M4Tn/GwGIKSsVbXXZohzwJEPNCTlEWcQEftLBK3FICI
6D4wSy8/BAi1rW8QWNI18faEtSLt5wr3GgF6e8jKwyxFoTFo6WdX9DSuy/MIn0YQ
`protect END_PROTECTED
