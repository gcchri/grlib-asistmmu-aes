`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
edExK5l7Pj8b4GkrZa5ActeQ9lGgZYeY1sk0YKlASTf4ufYtu6p7AxgD+2+31GLb
rYCkj+2ZcsKBx/cSjTQiK+CL+06S9ThdOUGaToFlyBeRoT2b23h9x1mcRcA0iqj/
2SQs5kA6Ufef7ufIExTR4krXM1RJCFU2YZd16T3GeElGCpeKW5I4XppcUEswrmdw
B/vrOOuySnsdqGM8g5yOWHGdb7d77M/haMLZkHNhOjRHU7iMu+qcZDpXSWx29uCR
7lj+aq2/rLgt/JGbrR9qo21lLxBo8NlQniqc/FTJbC62lY2vscwRpuUFX5U41kaG
YoSH1EPQn1LAx0gBUdwDzzQdI6sBuk65J8hmDQpqg5KQ4XtbYNiU5W7hvWeVqXr7
0i0BbH7aSpML4ZsMEz7BKubIlYcQm7KBUesTIj1tVWaVAaXCphPN4h6romXhVW2R
EBP3Ce1wv7LAIzxZeBviWd16edf2QsnIVi0pT+W4Id54dO4+lCkLW1VLOWnZfOK3
g40Gn81qZxpwcRklnr3epdPUaFtKzTV3P+LtnrXlks80UwO/IAVIRqE0feCVE+xr
`protect END_PROTECTED
