`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QzxRplyLn4OF9Zn2TURm9UYHbZb2Y7Kc1H1sWjXFET3OOqAlvjwtDH/HWc3fqO3o
E3STONNr+EMvGhXlM3kAslrYmrzqHIzZj/yCBfsERPEtVlvhKyANO5hY3D5hipGq
UyjqlOIsK3SCDsaZuKPxOHaUEltuFU9qZgcSZ65835YUbkQjRiYZQnaKgpES4QIb
QjwvPNKEyeORoxOpWbrdcGYe9bINGuSakw3pDIbqIeRKAFY6EPRk3rcbboBuwVMt
l9TBeTJsgfVDeBdfTmmWmRYSb49IkzZsI/ySxOABX48q3Wk4k2eXvcXxZsl882EJ
2x2LX/P4qEWGpqGzAgzEqbtAGqE0IhJfag8XvtHbTgb9hZ97PgRSpNrFv4GHFOCv
Jd/njrmPW8SiZIPWNgVxpejn3uXnMSp9Kl4tidbthhOwK0gM0Ge6/bpqa4DLeBQc
AAJTisaiQ/ARWF5uEe3L71eZpMScMiwi8dfTNwGzJ+Inko37i1G2XyZwTkrT1TuL
MoqGJU0mVlc9a40vhAAMCHvt05xdsu1nENgAI8lmsfAd/JRFRXaGaX57GlTYq3w6
iJto40sDktG0kdv1koAUENgM+U9DU7dP7KHTYhKjuetWSoms0IRZa4Bjduz8yvhF
thHMo9KzyPzpMV3Xd36qd/9DZCuiho5r1iTEXqUIo0qMO3DQZUSIGJDM81Sbh/1K
I6SYNz7VlBh5iRoZi/wmrt1YCUQjfVlX32LEcbeyqog+9TYoFGv1FFxsVPMXwlCa
xkDY7BffpZI079AafGGXnZ0BpkU6IF++WWZQf7xaKlK34SnRL2SSZk6LZMSwqzqd
BXv5RxImKWPf4q/LdhuIZtxYlyriuUX1TuYflXn8P6i/GZmgdWk46tb9HT3+XFPr
QubK/kQbiIPnGfxQ34lQrmI0J9t6L4ifmBCVLfTj2sn/N3NVIktSiLdhCAC8T2Nz
4NVBoRZSvIJyrVZtDMPL0gyxWrvq6E/4uRVgwdcVRQKwCPDxXJNw1VbzpWtfr3n6
LQjyFlRWrjq8+n5tP5srNU+wDlOqalngLcd75Lei7+OqI2sK3Z++HgdL3JBbWeFD
PE4nSqkjZWfviZ/QweIdNJBAH/7zUiIqgIkS22baQD6YiEEEqRY/qfomhQgSBJ8A
Mt0bcGim78v6XYev94jnmGRK7oI3dBIaRuWhm6rYJ92pnv3m0PTtVlbH9k43jsB7
LGTh7uJMzC7VtNUpC6Fu0rORt3aO7+WRe4ejgGETUem1c2atxhRBgw6ws1TcJKcv
Hh/w7TvIr6xBdj/1tnVka64LcHK1JE52qnSheWXTROuxnFJ/Inm9ivvq5ZKxNupq
mlU67KaQ2TiaoGtdnyIM7Z5/clHbcM7RvILmBvf1xJoPHiUpoxNqDSiPvw7egwho
0zl6DhKjOZ+8FtGjVuUpU4ko4KYl/xDicUBin0VdG8KOK2e8WvSnxRY6BkwThaCm
cae/DMKLDWYlIlIqcx+ttgP+M9AUNAIcpMm/0RXjYJIfyNeSsjDM6Net1dVH1s2Z
tzqBErLcsFfzShfSxcFJgmZy4usMOXd2M0ybI8ivT1RokvoF6NZvRS8Z0RXBWIc9
PMdJRMMUHhRkdQ6pp9LlxtYBczoCBO32s/vX+7WhHeUoBzxLuRqIi9xxwQZvfIIj
s4RAQM7rigO/GfQBokB6jjtVnNrmHPPw8c3bcBIy8ywF7OO8KGy88WccTWWuyHE8
2VXyf50vdM0TAw2PdQfbpZjbUD8JPzpEfx4JfdwfuYYKgDyM/uVZJ5c0dHoZCz5d
S0HZHvdxLhsREiIDqP2JOEsYFcSH12/EP/r8ZEAEJzZO/a5OnuUtTQLOEwvbGYxX
iRFt1X+mVyPP6WdjnOO7HpqBauDihaKP2/4SoCekJyeJ9Fi+SsJFlCR3v42OFLBH
fjcDjgXtCEV2nMFWrHCO+9Vfzzz+yoGIl5HY9vRPbZx89SEsVHD2EDFYx7UP9xbT
vbLY93YRoje21XCanGuQIbHAK614JfWZNGCKcLX0No7O48veqoHWYkEdaGZcuRhM
uHdQphC6g1aeIUWKCa451dFg2gSNO1mdCb2kyV/sDvYdiC9pHZKLL+ePW8+UlC5m
8YLguaxhbs5a7JG94LeBBbKo8Pj2EIO08+h3T7P70hs0uQrA3Gb4+e2yHJHjETcp
3AQn8Aic3g7LdSzPWaqz+v/YJwQrLeybqEO3iKAeCnxGJ4YvuNHA8w/uUF70x6Ov
LRkRzIT2eulYH3+3F+Mrb/VBXhSRsHmX0XML2idz/+U6jzhkvjXLK130lqbrtnR2
IEmxEsBMWmqhBECVe/5WtNlnu+47b6h+dVih7bIGJY2x1M5x+k1mP8mbfvZX4ZM4
FMdsoT+20cPdFsKJd5xTbITTK8lDSdV/fDUD+5WlN2eMxsD5c13Kblw0dfSXUuLX
GzJ9lmZlDpgdWZUrz/Z+g0OnGS2+4SHn22ZlI81Hocve6mjK6y3LJy3JReO2uRDo
joCBwW7x0lNBH7mwXRFe6KGDSqQ2MFqO3eCoDEhH0gDr5PTMz0pi5NQISVMtoP3R
l9RDudz9RuT2iXSrAtYaPRJM3CHk44GQ3TF1l7onXNgODZlXSy9SdGMsZWVZDbpH
fzdrKRBAEChdErvpkndjgwcwGnwYg2D0iP77SwXX3rWZWZ7CjkimUHLyslkKhaMb
37bT2BfOFU3IZBDz+BJxIU0GMovYaNtYz/OnIi5Q1qkVfcX8AqXnlizuPynkJetw
oHo4GfmjoZc3dzHPRD+tpvOw+C3U3sOtGvT08wJVMBD4R1w6ZbvpQjCU39nka684
R0oM6q01oukP2pW+tPWyhH7WJEATNKQZYmilqsEWB52cu41tNDw+gDZBCY/8CXhk
5XQxFr/GtQ0406jNnhoWrL9lgnN8l/HI/0cCCemRwzeYKBkfFSYSnIcL3ugqEr0m
yBB8DS3Es+vNeRZTI8vQLAdsYdjLrYs5lxY5P7aUoofD+fuamdV/wQMFC3bROz/9
4RIpYsGeNI1HG0kefRkhRPEPQrLM0kx6EUZuF9OGjcEbvK0QbFawY+qlYA+cf/T7
S7LJB08hrm5l9vSIJKubdFsgsAK/BfT3ZpfcPoRvsWwO9k+mfzuzDff2oJ357v07
9XDkmmaKoPBwG/eJq7LYx+6zuyMT/HvX95DMWLZAudAd8as1yQsWZGfrFbe7K0jt
A+77715D8rCtsPSWuIEprD4bOgQhdYAwQrsitnsHUDcPNIicW1GmwzLzcDnc2hQm
VRok4TAWm6Jg0FnaYbWIViNcAGlSoOsI8sDuWruR3Ncz/Ao/9W/kzSY/kl+QLoAn
BdZALDWSr7qI4026dDBc4bfTQOCGJrVur/gean+K1p7Ts7CrtnvWjzkW6pu4F1OO
bbf4LijrSlt3b44lAitfCkS4czB+Cvg5LECQZ8wKlETZ0i42tSbuWlduZ7XCdYcz
WEnWZtH7v9fgaA6/gcr/0vNlO4/PXSOZNXMu0ZwZs/BP5Z/P1MPLM/KtCMpuEu3N
dbAbrNN7R7q/tDTUIiwj0iQkJpf9+nAcPs2ovx9T2hnfzHw8cn3u2oYFr0O62sYk
1t4GKe4D+jUOSkVdmneFtoCZXGx1o4X4GRlt2h/zhssXhWRG7rHbH9in02VXCUu0
GBI/xdmp/6BFlPA+fN2gbQKiM4wkGKQO6fCjHksjTO19nv0v08GipsY/IJ06oBuJ
u5FyTpeK3rxy41xJ7blKW/iN8X0B0uyRn1h3+S/IFVdUTz3fPVrNHoliD5ayu+0c
lfUUFNsoc+QXwi5DmeF4M2RAUJqJoh0VZO8GRu6cnIot+iP0L3L8C1d5Mwbvp9na
A/7L0mT+aCHxod2pLiR3sk5okkEM3gIwOpFg3NYC9iX+MzF85vpN/0wX901XWf2J
7PYzcW+uwFQlxgCEI6eNnxOEIcLeMYRk6V4cOcKl7BfTu1yuE12dDjtZRRlgsj4H
0mv9r2AQaGWqeiFuPdskuczE9PwhzFb+7RSD/1Iyew8XLq6qyC2FonwcF8G6hr3W
4jVDsQqoxvPam4rKj/mG9wCskS7pFK5i+fQKqpPB82hLPOrKVHzr7Sl7ZWgTLpd5
vhEd+dQUm5pJfQ0UM+5ZCpEULHjOgPqzXzqOtlwWoDEMW4Z50+9spzDkwrYirnf2
ux+zCg7U3bCeQzmwE30TY7NkI8+03R9B2F5DIbZMLI7EuSrKCrAjKSYsIBo8+yaf
j9BNj/mzKkW0pt3NRCPOWm4xI/wMHUTppMfB5SMBiDg3Rbf3vQ0f6j+HGAuEU9c9
SOmtJeI7QJ3yGkLIkJwoFNMUMelroZsmd4iE4wBG5eiHQoJXT2xwKNe7Y+5r4MyL
UMbymerWUus4WZ7Gw1lgOJbyrVTba5a8ZtlQGhdkDbZQxe1gEvYU4K9+pmgYQiop
zmFYlfIRTjrwHC+eBl2OQ287uSK1apqkmcHLAyJXFUnsksGn3ttno3UZojGMQg3h
bQn1lo3WizW9u/W0T05ew1/pBwKNrZjbDtkeLRe6bcH/a/GUwPa2Z+XaUN9AddkQ
/QBaLUWkL3WEoCUdMuxTvu1I6hWmZXuVQu2NDl58m4ZbuDyICZ4pHG0nIoMKeVs9
VU6OlZAmpEAgVnGWADqzzC7ONtrJ88CCxQM494fQLyYd2lqCEPvp3fK7UPXtRaid
Mk4sIzUQ4M/mW5sZJayMz051rrYegQ8fpm+u3ZN0roJIFYFUWm6RbueO35aGrort
VJJ52D4BcITWoMugQz8x4jPAfroYEViV9MS6xZHDDTVM8EgDFEF3naGCWH7VAOQI
3jo8avTAdTcazP19cQwKIhChn3Dam9X5C0l4/Y3QFE5xAcE/fJrdeX2Atona5ys9
l3u1JZWJsfFk/yBqB5zL0DYNjC8NF+7U+UFXAvYtzDobtL5TCpqHD3XYto/MSu5I
Tar1832Et/FNoVzaJxK9vhU7m3JSIaDljdBupWSZ8LmPz0pPheFo5qOaDgi0ij48
S0auIL4O4CIvfBHydHkqROPudrmy9w9Md4r5R1BPOeZUQ3yRzKFGcnIXZi5myCYb
64YJPY+CgEC1+a/r6tsMtaA/84Nj7daaF1cpv9MX8Vofx5V3LOpHhODMy5+1/NWu
VgPRxaAyF64ywhY2iFH4WkYU6dyFE3XGMsho4zPEoI+EpV7p+HhESo+/Trk3Bu/l
yhD4yURTaVPZs+WckCzQs22p2EmC4Tr0S4XVoDzNgPJYLhHjR5whlaJ+bz/NOqpP
lf/UfKO+QqXUNLFB97zlhtGEAlZJ8oFBggTkwEeYw+IRH3ihAYr4MPDo3Xwkeylz
eKuJMF+BanEO626DnsTQqH2Yi87XuC05Syxij+XuA+dP1ktFFoVjfSu3hpetIl/3
nGj+qzimSSWSTdkrrQHW0fnidD2D9fzKTD4NbHoilEHqSyM/1CwqGaIFqWZeauu6
Q+zhrENqGcIOB0OctmzGGtW1/dNiXINyn+QQuStI9oJgHQoyUJaioNxAFGQ8jY75
pwiAZ9siPrkDKaJQeydOoewlaqBJIesw4VK6LvjDCD+sHG6XV45CoKHzi94l0jaK
ZjK/bqgvVPEYSFjgdIU0zgkyGe3D6MNJfSuI9SuHIkyuBtRMJ1K+o8XMIQrbcXDO
t/Sg24Q7QD9XkZvU4Fzu12QGbIhbM9R1UtAzUsegnNsKsNNyiHqj6DTRuzBfKWke
fPeo5FhwpUKui/jdRsMtlD5VlLgDi5g3nkB/ebimq3wfJ2zjdaF1YwX47SzR1HkJ
dKXOhz49qCrEQMSaEJtAUMGk2Y0anihKRhE/8c89kAZjcsCVf5o0gVP0rNJqRhnB
ZTNF2sJjRMEbeHeU1b8EP287PFbdr8oBX+b/3ZBVP6JBPQkwS8Sjr6eF+owLvMcG
Q5BWwqjdy7yrM30IoiezVTw8bWkQxP45eb1kmwuBvU20opkePGzYd69exyE0/Bxl
TU2S/vwVBJZJHkp+bjtrzGDFxS5wyDZNkgQNzYcx+SFYUr7NCwhljMFS5u9F9qDL
b4v5ze9RU5Ubmt+o1GzZzt6atKCilOtw28GOVHrwpvXtnS+iBISO6PvnS6kw2Dss
bJTYKIqQ3c4FwbI5R0AxcgTX8P3WvGScsmEg1hRj7PWRYKxsA0+N6Y/d6U/PeUl+
TLtWsQBUoSREtjcCgdusf85keOy6CmAuDuadgPfzBFOpW/6tRc5Dec6KYj8R7suo
9I7gAIeCLWAzdwYkss120utj2ZegPKEUvYyhSDYikJCrZykUjHWfmvh6MIOMjq+h
t64F6tswE3jtE4tbDVA92WOsnKXaYQagcq7suI9XyF+QxVwFSfAvp1xJWJo3K2Tz
2S18W7ZV7tB37k7X1agsJgabW8+/PiEwVcKYiucmzH4YzhEsRt862DvhkkTTQdiP
oxVufXAmMqgF/Bc70UADRbpUJe4FCDga85qG7zo0OLILqckI5RFlJewaDy1lRxXD
p2YX5Jx0K1MIw7yYHW6JgapILK8e1GM3Gqhm9PFPhnrD9AQ/+v2N8S0NP/dy/7tZ
rzfBZEd6Tbbmx6LHqKAyEscXUbBj69w/PXBIG79Tr86HskvoqYA3KT3fpatWKCOm
xoIkAqHTnmRRQHBgJ5ktL7HwSqBhf9KxenRvmrqNb3ApqyreA4cCINCjzr6oo4pn
89tHqGZNoXISjlOeLnR4lBz1LHpy5AD9aemUY88RTNnQRsacEolRsOFbY4xgrYo8
I6J9sLcI48X92lTfTNVgq+31E6bhoIzY5xfRPvRwsuEtKOy7kIxIb2tSc7qLwiuh
dzpRjmS5ydJrTdkVUURQvqaux4sWJ/gCl4YdsA1bofJMPJtVUCqH8MD75oVZQTqr
XLfj1pA0vlWA8UqsPYmU5G+lsjaZhh7MEEeieWTnSmPpLXsRZ5ZBeOsn+u0RCZDI
c2lcIzydH/xLxTEbuhxZ3h/e3ZDw6hCvnnfOzogIUPVWLUj1aCuJ38Q7DhtLOaIX
kV6BOu4cyQTFrWzLTp1Cve7cFsbARoaalJqT4vIBo1vxjp80XNuIfGbqsYWPONpQ
bQRaQ737Jp6BQzu/m+fwkw9TIzPZ4jZe1XQ2fpQXe5yMbPi3Lldy5xfkwUEAYU6/
v81T/CRAXTu+3M4bZuAjaDmMpWAUP5rTTsb+m2xl0C4NPxAkknNzF9VVZLrThr/P
ZoBvBkSGOS79/q3GQupUJOImIOWIR6SXgaQ16bn1hlZNAZxvyaUi/MuG4Ta8ipmr
5I9o6lxgQSRBwScZSOLjViPF4bI6QwnErh/Yy5tLoP57FOMguyC2z8nA3KUA6vIT
wmbTbGfXe2UXbckuq7Y5Tz5wnCNBwHutVdPs9v6+oO9zS1g2LnW6GgSVzgCO6HpQ
GPPv2piFl2BMUvO/2woVQPWsjVigNKXZ5fzz3BR+mlunDMq4CO2hPkhBrS+eliag
Vldf7qFFaoxLy9v3Z4dujSxuMDBW19iqOad9Ir0VR65mep6UTTzxGBy+TfTzlhYV
bHkI5fQcCNcJj+XRB1784eaAnYSsGrW+6zdytBijMcljGR3JtZ7tv2fRAts9fcjx
stHEMQBM+LymEd6JrYyAb0wggQff9WudvMrEa5rx0grcOHQlzVD7FA9KQo+T0JSf
x7emYOdzziXVPpw2ucp6xz9rCXUNlUwleyzBYzbfHOYM7mxeO99WfE01aqXWmM5+
nuQ8C+DQbYJSlXtd89cRr9CqAFXy2sOjdvOX++qA6/0PeU3nVR8EnOLFcBqh1z8X
kjKaNYkAkS4PhxqoUYVVf9tD6DryGXoT8mTMh8WrnAWgLh/sv7/P/MuJSxOlHGru
InfBWUox5Mkz4LKrNJbwTQUAcRbg1rZkTiXpCg1ltF3JAsoQ8NkW0Tf5M/DRHlwf
F31RSjmCrGhT1vb82cfRddZuN9HAntj3RTboz2E2fXeRBUUXaSJYaW9PXP1iEv/U
iH4Mb5ee2PL+2TwIakP6EQTrTWca1I3yn1e0dH+zJPD0GAg9hYHHIn3Wq3KGlah0
tCPAOEy/NG7viMhG/mo+kYEEDzUHiJBx6ZsAmXHR2H+IeONo5MyEZ+8XF4bx7/aY
ZF0sjVPMRET9FAsBGSgo/+LIVBl2o/UpHAxrNfoSaqA3N0Ie0LEvz4vIU6SvRk+R
nlhEbvL0GDv2mCH0znhuh5jqtPkFEfekrchFFOn5KCYMw3gbQt99DYKy60j89SQt
K7n1u3Kf0bMwtqrF8wg8it1Fb0AYYiK0R7P3XxXldvM2Ipx8oGwWxBU1xNGbIurY
nDVynn3EYk5rTYr2YjbEjTxpqLcvXR1+69VJHbiamlyPt5IT4W6wGa225qA1cIaV
bmSAeNeiFj6YYuR48jYAwhKPJHhHnkxhnNOl3touqY7W9CK67kFlEvhU7Khh2+5v
71v/X0H3+cnEq+Jc/vOo1/PrrdanpHtWtv6I3joCHYc85cdUhLkBOWEV7w1XdG4H
yAeTsUZkO1n5gMxSY/qxDd7p7EX7zvYGdwnmAIbFRoB18eX3MNRGipUojGXl+f86
0iLtWGYDZFXHuQKFKVh2yfF1Qtqlz6hdYIL7KYmfG4k0MGrHesr3dB+dfhFnLaZx
8Ou+mt4/3IIj1Pp8VRAVPpXIiqyVeyFrVp+WoAQyYl9sqF2XSjOvPQVS+lREanrD
xgWn6auYaID9lDBUzqhgSafKnEBWZPi09N4Mk7fUwyCnbQdUX44AZPHcYNE52jM5
wgdR7eEp/Dv3zEwO3rJD8JYpSZ4LCkB9LH0UK/Dh6iAP0tUs1ExBxyz/IBAru1C/
KswMrIoicN0+uuTtJp+cFyDu7wgHudwlxrvbjy/Z2aCBRJlcQb/VcEPitpMw2BHk
8eYlvKemA8EHM2iy26mJME4srvcWm1+dsvOqWnOAdq2fvwKvKjYHrRLqIxnvwpHT
eWl25S6J2M0bdav0VvffEIbEkLpWlL/trFNXLCcembSuuX05HJOjMddhjpIF6zW8
GKdrXvV/XXeUlbZsT9JddJK1Yy2F1ksTyuw5gAzacfEXYXGlRKE9xunKT3XuPDd4
M0d+eg+0VHRg4sObKjrrjrhyTjjfjzlglsi7j8KV2h7bk8xyPvG/4HLFKZ4dF1dF
YPVN/VRoA7hpusRtsF0IGvHcV+HwvV3OJbMJ3TwmfVaBl26IwSLOPY0m2SzSoZyG
yrpEJtjXYK5mWmorLDt+WVtERmx5iOcc3dwNKg7E5osjgVFZPPTp1m9K9Tk21iZg
waZqNQELrSj3SrcB/izYulKMGRMzKqGs8BdAFRSKYA0QypKqvpPX/tkhWkObQ0Fs
yU2dNpHzdOX5V6Qwx0g8UbDZdRyo0Wflkgsq3I9CRMfI5EC1+jpflOFPFh8XFpoR
NiFvid8FskjsHtGZGbhvNEpLJ+KIBWPg0V0OLxtQVRLpMHPdy9wWEXLabrkOImm/
1xPy/7iwyLFw/+2lq48q1j12tdJXsUHkKHsoJX9FNWMcekaaJo3Ure5fIZNhIYFV
Rj4pvdnKz4rj3vdamYnFc02UQSigSZGNrLtg0Klhk6oxalOA+qUgMPRRpSuZEki3
2MiXI8HqVivHKSeorSvIfyKe1x3Mi3ka2WjDP626vsRCJncmu2cnFt7TDUVvDq1B
UTDIKxJFV/ma6BeNdEL6yjbEHkjdmJYkdRSNXAB9GJEDNa4B+G/iiFHqk4ho2rW2
N5toegMBwwRGaHP2ewPKeZbUHXlh7+m/ZtL8ScfimjLcVQBoSvqMyuaz62ybA092
Yz1EdP9X067cR6yAE0d7QIvzxw6zzkmgs1Z1WAeoz6mu9zEmjieqOWI+rWVDSiNO
aFYz83nv0H2B0blVeJYcJo7/jQMo/nUC2tfff5Kymwrfv6RanvRGiWKExpcRZwFP
7wC8T9k43xc7Rvrpjodh5gL8SfLjk2u1+orTOLOspSSrxBupcyOXnt6+Jxw/Lr5p
ZsFFAZQTiiaVoKRJcHBIJf2VNiK65gzJE7nKK7TbeKdEI5nXywQlz1Xyh/eJIUBV
1wzi3kbswZJbxeXV8HQvw2UsTZUAgHpav11SYlN7XVtGdVr6pOGaBIVPpXxpGRWv
DA0IiHuMSabSffQUVsndbgo1w9U/pGwszC9Zy5/wwdj1ZgA2jtoRcfY0luzRGtYv
ayXbeVXsbPQ0qTse/jstOdvg6KphBqP21z23Hv+XIcvwk7/Dw4IHyMwbG6KJt7Mv
LinzmfCG9HcOTEnr7UXNZm4HQHYgMQ3N/GWn8WOCEQcV09j82ZFvdsGPbug06LRG
lGs0U7hn2QiGXCVQ4uotEHnL57cyjFw9PvjnusOS2iKCxa+aBoRKnqnlUFCONlpV
G47MnGNnPURwX+y5Rk+hFtmEM7Iy6i70e6Z8AzB+zBlfab9qJDYHW5F+eYCQsWvl
L7HyKsn7awToDLdGLU0XAQg/y+WXUd0XsLXkajHk5kigwfr6L0zNcffD4RyxOmC0
N2PWt1vSciATmo29dVuHtNzzcPvikqflFRAO1R7UP/bgQeNTVw4R1gTCHNyBRglC
0Jt6+a73Kn6mjTR28XzSKLL4ywQdEwddxzbUZabHdM64cXb7pFQMiCjUx01DMfUL
5GToI33ZvTkm6GCa2uFRGtIhaEqh3bpgIdWBX/x51WXP5B5ZzOKWff04ZCCwvCbh
HIl8QKF/L6VjitTuM1Zq4t6pOx2j8ec/ZlF3BR8mAeSOF9pux4tNXk/TyhVlu53c
PLhw2MbnczgtzN3Rvn3JchvpQY7hWGzw7xN7un7sm8LzAaG6Ac9T87YmCQZXjPGE
qFhYfRQELzmOSKlXnNLBW5rd5nMRYJxyN3xTTgSuJ9xHZMbMXqhBAU6Y+WpdyFqf
c5OGkactjQMMEH2K3LhxgjqyLsR9AUqsyKnuST/yV7V0iNKJlj32IJ0RWoALB+sc
h1BkJHEn8DxwBPJD/GkAiVdzCEpUmJV3PqZRz9iGnFMSrpk2jH0v5kM4586/zfWk
Or34Ax23WKLdrssuvvrdhYfjAy3Xa4SQUbXMfYt7r4RPD5UmzcGfaf5assShMi/M
y5H0HCYiNkS3/dcAnuOBzGvV6KydfKTpBqkiAw9O+Kr4frGo+xSKiHpBAbDfP4oK
OGege5ipvnWhfesRz0AdF+3jlwDlzUVpnG1WUnzKJnextYs2+SX4c4zJzTQs/9x+
lRUjf2/PIVzQIDqXbIAVNXB0kLBBd99BNf91+NnehSyQmdJn4Mru5D07jQu0uCTv
jhOpZ61tlbSParS8V8fuIi8xk9dCDBt4U7bRMCXwRMM9F3HghdpgxXJXkD9hBsYF
cSBpcRfaarF2pDoH3PknN/0xr6oO1q/9QP+FacwdqC0hFkGbIVlHq9Izg54YPt+e
lMDhKKfC/4Nap7+97D7lWdGhVjdQMK5MMVFGL4g8Ia3zN9EJpWVG4tjxTqd3ekD6
SG0DR7BOZWd/yeGywRDAnaghL1eqn2/eRk8XIBeSi0OFrDOcrPH43qnJIVG8qTHJ
6XtjKdHhuEde9ehS63uPtnY7wCOIieaQGFKD25qoIk1JQleb4dwoA8X4p83YKg92
oos1KI1JwCglqkU5PkEALQhl/jNyL/c45L4BBwCrChbwWPm3h2/27+Oecj++JRxN
5hNGSkvvSn/NDqeQEIOX7wHPV5hYvODhy21f+L9G6BlaSLZI5uWLqi78tj0V6k8B
+aizzbog1Yl00dvinUs3fXJEKlwTZnsshIPWhSpsf2qczt62GdXpZzhEZ08kG7xS
BB9BkDQp49GHj/QPxKiU1SwdrAPxbP0RGq1YYNAkRoLhumR+JPhNke3Rvbn99/hC
DCH7nXvtpl5/RkTfV/BMXX9pWzrzLA+GLFMZggLO05bQC/KYln/fmd3IGHPhomiM
/5QhM2FWxPQowHIr4vDjt1U+jJXZqlGnve44GmVQDt0SlibSN7HCcHKfqdvT+ktV
ol84lo9qSd9zZWlPT3sNJ6CKz1kIges9gx9UImljvh2mvykc7i/jJbvfTofGGAle
dy60r0tL/Jb3p/vUf3ggcDVOftg+ZGVAuWJXiMijYBgLN7HXqj9llgZtO0adOSvg
3EWzbdE3yH/P7yjeoJzXro6Ul0PDZiAerah+U2vVPmEpPbD/nd8iksylh1xgNcWZ
dIgOzHix/pnEu+lHnpm6vmcyukdL/JiCxpd5oQerSjneOCSnIbW4NO3pVOUK+7rA
ZkDXYJ+s8HYuVMwh3rjffLxukSplfjrU3xR75LuyG2RPbbfRjgGmgIPSdwIlrwdu
gFdqFmetWuPvNAMb4pQXa8GzeGgt0rOBAWA80TbB9rm5Upp1X1uiLJysWHpl+xHF
tvj/5jFTtvjbY928IcfbtJfxQB1cMYY5ZT07+ThWEVvW7AixhXafXz3hYv3llI4m
V+2dN+xP1aSNuU5y5XbVwtpIbgsr/1Z7MrkmDd/xXN/y5ZDO8xetKFTlVB9O9bS6
rlbnDKKRG/tRNnur1U4ZhX91iZmVKWTH1wto2wbyjm9+Q5Aw1U412xh/tKsn6XgT
PoLNfVEp7YhHDIUAEldlaNNZuGBC/9jhAEMjl1asoJL6qowXwkqXkmDvhn1wo0dt
mqO502lIgykFUCAlFhlinGvZzjMWZWCaiQGe0taIA0IIPPWLadKEqeo+vP3Num7M
yCw4b3tc3xhJp+plydrq8KzGiCvgZXLjMMQd0iC6rN2sGNfaO+xPWaSXC5T+1pU1
fkHByERix36LLtkSeG3opxWbrw73ad2eqlEEBix/9tKi4rrrs9qowI2hezSJTf9e
PPOOIPUj7Dt83VfaMNOZQQQQuUh6NzziIZjO/paXUmYUHM7oRLtmCp7bf/Upuw5r
HpBoEe7E1KtEyD1j3B03a7YaXW3fpYk8qytcwb+uI7zrHyvkOwndF8/7FGMteVbe
sFu5Tc/LWfONeRUBd2BIjk5dY7vuGWkPSc9gZZXq6nWvVORgCWELG/OLiHL9k0Tz
jttHyAuj1HYdm0uOkt21/Tt2gmEOCdm431J+6iXwx/fRGnLu6fdzBitqUYBPKnr/
udZ0C9W4DYk6hDwFFajIXb0nnXcirRru+MNMWPdXYdihNbzlRZ+rmRKOPeU7dirt
1dxSRM7BwvaC/Hd6nd+CIH1VNAvM927I0v4NMqiLAgWFBp8Eb1rOzJ1GVD5zxj+l
k0MaJkUNSDggc26G5AgwneBMdz3Tg4M8nGfnYt2ZUtw4rXRAGFkHpES2SzS5CScG
rwqD4mlodxp63wNeKQwEO1cT0gqO3RjqiBW+S3hS8ePXQOvgbJjAjChuI6//Abp8
2R2zyfdtBugbaqsC1edIIWOs5Ud9rWv3Vq3YId9nlDwPtSjIPHNdW9Nj3yIxhTdi
2I8R1ruXg+knU7Pbg58CQuv3N2SYBZOTU863wmPbbWoq1vudg4aXvvrm4B+Kv9qB
hXcCmgWy3aKtdvrP0WcKKkFfqveO8KnYr6Oe8LQdwW/eHSTlBtbGXYrzQ3pucZt9
1U+fIpRBRYs6621GbZPC2mWzLA+I9FNIYiUJJTcdX9OlWVjq57nhxcLX5BeZ0fXE
z3jRnRbR2Oau8TrLSZSiUw324byOu0hh5fGcVvDA/PTgfR1z5/rYBmAiVc8ZP1pR
c7/euTMg+Zwam5CXicwf98jBznaoCiXLb+/SyUA0WHpM43nDlsf+t/RG7Xk4gtgA
WJJG3Y+FaVGH+lSjj5l1wDOZE0PYfpGrwI19UcGdMsLc9dXJLsCJOWQyV76ycHmY
8O5A754Qb3g50vm5RKhJc44We5in+Y2lOvmwlhq67g/6R57zEzF+8iYtyDvMrL+b
4/m8VeetrtvKHF9RWn0XGnYiTeQZyOokxWZcaobYPRZ3tSK7k1SWNkCnbvCpsyiu
VcsE2GGD70TTLm4TQB+3vRHGBswguKw90RgiQTcUxy5mAUXVxZNAYw+JaePbU65k
bC2EJi18+zii3p5TiNGcbG6vizgE/qD3A3+XZkGCwHswD2t8AZ6VHPHKdKFWzQ+y
jvnY5E7yKE3C3RD3+8FFqP+Z3W77tga5Rbx5PYAySe4ABQF7BJTSJbp+jZgGZHFZ
5veQJq+ydrkPEN4/X3HngErSVE7W3F8t9j/zZaVItKuKzMVZ0zbw89OOeTJKU2mJ
MJRO9mASUjWPcBHF/10rUEHxRPjCq5y2B4fgkWqRsN33YkptHaVjGIkpKyTRcF1R
kuAIZjCaULlaAQ78IC4sX6cNM1wGRfVupMZCuojNcGKnn420USismWT+6t8ASlqt
w7jEk0iSHaYbEyu8F1G7THgPsWqmkmUQaBSaQ3E1FziX/r4sSm7Ra8DWdxZxDv2u
VB72Yc6oh4Tka+3rZHe2BYjneK3C0bnUPB9asw/k0LA8gQI2OjsuC3UP2syQo2W1
ON1gCaf2zblxzJAQdaFI9p18s2THctmxizXGskBY32rt8KLHUwZJiPKwTz2CRoT4
2cUaOdyYtdmQtGbREApLJq/iOfv/kzWk+hcRozsXPG95BFq3hEBn+ksDqQUyMVEZ
sBY+rohRIqgrHUL+yBgPaNOjsAjp836oJuC+xU/Ar3uynkM0FqhOaBdL/ZMZbTt8
GHsCzcj8bDlN4B01muQ9jSWBETZZN8BdDeP2/pav0YKdY9JzKIhSyaJ6VgsFH7S2
nd4MS5SiV2CFz6GtwOgGtKYxon0g7z8Kv/WMMcDJp/5tY4W0oPLWsvGsbc5scLX0
8/st24MOJLaJS65I3WEm7YIyPh3DweggEdCoFITw1IE54A3QSqPWHFocK50xjfUK
DQ7Zdn2jHFUZDIy9Vr4fKGIeUsqW9NFga3/4UhZInaANU0oJNw8B9CMf36OlMIq7
KX5O3g3l8Y0CvtalLli7VRTxk59LYZ3be1trTQbSzTPg791iMw84w+NDEaGSm24E
s553U5MbEUeWgI9eFeGP0186W2cSwMdMUAY0Pj0kOh26dVD4CGxdyK1WKo+Ic0DR
RWmzEL8+fNlcJcScmgFgxaPh0BOEo449zQZ8AsP3oaAyYuzmwe5ceQJSZmBuwWkc
1IJE/z6H8KKGNoE8jvtiCPCKQrByNStPlwYIqaToyoJgcE5a8Oo1EQO1BV9m0kzL
34XnS+7FaKsn97Wj+r2pOlp6y4EqCuqjVtxaOLIUvWDxskc4StQhR8Iy9+N5Rkt1
IET6EyscXaKb3Ung9oKlyt9hWGBg1Y7PpTo6heHqQG9XBpTb+oKN4ZaLawub07R+
ucHkd0qqIqOOvzK1HtGTTLEcrc8xQiXfkT8F04Wp+W92mme+ZidDcn0OQ46zrCHu
DnVBW+CFm494SiuBhZc3TkUQLZLHmJ8FcZ1b25CRQGubPy7hRbbobkNe8jw+129C
eo1Xu2aJlL9zDcC8Lxac0YD0HNp3oc7Sau+xAlcpwNtse3l+4fuflroI+XA59exX
Ag+0lyOsg0gQmv0uv0ueBZaIzhYhiouxsDiGPz4hm7raJIpxFSrGX3ir7Tr4FU+q
A63P5EkRQisWCjSiwsRa86BmVVMGw9sIjnROxrinYWqelajDGayHBfSIE+KluZAp
L4jBRqFbewxFLzaddIs4IdkDRbz/LC5Oi4+4AqxFGTMSjq0ihnwQkWQhBnejDg0N
EO6IttWvc5ue07HY9VTmyg6wOOBHY1SePZItg0KJ7evopgW8G0ZNzTXETpuD/4yu
uME7VrnEOI3elzHyOC2//jfYmSMcJyuyLXmh2lYHMm4YR0wndhuXBZiUsJgvAnSJ
zR+siBth9jj1kaT/hZGcv9ynVSq0VKAFq3fJOLN4Vv/sVMlQMTRbbnGU4cDqJOwc
tShUx6bO+G7cHzddtmhBQoxSut4lXIS7HPFtZtF35cCZeO63wWF0EeyR+K1S4/4Q
NNwA6WmMkEbeO7wTJ90bLgLUualC7POTsNVC6BNm/g6E9PRngnxeixlPSz+XSGY7
TJQVG8w9TXMPG6UpsdJxAmoOZkPO9a/Z6WkTnYsyVePM3EPQaE40t89AfAGCKQIS
KD4SH06qZPfOKe9WwmQ/lyxg2cEGVvcFppKrV78vHeOO+t9v7vgZJBB+y5SiW7dt
OXes0kPw2GzrdvfTUEOYVCtvAn5GsxPUxouyqJx/qXD2zlFX6iTuHTHZzNSGFpzj
qvJDJ/zCPLXnTcDYBTvzdkixmTs8QOFrAKJTqVtt1+/kmcx2qUJl/oolERt4QJBP
SDbmlSEW3PFKoo9qByuW7DKCfyE3FZ73Zswp/aAnCbKwPbpbOxqusN+ir8ni5+uL
Ram2LUNGZISCmdxOpc2wjWD3stZ1wO068k42tVe9bhAYdxUjBroN6yb4hWcLdHeE
tC/KvFzWr9l7Z7OTNRM3lNkceylRR2+ab6zznIkxOyS6ZIJQtZNEU+k5KWdq+Wj/
yHwWWvRQcn/fODi744aafH6n7KK3uo0/SzVzM07AK7oqLf4f8L8RMTZXdafWA/fj
cTURpYRqyd3E6YThnErdx3Dk65Io4t1SUqLe9je99cvxChuV/iqE/qyLOngqketY
J8ZxFU+Rgn5f1GY0UrkIY90hmnKwKZRTKmmb7KqQ6eYcFuFakIOZm6jGVG3tzGLV
A6D43W4+i05yldZwQqLT4TN4Px1VUWz7TGOvf76yajYsxxWDp6RSdiI4i9jeSsjU
8eNUfG+80HBxwdDrZ3JIIJ+4234aunkDqhM+vYNNBgAzPMKYngrVKxE2chtDA1vh
BwfGNyUsb6WRu9bW+gSrsf8pKXZ59Q+vvskTgqUFMHS3Xm4sQeD8wA5/tfbbjfJe
pYimViRXdml09cWtFm9B2XZhpd3g5MdTHDmNbV5F5IvvZ5heDGtAJzg7xfAVBAl9
xGOC1jRhNEjWua7XdlUrbP8vsdn7YzGH6eRp9kk0q9jBxA9htfOQcdo48eTn5ncv
qhXTklwXzgsUMddjo53Mqf4Auqo1cz5NPO7/FstAzmPWePDXxZo/caRr9L/m/X9A
xCizT29e/AJlyymq5N5eg+UKrQSVuy+CzI+Ke4tAvvQCI2ABTtQriidz/rHhPVs7
3zIydWu4jcE2zqT/vpBTSvK/Ma//+ljFyxBVlDpXddB8Xr3uhMTOVGBsRU5pzH12
7+uXxFCiA5Wx8dMUCwolAlDF4/ayt1X6BOfnYeP7GIUQLzWbK4rWZNBEHSHIS6KY
u9m9KG8dq9Ib5SEzLEQN5PEbjNKq+5C5ePaqcPesfJvCDcekfMKdLClSdgnZsBqb
HICGWJ12Ik4WFLMp9Aci4+QcjkQMXda+tKRUibUd7V6lkt0c7SWZFdQW0VsXgJ7H
WWhSD/OxHqtV/I5t+oVT5dnp8bjMnlFwpOStbbeOWa/qNDGplWSzjaXgQO7rrP8S
Bu6/AxUAPGavLhlorSNtgsN/R/Y4b6RTZiljE3bFfN1XB2xXnqwVWgd/cxNH4G7a
IHUwufMIt2pBlpKUYNUnG1mKkJHkG+CjD284zPBvCPZQi0h51YRKD783WmBpDD4o
eafkT8RAmysyzNWIKcsEbAx+YYzOecFLO2YZxIBdKjnzeFVI3l0gmWF2m6gw5ETE
/TmvsOSLPSQTj+74jTeNtUtkjj0+Ng+GiUoPh+U36MD0BEOrIN1ie5x2GQ6FvowL
52lMOxhWaPT+euXMBkrbeVBZPuYSnEN4BxOkKQt2Tu30q3Y6Fdei2J9S20rzGw0j
lNllw+JGIju+fmDneNKLiqs5noxbqlelmIKs4BvKmQedurVSwpLrueVhrX+NRXPG
CUjsfdDqAx0YjFyE8ITvD60MldFaElmxmcoSFXPAVvrQznNVAmqSYf59xS4rkEGC
elcrbZY1VOBdIl2owADERU3P69p98KEPloPnprh7GGGyMCoSklvzuGuT+HYvCif1
hu9b3Q8b0eYRBkuu3suzCxHBld3gz1OvDV+pyFdv6O002r67q8FRcJMh79drN4UP
ptrvXbu6OJGsUng1cDtdVw3ZXQfdp1dSfFP7nNy+9F6lrCnEGF9El+OR74kBEfw+
kDeT6LkZqWAbX6STnD9b33mYG37U03Kn4ZV4rrNPLWlCuWhAo/6fl15KJLUYTalC
bK7sv7KGEjs7jAwdKWfYVHT2u9xOpSQYZyBUzxIVSMvBllmsxJ7LyksGYlI8RHd4
l6+ZJikz+UGErkCtJEjTBNc9a2JX+07HPTrEgJ2Rdll78S5yZ2SWcCcWW4IKwWNL
dvHqVyHJEjxzekALeth6el7j9ll5BjEJ2sZ8YjL9Qs1ppGkxWOWIUqgGgVSndd+e
3YowNo5oPU4vMYeC9D6d53Ts8WPdDl6bwghmEE/t/pKThhvwsusqNSQT7aEUOL8a
lc/E/kbaTKJgnBAbqe9zwA==
`protect END_PROTECTED
