`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kFJxkAH5XqnD4mXEZuOwItj8Nz2Nj0RATY3lBFtz+DSD2XLRpK55od025HtAEj/D
F+O0zrpd6dA7G8g/SUWLk+K8ltQsgq+tFXRBa0DxgDz6ElupilTVZuk1FEPrWsA0
aACqxwQ0T4HcKSPHVdMi1kphn/m1we87xv+mvs3S7l/BpqAq0SeKubKPCvSab4Vr
Rs1RXCKiodOkeQ/gQ/wIg4qIp5OMNYIDmuvYqxpnGwHrcf9V/QUNzKgxKPPIHN/L
jLxyrpmPLtV/pRiI3vaJdta0i8ACpAGRwA4+dgiXTgRKnwonI+qxjzgCMzn332Gz
9ioIITU2Xg7AE9KKHPhre8Ld/exPPGHdbwq1usN0myd/USjPmda/XUFcggJce54Z
3ZF2enO67zxOzWXw7F8iufOwKe6ZsEFqE04521xRWokcezMh/TGGio1xruzW00Lj
quHKajIbB7EPcjWpOyqlnE6nZVZxCkgqYp5CqQOChC1XZJRTtVeZnC4bfi+1Ve7T
ayunEAj4ut/2FvKv46Qhty/mKqZ1Wpm+X4uc2gwoUSzO/uEOOJqAFegsZf6N/wiW
FpGdvNm2wZGR0wf1f1cXM2KenIKYP8ROYK9QC6MrbQfg4lk+xrphGr3/gJG2ZvvY
b4z9YJjSaz84SjEzblXR2vXdVLOdG6ZihHawPBGuI9sjHeahTj9xdWGWMP3bm90/
QRLAZDdiQHsQDpzccHBPf0gnbrEuh0oFz9Zkqx2sAOAYXFPR660vtDp9j6nP+G5v
IGrE+SmOSoFN7tmtOnHaTHrTtL5/HN26u69kfbNElZOLEBJ3PptMysUXCRB/9buT
MQRh4eVCJaopkSeiBnHafYiZ6TxPHNMEiUdSAxXGWWqsfJylSV9vyEGxTeE3/vUq
abF2bv2AQL1oIz1IjmNLeBKHOMRbZREXnLr5Wf6E/lybdGteJT1RdjHJqjInZa33
uTdXdx/1Q1xZbXI7kxMjfkGFEle+VEXBwTndcCOhbsU=
`protect END_PROTECTED
