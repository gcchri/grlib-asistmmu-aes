`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
14DA2qtW9Xciz6Dhc4q8r3HwJdKGp1OVS4qPxTE0Fh5c0Ys156G0DJ88Id23L+IV
DURBmcgODtvVSUpf3B/eV2FAJ6qF2mhRTCzKuc8tbwTi5yT4LbfXrZ0fk5D33vCM
SYsGIn64InmCffARUALcqp66/GkgVHyCcNysaCVvaQd14QMJKlqtaQ7iAcMFlwn1
Ca+F/zJWFx1+lFI+Ry+s7PtvzwSgVGHPh15KfWrJaKyZqkxw3oCk75DT0p+kPK1+
xWUaEyleYiE1NlqDiqxuMkhyrfTtkpirx2Cd7Fi9DWJd7lyukP4Gjq2GZGA3pWjA
xrYartajwTkeVVMo/XfuexGIHPXIzeHRzR6zfg30WWVpUFNbG/DJJNR1RPuQCSnW
jV/nTUoNDwz4teO6j0+QooQ9Y+rWXEi0e+/x0dNNAFE=
`protect END_PROTECTED
