`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sHkXtXNGvCx7PtyvtJC4lHLlmNRDJGJU3yiTRNKAc4gd/R7ES3NvhJMgzU8MW/MC
ft+Ssl8y86yZuSgzynebIVIXUgz1wH2lLjfmnY/E8m5ZJ0Nx0o5dOl1TeTIcEs3B
ls4qxyI9RY7LyVCQrq/VnqWV5E67BdHqAQCiVj0MtzJnvTDE60xTSH/gx9h9JrlZ
x7TezLnuRAXfLHEIhUUfq3d5IT2igd1/jLpaEoTJ2SUld+6DaIXSvbpVbgthH5K4
mVMQBuz/Jsfsg6mlcloz4WyQw/IO8I8sTgALfedfWQAYL9Zbq1b2G11N3XsnSmRT
ud3PUlWZ1It7aKm39PU/MsjLW6jJpaGt4izDS68KVuqUXNeSKLSAPk0BnApjrHW4
`protect END_PROTECTED
