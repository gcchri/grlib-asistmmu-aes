`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dNsgFMnWpBxeFJ7PJ5YUyVY6uPHAokAeSUTPs7++yRrqrORhzjvvqgMGs1p8bZxk
MoD/9cg4fHPM+i+j5K0hER3JD7mpxDQqDQ8FK7tbQjEHSp/TvWSnL8RlEjlJ/Rt4
tts1WXrH1FjjhIglcdjZpUudOwUx1o1d2TGlkliKHBu0XhIO6zwSfCfWiXOLRco0
u1lioRXj6dNl8U5Uj7NpEVElo/TD3odaVUjmSiqnGJrRanaDbnh2RDQydgQ+e9eB
L1JonAPDrRTELvxrjPO+OlaXPaPYCLGlOtdSguV06so7MM3Hv3bnUpHqMez8T1x1
6uRmO6734X8e3caUablUA1G/+ib9kjRFIQPBycq/2dW1zbxkK2rblNhiM+kgJ7Hh
`protect END_PROTECTED
