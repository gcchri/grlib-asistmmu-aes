`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C2Rlr4NJUtzo9Z3cUAWOkuJxanjjdRBzOcl0OJGzmMyvNOa+5ZKDOJhhAIvHxOfz
Q9v0eTkI0Bcd1ARW7TPOCgxFb4xi+l1BR5BdXAtW6ehdyuGTe7HzC1P5JCA3PT7k
H4PwWxk7Td/kTGWbaGvgpbpTAhlgYz4Oa+d2h/uZ1Pr0aDrUFhfrQvnRQSGShihN
o4hl6EapQep6oF0zCP+RPLdB0s2o+NzXr2yR42iBq0/gDh8Pz9CdDGZ6am451hYb
hF/qcN1CT+YQkd8eMMGXqg==
`protect END_PROTECTED
