`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/R8HAREWuwozMu2z8MC8FsMuSF/yANxiY66Xv+Ejy6tj6AxBme1qoQr5idS+60gv
NbFB6YsIKoQ/Vysvl5AesO7yFNC1o6sGcI7l4w5RxFRur+EwvlNYGw4V3TVgvyDl
mErwfoVF1WDkkNctxSRkKnUmtXVwv1Ni+sacFtqX/P+Xz2NVlYTjCM9seQKotZOP
rEVcS55sKIsZNxN3FAwy6g==
`protect END_PROTECTED
