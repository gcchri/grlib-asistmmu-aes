`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YHwjHZKke1V4ufheOgQGdhz8rZ8B5eoUnfQagyICt3NvYgh1svcB3K2fx3M39tRq
HaDJSxhUo92z5xnBzL1GFZ71u0Uk6Xo5tz9UAGvzxRb8AiGKEL7+MEGGuZIVK0yo
wj0E9KheJirk4E9gK4EYC0MtK8D48vhv6cpM2yNB1eklivs0p+TcG92MxKw+zet1
Sk+rndsFihVoxrligTcvyadbx5I0tBcBfyDCYL5U642blC0iMXXXE5NBSEL23SPM
WyS+TfVZekWsSVrldT/LulafIUDKwvDb3VNwHmADOICwcKEMmWQaP1DntrZZa/w2
Wg/5akiymXkGu3/3fi9sVa1IqWDnFHjrYLVGqsxg4MzDUiLNc9KuhrfA+xKKTFLP
1iyXtj/4PqfdEOa2ulqLwQ==
`protect END_PROTECTED
