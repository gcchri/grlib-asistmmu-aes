`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EkjITPkIt1JWyY4LXsAwQ7VARvmDMkQ7uPj/DfZ9tm9psj2oyQCBakoq1guWuenh
gD2ZX49sYibWGEWUXzwBqWn8X5CarKHkjuGsU22XabgJ5VZIef0XSxPzmZ02Wsu5
IK223i2b4SIHrL3+Inwia1JZEjLUn3OftmTOAf3uNT/ZxK8947VRqY52Kn+jssNx
e/KJSe3FjzpGGeH37kfazyibb3Uv+kpxYujaZCUdc4z1B9+EGzmbQ38l/hdzq2uU
g/29gkELuqJ9NbRO3B7Zyk82TjtXhLEiqjcySunHliE5g5GAw1jHWTlQ6pc42oCC
GXeH6IJyZ/lfEoOgFLI75XHA/nkMw/py7oeVZVanrVz5KAyAVKo8efwaQbhaSxOR
kuudPGkQRNzF3lJhr7MO1xJmOPpQtuYT1rL3O7c6N5U=
`protect END_PROTECTED
