`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fDsCgqles3Ef1UQLwnRChLdPFPZmyEDl2kIxL056t/v/hSxXkvbWtsDNlLJMpPwc
gG56F46EMLdBZhFAUho9f937uvmXPrRzz1l66GqPejdzdY3AsoKMdEH/A8ZrXlT/
Jy4tUqmReMyo+Vr9BVS1moaAfld4Y4apPWQWl8Yx2HlkvHjghSQ3/rrbheEeTXk5
inwU4QMn9SunYSYrLvAZLI+3U9c+1z5k2UNWhjIJ+v/WQ0xVZ5uHS94veSPxCZ9X
WgtkAMc5NK5DwQZ6Fnmt+Xl4+VEDbOLX/mApB9xQhQ/rX+TJrTvM2Y25qk3OU9Wl
wnH6jIacl/UwPsigjxJcdObEDsa62AWx20LziXkj2/HSudZCjpNaFewyIJtvuJ1w
UvFI8QcHt2NOGfYs++ni1IRTvrLG71OKaU10yQ9XwypuAtj79J4IG0Mbna78psSf
GVKjaEbdyKQlAx+vlq32JnFliQlhqUE68rWfiE/kjcmQfTg0CXYEt1G0x6akwwnm
bw1eAZEN6O2aPrcpv6wRK+y6lQxkki13KMHPzuDVI3SOT2voIP14Y6XVh1+KrnNr
vGsWH+WhxkoXwrX5oMIx1hleqRVdAz/dV29GmK3oVEReANwaKBCICvMtrvdrdahC
3NSkjjdGJe9hIBELgPtIabyk3s7NfR+Hf6GK3aAixwl9Aukpy0RyHL89PcUyR10d
FIEiKyTtIsVrnQT6FFPdJrDUL+EiQwdUqeLq8G3rqog=
`protect END_PROTECTED
