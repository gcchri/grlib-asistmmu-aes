`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pkSO2G2TC1XnUxhoRlxHQCJHPMHQxx6Fv4AZM53THBgcHKS6g73qlTKz+/Wfpi05
futsaoQJ5QGIomCSWL20etjAL2UB5WyCuWdMbiHecGRdsDC3zu2hPD/xr8FTqjLc
De1QOEbFwXiUzjm+XfuRsGtjjs5cWptT1xMQBlwO6Pa2ISzdjQaOSQEoLjHtb/uN
K+SPBnaxg4iEDiEBqveTd4B5i4ocA7iX4WEbG//WlZ4NmOumyEDEeiStKnnkx2w8
TXSyaLeTjg0J+RWVdANzConfXS/tnYVvwnSP84DhxZ3xS9zH6/zkOXnSyKpfGw4c
6vH72Wfbn3BHjo0go9KoCewGRpSqMcS6T7FtODocJBad89b0g/7p9LCkonH5ekEV
2/xdeTilKpG8TYeyvcwsEz3wya9qugeF7UuVPh0QBAwiY33gDMsaJQERWd31VjAy
lQzFeqNOVavFeuUdGT0k1jgzOn63F5O+jGk24JK/O6eKPIzOTrdQBeOEWbxzSt3V
cBJmScmpMaVaQ2ckhXOhekNLATL0bVcCU32RIyuxhKrPa49ckB7knHVcwopBL1q5
SklGkGFEjFGRpO+s3h8xQ7QYJ++B8AhU2wBgEKZUlPWCeukbT9GPCtWB5QJGCwXN
GP9dn+1z0HPrCNbchNj+Zw==
`protect END_PROTECTED
