`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P1MqUNnK3pFCNHeHt3Ryn3vd7om4V81J6vADp+78wYiN33xvyKgf2DaCmobyHKGu
cFCXE/iDSY440nU0rlz65vfzI2tb4w/C6kwC5sxQPhFbBalpKIZ0EsETEgveTp84
URbDExur8YfusO9R66E0In2hv7fiJWIY+mfx4KBYFfSRwaMbLEn6Ou7pTDLTlGag
IsQL0rZBIJP/xWqDwA/RINrtaUVGqV/Y+h9OWfdvlel8LVpDk+HJsxSRT43QQ+I5
Cg4I9lWaewX2Dsmuey2EmU/q0AWVM36Vde2cvWAY6vtxubymhrtYhx8PkVthNwaa
1RR27en5Lnd4mI7TKTZDANj9VmDdBK/pp22pZP+IGPIbP1BS14d76fEcStjomny4
3U2Wpksua0mJEIFr6DfmZesYDxU7MU6twvLA/aQEglphXuy08g8RnSbibWsBIxax
qk+ZjhR3WXKvOMRR8CHCKP3V/PK5FuFwsWsNR2mOdWPbAZhjSjmoP8kO8Y0EEcQR
`protect END_PROTECTED
