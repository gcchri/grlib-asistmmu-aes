`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vWSM4wtnzOh6MCZQ1VkPVgQrFe0gcTlNll6QnRbS9YlevUCVDRfGvbeMS5vE7G1f
H8JpXiEosp5ypjW0V9/WrbRWo13+TQow8Aycw/cIsVkL4tuYAP7CFd116WgMBX1B
q56dpXz0wiXMPCKMx+BEg1oNkwjrM3qmyd/SV/g/WbbqAIpKT5zuE4eHnkrwnTcl
xtBzpeszVuEQz6KeoDExC/Ch3agVMWutNB7od3KDDUWRoqLoTqU2qzTXiGdq6+Bx
vP8tYkSSHtp1kf1eDlSkxW6hEqsgQrjQIr4DFW7eCGPVqzlB/E0pZuhVw3XOMyKi
AEkEI0cBf8V52UjQO8hVbyKQVw/2F4nzxBAJT6m3/yLUQOlWENztoM64FMdnv3ne
cro0wpehYwXveDdCWHUf4orjL7/H39WTJBgb0RzAu3gSu9cF51sh4MZ34Nz6IgK5
/gTuUzHlUeMOLgqeWWdN5ZqU57fCNzqgtJ+8DQ60Uz7vFAbkajMPUpx6R1rxpe5K
CzsgD+YD54nFrlhwf716zuEbva9vfvqJcO7xpO6Oj1E=
`protect END_PROTECTED
