`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GKGUdb8KPiu7TItjI7/+hP7ERUjkalzZtDnAosUkEnUubK1jkGTYl+N5/e4smqxB
3+8f1F0LNxJ9iZZ94fbww4ScADzw6YetPGNc5iwR40YD7iP0RmVC3GuCB2BBwDbi
ed/a6Llr7zgoPxq51F+mRTF/78PkBjGVEfaHpzL6cQgMnmhMdEo+lHMg/2c/Ecw+
lFDMXheSp+TXqfICpns9nLhhtvfUmp9Fujax/qy+SpVjz3MBdlByNByGXSTySfzg
wgz2DU63J0fAa+2LcHo0C/NOKfw1djOmiNHyq/QXmDK0am4AuwngdZWpIcemfiPV
lp8ElKekPGPyXUEqVYWqZBM/D8w7+IfoEesnEgrGwQ62CMyMSbNVmpXhIxOQw3px
3s/S/OlJ1bHpm9rPggKxrvH7CYp19wYuXz5A1d7j28HqtModfDl0VFvhvukPUxQX
vh0p92iC0mdK36o8UAatdAFcKZv9A/3rSkDA6fh5MKEeQw9cKRbia/7Cndck4qAy
PmgqmTi/E4NDD8lzrmSlU1/KPMU/dgn4ezallUNE+/rJQYaBhQYUJbrBahDJAogm
7t9JO0Lvoc4p/EUHiZ4pACPMeMTXOerFvUuuG0IiDjM9a7F2w7qXXFVpU6auck2Q
AwtKVxVLA8Qw+Utj+0NELS1mcTdT79yKubvcvCg0iGJpKP6q+fgk/HaRzF1rfzDQ
Ec3MwNSS9PUOtUA6N6Dl8qGAFaFUHGysUIgrluGt3LoO8+2KS5CwsRKUw3a3TiDZ
QTR6S6y/qI5y1vaPLThDk0wApou01kwjRxl3UhUL2AoXA1v7d2FfEgRm3W4XUc8f
8fXheiI2GAaOXSuxgiTVZqR3FNqVOe4I99vSbyoOU0jNbs8KkC83w/S84da8yBjQ
6AbFbrEt6N2yCZGyu2ikFD7IACWBsRIBmfeja3WRQd+fwwiNxQvpYEfDyhe/FdrD
OKss+RJg6zH33+zey/rHAJK1UfmQqzMUEOZMnNNOz4761ZOu7SF838utuCFicPJ8
202bl7Rt7WNPzIMj6Bp3W1AFKOYA2c0ESSir8dYwOtpJYHC4rSc6MNlH8cQqz5Lb
YBcTzRcAybvdGrbHP3tdSikF+14EwYvD7HqZcuxLY4f91kYvHyXvU3Qy9seq0InV
vH64ZmfaYYpA3PVcMJAhqDeL4c5ozHUxMnp3vJjhBkRoPBDUIxHp+bkd/pG6BpBm
soXkhBKWvan45OL585//NAkiWyj7x8ns5RxkjNOujdIgRrVXfYPBJZ4qn0cFUey6
6c+ieDEfZN/oL5oaHDfThOrt9I7qUfmIQevy6lJPil1wz31ZdNzJS2vigH7uTdi4
794hcVARjv1CXZyfiBDLnU4TbSc27uUSSlXTEqd6h/QWN1echUwcrk0NS5fpvkNf
LGLgF86GcJQ3RDInO4nJzIT9tlGv/mBoz5npOEgua95StTfkbCaEPiPLwEuowcoq
`protect END_PROTECTED
