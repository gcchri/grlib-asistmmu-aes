`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
15soqA0MvnhOcuSf1uBPEeys4KSVIDNVbXLop1e8Z6PJk/Y7K/NCCQU1rr3YImxf
NdeXz1NJxoaCo2H0pl0dMUOhAzQt2WcCwU+4SPUjURClZF9BhEeht44/NWctjQNj
u4B8UQQE3sRQaZewdds6ku6gepASaHZG9Aee9VajswpBZCtWjBZ2DdoT9TXZl39h
NCtwAI7aB4GhaS3VpIwIOhHwKbywsLWCfijrUXcV1U8i1oaKOkvX79yrbThntap9
Tjb/iTJJEiFySNu3izvXWl+GUm3ivY+AoZ99fwGIWxGCxwCCRrcV/eHokhfkgYQH
xd3tkvwyVr9gOarL62VU61SRqAQtPwH9FsWbliL1uSFHdNSa8m1DZDEO+arhswxD
IuIEzGJZ7PkXCexDMk+a1T5kCcqH89DszAQTrjR62Ik6qmB9RE8NvuWXxQql218S
KE7URTDrPVIbgpjrnS9ixC1fDhVZ9DmbbMnuefRdAZvB62FDHIPdUNZKOnDeqWzu
9JO7tfvgxRFnF/B4AfqPeEHbuQbBWgTg9H/FXZNivcyErKirmu5YaLuxiCBduzhf
d4wkiNfjFC1MDV0xk+uu8QYhzWilZuARUYj6+6Tj5veLwUt3d/rQKsM7BGGFG8oa
A5oXRDmulvZ9WfJe3t9seZZxurO+KYme6su0CnSjGOsaN/JObcHweZM4Oq8tr1/4
w2t+CXQjI7iqJvN16S8VTJSnHEqp+e59XI5FwO85XB4lXboejt5/dhCOjQa8WzOY
aTkQ06k2Uw1IkySjRQxMwDOTG7bYIEnof4oHrf/vwkRRSf9rh8DNHO5MNmhoSlVU
jzs0dfXs4+icU1DymC9oNZfp+QnYbKi1xo71TO4mdcXs6dV8h3nTnuEOdZj5bhLe
ocuUXVgMCtQRgUj6W7EUyT9Z0FiXjLvQzfkxLC29FJVhC8IY5rhl9mlhkT0zCQJJ
hSSajPqJmL5L6qoLSWCMJ8nmuUH+5Y71dMl3ukf0+ydl0/VrZabEVIl5grvydHyh
Gmtn1Gh3fTKc0DNbDkM0WEk1wlHTYLLt2HWi44E89A5El8TFkHReVF6AE4xq3/Q3
tjM6Yx5UjCLDfpOYhI79gUqHqMeQq0Tti3uedE84n8Wal/fOUiykEwNjfLByoChl
jVMtcXVlhdyYwbNHz7Jxisx2VkjAJQ1DZXsCxfKUR5k8r8n9YEe6vx2pjVJYgPsL
hAicX/iUxXTUmklX+1+Jq2A8IRbSshl9SiASnkWUcXdMhkMFb+EuYKiYChGEQBau
YH03d1WKfLOAxMyOkW59t86DDY84gatnXI1KQEDZ3+VPnFcQAgGJvQALVwHj1lEy
LxxzhHI6qG9W59ujA3cNCbx6zE/gsBNFFQgXHmAP8bbNp63X1AufYaZCcZxxYr95
yZaHd7SBTMtHLBK3oPPqnV0Mi7o3O+kTQh+uEaEtSfRcDiRzpJb/EMs/qvrXP6vG
cUh2vaxiGR9jMk9PYPvF/r8XMB+e8nEr1nUE9Yxe6LpKjvkJeKG0k60Jr2i9gfk8
Cdy43JmpQL4olS44yPEa+NLgAGFWTMBbBykGzKZsDPxF0vCXRYCAH+8rpNZ2c3/E
xsZwlmH+fDkKprOzl5IzxXX3DtZ4BY8m/ynLvYninvDJviE7ImjvqZTPCQZ6mmgm
8QP4+c1dR0AbZH4UCocjz2sPD+PdIqSCdEkuGj6geACww1YEKzulTQSGDR29pXcv
8oHwyRkxImRHVC2puYs6tI/a1OmfGus7bzZLd2WPEP3n+uXfe4wqMtQaenTLsqj2
BfqkZkX1rZyf9sxNXht80XIBa/WQuIa6ylSv7NmZH6NWrqboztnDMrU6HkLjScS7
Cy3ajkWUMVu67pS9YcvOOqKUT/Gh41DAJuDyTZ7dc+Y33P9rwq/zfbFyqEtpwnKS
QOhJxOVy8GVMqGGAN22RKfa3EVvdqZ7RqfWzlxE89bpN7NHhzhkjpCmlsxEobzcw
Yjta36NB7TWNCsK0oIhPFFJI6HV7L/b57M7WuiEt+T3pT4JAaJJAytjASNVw5ut8
Rynh1X5+gpFXLE8kHtSeI0Ymv9IjfFTwZKUTy/jk3vMqXMdy6zlzxx8LFzQLptSt
pYIfiPhx57F9L78W/9gDPZxdi5RMdLFfBW6IKJRYRvHkYlFdUdaipeSQzUfUVBl3
7m3QnwzZenLD4Yt4uH7Grq67SueEAgk3y0AuYa8m6Y1SzKDyR7irkgDwZ3KS7wbW
ecxfYvNP8Ud1IaZopWWR/ICpfah7mnhwrKu8KsmVIayxbhsvgMMoY3DpoKtSiWul
69wd3cUuindsgvuGCWMRlpDk3KTeo0Pq6bmihnPuvryMD0VZRS9u4VNTCkeXX8eQ
2/KZo/oCHjDVMCNNAxa6UOItYTHEvdvpCXPZVQ/z9f11lszRfG7UROujQRAtGjyk
k2q65CO7f8NqiDSp3aB2T0qi2H6FE8umsymzszPwxqBwKW5P5omh3G3yEKiOaDco
hZ2zjZcstPTuALeFTBvw9ri35APn19RD2c8XP2hp4qtTmNlmZ2pRd382wH9knRgm
HbRPmDDq5xMMYP6VQTSD+5/I6FZGc0lbVSIDdaQjzbInQE8QnYyxEu/l+1pgqPED
ZNP2iRvxgtF0J09RgZ9/HuNXv9fdYwbfraUswdqXscIkGPvtLA9ds54O1Sf7kdHd
deKGzw0xxfO6TyH3tOPzsxDxe7qKJUSgKxziqJrHMGMyABQaGlN5bgxcMELwR4Us
/9IDXmVsxuzijtz2BA9sKD3j8QVV85b9PpAuxNw6bnp1s9m8PfF0wQExzOQpJXB7
a06O1kwuu0hQcYZm7t2RFakXexP0sDLYWup5y9UkN0W6uGApHRfPW17RcfqSj8BP
WBi7t59Q61SDkp+Q0Bu448+3CQdHIqUUewuNsYavMFs4OcsPNO/pnJYBWRJB5Qf6
l8P9IH0AiUM5bx6ix5ZISbwqHJEebZZi0DenM4esOLsj3K9HzaBGwTrSLtFjn6o/
X6IQ++OpjUf8cSJOw+Rx31HKH/GMtAR8uo+XpL0kIFHUd9vdCAVwv/ApzxVLsjXi
XYCvzd3OpMj24clRsZ4r28j0+J5oUR+j9Xe8EYLtFIhz5EYv+hm2yxgL899axCK4
91CKTEzlk0OihjMx92Yn2IpT07AFYKqfJJVXyHbX7qLZ9CZGWbxZZd+g5O+JFrBe
SxunT2wWo+NK2Oz3BBtsGZzkjYS5xD9KPbv5mr2pEVTi7We0Yw2KsfJifTcBizYv
Lwxani2kHDxKsaV6h8gV/XktWGgpVJdJE8H4NfQG2inW03akYxYr3b7wBtihOhKR
FUhgj4+SINFnYrB0gU9j5boPC/20M+q7dPhAkAatzJmiIQ03mRNo8K8PS0djPOhY
vq9UdhuJ6lvkwMd0A9b03JoIV9wZn11nduP7d1ecQoRQ67BCBPzqgAtH7gC1aBHI
KRZBKMA9gFRHHG0uEMuuacKREc2bEyAagy9KnxFFyDY9mHn9QnqDfJjXGBBLUnbS
V5ZQL9d7gRf1AeVWrC8ofGj8EUctFbdL/iNS1iiNCHKbHVMkUyJ/UESaPEfMh5EO
4xQl1IxQ1lOuu9lJfZw+K6uScEe+97h06LDCJcWoT9gIvoVQXclRa91eRkNIrG8e
Blgrbtytf+stBqDhTd5ZMwuc5xYBnbe85UmKCKQzFu+O935mTKHRu+gSvfWtUWLD
djl2wr+NkYHDNdnsAQyVLCP0NXH6MD1jiUgigDMQFY2FASeza26tXB2vg9XGzwqu
DHciTezxA/Djq0JR+zd5fynlciepkPfNQe2w3wWeXXqfIZSK3B1AI8lBJDMAULZL
ANnPN5sPQDyti+rj0/HylI9caPHCz+tAYiQ2CUnXjFC/BmQ7xp40XgudcP91lKON
+63Dy0QTyh3ZjJfhy0sV8L5yPyf3KgSQthJSO+X6RjOXNuLj50pfIhuWW23OLyy5
WCrJZ7rCH2dO4kxc4kih20shkKHmgFi2oE04K7STmfaS0DqNj/11cP/7mQ97kXn5
vQbr1z/LYJfLTIU7XuD2bkD6MoPydQ59YCL1i6fy5dbR2G01W3kVUqC4mKsMeu9g
l0vE+dC1sjp1PudZHDd73agROeW+w0UEEBehV3CP57lqClZCQqKZ4uTKpAilnZ5c
7jOBhAPXS3jZ4QBtf0n//bGOP/Um0jC7Wwg374Gwn72HxeL+FSoW3BVCgMc0Xc8R
0eTpNAQlYZChh7nsItfMqVks4eEvrZfi5Q0MhHSFPGVwVhz4j5mHhmw9Rltpgy0p
Fq7qOXf/gDCBhZEAC27lYtnknusM88pevrSjIGqTstZNMGV7Rp9lmoPhZfoUW/GX
+S5+SaZIIP0LHEqFRBaAGiQ+JxI9rcd+YpeMilTFSPGFY32BioP3FWY20vRfDx38
O8OcYbe7b13Hbyn09Z9eHoA/BRiXCZAdBFtZcKHWY7NMJw67PAp93SykTLAk5tQ9
GZGBydAM2OvlX3SIyo6OFFtrkqLKUxzZhZtaK2iH06AHKw0Gp7JCL6XKNFTSVYmb
CpYHLDclcH2q8nXP+bsFTEAnQXbBX0jIB+KLAAHWI1jjcsxwS+I7Mi/nZCj4ATCp
fgwjA0yNsIIGGRe2RiyRKrThOlsXIsVx1nuvCx4LNuXfiHRlqaq2GwMorxYmVcAu
OHqksFq7WTQxoBD4G+vmGDYfFRbv0SpWzFrK6OQoCISR8ePciP99bdfYiivSs69A
ySL1FY535bNcNc2KNZM4HS7kgN59Cp0O8hdSYGoiVg2H+x3QhRhN7tC8FmF9LyNu
AO/0WfEH36jMSjPHRPmwVp6MaNdfrZgzls1KUahRlDAGDtAOhwgKk+Rnc3dDt0qv
UODgGNnRVTUGQ4EXWvaMu9RihfzKKGnFRNvKz5BmcR4ratCQMkO/9PLaPAofSaEA
f/xwtkcOk1WEovmMObMxXTJJerHBx9wj9DEzsnBbTK9BgHLXHgpQvTNqUdlM+Bj1
2sw08hsTXolPGUJS63ttw1yVZ6LOIqBLT9Q0TMaq/VCno5J5UyzRIyFUMWHJQDCE
zJ40k3ZZ3CpnxYsLIb0QuJQl+CfVsT2uQmAC90nj5dPVOxwd6z87B/aX5U6NDfau
OE1o4Gqv8eeFPZVPaExdtNmhJC9G8ZevPMDFw1l8KalCc3fv5V5GH61ol3x4AzpD
ARjiSSYZZtxtBXG4MLzXq5N5U9z36idK8zCKjBh18mmUAjElMXI1zs4BQ4xV9Vz2
A5uoYv/NCFw1is5uHKWVOWanq4pHO1U/fLW9b8hCGUcQI2yJfLBNZ+LMsVINlIpY
M5aUb0Ahng0Gabq43fnp5x0QV7Hm5YUvV177v9h7sYgPatWYGJPZ7AblR4xSu71l
3P7TyJWUa6ss1Vkij5Du1+g2tDYPxbEKmvzGeFG+MmUK1wD3w87/jHAwhnvzIYOz
7M3l1f06c8hO68buawlAzydnjHGhAqmFYvCyydaqLwjNq+q1UOjnUlODppN0TKZ3
Pz8mTyAe9CejQkuLJWppAxMikU1dwAWHHpgfq38xre8gI/B/IOdOnEuaHxNI9Vto
vZ6k9pgTztY/dGIN4LGi1sUmMn+uB4vpef4/FJL+5sPxBX3vjMLVxcAj1auVJxhD
KJQasrdKzysdXw89i/g8h4cGHaKPa0i0y4I0OyBfG21hzEC0vswfDqBlLahUmJ9e
hllLcFwiqA9Po7If/irMXG2L+Fg0W4Du/xebE7PS/e8F8FDvpWWVHvkpeF/+qYPz
VgwYwu/76TL/7locaOJvA6UiPaypq3XrQaRP1/4FAM9Q8u5YWlQBCe8vwKVWXDF+
SWBvWX1jnmryewM9PUOWhU+RuwOhDJsRDhDEZVtHMvyoI8JrrKZBI5Cl4oL82nsY
lZu8Yf/dodLJ+JjPAYVFeLXzLd8YVT8+kFf5KlzNF99C+6XZ123dPzeIPzFKfOX6
QJu28yh21JRmxqdLGxUtpHI1/hQ9SC99lZYtgcEjE0buoDF3jjJCp0mkGQlMKw/y
KUvsrLzhk6aWxvEniL4VjLO6uwLgeTlU4vUjgtv+mLL4UbPQ/lgeXzbxAppyexHw
0XBnGG9Xv3rcaCpIg13frKthAQt+dMkLAKpGcZKRR9q7usWlPusFftcmOL0UZLLq
8iykj8ezHzI1hYGe8B2hZMKY+LsMNiTkjY/YBVEDICWk4drcgLIkUJg3+3uwETs9
gUVkMqyiX245vMmpv2902tCyZv3rFDObiiEyJI70V7Thw/nrKgbQ3ocaoAorv6tQ
bVvvaXvTli3b037zjJeYw4J++xDsPlKQPmvJ5X4zNs8=
`protect END_PROTECTED
