`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qxGm4h7UiNaOTTEstVFS2a586MT81Qpz2uHXFxHFsbiOT5j7Monib9j6scUvyfy4
x1IYydUpPni+biLW/0mdPECtMTymUq6wV7w+gk8ENvqrZU3wN+PQpgXKzorVbfhZ
W8nPRWnazVSfhJTLpOLbUjE6CAyz1/yHa4g5acPI5hjB8yFkkMYLjqu1qajPPGTw
1FTt6w4YjtR2vvGuJQydKHAcQKaNeNsWMslGv1qSlBtcistoeUA6oGdmvaO9OxT3
rONcVeSySxWrjah7GXGD69NQAUaDHG9nnbuzO2YPc6tD3Uo9WmFsuTEJoUi/LXUM
f7Dm3DdyIhU5S7MkZpe8iNfnIMBUq6rr3baNGqaNiE8buA6iLkSUQg3cP1b+9s8P
ZtCuZA2p3RzEsrUu+e3b9FRmBp7q5Kh6caZdnQV3RBukFXJAvvDk9YpDSH6y3wSO
ocSZ8UXtzdGYljYVybPKjOuOfNVz1QocwsMPS6xgXzQDqOK8ogfmp4K9MEf0THXe
I7/nbmYGt/sXQLqtw52lZU/Q3i/SFK/smsiLII+5d5lZ39EZch8zJShTKEvYB9cf
CKKMPvSL2+YmktLE6Ixqz0M+xQdgxc8iyEEI+afdQUXfEEnP76/YKKn0xzllvVZg
dUQRI7EdSlGUs00XYvQQLA+mxOtoyzYf8zYmmJYiY6mF0EnyOO9z8rRcRBPwLsDO
WinHR/i2mz02Z4rc0U9y22TrZZDx1s1dIeB3Lii3pQrU8cqyUjyStfqxllZOO7zt
DWrc6nUbA7UNbgY6B568tcUdIaAPEisjvItcX1NBiwU/4Dt9IZe7xKheEnouUd3W
D2I+jAgnoqZCzgwbfr+l/Wf4gK1xu8HUle1BNidNeJxsSttTWxY1uvXJHI0vl2Qn
+O4c/+kL6cncmHxmqijFrbx0p/KzC9nVGsyqeqzQP9vLJ/tSGGHzTqrSwfzb7Jxh
Y321tu6/rysuLer1Igl3KwIuLN+sgXk3NnQ949UVrj5n2tVIPL1LUj7sIBSpw5CM
MSjj+9VBGwsxToHMzfUiJF9Dd4alioeCf2N0aOs0/SIFwhxiO/MdgW0Am96EuUaa
LwnQqY2VhYwM2fls3YklQRap8sV5n6VfqrCP3TtGyxn66knQEDHaQaJJ7X7F/Fzb
`protect END_PROTECTED
