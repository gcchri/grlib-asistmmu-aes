`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D1dvFy3lu7WvEbvdve4ijr0DU8rBPKYD+GB+HjHHX0WkGsmvblk8e/ZWKu9qyY75
WbQ+ci/2wyTqrqyQfXuoDlK3YbSuyjesgRWBHuQwEEjneHVew0lUOz2s4Tb8qNqA
gG6snROBCoyCyf4VWMvkj2+WFZUEJhHL3aZTlLuXFOQJRqZNurxpHut2thwLE715
53He2sU1+YaTAm4wQ+aDWRwCqrONR+3e0eVaMet7U/OphlyMsKEP7fwDdoUlqLn6
ai772Hr3vrovrDK9ZypGomzxNLTNL0Q6hqyaTlpnSqf+2Ibp4HeK5JABiGm1w9TM
jTVwQKj3BYCnSiIIn9JrGVJCitj+EBuK0X6p9CXvAXEAlEIZwxGaVaTdsiV7mJa8
jZxCRXtwtXvY943bgiBiscenRHnjhREoYBKh7XfpAiLZcPt293+idp7PsZV42ZQC
IC3Qx7krWW+Ko1WFiBn6q9AJ2fdKxq0X3pYjcOVa7uZxtiVbc0Bww3pFToOHD8xl
CjN1yB3rf8brwdpXZUWrpg==
`protect END_PROTECTED
