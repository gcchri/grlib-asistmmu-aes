`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rT+DsTSaRqlK0Hc5CwzYnubhAVkG2ekekVQMMAB9u03DAd81cJNsmNcerbKdjGNr
2WV3u+a+PMyeBDLHCc560bbOYwniKF8xj+H463CQw6rr6YE2x4xpftMLsw72Ff+q
mwH8mGVgPS47T8mP9wPFZqimjYZ09uEUv1G9zTgxjh3BYdMgGpn9UD5hq53+b064
yuGylfkzH1M13Kq/pEbk9+y1vjKD0An6U5nVnDGR68eWr+RjpHXSO4UxIpFJY5dN
5ViXc7aFRPItX0pslGNPR++Wz6OAlUpHQUTB6YkmRgrs6XRgfmCBSnEv7ZN6biQn
+JRXaYFINW/slSEZRzsztY0mcafi6RrkotfwViuteRvdK2lVenp96f0yd8A7JSBY
qVkYvCh/h3Cz3Bw6xAmseA==
`protect END_PROTECTED
