`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B8acVQepC4vcqSBFtVsIUCVUk5kVGOkcf4zdfPnjKL/wNZULj0I29YRteL6tr7ip
DKP+twZRS3quLZEyQyDeHBCdvOrG4nK+feDDGfsDsUi4dmN9g34FSdz4CWGnkcVE
bR5yiW/r8rZ5g/yARZZHF7Z3YddPQTNdTbXUCIHeO++S7Q2hgDMJOgc6QNRUsQq2
vBRxBNgNNA7T5/YUKV/2CgX+bYv5DJRG2OMEPJ8XoiQA1tnySi2qXAcSMF7iRzXa
ecmX5yVO0vQcmYlBxqKwcLg8Kx+ofHhpEQB7iEQHfDMOg6Ud9Agg/bfScKuxJfH6
8nRS4rOcj9Jd8QlSc18u97lJBzu1l5npGd8mpzZ9u9F+dI9PnLq5jjqVBhsYZD0V
auv+QlAw3eZxntI6p8pexoPAcOCuuqnnaVQpxcWpGVpZLalcOXZUsO/hpS/7E4zm
ssi8V5DM6lkdnTueH7tzbUmerzFFsBG9frV2RqoCVpG8lz4aPUrKaGg9HJd1m8Zt
`protect END_PROTECTED
