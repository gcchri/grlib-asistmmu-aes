`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
juxdOzGyzG0MNO0PdTdaWFP3i9Hw/rjROEQM5kQVmJdkDtTpBIiaPdJKvu0Iaalz
WmcFh4srqWxfzjLCx4V3Gu6OOGuwPPuGDxZiV8fvC8AE3eEBF83GbyUjCcQa/fZE
WKa1nr0lppxsRNXFAARKhiPbsXpVzjnLi2ahmB6i+08Kjt3ODRXu4B/SmlXXBF9i
GSagy8F6BRTyrw0+3WBXYHeMV1O47XlQrnsM9Ww5eR5cilWNP9aj9KgHTEU2k5F1
fUNvhbv4jnD6zIGMdc6SEEcPFsVqSa3BaiST1g5nOUpNTjXDa3l/0yq6HPQuYkDv
ulsT2jt7rZqb7IZSbfa70DuHM+ksUTy2NiKdl7dd+93WH9KrE1ACyHpEQgPkzBig
GmI6HzvU7rXqilCkovfCEOb/mK+YIEzCjf+lxl96ANjgEUkIHhdnBcz9xxEFxfJ6
J/j4rhTRPFtuVNjPEnIKoMnxlFDzImsCVxNB0plPTohSPN/sg8U4gmMa9gmcZ/JG
M0Y+hZVGNRJsOZ30yUSxQmL/ZiEVGY0dzVORbQTdgQ7yoF5t/rUQ6GjA3NZKGFh2
YuneiA9edlQ8OWsIlP8WwbW9tvEZLefO/9a/xDzlB/hhDJiBKZNXmO+q3AZqlxAH
V3VMh33fau+1+g53+RSdVNW6TzNMSM9drE8WLDcSXO9w1U1jgQzfcrx2s1Rw3Uc/
GlKAy8bbn6ojHNWoW5kISzjx3yyEKRAelfaArVPfVZ2v1zK4NMXQgjxrliEAL5SD
z2htH5Okxu2CMRNxSFBpiC1M7YjkKRh0DdPnfzahsN3A8cZfEZSoeWufgDeQv9dd
E5wzz5E90VHy/pawlV0404u4skCU17jsN+QpfymtBuhvAetD40dQj+F0QN9i0J4C
ZdGF1rcne/HHAFtNIL8ScWrVQ1+OVnJxMDtAN20Z/L6VHngnWSupaH+FieUXoWda
XEqudUYRsdwzNz38tl/raFF3JmrqocPZsMl3QmfjX8t/0u77wQVXd3Mw3Czf1tKM
V8hGidK1eGR1qhvJCIDxUbapzCIf8G2Z41UUFw5sgiKrSal5VQbeCTQ+FLR67q8F
UhQV9i0ful0Bg+XZgmvLojtEaK1Npqj03xIx5rUVRfPRRSlImmwC4DJLkLKhYyz7
fLf9cVd9mZr2F5pVtfqdP+7RJA47NbAYmddAqHRIdosj7SVrnktXNE3rexru5Q8q
16YT6QAZCD58gZnYBpYqtoJmU7Y85OS9XFq5HsFLifLvv2Q1p++FcxN65c1E94yo
YJaCNgx/0aBD+SPyEJG7oHg06jnv5kKT80PSmeB+tNYKR7tdukfMYHK05f3f2jE4
TJQdLVg7uWNSWuJihWoxQBEpTL/uNJBRJbO1BJMaN60TFumOqiuIks1574zsvmKu
Vm1atS9bHvj7Wc7wUcBPBPVQmFHkP7KtVDaaUhiQuB+yAIgB7TmTjk0VjjqTmez/
WbCoYXvetgtITn2acNAt7bDVyW/EYtziUSabEGQNW5Tr2MdKcjycBOZxLfWAec/U
VYT/lhdzM0oubQQrRQQhKlxk2SYLsUgLZeiGdZ4u9T7NGM7GBXieUUHcvxJ6tcpb
f9XKZXFUj3twqliegwPH+EntFLfmzUTeBQg+G5Xrw9Pzbn5QE9cEcA6ZiwWMfvKa
yj8uyG1u9UFYtS9lwdjdrwwyzlH3ISS+PFTFDep0/R5i2JkCd24n8Fn+F+YrHLe/
cFhIBuklzcBk3Uq+yFjLmrHW3//8tnasH8sZuzrwJdyuq0gKsnJARxTBoxsxDrld
S/sKyQWxkYkpngckH3+qFNWPY17Bq0cRIG1LJ58lUlc82MN37hVlregSuNDoxvor
3ALelz+LgU66Qnlx1t7dDT+blVhQbBlR0z85AOb+gt1jO68UZfWq2UWgPQcTnR7E
1JSoCMEcLoWHOGKZARlmCN/CUZ90ry3Z7BlnVCWsCP6fxcroeoH8jaWDuYZSSfmL
sByk2QUla85pj1BYHIUT+qeij4OIojyo+KD8/+4LXtqRTVPdPiCY1TaMOshWuTI6
`protect END_PROTECTED
