`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rs5W044VMcxR0b3RGB9UuwMlhq2ywiOKa1cpHw4tWsRis+kFwfzXzolvRKZRzwJg
B8yBFFCbC8bC7PdnaZCVryULhTkE63keM8qOgmj/wh1osmI0Io79zl6xtS8/EMv+
9Jyd1amAckpRAFLSDIEVfaldF8an1EJ3aG+K1+q+YC4Te+MQq+jogHBy52nfBNr1
0s3whHX0Tdmw6g8rzEg1HxLfebl+MapwjUstDu0GR9hyGU/xvEiNAyYnTsFGKhUx
4om66VxBVGUtVFT+ahuZiTqY9IeNYd4LtKWoqi6xc9rVdNUOE9TSYrNTsWu0nSo8
/jessKO2v2LLnL2xe8U41CzwBcHS8lGxaaxwOVSEv5ac8C5pUUI2t9h6UW3G9OFj
8gPSjF8275f7o50j8J/KQ6kSDmimULhfs0croReURsUfZfSO0zExxlL1hp5mxMDl
XYfVM0cFDyCnhKrbU5TFWHi2egkZ3S2Df8uOHqL5taAa53Bx2BP5foxImJuQRiel
vrD2sM4wQrp0SU/cetUp03KbM7mORIjJEsXmf6+byCpLsTyQ853bZWH82hNaFjMe
LgNEto+FK3UpOr30Vp6+k2L8IqckcIf0W4PnzdX/s5qnn/hG1vYmzTUqRxVccDil
k6b/g7MRpf9VExwbzsXmnenyjgvXL9482sVQ6k/gzKs6GibTGUcxwAl6kKUvtAgB
1G3Hb6o7BQGMMomaVUc+RRPNoTeBNpWM9Ctmygg3Sz7UXk/11hkBWCmrsU1EWeQZ
KaMoNFgdoylx15d4YgHUUdExHSfNJo6fRIPOMVjyqsgSedLaO5iJTcKleeagUqVv
sv6hRzMXmSOPlTVBWiMhwnhZOwdveoAB7rBp1hZ814+gGPC60IHPVR+LxH69AeVa
5F4VJ84hiAK6j7vPX66huJaMLgJPIy8mHb3nJj2Asx89x+geuoistzZkBHX5zIlW
sXyV4724ulCAktqpBC+LJ7gtf0j+aVKs5tGwWIqbhfE2kYYdCtybZPJROx9YWUvO
Nms+roN8WWW94xHFU9HfhLkVoRbwZkc0po9NTkkHQg4=
`protect END_PROTECTED
