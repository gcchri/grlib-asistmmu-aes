`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IIHWFB4kOnXcTc6nw+UalfS2Cz0y02WShgTPb3/GKXPgp+heFR2HftqxCmD59CHc
CjEbIWbJ3vA4mcdlXx8G1S755H3zUNoIEdvmzH0tYqnmBbvAEula5sKChzFGZwei
6XmGt/onTkXkKr1J2j61AHHe1ZhpDQ19EDibwAcsZZ6aeDN7Uyao8jYVCC7JdMEm
d70/tEHzkPynPkbOblIAQR+kXcRm4sBmdIiDBSf54o2lXlkaRW4MfBhAmER2EUh+
iStsP7VXFtjkmpgsbSqyicZ0SumT/F6VmzYhAs4mBSpqs8+WLAyCgUXrYY0ETKz0
4XkXx0B1XxZCARUr4bSMdg1d96v1Ws46FY+1i6vR57CqZ+PilRFhtdL53vTEZqFj
0y6cMP1Z6In8QJG4XftLusDU1X/w98KeYtSjCkvvrbwmuomfgAGGEprt7QILzKKW
`protect END_PROTECTED
