`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ltH4TtVhgMOz3WnnOhCUpxb9N4U3T/37BnD+txOsVQEV7R1SMCzuh3hNgAAwJ+Zr
npF6ROFKQH99aPicyNVemmO0Ga4ehq8MYh4VyqNQIXd3UQvI0W+bdYKvbRBsLjTS
ugBH5JlKtyebrTSzD3uKM1tWZiuMyAY/FOlc171c0rdBTtyQLBudhLKOGpmiD5ez
2+rJkqCi4nSO3eF5AbWOWsWnmerMNhMf2WCtO3IexVkDgfDjAkhLcqzAgUuWImIg
VVpZn942DPTkZWxOI4sp2SRy8Gy7DoM8qTksuFODzBuC/d3N8y75/Avan1peDeIs
R8blP1QJ6hu4LJDdhd3FpjEZ1z26HGp5q3ArTMd/rmGZFMdENKNs2jsx1u1S1wQM
fqZQX5lqpGkWKpM9sCWXZ6cj6QPa9R2IRzjea4rnMGuP/Ln6BoNtoZfb6St8oUjY
Pv5i/YDSJD8M9oxrk309oeINttVHobVgas5xPA3VFLGosE3bSYeo26KGbmsn4AFx
Cxb+l8R+fMZeT0Z3Fz+22zRSMGlX7IBpGVpJAJxORrN0grhzKHye6xqGMetJ+ezW
kaw5D7O/E+6MYBWKiQk+4ZKc/JzRlUJFO5/s5Bm/LkceYsZdwVYzqsvy+bQ/PFoq
T0MSmNSq+3YOj3NsATbJ2PfL7k92PLpBgCIuySznIfZDjt/EbFvzYLia63zEI5X7
BoObH+eNi8oyoWeKXc8hqhhekAUfAWuxL613A/s9eeu657kQUfXx7aGNrGADgv+d
rL3FsgOzFGCx4hdqq/54Zb5ShnR5Gf+Q+7/lP6dItwfp5H94PbOuktEZ2YZhs7V2
CBI5ww8T9e+H+X0+U7lReMYam5eI318co1QWwV3AUmo6ByQ4ahPuwPvu0AwRIyy5
UOHESDvrSBMr13xP+fb75N0AMo6z3UMk5UunXhU70dgcb+i0TtQvAuPjiBR5Yfub
KbTt7BRmYnSQzz+H7QHM9DYKF1M+OuSTuD4CA3fJARjD/NVdwCjRB7Iw7/Fs1wMK
2QpFsLq4UJk6H2hl/DYNCb8snyaMFXYTSmwlBioysL8wdqBRLqL3dCQNq8KRR6WD
t5PLlureNT2lOJQXpoMsfD87vN0qFMawRxxlqktUi8qJ4YQn+RdelSHxVlrM5NRy
rOW4w6EP70Ppm5MKavLjvZZmMk0lk63LSdCI6ayR9fPV3Jl3TEUkC4CiohmNP1Wl
yil6GZClRwNs0dYwHty+5OC1axuzywQC/MozpkWQYFzYF/mPKABKsCqNUEF1O3Nu
bltQmmOSe+CGd6nv+NiDmKLYq+nKam9IXtmabht+Ddk13VodeGmBwsiB10mO8vp/
OUp5KqMFN5sQhTefwyM2o6q1Z0IzdxzCfb86t2Y38+adJssOa3prHjrjVCtYlaYL
r+rNclwoiMRqnptaKFspnliaNtkfwAlK4wB3ECs52tguHnBVO0IxFXArLeQuWid9
eSIAX4EZggT7hU8ZLd4Hjotf/6C1CautWDd89OfxcnqOF9mcqHGUSWMtq8nOWp4g
YHuvRgvwSXlvwutYTv9GRfpRhg2nRu5a6BNu/yBrfQ7ACEBH2lzUxi07Rt/EBRg3
MZnMSojGB7uVme1N2+8W0eZOytG6TMvcO/QoGpiLfdwIwfJN9t3y9Epsnei614NJ
kgctTvZFXj/CxF7H7YGZKxUNtYGCvFnWwOsqyg7WpBVKaj1KPaBesdCPyqfsRcof
WzHPPs8GsF2fIh7H4IEFXTWCxG8ORnsnUFKOaV3eEBA2RE57pNsGgj4Awldjh2Dm
Wz5IFA1nBdvW2SDVHxnV1YWak8olB2Wf712RwuHcY0Ex1CbrQ+c9JC2pBlYNUjiL
zWl7QUAX6V1SjBVG0sjNxgMB/NqTTcJyo2Nc9LoRqW+53fa+uSTgOVlHsfQn8WYN
9RyyJ+YiK7QKPCqLls1NQrDMYrY9uFg1Cs3Y2kpqpI2yR39TmB2+DQibhhwF/aCQ
3XPOtgy6Fa8i6w4WqK3KygqUTJr5Jx7INwP/gKvXOFGetMsIE3qthatpaJK71xy9
BaWKyEPvsUoq8GvkuX1il2DUpbz0UnNHvaBTkLeYRLZz7xQYYRLwiJ65QfxrlHum
isR05OpzEgRf/Lta+59W5i4hj5CZ7vrdSs7ob9x83o6w0yQOGcyH49rKDDiDnWZ4
Gseb7SVcHF+jLGGcFdbkpOUvjOdBn3Ig6ZMjq0lESOWzlFnFimpgm2S0N8UiKVWg
dlu9bPOCZ1K87c6RUXci5/HoeXicuu3gHw64C8lwsS4hPu2HCkTJlGxuakA33GwE
vL72E5WRo0/gArOhf4ZNKxucdsC4eTVZC+hOeUMKrIMguY7P6IwtyGCbaXcH0fwL
XxjjXyylhjZRXUPc9iwPWWR3O/d2GeVRd9Oepc6+OQftonMNCMlu4996gXB/BGUs
tlD3H5Ne4lCufVNgbf1/ve3K+dAkaeBhn4/2q05RdWh9NJRTA+WmCBl1HgwswxYX
rzLZ4WM38uTKqAOciJhpqay1ByglgGVQo0eeSDxd5ae8lusVjQCIj3er7FkOxRim
gAK5WpP7fsbrJmz/8ViaNWAunET5X69rML6/xLFeDCMmVXXSugvzftYFv/0BmzVx
abe9HKv0T+VwtbgF8S+FzjjA/+C+ULcc30I5N4soVf6YZ9ldjN9zY/scgr/M+uvR
4V6cpIuBHfyrXE7BE2QRdPOYHuDyASlJcEc/AiT97v6N9aFREwT6uEpQOCRH+5/c
fKJ/AxKgsjlCNsrrnMxoypCWQ7LaABYbawAxRXWWXj41xPgge+2XmQ0Y4Yio2hS1
omr4LsS41k2OwMu1WLPCyuq1h48b6SG6l8ISi3xtiExnIuw5Z7gg0jkV3kbmWhKE
9/w8Nhh5YGlf7HZINxla6DoUnp5btIktPqJCy6DCM0409cHMwpyBnuR0eRxL8DeN
cGqKuuRcsWiDNpoHN2HVjqyzEEUh0mjD3NAA2jaSPD3+k/0Geuuk7JXO4JoD/sQz
XYX/ZK5kAkAHVhfcHAypOeK1DNKkbEVYpH0d/koSzuka2teTNclUL8ZW40m1QJP9
sY7ip0eipSIHa8nXoMTtMoyuUcGdGBmQKv+pXP6R5R+pmPOboEBZiMsOqAuRAVhd
ipMl5MvI+snEDibTdtMnKs1xvyYyWCqqjs8KVzmIP2oCN4qgyeoyViT/HrcyLz0Q
iHzUAfIi9m63WysdptMsoVx4ivO7iFNTt29FNdwGn4mpOLUVJw9rBL++BXVxlvYu
18zxspjdoxQq67wGN9QBy7sxkQMf/C4EoKjo5J/Uj2KVHb82zB/YCq1BpPFRZWj6
CAWd6E6Hv1jShnaoikMMDqYz9eMyQYIkdNDhXEq/rt13xxHA8lvsOTr9NrPfB393
IKGbU0PsjG1YIYoQaDqjcABjAtjH52bKIyzWznA4yrjIkdf19sRxlx9iJLX7eueJ
AJHKF3DAkI8xVmW3jkFF963bSp6PoKzBuDIxi8JvHj365t3CRjmA9dcv9Az7NaBE
ZB3OYZPCQ28uBtbtkQ64BgGn03Z06RddUXwa+qdPCYh3oVuPS27kw9HrpOUbshJ2
LxXMDQ9Fzon38RyTEI6Tpjf8cmupB2PW1ZHRLCaPLScYxXnY21UyAW4rw4qbKCHJ
2jfSz+Le3CpyM1cYeuJwsWIF8Dj4NPPcT7M/D+ULbpf/8U9Xvu9FRyflOMi5aHfe
xP0dJwkxWHc6c1tgwtmvFNR6N08MaxApO3cumrppBcn8dIJmE2b6ytUHJcQdcVTb
ch7sxjVYfOu/wdKQEZAEs873OY69u1VcvxIXcIHqd/gFpd8USr+iqV8jJeBTH8bN
18A8XmVMiauF3axXdBWDZL/jYDBNRelt8sNQxADQ2/V6G4wCREXJ3LgmwfyCBTup
eBE0DGzEK6am8P+c25wFBGqqGC5vbPEONnxz3gGo14dcR15aNg0DHlJF5vc9CIIh
JsKLBLh7MEzWhVRDWVplrCygyguKUKZyPhVb4aQN/dzuOw3ymDZhsmY/s3uy3T1v
N3w0tTGYGKVZDGo+MYogFKe3DyxxKGvSJwvzYaTQjre2D2LxXkgc1znoBI9VRRgX
arhFBhjbKNOC8dvOeEvcD90TESvZf/lOHCjorQc6wrNHhBttsckxGCXqDp2usU+j
R/4LkQcmGmF2qX4xddyJdPgjKZOd5r63S5RtBFQCaAidz+TozFvHEDBKNiTg/uwY
sFr/cfxPfGH3vZHnbawremj20p16B+nXJZmUF/eJ2+poqEDbral4S/xFzIwZkac4
t1la1jQmHLtBPMWPt/fm16dMobtG0vtWwxwcjBq9Y7nsde+OicS7to0yhPvbCQUy
2oSEvWSG2yDABfig7MJZjiqAtPVWDnbWsV3aA60vYGuuQpOeiAyTafigRZU3d27k
/kqoZ53ns3svuoYk5ZoZPfa2Bks2VYHi0dO4iAL+g9JiHkcsGZyJQiWfveOKVKLI
X2o7NgoPO1kGPqRPoKBT80e/8LJQ66kIf62IPrPg8WRj0xFPcSXPpHH68dB0Fh/C
3NSOrIUUSSrszvBC9/AvUjmivy2AsbnFOEw1Gz5M91v9q7rquFDRPIPP7+uUgxuY
RyKkOTroNZoL/BzXvPlzQK/djtQHd4ztC4fBu/zr9LHp9XzV68VeE5tIJFCbFu5v
IE8YWwy0+YP+F6zOIVHvm4SqLWJavd41O0Cb70KPoiWeKlbySH9iFw/ZqQAWDtKW
MKn2Pjgqoy0g+CG4OGscRjkxEJz87m47ZJ7qcr5Doh2wm3x4pswTzdmKCmW2l2xR
mKgaA7g1SS4MlcLOPkWimN5b6e3YalAOn12YsAEU5H7hIWkGRigz7KJE21VkKVtg
+TlG7Icf4UvGiuMmowYvZIaPrHyZo7LwbhnhnxhDSg/LoWKJzBEcbiTkpU6k+mYR
ZVRAw+1O3KzPRtgvvRrhfMDCatdcGOzF6h5+sP2SW8/ZdCinh/StvlGC6VgMXcdZ
OHERL4Y+urQ33JOariEkArqlLouzSeHsLJuQG0rgEIqJliZo9Ir1rihvU03QSqVN
HxxsmDct0aJcqRPYy51EbO9axnozSyGYJhgNgSTfzTCk34d51wXygwkCZBKiXNPM
BqG9PMR5xysjTYA+1bw4LedX+qvFavvOhLII7bZqeCdQfZ6NVf1t+ff/6Dh01QAg
s0XnUOjZZFXsuVxKswPxGxZv2tasQNsKprt6b1+7KERBTGk7qXgyYQxXVKkh7G/i
NuDdW9sHSKnQsA7fJ9MjS/0T6A3DTSUV680vKPKSj0ZRR7Ue5B/wirkec1m8BSoI
ISu2KW3PWerL6g1RSPLEVI9AETgEUZie5dVRmFRfZud7Vmoa7dLWCvkWz+axRUo9
qgoXOgN1opyCYzSgHbJR8nQPjlIlfK7hBn2WPOb+7DeBnaZY3IbMpq5GNAkegmJ0
0GlHTmh8RqrKQIjfJDll3JQ0GGjWUkIxcvbKlvxoOUWgApKM4j2PZXAUVjExlx3a
NhHKXNn3WYDtcQretH8//Wsh1RgaU2pKX/biLeqGJ/vbc3rQzSQ7DLPWyBapCIfR
gdq+rDLcSEH6DRn33pNuH1JCAtOwtFo36trOtv4ZTsN5pSP3xa599kheL3psSyYw
tmhgosU9xyxmjAAwpvlFG528B93OLyZ1KIAaBfMbwW8jeSmvUNGMnK0Uxd9dHytC
2k/+DfxNouWnHhxVXAz5XVGFdqrke1p8Jhvj3wv73Is5eq/YKSmRXdbOK5x6nbRG
SHSST4kbAwe905gdTWH3DzQzEIYmxfWWi1/hM989ad0PROyzx7pJhaOd4Bo0+kOj
iv1/5E1xaxuSoTeAe37RtSVAqsZtl3SxKl9aemFbp9MQPNgGk3jPW6Vs3F7mZQuc
LCksyBrcbJpWtKY0cnP1q1SX6hZBfW3YFsYdGdr2nT7liMfMIgQSspcTwpRS14oI
lgUie7YRaOLlPnHJa8+bEv6boJ/DHqLmfI00RSSvanYAzvJPbyHg6cw+1OjuS99J
doBk9UM23mzzhcq95OzYgD8tEyubp4KHnN/JbVYKomIOi6w37ndgkHVMi7eVBuu8
LE2wERBbJ+MO3bJ/oJ0SelXh2DDv6bCeEEVyvYkLrJ76JAr5U46iyEhJZIgkwW+U
UVcpTxSn5oRmbakNI/CZdcGM9fDHBm76H5BSBA+yYui2+ExFBRwCNZ7SJ+ooCFvW
ZgQ2BRWgdrsvfFixoiQkUg62YemSCtWSymVeA1+FaGZHM/uLe9n9h3VdqFxgzxSJ
Xh5bnQSroz2voaskhAdpeAAyzOKPtyc7hwt4861opVfeIo4OoKl6+GkhaOyTzveH
vwpiDSHzYtGROhXtl87ya6VQv69J5pAJVqMtGDWXGaiBpapqPE280Hk6Y+GG+gIR
0fkM0s84lbH4XLXlsxM31veqUFrYfyGkLPj5LvpeqS81VmmZkheIVRzoHSQFRMOR
RvsJfLWTfeUFmSSQ3kb94AHYWelUbTTlvRsx34+GkMZL8YHWhyRPske4ofxhidrG
I3MGL1XM120DwoZF2up9OjsaKKQnu5aDr09bBgMDKW0aiv5O44ZydtkHBuAfgHlX
jcLewyl2+aNHEFW/qC82zb4/0ZZG0ihIszyQk47vAerUR6zYLcyGkUOkiTtJHxoT
vg3D4aHovIdEVv6ZNgHmeE+FaGRqqPlH8HVPdk02JYooawebz1iBJQZUjzevhG+f
hW5JRzxOr3exojPUTQnSxFhlxhHqZKTiyNnIFX44Q5NQkv2tYSlsUO0DK7sdykCM
imkSIVmKeJx9SJ+6SXfeCCg8XthIhwNVUBrDQ1toq9UhWfJyCrSYMDcK9iq+79dK
CIodKWqe1cMl8Typ6wek7CzQMoKWxgxkMOwuWYy0qjEC/vMrTnBOSH11TN61p6eX
t9UyuUwcDrvtDrTbfyOByjS/SPsCLBQ9dS48/bbEMqYafz1zHX9Ln8MEjBJQDdOr
kgUDwYtdDw3nc5Fd+7p0Ee0b9HpcvEKcP2ja4VlRdDWHIVyTekoWzPAlegQ6pxkS
Mq551wgoDc+/VdgoYwIp8xiTcmqN0NwHGzuK5qkArsT0wtXhgUvl/hqy8LIYkQnS
HBiZDgq/hQvG1ScJUPDtY6KVEuSG3YlO9Czv9yhVNwZeNeMlEzEbmcUaMsEJchE0
ZYpDLFUhhdjppcYoQ6FoHzRikn0HFQvjJ53McdgYtSuqDAvWXfZ52j9HzWzd+lFt
mIrPZJX7fFvSFk7xQg2SJ8EZoInubwiDEiARnFCeDpxcP4UQYYz+PiQGmpHUK2vG
LbWqi//8GNvzzCR+1kL8P1rjcjdQoF4gaxUcRfvIKyvioI1uDe1XyKVsgQ3yjOEj
Qo7rR1I4cem3dvUB+IdPvvWW9NLqGi+SJ8ubpUwcLZ47gEIfDeqZA3/FzZfF2Op+
rqpsPJy+6DKkNxyIoWumfj/q8jFpVBA7ULXwMOZb8xoX2+CNTL8aHpRHb8f82C09
Zh673cuvPf2I16mqWhBUKMDZFueXiJRNv8gyF89T+dkz5wfteEZA441QN4UdDWwZ
Ca5M1/WuZB7J5UCjz6NfRrQs064+Lh0fvusyqAzQyl7WJNRAPNHmToaHNNW3q6BC
O5z4Xnh2tGg8QPsDS0qRgmDCOo9+rLiIiHrslcgXg1GKlbgVSIBf0ppW3XcPyrTm
vnX/pNoUAfaJ0bxPD4IfEsXyI8ALsojhWH5cZHtcVqo8RZUv0JGbHjrjhYm70vc2
yD5NDTuN08KBDwq3eoBKMVizFmnxBfkpDX4ffjse8LOAFuZeUg/fTScAnzrZhdaQ
vOD31+dV3gkDXZWXNm3GgvXde4SuueymV5SOv+VyIxfpqGPtzQB+c1KVE+xulhUK
6KL2ECDQcukt/6tDEgU+n4iPrSX8XudPk89DAhI/PvHGfK6om9ZBfcZSvmLSgYy1
tRNbXFEQYLPOu7qKUwgQ41AavGW3HixJrCRRVXuQGAu74O6K7E66mmXCZyn1kWdg
f1xhNEInc//e4kW3E+tUPZ/luswiI6e5dr1JHghYo/sk9PAR4pwpnBHkovJiAlbW
QP/ITrg0OZCCnpNkefX5iRVRtarRCuGEc4qS7ykbPSTuF25MO44uASaQ+vpV+6vf
d0Fc1gd0IjXdV4vL0M6oONxI05Cx0hVzv5HsYZ9t5xFje9LPG/VkIZ4E1XZe6YZu
uPFYbemZHvKcRWJLdRNEQ8h1926v6rd5+yvK+3qLyplU1ba6G7wLvDjY6whccKXn
CRNMZVRvw6hPj2OyiNycP9sDv5sxH7t4ehkv89hrTNbY2o3eAJFbX13B2ahBgnQc
EOutkCCTbcI6SU4WoRxbRXj+CXRJi9YuFCC2twEAF3PW1SnTlvI6Ay7lx+nB4dPX
z2QTn5jrTt79Ir/lI5uizmYKx7lW+WnoHh/XJT3U6HcbIFbGYe6vlvwga6xDPd7d
uP7uZ9Rgba9OPxzExm4AIMqN5lAcwwO4VXG2JAbUuXhQuj4WX2UodZtA8oRRUOXr
hMAsCtTg6Ll+fvisdExEoXdKRjZQk8AY9orEFU4NQPUxzeEUCP9JTEi2sT5FbicI
U3QPawx5IlxSiZXPMAX2LMY5MBuk/RPgyuAkMhD0/x7f63AvzCernN1y7O5DWeRq
B5/l8XsoErdn/FhsBYcl+2TI9AcR+sbqiNKv8D/l0k6FxeSHJgsKcV6DcIZkqA3c
NXmeVffYQ/ZCKRAEvOHEnA18gW3IQ7hPcmjzUB790ueirjK9SC3FejaIZVL5Ivk4
V/LdoApGfz6e+YpN4MClx0SS8Zm1Xxs4MjlFlCgjmrEAzHYvtxD2gr/DWya0V8SH
Dbmwit9jd3/n4tYJShSLlHVBAxOtB1LISu7gm3uohW2IMxzxm3rhsXehk+dbX1hC
j8TvHdyo+mE/cbPzljzMwAIkyPauu9eo9JGWlSxZARJjQ2qY6oH9Au6a6PMywm1T
7MeNP8IHfGpNQTevAq1bqJGxIB03XChiUQHS4BcGxvp7IR6prwnOKRxmfr04pMmo
zfEPqhBg7HHAK9wTLF5Bk6MRHwCIoiKl+/OkG2zxyWBewQoCJGBo8yJ53rbq+5td
9PYk+8nXWka7hHXUazNbZdc31RxXcryJsr2DRF2P9N5BSpPjkcr2xgTHV3H4863c
dUB4V1c5PVcnnuu7nthCwmxMtRVIgJeZHG2KnHUFCVRVVGzneM+g88DNlo0NUhI1
CS6jvmvWNPzEWTnoCXewmlWyhEW8Kq9LIWAfX9CFnhTVAQcVQ1CcYeAdHvCDAw8Y
JelYSCvpivFt2hFXbvMLiMf6cXS0uggrehZ3adCcx6qoJXJEFwygS31n1KNvhkba
onwPztkFQKzzbS4S1zQ4vIKQHenHdQ6uap2/CNyV4insIcNCD2tVL1DaPZ90/5pb
QbFj+za4pmum/OAEuk0ZcSyV8oqfsQjEdV+EL8+VwmOAyRMa6kIfHDUe+FEk/8lw
emUsGI3UB16Hx83mKcoSB2lG/lIua4g3UfSYkNrbpIk2C29rNs0sZgQ0wrFRPoYy
Lc7zAr6wwlWwajpBUuzJ2+SNCx1UQ/kZTpDJh2uYsQWHuZ3t/WOvSSkuTc6pVkj8
x5feDYXnUzHFZobj1IzpWohGrT/wGCcoAxXHKr97nHBZXFcdRNNa5zAnGaXLMUyy
o3NczcCNuc6aE+OClETsE1aDg7RZnkbxg2KWGkP9M7HsMkz2QUguZ/DW6cICSVTl
WZ1CjHUI1/gQcDPWHLtQmqiCkLdY0gpWwHEDHKN6jIh/D9DuX/+b5qpjBzlZjICG
xWxHLFvvJ2d7OsoFY4tqAHIK8zzh2R/QK4SAXjGMC8GaiiXjtMAFxHnJVXD3Hxts
xSNF/Zwod5eH8HHKBRSPd9uTqcNqRINKiT+R6zJjCK6ZULgD/8WaM53aLy/bEjQq
pLuxQ0neT+PB04hLK+v1EL2WcRchVox5rZq6H0G/rchSmLnV+63WhO/HxzGQNMbH
OD/WYlMBM7j3ezdGBxey6JKsm5SC+/CtAesxrDRo1p8GluCglZCgENMY0Ltu0YnC
OHivSj94vIZwT+ld4v5LcbloocxwkTsVzhkIJhpWeaUpoJe9zazERlp9IVXKmYpK
LGdy6Jx2xCqYYlYzvdmf4+ccQNwSeG902k9T/w90fHa2VMAab+6qtI5EsP6UDrq+
UHUPbeSoo/j7nO8IY2dz0EufuGNSyJzNKvzfNjTpKTO2JJGRtIyUtaB42+UGxy2E
q8XbwhvorH32BQpsXfx3JrB+kRn/+3CSQod3pBbhjgCIJ6Yi1Bo9seL/BUTm2A/L
2dkonxmXkUCpRNuPQxNrguyFb+eDzz19anudb7AEq2NSM6nUMIj3EFSsJsKpA/05
se5RbiFdFqT9f2PX8OawHfQldMYLfPeUw92wHzy6TGUf3/2e9qm9EhVZSJC+2f7s
fCTqTz/t1gW3aGP+WTpSVU/pdKwN/AsjbcVz+8PtyO0Yh/HR28exPmA9AdLhKMTL
tf7dQ1BF0up2VQo26R07QXzCxX6rUDeKHo0SftLg8vpKQMqXuNA6fVCMVsyO52u9
PEcBmfwOhyUKNR1ZV5FcEx23mj/7Hkxah4mreq1VM4+5TtRyB4zOnrlTcVB3R2It
NUgxkYkBY6AZetyVbyNIs5pyZaBc7Z07+2uG0RKoQcx7f34uQiwS49Eql+qCeTz8
75kbIv+ZnOjC0OI1RQFP+rFys26YPmDGUW5Gh/Ia4lvYxKI41/5Otvu142IBjZBk
34v8+GzgdT0WP/iXWYZ8Z3xiEw0eLW/ALtPuTNTydZw9vqDAuspTsveRJ6LRfxLb
oqLF4iyCEKLtSFv40eJYvIRWS0lGcm2mbS1kIHHgNpyT8crFw/x0hSLcd0jWksIc
w2Ry0ySkKDcA9aYGjkP/xdvPbbyQwh8dIIsA8IPNu2a7Wr/KlR9r+j+hRgzJiO6Z
x2pvIw9uR7pMPZKmfikLQD4kVssceQT39zjVWVvoxEvhANanQh3dZGi+qFj2rGQm
ZrWjfr6wHkXrjw12O4lbMVpZmQQkbcpRsmtt7Gtvh+gZ6JYcgOOKBb1Ygs8wJwtl
KoPPGt2okqB9AYuXkcwBOn90xKuc/umZl112o6Qmf9e+WpWn+cW6xphLQZBozUVW
Y6MQdHbbgIcxT/DIf68hP1pFOX3eLKvdmE0rTjHxjC99tTwpTfxv7FwLvhE0G2+6
HbPhbaOn2bDxnWIf9xqbVP9nEN/p2BC0eabNECXTvezG4GZd8RPvytiMlZKhZPk2
ZKeu3Q6NqZIqpzj30cHy5SPbYrHLIDxvJiOanIxHpzqOKPDlHTxbFEmS0ZThG+Dl
vnJDbm8BxDUuQyMKdfPX4ASaKvw3cpmgr33OIKzHAv0FTg6RZ7vS5Uq9vTSPi7Bu
k63InLvaYSdP5HNkAuM//X3OJyGXg+LY7b7VrCMAwvyM4YhymKvvWHokLSDptqfa
83E5fFtn8C6I/UQK0yJGdklkRJy4/Z83uwdW4DkZjeliTKuXozo3C7wWjQa1S2TP
DI90dUPATqSsU9Jmc7ZNKZe//waniqho2LsaVx0MJRcbg9iMPJgXoGIa1EKEoEEF
NDidGpraKXSUrjAjNZYAEmNuKiI+Rk6N+onEA7FurYhi52ZZHQk9cGLDyR5xG7z8
xn9iLWuR/62HFz0bbVXL7ILv/i6M1Zrbv+KOyOQ3lUKNvk+juq+XgXq2lzSHZfN7
vHEGMJwYCtKSfd8YXevEh4BzZzNSPYthP0z46g8Gg1YJKA9YrVvyWhd4E1BEKCdd
cBE2dScpi2JKvzoQqPYfe/QP0lnVO9kY8lXdRNMb4fEVlBxHhNflwAPblTlNeh5c
ku9l3aoVkBxaBtxSIqMDk7ceqCzGyGCTNuJ6S8IiJLo9HQe9DoJ1MJIZb9BGbEFh
Y4rI5ezLR1/XPhhTtCoZBZE+7mju06WkbwEcHpHg3LHLY+STiByPzFfRJw+0xChR
W+QQkNN79oO/GNyXKkr29DpOd91w7hsQog2lPMU1qpEPBPu3Nq1Tpsaq4e7dilyM
XfoU/1pnx/Mba1jYl7jexLHL+LHdeSH8DWSFDzyMqah8qT/yXTwVYuhLx5xhLyDA
2RUNBTFjTTBYRNGlGbTZRG3GQceRAtetSCCdSUHUbrW8Ox3VkqQblbYZVKlySQoD
/SMFwEI8m9EgVC98+eC5wa3vHZdpv3zwr8Lj5YaJAgzHMRxV8GjQs+QKx2gqdhiQ
GR7IUxpZJz/Blt7Ra32KeA2/16bYqRP+HJkAsKC/ycYjct2ZQj4338UmYT2u15Jb
WpChtMpXLe4kJtpC9tsBbwfVL3n2xrels+tjCwHTDV6WSepN4uOm7rss6L0KbJN9
wp4kdXn8soxj3lYljtGxxxZ/8WEb0Yur2jNFEaW9iOKzbKASadAC1ANHSUuSiJXj
tNQCvNQwuc0N29ZKk/aU0IokYB4/Yr7UetN3gV6UB6jE0Hiu4MAn5YtfC/cwhpB+
fYNbFsmsOYE9TNSW8IJSXtMZgNL+ZXBCKbEYJOY3sLnONXQF49bHA6M5I0Cjuge+
q2B1m28CBUgpVQ9O/MpXHWsFN8UU1snClwOvL/MGpE2U//ChEj94aOYmsQqfQjEs
Wo4xDa7vKvBTqwk05C29e5ZJBOMKakf3JqKJxNZF4MmXNYfXhqkaVa5vtP/7SFN1
/LU6wwrSpD+o0tSdlVtAAB9WhhIT3TClCWQ8JZhjhcPdnMhqGAN0G5l3od0pk4xJ
C3zAJlouPv/5i8kwhSPDgspyCMce9TW3gZ5GLFL1lYwFktS5wwQqAGoGxHg8YD3i
1Ww/1lWC205f1X3U3VfbYjEIxClDyIWIy0noaVg3I76QdbjLU5ycy+/NO94Mp/q4
66G2UHwnxovpIs92Fu3UC1Xk0SNyiURR4qHr0oCONe7talroJD6LSDOS5PHNvvcz
d5RsMz//Rq3rmLUlVQ8UQjnYz951i24hXwYtU0jmS+SlJV6/95bnAzQduXURsp/h
k8yIshFNSYop1XKb0Eo+xIMBbEfAlgaPhK+Wnu2wuXR1ySm+c0kzKBOhIpVDuyQC
8hU5JlOoI1i2Rc1bu2npeVthBb/07Ovp+76zoeM1pQhaetJnYccMfhZ2/mAIe+7W
nGMvfFFKuBCAXbayqlQQtk4yyueDSpXs3g54R+62AJhSw9DxtOvhVF/1CEqDt4C3
09a3ODi8/8exzJoUE7NsWQFMVS1eswz+Y+tzhuYc0keG17V6qKiGeoLXSZ68ng3Z
rVt/Ob6bfF2v9VCgRZbh5s66oXeuA101V0Gy5yeu3W8s6okcC15NWhstGTKNZGXj
X6+wtIjrdSlHJHbAq42J8vbHc9I21nDphkwRftXuoyaXgIhYO8rYbPAD8ZYui/dN
nXkDrz/UoUZJy/hcD+MfY+7NL6nQ1cdaI1GxdIbodwannIH8SNkHTizEiQ8B3YCf
mfL+jO3/xRvVaxFf35x/r+kwS59ElRImhJuDRV7L6MvK9L7u1KOQ6xvGe1c7f5n4
p1yp+5JUaV+wKwDg6AoA+QCDC/JzZxlg0hlfzCVggOzR15Phkx9JIJjIK60eEQTy
nlR0wcO9s+aA/biEhxxx6BBPWDSsbQ26vtW9m7L8oTr7RvsyHQuEAxFR+Pl5iPIF
vlISPtBp08tI7MH2Rrz3kL3fPCGVEiEW5cZQOHbRkLj5K+JcANmgVqbvMd9lDBDi
C9IpEdIVAI9NTfN0E/BhXpcryZ96Q9sUEuVFaDUXU2+rG+xLafN9M1KqGu9YGPeX
a8kM6neA3EbrI6tsW9mJTcggpbpRyfOlbM9tAHEBmGvehkMya216YxaE1dLZQGgS
OK0UGVPhLVy00lFCi3CgGqEyolEb+Ki3OBJXWHSeUEbOzT7s77NZMNHklXvUT962
MMXEIWBZvuVNxgqT/6ZB3w5td+PNTWfXPCRLQt7WcI/IWDDbagLSttbXkMqVBCHC
Y8EmuIGezBJTqAsGoKFGHNsTnlVY+k2Brh3fJ0NYiQi1d+SP70LwF/wV+JPRRtl3
yxQPT+SUJkt4zhLEqo+cv1cCI06UcKEfgI7+bxUqUDTzdqQwChgxn8FjjZgVwI2q
/+yh0ynRFAt4heNy7cz7i1DNZDrlLkKrEHGz3lLzYVpnjODetWJx+9eJeNBqSa4r
2cv6l07WzFsy+QbWWiRLChETpVObRePa7YUwmVpSohNCkEivwm1kEVN080xk++1T
iKA6keDyshSwfXM6J2QS36QurpWj3fF8grOiNFknuiHi9GS8FJ407N7nhuG3g9P1
I03BooZR9WKRMbgnEgGwmZdbWFIwoZBF85DrCsvcpQQty9wDzyPi9/g+q/qsfUFa
kEct+0mPzCMbmXekHXnNMeYITPnMnNUTtdUu7bmkEp5Dx1rsF9pZlPQaqzcEehUl
PfQ5ED7+eKxyfMxqbb3lEjU3Cs3XANT7maTOGSaBYYgLro+MBQ18dCb++wDa9f8r
YhRXCgU4+sJVD6ZgpbbkkIP6fHU0+bboGpfSmv/AXjLtbZ46H3NQf7+8AqV/vUYH
ncfkPQtLb4J44T+eQ+sPKuNryPlSnqq507SwCuujCWfmRi/+UZYtSgoTX4PMgDeP
5LWNzxSqeE4ybfBwmlCzfNj18iS6u0WcS5lI6M59fYJ2zsBqRx/+1crLIk7RO9uJ
jGllgXzWLooQewVE+ko+sY+ZXvYjGwr80As+TRgDgilHOy/NoSwH1oGqzhuAZCtL
Cnplkd16W1Ee0L+Ej/CxPSWoYIrtYU9k6znXy5FP05YG6xyZxlUJDh6ruWjD7PWw
PGch/Z9YUBkcqzplbmcvqLMzHoW575PpnYoqZX8n0BMGRy0kGLcTOQ3lgfB+Lvxx
Up5K1NkJANASXZFTVI9uwm1MwUoKTJaRbtFqkDD5x8MTF5eKe4uCr9ikIXaC0UKw
YxYyHcK8h878sQgZRw7s4QHaB+Rj5wibu/8rtQBF7QkOdSH4yeSKVLJPvrWnzrjU
kXWNnJ9zNes5Td1tqIdMblxu28aHz9gd8l3cq8LMw4d8ObVQ9qzY7CFYaY1LyV5x
1sBL5C81NVNEExQSlLsS19HxQlrcV7JPDEDq0xxAO+NUPyD+U4bZyS4byW1yI3rt
WLberzk1BNKuB2rtDK77+3i5L05BIQ4diDinBXHi79D5/oOFx6taJ926V0Mz+Cy6
OW0eAakwbs4dOuhTvS0Rav1tkSeVswOZMJ2GbT0IGYM1uvljvwlYhsZS6GT26y0R
e8CNEe+3wNtmcrUOliENb+WU0lX+MgUdAk6MugYSWjDmrvDflBsJr0QZ2/pFvswf
zMLoM6nE6mtsh/QGU4Atg4UiRb/9goJD78sN7d27ZxAj/jlFpaHAoDgsjQn5/Xji
`protect END_PROTECTED
