`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PHUtTU9m5Gbbh2N/cAcW4mAYJFuANJ4kW/xHubsA+2qpIH7Yli1W6aVXm8KsLANQ
Tmz5JwvrJFBWTIj82fKzsOCvebHsoQ7by3XJaOk4FEAyXGELUh0wa4P+PxSf2qRY
GWi7S1/l+WCzRpw3l1aZkQy7mvs5btMbRwBxGGsUkWXNt9iadSb1DjhvJFd7AWRj
PjrzP+vEsohR2oXQGWJqIgVJSQX0Dt1Sby9JSnOANU0hfLtssbAqtgc+YV763nhg
/Mdx6tLtyvODrhWCeKGX3Tq72XoRjNljvuzUAce0I7HKXrT5QxxmAydfPjCXYWw5
XN8b/SHve5FeDVQaSYdHmr9v4rF8Puc9kfg36Lyb+xpRhpRrgjoiHHet5ydPqRig
jWxSS2A5L9qHNW0wWYPExXu6uuqkXNNahL+FtBWHp2WeYQmrMF9ft8j1Bc/XNcEb
0InvDGvyez4uvGd536KA7G1onMiHA8WUqyVJ0AONUigd4kSTdv4U+r1MVR84yx1t
`protect END_PROTECTED
