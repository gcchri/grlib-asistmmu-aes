`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qMYqbHD7Ra2ogCGgw6onMHSr9PsnMaV8mJsJEMrPeiMQOAPgDu5FUJbllg0vtqcz
5JGV+IvMsRDfSOjFmRLL7ggHii/OyVb39pCkwL2Cns5goMwGQ+MI3Wd/SHBhAKBd
ZffQghAbaYbGmfcHCh6V2SGQ1PY9c6679U2Qg1SHhJKtZEaFLumgGd+CH/+zwxCg
qO0Kwi1Ekke4luShsfq2UQU48RZCg4Cf/u0kHrm4UCSOzIpq2DgdNdbEXun+jYLM
zYFF9QpLbgR6LkcG0m5VrvrvqNWVlyS9XtwT55M2oJmm//xFBLRaSh3YeoCPu6rg
Yn/jln8abAOA1azrO7mGYds1++yKrCPeN0XdzpEHar/DenZYGlcFBa1lin1fcjSu
6Mwkbns7o346sFbYOjAPXgTJ3SdNkGUyC5W5WZOqD2+Dsus1gGcGXUdrE5uaM4U4
G/lN5DPN02M+17YKyxM1UfxV0G/93N1+zxPBttj/DIQX+vWMXb2r+YOglwwRHThH
7m89fCQw02Bx6D1R6V9VvKM9961AJ6yvLKajeMInVnER88oO91t9jpoUdLBQgIpj
np3bVX7yLntI2miFbsblWQjqNsNq6DRQLc4x2Z/yhn7uWLmnd8h8+3rAZLNijjE1
iZxjRhARhCATHO2xfeXk0Y1jHiWY+hYFFZBUx85zEbsoQKcKuWAsXXZEMQWQuFWZ
nZqOjx7wC4gvZt0lGwfZ4RbsdHCTkIXId6lTzyyWQ8MH9201YDK8GR/dNZf18zEx
mAkIbqKkHTLKbxfpvxmx12wVkhDv+/r1ort2g2f+eNF+rLgX9UO5U1XYiu9ygrqq
Au9quJ/XYfgrUM35nBiq/QyCLIHTRhSq29LJKlW0lBhCgAoCE32EVkDoWEZ3AOvs
iOkzRXdIjZL7GEb1cYOXQH8rzyHn8nzjz0MiLE2dx2jHVUEt1zqFoNbqdP5HF7vy
lHP6FVbQCDD0i+s4nbwT5epcMdp8TOOQo3I3QAjyeEM=
`protect END_PROTECTED
