`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UzPjd7By9myjsirCNsuVWgUdV0ywfgNfR1VqyjruqYIbllPJwG4V4hF5mGdzAaTf
8OqYzKagFpz2LTH1lhFdiap3ttmiLbtmlIwsyIzqqMYWZHeEVFNqp7abr9zXYVaS
vwMGHLSIpwgx+BINv7qQjHFA+K9c/20kVL8bPq/mtBXO6OKo3JsXs5sZad73hcLk
KvP1RoYm04JsERouyx62z1J8WE0oMf6fPZAOqAlUJnrQzEsPIdUL6WfoudvA3fT4
I/8xoGR4WPeagP0KtTgYWnUFUdSrctBqy3TH6+udm60aW07JxUOqUeAfJcVIWIGE
G2JrhQBs+DOyH9360k/AZGCfTQHARxBqJmUpjpTTVO18Zbio0n+JYqTf50TNkxRm
LATFAJyYjnseVSpo3EfU2GYXTBXdbcRD4WN4PumahRqEk8mAmW197W1hmAS9zh7I
HlfIBbOCnT9UwHHX2i5IQI6EqnCAgm9X777DA+H6++jn9rpg5RRpnHWteICsTBIm
Mf9r9ZxCvLv7J7aZEXEB37ddTLtc5By3FDoWj6xL/tSHJdf6Qam3sTHfTxJFCqVU
ttN0yPACbmUjaxBvf4oYZg==
`protect END_PROTECTED
