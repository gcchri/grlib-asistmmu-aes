`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7q0zGDyPY6xXzzgctHye5Cs8l+GpNgVfWTQmmvEXnO9phUHGao6eHKNfDfKuRYTP
Fcsy4JY7R63SmCuusp1gu6o2Uut46IWsAZf9NRNYsZw99zuy82/mfWT/l6CqX/wm
s/ojSCIsEnL3mYcw9muD2vG/mYARcNchpncSZgtwverjPW+QSDCzP8i4ZcEZd2WD
igmT5bDjpqMxWkPa/NkzorytHd+jgXwKXTeZlKsXxu+T1MIvsjBBWmiYOY5YjASP
CUbTly2kNs6IzsiuiLK77xALhgGenh2Z+kTxhPF3JUEXgxcHLHby3zp5rX5XoY9X
6RAASOAEpJL/YXPXlETjpRWRPZ5gPzLpAdlxEfB39HJJ/ojcm2pf0vJKAk8sL9qd
oyOeFpybtKOA4O7S+s7D41RVHh/bOMtnMMZjefkDypfW/eFZz1stZrlMaGnyGCc6
lUbwYm7CtZH21+Jpqbqn7ms1g2j6Ng4stlDMe6SzU4B1WZxQjy0TrtSoqOflZCTd
UO386jfuScObZ4aHw7aAXgyAKJVJtvfAnV9W2jN9+0aVfDaoUgeWXrpingCiBZCq
d7yEKcfmMmBdHXQOOrYraODFBDx8jwnt+8zVTQQyMtRxNT5MjG09PfzBxpwNpR2u
Bx2v8mFksWykdEH+/84QuXzMrZA1bLWPRpiGU9Y4hf6tg1d7DcvKgCF/XLzEdWej
s2mNdXMrCfqf9tQuJrWlp4Ucsg9wi1Ohbcwa4Qsk2Ug+8RZx/OPa3NUdVJIcx8Ml
EiSEu9QQvcju6BS9pBK0cUKxOtxtfit3CiCnePCBiBI3cZJLSSmOaytzLtN9mJEQ
TfjkVquD3KZAkDnjMyUerrcAZ5pEWZvNBGu7pjzvotfJ1kXwobXgCS+PTeKN66vM
YYtHTVTcsih4m5GeJyonUUMmkiJYqvOJ1ra/xPw4pCNM9sQFItD8D48W9OrG9VvO
zH2z3vUE2ihs4UyKrgyyt/43npWs5vVLTkOIjcgOK0WMSqboYIrzCwolgXcVxqAF
5RXl1AB2CSe9CkYLVdMSugfN/1N3976P2CJtsBgSWGCjXKbIDKzZx9hvdAesS3+q
1xAZqFNzXuIulA6uZRYVYXbxQ2VBeSnpALUpKAjT3HxFA506P/QHx6gu8M0jpfhw
Mkz9HQqvd0zjNoV59g1HxmgP8JhiyoDQBOaDKaA5gz+rtH24JBNJbjRXjpRIMayj
e95g9pCPhaW787hio9Nty6U1J3Jo7ALcO4DUarW2/wymiuMSWBFrBmhyzG2PNogL
8G/nDoszNQI7X52ZzxWsNWDAa4foQg6StfvxpgArpcnOgjCKwGKRhXzyc/fKJeLv
v8rwaGBxJHxc+0DQxQDR9RXxuuWazfocgPta6igWt52AKNChVBJV4aGfdaDKgRr4
bNNONxPGiUhwacEImGfbXZjl/XSQ4jlBPHVsam6tZkfY5EjBn5Brwetz+v2ZMiPj
M5gocHrTICXur7HRxFf/7iO+UY79cL590ynLVn5VsXjxGV+dS6Yi6UmMRfFnIjTa
kX4lv8YyzzrHADajNhuWEKbbd8GeJKZiJmpj33sawPh6WVOLuYMgaeVUI9J9TCW2
b2tsrfpZ0tpYzE6RvKY4Do/KdWHmAOPVY8l07LEl3ax0H9xrrsa/x/oSUrBJ48bO
nTml2cLrSBB9DgwfP5r5wEaRYlYsEjoK8QJNL7riprERGhBS6tyBErdj9sWyFilu
fhsRnqBaWhB0tLt2foeNJgQt4jZG3AeFdkNB2VmsjXDZtBBgxagEGOww1VsC/eoP
EK4o91O6Ket6whtki8aGVs/KfJ+Y+STx+Oz9BmoC5ZVXXJL6OnvRGedEX92zGAXw
YCjLKybTG/JpT3Fb8YSxclOkT5ksgORmY27LvLTXISr/01R1I119O6CaUhmiz3o0
TqFvAHQEoRRj1F0qWi7o+rl32nbKTXcTzKvI65EBIwOmH4pWl4JcBvhV/svRfMb1
gw3zUCVpoclkuUdsqkbU5urqVdewT0C3zUEJUzA2MOm0qcLHqtL7hSywvijXGkBZ
iCr0F1NgDibOnEg7kwszLwYFCMcJTCgX+PCgc1J8UVA96Gz/tEdw4dOBtL17dVWq
ZRQneCbBeJDygLwi5SHKe+ssh/RGpZdQ/uJA2TQyCVMOY9BS7Mb97beIlkvJsGlV
L45elGOmNmpUzDapDY6BOWZzUd/28bVhjNDAS0/fLYQu4Qslg7qbSYZYaP9S0ldE
Ca0QV8W4S+WWpNP13zIKKlNu5NiRb1+MF0Di24mnpdv6z3GHDP55Gn15OVVaqTGs
7AnY03EEKkyUv8yA24G1uiOjCePwW1k5iwHbnJKKNoIA2tPQ3S3YN5YqjxgnCtAB
1gp1QfIcLy3/L6lPSyYBF6iR/htlmrk8s7fhVyM+tqZeLPnLqIuoCI31pXWK8Reu
Bg7yibqkIkNpBfewgb0dvKqueErFCx6ay3NWkc17jUq9e+uXOKTyKAfbbmka6eu8
/0/2PCtlg1Y5nWiEownmwxj/5zcl1lLYbW3oT4iIfQ0WIOc4+nyHkMRoDCJnku1n
OKI5L9r+XupXEPysdmU7gnf1vTTQkNGKYwry4vAaIVYJc1CZ02FVV6Q8x25nYX0V
shxbbzPJGD0s8NuGvDW/Rasc1ZNX9GN7aEBAiqWNFtYuqq8EY065QaqcQkz95OAW
8GLpHVMgCzrzfuHN6GyhrlKeAtjPS5Cm4EuzFkSplfYV+e0i9gZ38hJyVRdtOfz3
nMiw7uCVMfnlVLERz/GGEwqJaiJYwH+2E+gc6tADL8/AIOAyeyp4QIHk0amkxucl
4uiE98KCNMixZ7I0XwLuHJJ+MXJ8DDzWgHtW2OTC4YEKSBN2eNn2H2Bx57zuwnLJ
WYeQdCW6WkonConTE/SbneGGE/Q52sLAL9/oslU9UAKJmyfbPMsGz04t0jb5xEFU
2en0+gag8W/Vx1ZXxnqUMpFj71WGJyL7YA+KXNamlSlo2gyYMqajHafj8IeT6Sz8
BzeWurbQPaBwpjnnyj1lBp1aWMp+yZw4agp95SAW4U2beuhYuhPIUIs3yl7rcsBE
Ocs4EJ6UfYZD9EEPRR3Q7bsGsc3SdZduNbwg+JDKWo+W+Dsp9pmmZ7/V71hOCLEt
yh8eB5MkV/kLOtmlfdDgw4kBSzdK8BgJ2ICRT5TMwYno0NAokF8rwfGYlPABm1DV
qZFNUcJ7cfsiTjpe/mVn7hhRqeUyJNrjXSXNkRMJsH9ThQ+mb1Cg5oAmIDVuAS/H
X+OD1HoCow3Rqzya1wEwvLIPCtm4QX66VP1we4+GLMuQkFjb++2d4jNLpjaP7Sto
`protect END_PROTECTED
