`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GE8UWzdYc/WrH4KiZnCmuh1cqhmOcu1xVrRVadrcVkwWMTpQPyRH/aW+l1tGE8wM
/4aACVaMPA+F1nhNswUv7UcxnVGAgEVSj3GVC2Ih7AL71IdXHL1Nu5idlAFUVAIQ
MpyxdKFOqVm58mJo7WOn70zvndH2SNdcyhu0+X2jaIrzhVM8MmWg7TfVPQZHl90U
xFXsEvhYHFEV933MPQ+uX4MaOZ5ijE0hGCJBqzdfVLSXgqZo7gPVu+uloWCsx1JB
uFP5qUzFBeUDFsNh6K0QuoCt1ab3L221GYjeN66HVIntNKiuRvq3K0/sEUmAPD3h
a1lhueGcus8BcllU9Cc79Ms7Nt8QTjLsTg8UxphbKZE68F7FwNrDV9XYnd1LpO7Y
ghO6pko1IV3DIbp8DUIY58UXfhwcUsskYRJCN5AU6gT7ZWplMfzfxiXQELIPgL1D
Cy0hcn+Lh7OI9KQbHiR6a8n48YH/9LkQoWTzGyI4X+9fPdHKybDHdxf3cpm70DHQ
ASBFqAU8iPi5YJfLGqt/1ws6bSYokGjizBMtzVQ5LGaTlYo1yi7tmPn29dpzv2Ym
`protect END_PROTECTED
