`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pg2G7jlxvWL0dJtw2UdwuRlXJK3bTuNqN3lAu/C5ORHzoA58hy85eZv7u47sw4iP
l7lA20XzavpZKAgIeGHRHxjM+QBU0NAgnDLwGSyC4Q21dPokWSqcm5hL57YSS62w
wMJdZV6TQQC6dXAJID6X3t0p+6/kFubL0dOfCu9TVfh+mY7y0+Iymfftq20/usYq
omG92R83lwets5g7aGbvxIAfkp2hPdxZOUlEyWpxHLUvnmj3496c8icB8tUY3qu8
1RnxcaADjS0aUq3eowZYeZqxmV0MKpJYU8v8bZZI5ynBKeje4yGgNb6H0DY7oChP
mPdS+Z1BuClZEuyJ1I6LGnZ22eXH2j+XMm3CI/vHApYDrf9BhvsD+5IlluWMoLOe
sU/JuaNMbSXSqR40VWANyTq1YqemvT1B6oTx5kz4oiZzXvSYKQf3KlppA7ADuaPD
tJi3oRQfb4rv/S+KT/4eT+G9DiZawIUApzSIqL/K4F1S/f4+bIA7aKrAq0/R5W6O
vOv4NEodlbRPodIzKN54QCiM2LTMqKklblDAfkhTU/ra3FOxqzLGh6fF/iuJpP2c
A7tv1Fm2QSspXwAW0oZdhw==
`protect END_PROTECTED
