`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gYfJqnOj/0L5jFwUv4JD+XDnSjDh0j/XpFkYTZHXPvF2T1mFimd9J83/gCID9TH8
1DacSMOtB3dYgTeA1WU7qIDs53xlmTcTw9gAQ2GJRudHibjT1w8YNn802fs/GupF
1YiWESGjXJvXYT8B0H2HfWlS2yc0eQxGUYxh2mh/6ZLC9/u1rSN8e/icaKyotmVX
N9brCs4GDwhlGH5w0qahcDbaN6l7xpIF0Q5yohcm5qIqzAE3EzOo5hJrOrrZyNQ0
LkyH3dksA2t+ufUFM02fozqFFVdaPpKjlodJbk5spOo7vxU3AXn452QN0oezMfgn
QKqn++KnsqkxIOEsSqlDIJn5y4HgteceQBNs8ADePIfq6ona1ZCaFkOK75Q3gdVf
keQL053lsG/HV6EJHznovhJBOqTzwBRDMgD+No/TVNwLBimR9kAYht+OaPCb91bb
RSq7fAWZxm9GHQgoYxcy/wlV3JiFDpow/xMCdgCDN+b8k1+0Aee2Rdk38y6CJetV
J0VG66rPdQO/Bplf5rRCLvJcTKCjW16W4hbDGkLuvcCrYcUFuELeW7asebVr2bRE
ECQVPO3T8Z92dbp0e+oc/i5+fOIcUtMKMZBYf5K/xcQ=
`protect END_PROTECTED
