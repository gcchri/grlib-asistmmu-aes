`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LSQ8TcdqDZBVI99Kf+Dn/q6iPH3yDwXSDstKcqhdTOBSqngvj66pUpPKOvp64iw6
zXs5zzzlTfspCLoUwtt/Lw7PG/E0Eg8vfwY6rNPzDXJxMFDu4bzj5ff9CjVqgXPu
aObR5x1ATfjCP2dPs756IjEymfe92NkXkTzMk/meEL0G50IF9kMHfXOzig4y5CZU
vOL0QHwCn4ng4Uqnd1fLdhGwL3+/tovfPHRjy6DqQscm0fZHrkFzWW5YscbHZHXM
5jifZuxm/V20xa9yi5wTBJMs4hqhIlOGpUpWOxnhfgiy5nSkK1hh+uY3o36Zp17i
DuwUPnUe6WR5ohoExvwaqA7eBa5HgVItWO8P+o9wT2yFDkSW6GjmQd0r7oM+fumW
hXm6X04HS2NzfjlO7lZq802CqsPBQVTa6n8svEQbigIA8/U4YZkhmgda11G0Tpmb
NLmntUI3+4n25XgpLggNp13qXIyeRX73BG+igBtI7kEhlpDNiHZsfKNQUL/Ps9l0
jbUUZBmYFN12O6Sjsy5v9OqdtjwzicrRuzRE2DCIGx48Pp1XcEXGztBv1FkUZQYm
TWcbHM6b9iLoYAJGPkUVBoy+t31Ae/P2uTlpCkZoc5Iee8DMIR7uyvZkpgs+Oe1X
UtXoYyZvaJwbv81iZE2hfAq81i+OVYO12dqBia87bV4NtCXJXbcrJAPPa4edPLWi
/fQAvBdgyP/0WD3279xm0kij+8ld4hK9UXD7BINbOcjAvwzpq0Xg3BMjMsr+XxUq
xTXFlw9LzcFMDpsTFWT0LbCfJmQ4ckK2U/AcS5lVKvtDxfNnnwIO4i25vrkuO0B9
KuBjm9g78RLDFgVaiAv/kvTfXMC3bwh4kFPf/TFA450V8djJqWrMHJcFMK2zkitg
hTdOnGHtjklqXj+f4diuBOSRjLXJUetulb7GbzYt66MFRF/Fy56F/bmzLj56lZBB
KJwxSNjYGMnItSMf3bMR5YxL1mT7hOk6DTEUrPCv3USN/P51run1o+4EHjEu0YaW
/GZdUGSGTS5YzZ+Om7uKoMg2lCs3KbVX5ohSJYL4bI9JjkLpn4WHAI84TcjDwDTK
uy3vSMn+CttIDuOJApZUV9gme+hHTRUy1pYaPOrsdqgO+6mAPHUh2hEhQESex/It
Ou7cmh1yI7Yd1Gw44MSJVrE+b+eEJo/6ZlBeLboNipnlqo5esKh7dadP6A1Zx2zr
UOc55m7j59BdLrDmwo7iRH9m15828/qdlgVWljLZl8dVz+v1ayN3trBt8BfGRTDz
Ho/q4lou3+lbq5i1zGZktRf0t+EDy/f4oqCwgWXjjoBg+ooGjuv9cDmqzsixXz6b
iDcdcrYbOslVsvJN21jjVoCxmh+WSpKoWc0QwiaaTmhZ/q6SwExkozK2YDUyCZJY
VrdKXkVTNBBrPwbQxDa/hrEC6BuI0sL9Mbo+AjWIdkIQwNiGhgYU3B8CdO6RbBaH
TsPJSWAU8YYet/udCg7yWHeWQee/JamJWGXXGbBFuMz4XK4ztt0PT143pI+etKij
4o3MINZvFl2ljNSk0G3OCvjJPREhzRwXRdbQmPLXrOwDUovf23G+th8KzfdNihjS
1LH1LS1roSIRV9hIRJzOg158M58MLUim0D2i3Ni638Yts3af0Cojta1sXspGJNyZ
IoCqkCAJvfb79EZLNmp1Mww93pZddeV4v8ikB6JEXN+vwCAqNIuPHso9Z1WWGDMk
SIC4dWA7SbF/CM+G9kIp6SicRkbEp49mjxaI+9Pi3/P6cOSZalBBceRn0LAdwR89
yfOj1B9ww4QHyfm7P/e0j+/pysN0sQl4pPk7GDxDZNZBDLn0T3qg9A3EOUDlm/mb
Zi3agBPuHCA+E7DCErk4H0naLsSkRAoz3iDX0lqge+dCYowU4xpBHnMBvRiy3lWU
7o1vZ3LYyHCSIRtwpH07hY2GYT214DLf/WPEurHx8171YEjGn8oKJPxjjkwz36sa
URrdimHfsx2v3HWRs5Z7xx4gfML1OnutoIVY5S4s1xWHGLwwpcfYj4hql/xbWJDS
r0/NGkyurLAl4QHaWj7TnuGf+FiCIa6k6HEXYIx16yv/p8DUERt2rdDAv0d02DFD
ajNLHVtiISJgZsKhRxJ/zSm2ZSjL+B3NJXfsgYB4GpeBlAYNad+/ewH860c3v/c2
f+pP+l5ARsgtsHbRkW+OWbdxY/2bMxgzCFVimhxpV4dX5PDhhgvl6WVIJW3ASuAj
/0iRPqebNAae/uoGtfZsbBIPZbgzSaXb0RBtYpeQJAMY9yTbPgXBFPZgGNMpweTJ
9XMN4NmlM9xGOrEFzSKiQ0UPlwajCif0oXxzHnQ9SPKzcuL7MyJEWwTMU0tp60ya
Whh0AKEZlfU/J5cqU41x2XeM6nld6bkFgFfXjEQ/6DdEi1AubAzO8D0OVh+rIAYJ
Hg32UDIOfKZt1RYxdHOqDIsFE3+ln1JODhScj0CN19MEpAa7Jf0gLZ82iVKjEqyQ
05F5KzwVSblrgxWUa+x1WtcWmDnTZgh2ny76F019WcdPcS6WmVCbA/jXk5E9fBqs
Bx+yyseNpnxvIv4RwQ6kB0ukHPyHLnwWR9Y8w5ZyFM95CW4ccvGyxMVxX+05v4+4
`protect END_PROTECTED
