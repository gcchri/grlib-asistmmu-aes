`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R4zVA5VmFf74FXt9LEMnXCNbArCmV/Y42dp72wLfqfcKuVMrXgaqtaqAqVwioruV
NZ3KpjXkZWopjZkCPbCK8dSxr9JxDpDymSbFHDnJDCv+6pfNGTXWuSkof2RNT3X+
+yuUw6QJeETS1d1QPzVNL+8bTKQyGubxn/vDerAzPqG3WUNdQ07BtSgShBxO6APP
6L4EbK17UNvs9mbm1i+RorSen96H7FrQpXjY56+dYhaZGYWTQ5K71hfwvOvnK49L
FwcCGSoMAe4utCUKfTIdtt1fNUdoI0UcresnoqFSsqkuD1KTNTD/QNRvxxa/TIFV
nW13F76SV1EkPmefijmvimDZQfc0ur1XVMa0bOxLnBADr0mJUOkrckIHQsqntBWk
tDPVqM3EcyQP+xpvb2vf4r5FqzljihsG+zK+LSr+Dsh4ZLta0Toad3FkujIGlgDl
J/IzOlA7VGZns0qRAZOFeJoBF61o1pmL09BMhguyOwFaevGrlo3wWQ4qIgmatkNo
pDSnjJ5gfVeVu0LAhBB2G644y0gDzljdQfs+EAaJ8dDRN1IROFV765wCCfbZiTim
D7Xucyq2E3t28QfRe0hZfAY4qUz99wdtj/PdP+qSl8G4CdWPwv7B+pOHuhBi/VhA
YlHMaTYvOHUDs2s0h5IKnKUNxQIa3m73ADv757bE31fI2CagIoYBwSz+z5HjjRTA
vFFX49R4LxjBJo2YFnk6PEQguJBb7p4CiL0OgCcSPfc=
`protect END_PROTECTED
