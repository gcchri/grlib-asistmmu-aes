`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RcVOfwIQCaUIbmTyfv8XSm/OPBTEX40ViuP/VV2Lv+QFI6t+8K8TwDM6SiQc6WHB
YfiS5wpkGcCJEfEriIIBhw5hg0TAHzqVhHULdCYypMWZSFoD44cjoJqkC4URDHfv
DO1vXRCTCROFptsCOgUM/c9izQkcUOYo3NwB4yqs8VRJIQR5aKbZPBXbBBz4rwc3
sFKk7M4LfQNDR4TAK/2L88VosWye7JXTF1AxeG/TTGc3owclxPZAmFeNOKIt5U5F
uvdGNWfdSBAjYiJmgxmo4dWE0VesVa5bS8A2G55AtJuOmIMqpT1LIqO4e+j7TNDu
anQ3cBPM9gjmlJpsNzcUhF2w4eUgjcf4XoxH/0hL0fb3yv9OZx/XQwB4THz/gpqN
5a5yP5ZMO+yT4a/gNpcWZVEBwHNjpxPSoyEsAr06XE4BuY3XfYtoDJwXFL7CsJtD
GPO6ra2Qzt6oc6FQHqXT7xI2Ya+7QupK+GBnijr05mqohjelR9R+rG3Xj4TmaCj/
KxyOMZ8wCvZA2Lb+wiSbA7IQgtDxTJILsIZmCpFMRztXMAOX9qiz3TTO2lwBT2ur
frkw4UqA+y543oyhvxrQcbD2pD63qz1MWt/cxWsjZpByVIo38npDOcsic8gCboAj
CWctCX65PpV9BUDhvmavkzBoNN8bVe8Z8BOIS95q4kZjz0MDaCpqLu29FWtMP7rD
EYcQk5zxsmMrgPZ3H63WaA9aWub7aVNEpSAcazaYC/LBF79hvghGg4mKT2ctyBpa
fNeusHSZxgLNWeCBR/2s5oYBkqXAFJ8F0LfQiHgDMNe8sjbKmVVVdKsuu4V4hB9B
TctkPHhZmhUOEjfyD787uU1gBEpz7f3ehbTr9P0cULZ36XnuKVNRMLkSlyc+Vam7
WSt1MPKO4yURWBcyT7GPb/lfm2SbNOg7X5D+wPPuGNY8aMUgKRkQHm+HigNoLj3J
hm+LXDKax2wJMBRAJhijmpZLKHlgtFDMhUrerY4XCFelHqD5NXn4YqQ0WiSZ+QDc
MRrKzFBbWF1oi4jyGNrWwohCv2IpIjXBaiPn6FdtA6czSID+mFeAgxSYGiDWXvmd
ln+C5O8R88GD74/SsBySd2Au0+SGt0dRrYIHo9g/qZ3YuYjGZDEfVXTbQYGEiAoC
11rnz9r0P1SFgZIYmNnSddPku6IsYNh0MU4gNlZQq9PpMgTp/zFt3KZh6gsjTe8A
`protect END_PROTECTED
