`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QSazM8Qz3wnnaIDtnmoezJvUtF+YhEHe1HYitH+zvVrnclx638VXhwP6FK2x+nCx
CtiVZZhkO8MmtCV5SmXtCLmvFEMYFfCxKR7lCWNn2cuF/IsjoomwkCBYR/6TaaNg
64nnly2Vs2vnsy9boKcE4c6DUA9vfuemKrSPcEaSkzYXN4WtmlE6qP+Um0W71JPQ
WkabPO9+V8XbbHVH20KbjcJEqTBj6cgYWWR3H/Rv8qE12TS8idv821lCjnQJipJ2
9vxDpS8LSQRbRePTR6idgwTsy9sl46vl1fUJWVD/WPQkQCxC4D6sV2YVMN1ZfATT
dZ9OfiVWosly2mLp2XY+fAKz7b8y18MvjE1Px3bVBVLUKbOHdFxT826PV9Lbkv3F
ijFfo0/5YVNFZ0Nvhe1ggw==
`protect END_PROTECTED
