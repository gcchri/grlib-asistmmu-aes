`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WTBA48WjlO2RJp9rYTNYKGAsqFhef9uj5CpUFZ3NCp/KmKsZsIhJm+AqDoN/KaaP
N7iHQTEvJbLZKDmjqilE6+emkkUSJimmp4QVMZTuEHlW1LCw+PEPDu5aYdemeiwS
knYTn4vclko6Ck65sQncD2LiIgLwiv1wVVIV61vgMvBajf0w2TedN30WOxKY5gKi
COJZb1FRgy0vWdxY0PvquEW8evAoDNXQpb9h1KM725jfMgUlH7GI9sW+l7PMr/wN
rCtsXSnaNsxiZYR/3Wr8zUvq8wqXYSi3sBmpVC4JM09hglwxgoVFA+e66h7gk9zs
Zf0dnuJlG0Wb8B5sW+2uEALEAH8IugT6tFXFVu1YYjzuqaU8YsP+Toh2vSfM2lPB
urkgwYCYlqWpc3+wQ/9FpmAQYEoxzsvhmL+0p0arQJFmAF1Lz47SIjNVmz90Jiol
ryX21WJlO5Vqc6FV53L2HAObU5rUdjcXXFO6/vrNwAXu/JzYjJhM6svLU0npI9tI
LkYhSbbvwrSjfgiRWiJhsSAjX7fp1grsY9eUc6ptdE75x98M1Ld0sTMg7PzqtfyB
D9TCw6NmSHj+Sgw+OHQgqlW5nIq+wqgloB9TF9MGcZV7jRYcf433zheBvawf6tm3
F/tNAqCbk+ad53MgxLD+nSk/XyzYy4N++UOyZrvhrf33NQNYnf8jeCAdNng1ryWq
6LwwK+fpVTAAZuZOmHiDdwRRqVdDnr3aPVCPT+pkOlclbACxSMmrjbhHp9kusoYK
xTzK+P2p7z+hSwiErZf80pQY8ZF3VQHdlk1cPhPGCCkU21+MjunQRYYwyfICul6z
CiIgaUef7vctmOKy0ySQOrFrkho0djeJ8WpJcagbn37aZrD8dGsZzfYL4a3tjyUc
YQeyK+MBulS3CdCKWiEUKW6fY7kf5SMwntj4Vz8n8JGBLUuDJJ0I6SoggP8Ugyt3
iPqk77pQnfJlTPKLGCk4Sj6qbD8n5vL/emWPRQ4fDl5g5AlWsdzC1xW9GCig5k5i
06kxRZNwHwrYaum8avA+le1TDOnnTluf4Fncc1PMh+EWxYT3XoeEZM6HyOw9ecOg
83IDe873a7Poh2bvBT65Lf1k23Iwq4l4qdmX81O82N4mJy8XG/ZAhhehfvJzWj/Z
L7xwelb65XvgdDbbqa5ai5Qja/DM75e7pxkkX+YbOuYgOGOPVJFeiA7eQxHDC9Y5
LZgX+BvH+tKrSXgJpXc+FqY/j4tZ1QPrpiEUCWs6Yo+IFrIqxVZCqwwps7zCoqwk
eHS2OwDNghMHzPDuyWkJnbtC2wWN1Vouwb9hgT0fild9+1w+sPtY3T3OdCl1ZQHe
D7gdS4CddFGauToheJYp0epGTfH/ktpWtS+bf40gnVuHiA6dT6ZLshIL0R+tqx09
+pkTU8VLEEMq4BvFVdmdXFMZBgMf7q6xmu8Ormdo6twLUc0ZbN0cC/VveAU0CnPL
sn8qkbTqQFaaQwALhgaOC2LU8IdoDYumF1ySWiGbPIqc5UQ7TXIAQoHFc22z+ci7
HJCGXUXR2K0+0LiORnEhEvbkZ+1J/+lvmdmANxMg7hmv3Pi+oytcVYbbAiAoN0+T
T80U0t6HC9mudgB4Kiz36w8vuxJb36VTK0OT43U+tdNckQ/JHzbVgIeBZCJut3FI
RxAffs40KvySdTiQl9o65F0y+xqsWoioGTnMFntpC8g87C7mOf9929T2sjKerDFd
rhWbUDB8pHDBkMxkoBHZK3rHxunUqWY1t+keWtO1Sj3V2DEvSpqb+s1WNIkzFinm
nFsboqKdfqlXaq15lLqkmokmTPHqn3rU9m5BQLss6w+sPP+5NE10hURbT8vfsrw8
iaGxIX2WstzMS1zo8ueiM3r3ESJhCtZMGLpwjzhQPGuqvC9a3J43awR2mdCDihOw
0dk7K57TDUPdBxN5FW/xCnTQ7xIlXA4CoxY5gjP+ngl/7E2wMKrBsThMvg3kRLYY
Fmc1raQ8O6x8Pzkd/1qIAooq/Yp6bjFL6ku2DWmq6W8SN1yJBnPQSGDazTwxNkAQ
SKukHt9Q9p/TUFQJVs2TwYFHFI6IvTpS5GwjIYWWIGAztCToUTdSi1JGQkj0Wao5
vclxYMrn5saB37kfJPsaha4pWY8pXFkiQtDp+Lxps5fmdQjpGJt2BFSu/fSK4YyF
spHQV/VGmwjC+aKptD7YB6cPmdHzSjT+iOdQv7FT37FLWFNSrzbnGtAqFqz1eHl2
1O2nI908UMnpybpzJbdjHT8Zj4uiDj4x83gozhl1flml07+DEZNYxeZFeq2nVeDQ
IuNZyJb61deOQHI0zs+InF7TzVjQ2rMBY1SynuyL6FYa87SMRpRhV87chcY8yozX
Xpi1ZXQZH2aJ2Lg+HkVhavt/muNJDExTKSzIMRdqCnvnfcXCWEVl29Qq65irP/65
WlY0YCmiDy4iQ123DVix3OAFfaGlI1sj6unqaqdY3ONrYHj5t1+Hiyg+hq+TR8Qp
xKhM2fI9TrN86rfMgfMzQRIo5I984MKPNr5kg0+tFffloTFS5ainia2woR3cJoFN
1NkUbn8n2w4SBWPwwvPZktSrB/61Ci/u1eB0S+7Dh1KYR+dDyBk12DAVZQkw62+W
aV/XtQlez6uShBhde6aWTiwD1Rdep8+CH2RfI89Udc1pwdZJKYtdzB33TRS4TWUt
6EeE1biPsTOs7ST+TZ6cnj6XnwyApj7F8ZEskcWEPKxz4dF1EnjJeAduMwNPln25
UU/IafxhUQ4W0CC5Vr3d+RUlCPHahDo8xt4uuumKYAOauld1ruo2p8+UpM1eU+oI
uFbCrDtAYzvSht65fkJCJHzh93S1tm3Y9xODKGT/ENcCC+088idUSWr9T0+7K3d0
Q8LNiWjsaFxojqZtL9jsYCKeWmijWYdudt7Q7m5sncwFNjku1htrZW2RJVzVOgxh
UIsKb40fbeGGA2UaGHb+UtyBwoLiI0NSPxbothjnT10yXszVrDPAeYei5eyNqRL6
VbBKKAkTlUk6/NWRvMU9+Hg12BVlOLOyQhzZBiFi7KLA6csNX6pGYX5hdRYkCos/
J6ApyoKrzPzMpw4RK9Q2dd8xgpe2BX6LN24fitBG/pmOWYsfXx3ZEtbcKJ9+9HVc
vgoLzlAmSQzNdsHvx/n8r2hQWRiTrB4ncPVNFR3eFRF52ml68P4FIgb8hGXm7AQP
/obiwPz5cdPGqxLlJk/su4Zyal7G6P5Y+qJ2VjI6HlavGXogRwDNgo4ydnZcNgiz
BjQJeqlEqYbPznb4NLQGWcCHxZ/Guodc79xd07uRHucHL3IqnW+Q5rNaiBQf4IdU
DgJyJ/rCXbIThL552Fk1aBnv0qEqb6PykIwH5jFOBfAIHvsbtCEYFOaZWo8zDewo
S5aqsREa9m29WOeqjfjVNXZdnpzysw/D3d48b6iWeYsTf/M21snXjCTcoLuvT2ek
ouSpTEibHc9FuWzv6AiH8nx8lEnHxEAq4H9ne7TXm0+cz/HoN7cUSVEY0oNr5Tph
zyyhrVoCYnEM8vchGiQqxfVaFU+uSbKwzbJ78rVyyyIwdDJsjUOFheVo0saas9vT
pbCmZc55TVfmtFjglmByde3t6fFA+NHQ0GorJrjz+0lYkb52i/W3oRC5xPpahpIT
KsGNxxY8jsH7MiNUvRvH3RPqYkAQGszOcn1ccsGsSqJSM3liDCghb0GE7wwqu/+R
dC9p+6qAMxLr5F3NE1DXCSSBczrAtMqboKXYaeXqkayitHEkrB001tTWSpshXav3
b8zPfTFs4eOVbDaJb0jE6EqdPKTY/CPKY0te3arFjEXwlI0MFJgYKTjwdOmNCJ2P
Tz1qTJgJ30/niA4AB6M6TOGHFhmfzjF8AdIZN7MtjuNBUN3dAKBk1YTVAZZp/37U
V+NY4cuNcWQS/hwGQgpvZbqA6Zvuw834aMWL4/N8JPgZen0bPX1aLH77Pty2kBsv
Z4shGjihZEj82iQPeUwSscxnep4HD+cNPUn88lS00dKaF5WcCC6YBK1CehWjWe8U
sby60sbtdEp/LfN1AO8CP/bIOyN1Uxhpl3HqP1yzr1x5HnGEYqiI87rWzTgjs73I
NsDaGaS/nTzoNxt5ywNT2SDB2trVQTX/nVOS20OFjVeWUWzXvhSvfESHh/x8TEhX
tCmR8fdhc1FsagMN+h+ef2HIj5KiOvJ0u8QRrxWhfaxuoP6FI1QkdlrdRE/Me+nC
6NkoNX2+9HKRTHyN9WHNu2xT5X1U4r6qMSTB6cCSx0Y76PxM0dA0Aj2vLoIRHYAx
+xIKz/kaeSirLWGnqf5Xp/Ccu7b6ekKil2W1u/ydK7wwNvFQmtrBeQcgvjzZqaxy
Y3s56LoZuKffulKEE0LgEZp/i3Xn746D/Pv9X7M6TCYiyKdrR++WwfQZg1nW6u0r
onvlow+wSZK4kJTgddfetxnqmTuhtCLuVosczXYCYPqXzhkxn2zXyjuDMBheHbBx
H7anGaaYgv0noEQE59nRaViP4hYGN93WWZSKmM97qYNvV0r69wemx1wE5JMgQqr4
vPz//zzIx4xZTlD60Kg/xwkNPVDmlw5Kq9z+m4W9eH7J+LvamqC5z4Ne/F0es5Ef
h00/OjhZP4iXx3oKrLbourJJ7eSHSwhiaxLfxuTmnAHg+79d05XPpdnCk2nigB0l
WHwZgk7297whmfZdse3wgAkaGCdTezfBZKEoSBDYNLIha2pDN5XbUnDLe+slM/OQ
kMy5TcyWjYHZ7RniDqL0LJCQH58xqgLJqBf48q4SmlYQCsOVwXoCWtr1OWgw62oH
6/DZJ9YxzIKa3EILIjKXcjZWeW2tesPDN3ssjpzo6y6RyAKU7CkIBivnAu5EkhWA
DA7LLSCSdiTdEz1eXTMIcuYj8m/jOqC/sHbGOXZw12fcEB4lUNt4t8Y70Eh20ezf
pt9LcLkbC6s6FCex+KdBPXczDU32SQuesFvnyDeQWtgYB9tvg8lU8ygzPu1Ba38N
uxbiQLWpUNtG/yWH+DvWG2DV6EufBiXYtNgv9urZky8o5nv4AwgVw3zUSfcvtnns
XmmuBnSE420Q6FoaAvkKj05HiARHdV+W35ZK/6+pwYLn5F0oGx/likDCQS8dG68w
7Y9Zt25okXdtMnv4AWngABfcXLDA+pT/G443VjnbyxcHihjODV2515ngNTDWBhfY
mlYWkuN8LMkHLXTSBbF3sGo/LTJmbk3vGvXvK2Nej5Z6gGpd3JdBvaq2FuaA5Pko
1sL93xsoJXX6wbcsjPpnGaIP5sFDpcauPPsJ7r9XxP6G8mZ9N1TG0XwXuYcWDMNz
470F3G/1PnMug1ebrkHqS6OW8YzpLDxFmA9um5ClN8NvPwwSa7MkYHL5pZ3aIaRX
8/OPvbouDvmTHnnG1QaRW3F+v+a9CneIrxVl5li85u77x05u5uOeLsWOde9AIe16
hp1xgtG6UHzTazi5LlCHFee9leKp2LtCqTWFjhn6sVg/VWlDuDT1BityJKTJpiAa
Cf8gYkXjUaK/STixAm+kB3bFWxrscHRUecQyOtSLuYUopd6dghfBnOzBeGjmeWF5
jk5B5dwQqONfvScN52Etskx+xZbZ72oxeh0L6q04NQsctZ36vUhnWEkHgdXGvYJd
TK/14pR92NKK/RW8TzEs6NrwhmFFkMiNfGN/2JZsM07eVUZUfCxe48TgfYZvFMli
tCokaQMVLwNuEzq7eFZwjJYN61w9a8QpYlPSJ2XddjOLGIo+3fX8tmUWUPreFj2R
uw/KodaLjovuDYyuHH/3Rih9UE0cWPu/1cotnYOUpzYXTmje4XehTCgn9gdwudM7
KX1Fvni6tUMPjOgZ6l5hVLNnICP/GATPkADr1OD8eflJmz9HFJVjt9iqSs5UPKQN
+SjVSO20c6WeUnOgpJWhHzF7tyAAWVtRdqc7juz1FJB4dSN3Kdh40tCfcR1uY/XF
oT3Ce09G4ojNF486sL3S7bbEfK0klsZJSO+PMbe24XnymcbzkwdKmmrvwL9r1bWR
jquifX0lRMsJR/49V8QoQYIbFxPlfsleQ4UKnohXz5eWpCWJGBNocSamzs+t/uGT
nSiQaUx0HRV8q0XYCDo1J0ZQcVCgC+0KHICYuByFaU7SaNSw1H0ow/2At+N0IlOR
T09j3nQRV3pP0DJMhXDQK0SulpGMfzUbydnB9AdFB4wHXFQvLIJblGhlwHTU1lkq
uKROFBq9mQtPnMsmH7V6XE8spXgezkDxuKk/BOrjXJ01XdRW3YkE/+AIKRJsuhWR
k0smjA8keiB/IltXOdaZuiGytIorDMiaDYzdr6+LeFV9MEV5v+pDr7cmHXFZhreF
HfalUutLDfD9pRuL9FmgS8dZ/WLkPLHcrvC7ln+UIrqdz1nvTGg7lFp+nOkn7tHY
p9xAPd+P5Uz01di8W2MwNrHjvA5DndbBq/LGuWt0A9qG7QGCdRwgHpdJs0mY207J
xJL3C7do2LM/FOL6bPnMvvbyS/g8fga9EuE5Rd/Iz1mD8+vB1KnKUUNbfPpmoR3J
RMgLtI5d3TlSVmZ4EqM5jnJXy6NO4WHGWyteNA45rI4SaNivVX3MFo8r99vSX2bz
elcxxhkYKBO+M2EJbbvbfELCtuSpk086Le8Hu0hW17DR6seqy66NmT0bLSEdjDaM
JM/CNPai36Gaol0gpOeJEIGNIvvNbQmcRsq8XJSktJvoQ6L5pkIGj9qfra/NKAde
qq6FMutaJaX9vC2PTV6GUcnKGkgphiK3iZhqx0sV4NDr8CZrMto/6t/lc831CjiO
gbv4ppt45nQzDaKajwmxq5VPkX+eHouWLA0KzkDYbFsxonS7yHwO0MkaDOvKMBU3
gbcgaUlbQCKIE+nJ5xXfYuM+GLts1QOpCkHn8eEnVsWin25dRpknu9Fruo/SN2Aw
zn2LjGwqEi0NdCPTs02BQ1GsP803Mr9nUtNbEnl+tMB+CG7zFn0qTVji6xL/pirs
ASEIRt3eyhuIBzqZWoYcdHlAFsytT9+ZlyZAPIQkbUCHQutBIDso39V2nTs6GThB
2n2OW01eklUz5BHR7JyTQoJLYm+nUhwpl9kFj8rbeNAoLI9nUaPeHWV14EoEh50U
57NummHqW69karguVjp9cRbR8+HLkNd4u9DuurM9DbE7gpyansdENHYhwn7MF4My
WGFeFd7XoyrddMvKyCLaJzC8Wl2qZBjmyu9++GIJidKZtspFBzAV/72WV0s/TOrm
IJ12ntXHBNzVgxYUFdnqnT6VwWADaNcYwtFl8jcV1IrxH8wkB+oggavQpYkJokJ7
3UAeJnLcZoAv6XWt+KwLUuUDcD81xF8tPEUU7s5XM8VTfO68JSLeJZKK8ZyFqGR0
+nm5kCQsVNqyHlI8GaRRapKoi7spUpZltSPcgNYCKIL6kh+RZhbGjWvfgyowolVQ
aLLswpr0i+fCeqzWTbZmQj5aDLDTrJJyhl4H23BImy7AVOR81MVz8Ah5dA20efuE
bOAq9Gp1kyq4R7zFfTkzUj43GCc+Vstr13FPY2ZSnnFEytYAvyoLcUK9WNlu/Sux
jTPb+BMjmR1QGr0cBaqI3J6RVgD6O7PEiYJYd8W/BUz+DQ2uxtwWnah+9RekjAFh
x0ohPzzYpVLkokTk13PT+TpgQTSHaOjgn3b0w2B6PXdo1GFaeH20jfpPhZDim8Gi
ANkrx/2IgicS/WqJMNSDMeMVCYwY+qzXQ5OmKIQ95ARaD/N4m4FVdKjHdqDOE9i1
rLKfAki7BlYFDlv0QBajxWArjOqpXuxdBONvyos9+vRr3ZCmLlXqtkVlZ00M59PL
MldLPQdyG6b6QmLS39ERL494foKV85OOvZm9EKeOdRew3m/nd696ln7F4qLbL6JX
2spg23j77UEld0rl3xA/C3s+43lU58o6yosFuqtl5/8//mOVl17fGpY/hUkFKaMp
NhimLUhv+qU8w6m+AeGLd6p+gAcVM3Tf/2NhEufvqcPVd9dAojXu99nue3x5LPGo
ClAw3YyyDuc/hHUFnrZlb9eytLuMI7tLv3JlOoMQHfT7GVfnLbMlquGtwNZf3OhU
sw7bcgzXFm0RR6tEV9SVBqb2m75/aKiwdDVg4DnWnHzG4Z1beqpiWGoTkPS3JJRT
a3zcpw0nZa6ly8u7HJQwu1f9oGmXNrLFegTA36Hk/xjn4Bj7pApArsRSM+BJxjqs
deFKbPiaBVYeRz3VoWmkVSXkMSDZMCnof4g5g4A902kMlHukLmcVV1A0mIkro5iZ
hmRtfpGQEprjni4imVrbrBP6oFWk1DAnbxIihYwrmcPmh/NiNowcgeR29o2kkiMT
eRuUU++tUdtfG75J8CvvmvM9V+Nmhg6okfFobw7X3VirAqySAyBKAw4lFSWkoRwj
Kilr9MxhDUcy1pRiyElYSh4Q5YBHzUsCKqM67dSyYLHtyNh+pkTjibbTpz8CatuD
UvaCojqDKcvSAPJjpdBMgEnD57DLn/qGs6etHn9JhgvO9Z/o02nsnJMysN/+g8C1
fJJaiXm+DRfSBEclSZsumD+ZSHLGS9W5pKxOJRPcv+nR0FIy19pdvc7lEX848QeL
BIQNUDXUkX9gvhX89J3y1YBgUNABy/aPU2NjbslZ/wdFJUpUwtbPIgRxW7Zwp0Eb
8eNNQrXAIb944TxFS34zkToSnFuW0vmZORszJnhdvrJhH4dc8N1HeZSc/xgDPjux
hu4AAacEXdIhlAOPMahsUODErr3AiS3ULzaOK0+FyacUow9RS7Q/DacBCRMbehdz
+icgmv0y6MooxtGJOtAluA85Z3GN4Yv241zstVVDeoG2UpCHe417O7dNgZOLuGO1
hbv/WJPWJPxu8zf2umGe3gt9GUjxpjUK9HUfQCjXI0DqYLK/XOIog2yukVLzJeqZ
auJJdBIlMIpXcV/2feMxRMFZKW1L/oW2wydP7Nt8Yu1sMdjuchmh1ZhwqQzdwKuV
dGrvHHlv4bcSVIGUR4XWNLcsRqE1xDn2BWTl1FwdPlvRaJW44Ggd7xzLulT6t9XG
Ge25oqOwM/sbJTvtGp2YTZdJgFoLD8Z7FRq0St/aK77QbuL4vZT+X+i8iE453i5N
WPYMDvqf9f+7WpagPQtufcNEp5Xl39Ar9pGyjN3j83vcKkCsQylXHi+rXVzU1qbK
mQxdsr8e5iMr+VuxpYiS58CvLdBW+yhlihKVjeWshbLUUlHe5iyvSPdLLT5ONmH0
EuNP4lrcQqwl282p0uW7D+MSjEGd7gCQ+RfT6N9LdjRx4oQ4PZWw+WfgP0bdyd1M
VNaxk53SIBiks3b5H8xJmcOd58PIJgOeOYA3LTV3PbcA3h7oRGlkKSV/zbKgcyYf
ThHDxPPOxqbHxqdIPArs9OBX0KwwQvJLBQD3hQ0tCVFHkb8lM63X+qUUl8rUghsx
FFPAkNDL5qfDdjPOl5DeBoG9BC3aOgjShPHnz1ADGXcBh+Q5efFMCml3TfNIgsZn
Bj1oesyhaPPfbolHRWySH39Id0ldsyw7DtAcV53bhhfMPI7E39IJlmGI9ZuGFa2I
cWYzemI8RPYNIM1fDZwRK99znkCCA4kxlbe/RYXnmkZkw9WTPuXlARHsIXIfyLpS
xRoG6GVgiP+8TW4xVCYVii0QSg6TmWI3AD2HjmF9bDRi1JEZpGScB/nrYZ4zM7sZ
8FsZFWyQLHSsDjuuuiFwc3tyv+NWSyP2pOHlEsDn7wsK5frOyyg0oPvDzvain4nS
348rGGXFxwcX/gFjPcOh3ryPApqhq/hMzYiFkbJH2vwHW1AAXKo2hGv2/oH0dsp1
W8Plxga2eV8rFq8PG+40ruLXbIy1dHG1WWZ09Dzy3fPQRh6MWQb5Ak+J9iqn25ER
YbY24uEn7jtkSUQAp9Fm0ombxYOLuxvBsmI/h2oL08UpBSXC+trg/VAIww5jRGWI
+TlXjvU08xIgLsGg4ebOIW9CZeTD36R0d7amD3FtkaB45VGpQ4J+Wq+wk5YxMW1Q
WMjuyvmhe9YB917g2cAM0FIE+QNOUtXZfAqmwoLF8VwjnZ1mm0c8WT4K0q2WULaw
AtgMZ99vnnbC+yM/yv4FGEaUm91TksdDetfF1+Wo8xV6Kkbw4Fd2K68xSOA53ZB6
N5v183mdfag4zIhrRkQ+cy1uI7aGH398qaTQuOFbb7fKB4eDEbrJMYriZcbOyhTb
HWGfVKoK3tprMRsqytaku/xUGY50D9c5rb+dD1Ejauu/B0kacoglmrdtTl5yKpUB
3dOk3g1SGY3wQe3XfU+4sh1q8pnRBH+TC66vyJTHVJbBA6lyCwgH+H++cPKgQDu6
Ah18PTAkWqJzn1VLQ5xjnlqu3MAbKe2Pv8Nlpyd80x7mClR+1q3AYcSkPOAlQJvf
ueu/4L7kXl9FrCyc34MZYy4tS994sDlEyauwwQ/0wVWHrl7xB8wJ3Wed0AhHVZUi
FaGt9lGVQEf9Ft4h4Ddko/dVlF8FcBjA7c0PWK1S5h/7oUu/YfuGvv9+lMwsUqWd
rfunA5Y9UAO3RH+b8cvq1BUpfa7ajPzVgBa2uTaJ7clOEDPXZrbzBRN7zRhfCN5B
QNFv7vNtQdA7ANreYfdFEWuCLmcTaP6utjuQfRazoCRQ177+Lhp8yA9+e2jSZy6C
rUpfAu9TGoTa/YFKZzeJjfygDH22XXNXgQzxgZyyh5hHCkQPOjMT7WyECHHiThWm
pCu4fKRLSEWQTBL17Jy8T6Ayl0CqTvnUacLVfAb2WGhV5uQrPcKboacPwBRabhnQ
ebAln9hVwKBVAUNxs3hx/VEx8bZSUeFOeKmTyHNaeKHar0OFUnuS+tnwjMrrQkT8
QDcX0vFYRDd1r3N7PSY9ytHJIo/QEs87nxxh+MLKEROWNm0Nikr/PI6qhxW1Ruwq
akUPvdeXcMXTJbFq4as2aIkMDRsdg085HkJ7TRtpG85Qz8aVjbGOD9NOPWuAAai3
QJUJQSq6bj+uQEDh0p7SVyT/AqgK2IxLxqnVaxICYZVdObZKbFq9dVs0kAirEdz+
5IoXYG2QQOT391Jguawqx0/he6qzv80pFf0/nMK5RuOnYzl+p4gOY0EEdooWxEUS
OHgI9nA1C6AOnkaO37JypglHsE4wPP1Ow3ue9jSfi5cYuNCzLONXg44OyH35mxS7
JUky8MfG4DCMEIkJLCKNej83r27/QRDUzQPCCvwEOJXN86lpBG9arlgwURP7ZBxA
S/oiRh7LTur02pbtCh4Dp15kvJr0CbpkV/cFzq7U6Qe4mg67VVOMHQjXktoVTXfi
4iHh3qav3wFwYCeUKcY6XUApVjMVRzBulLeKB3y2ot1arqUJqt+3utdvMAa5tT/+
VuszmmdOfr6vzopSqVDXCILSiFYJ6iVsQsLJshAIzAtSKEzZPCq1vbADz+SK84bO
iy9GTFDx6sPDAd3TIXTHhk6zFJa2JRXbnf3MV6p4syxYE3N1jxxVab8S6HmR9nrZ
UCm8BbZACrTmd1Js6/LUCkKEp6D/drwk1R7zg+CnayxTubGBiROy80+BswAcsJRo
mLNWCHrMxXdz4JPwW06AdPL0/HYEcOQB3B8A3fMGrLhuZitVdUmhYxzLmKhnNndS
EUaGeNU7VRs6PYx/ZzcMSb19TktUeLOae8XXqqKeZ/lswNcrJPyTjqJCAFGB1EzI
/CAU9rtcfhhmoDnqVJ08nsTdSQ3OQppJOtg4DNdx6171T31vWM6aCyEs274SGIIJ
BJacna7ySxoLv4OeOwoqI3PDIJtH2qebaHjWi3MWqlII/BMb3mQtRVJbzz5yw1n9
KR0jU3nvrv//EwzSmvvNGEbaK/DU/1LwE0JQSXNWlDB/Avg1Y88nEfxlgb7p/GRy
cScjPSRGO9wZAsPgTBDUHv+xIQF/TPR88B3ccfEcdmk2z6SprvcNqRG6SPRMZIfc
EX2Pg7vIWZ0pQ2WwVTDNjIFRe8eXObVV184AS2OtEjNtny4LOqT8lBOLqpg316bC
Kl/14Z56eeJEt7itJbo7WvIeexbxUsUuWilUwOmku3NoSXiKOH0iynYku6UMmpUw
C5mMcn4X2k6Hz90b4U7ZbRAy5P/UStdkhBoSHkHlXdNwxgPeo/j2I5Qhk5WOAgGS
n6V9gno/oeCU42CSUDdVycejS+DSERCxjMBkMwhgerTGBiAL5ETx6vNmAMrJuYXX
+zHu3xP5nJP53419z+rcRpBw2ZwymhMgkc6DIgLXmPHm5ypaMRuFGjxmGR72hgXd
PSgI5d9v+MHdTHdRwSFd5COJnmFcT6kxTgyipm0mbe1YLK9aNs+Ls6drgqi4+tV6
w00dubRgcw/8doZB7abe6Ap7JfBkhIamYkrPqSWzF6AGrHRhKBQcYbWqDS+z+1yU
RuxccX5hgEhUi5e4YQD2QicTgWcZ9225qOgYJ6ThUMe7F7xQZBtKhko3Sg8e2x0G
+zCKwGU92GvHQFZLMrMrCMK3ZzBd3bQC1d3DVO8G0H9CiZnLh+88qo6nWXaT0cFX
Xv1qTTPkMvOGzjbHzTcxz9595fJSpY6PiUxs8g14cSYpNFCcvvCSVuZFMHRntsBA
K16L6sn7rDdNfN2hJpSkEd2dbYPZAPQkNuaL7bjAlV45gsJumfcpV0VP7njRxMBE
GiTSA9BgYmWE9cPoac9xLV3v2OMDfh9JD6cPzPtCzB6FQ9lFZYZOAXQhBuqPYaOD
zROxLh4GGZecsn4pNGdCMZ2Y4uPoHiLHR7l88u3UUP4RdtcHiFeI82QpIVk3hJ8b
LwVMZ/Z5XAvDzrae9cFDbPu+laJOH1YmXT+uOZyyCe7QF/k/jQQe4UGGQAtlxld5
EJLd07yThA2GgjnYQCK760Ft05GHGM+IL/GJQxQ2ll8jOfu+tPU/f5xjPZ/4zf6k
Tsr5smjziUkjmmbXvqLHyzAli7FWWPR9EbtPoLUuCuG2F9cCxwe7E9XlL3XSi0ls
WvojcUjpygZaDkJ50nYY1oGRjobnE87djsSwV6DmHOBuIq5Wbsf8G2ED+FcOpJkt
N2zIhTKjKZLboWh2EqrQuK1KHGU6umQV7ujdqCOyj1dIm0d7G1fEXltT92ph8Fcx
htJtvmyLTnug1sAutkR5/6o9BPqCHOhOpQ2yzB5jhx6bITz9ueWVRCoTD1iNZUz+
keDQdrGpMu9lFNsjLZU34fVfijzuOWhMW81vZbgqDdk0hQcx0jRquAGMK1J3dajd
9WjOZ2V261ZLqn/iF87k7qsgIEf4nYjEMLMYA9gtyaOHG7nldl+kcWX1C7i0Ocf0
DxTY41MpXBiV5rs/it9Wt2eIJB7n/BCf5xSNpO/8sZ4gWUk3QC3/AndWEHHQBsfG
KmgFX2fZXRxiBQjb8yDdzA==
`protect END_PROTECTED
