`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uspWHGQSdYmOl9HMHZiOMK3hgglAo56cxRpnRekByizUagQbSW7lZVQj/ub0zme9
D+siqVGIfFsj4569fWx2nhnfJ/Wg0Bykzb+8UqQF45P2T/Og3DP32OeGUBdQslAp
oJ0p1/TqnRhIei6kWTE1hsMme+EYEzR7ICOJ2AeJTKWjWXryXQ3MvK0VfDebIvx5
VCP90U94BXv6X8DIkaFCVrRbacq5YKjNSWpwkmvpieI+HU7afdjLqdzQ4KTVWoUc
f2eGWNuo/9jiZZy9TH9i3lxYCwn+MFV+eFrny8SjSnwVL5nF2x5A1RreSdMP0cDk
q6aTkbjoIQ8xLgfBvWLSb/w3DIh9jvBZDhRBHyvcfrhruhSqZ4ZuHrKBcFyFbX4C
m/hZVNtS7mTnuCWVJecvs9Pwve7UcSMvioirEcsVNNzmkZruJEMJUHklpztkm1ub
W3PKN6MEgGppwG7pGVJQyga96V86CHr9WwxdHxEOlvH2VWMGdmlwjI5RyVU52fxn
S70JGDFgOJWiK2nG1wOD1hm2B6Zi5oUymU1LDAo5l0NVGtbyWw489pWkc8iN8CPn
8MedJL3Tns7CmFrek6rlPUNjnaD/4B3I279q1nBNn7nlW3zOqKpH1BlSnNldbAAV
InTHK1QTH7f9kvqqcaK9W0dw2XsZb/XIaJI10dT4SapNMGubScmi2nQOHmi4j6Qf
uWWBReaAsZ9JXw3pmjk2HvgDXDLrWsJpQB/HciuHCWwt5Nag7bXvksrKaKndX5PG
XODMs33ZLf5t6L/R+Y4ZjU1lqahtTS5CSq4JCLNgDFmp8k/LmUGAr0UxNUvxMIIn
yTlxa3061y6WgV6NKecJHCzfeCZrdQBUw9xNEmsCBGtwB9IsWWn+0POR0l0RB1XG
MCfuFcpErYUYJi8M6fzKgjuuO9alusR+QQnhV+hZRqFfNN47hJnamnVjdM2rxLpC
hxYOsDzS2zLZeEhw4prdy9BnejUVvc79jy+jw0YHb0aG2ozSvsnlehLuaD2xXlEF
Ylpjx6llI/g99wYG3wqT+eb76QbODzDbjdf9L8ann7TMRlDTts7ghVkZMc3y2inL
yDQliwEr3cMErux1jCHEkc7HaTXViSvQiY8ZDUbvcXoCSRDILegynPHGqw2Uyj9n
jWrDwatRlAnhOGqbJ64FNVOdhtjoigCbK7EewDw2ocPKe4lFNoCWjn+TgWLG64/r
kbslbZ1lqwtG4lNN/BKCP5DUWPC2bq3xxAVI4C3Ld1030Z5EY1czawESjwtvYAnR
`protect END_PROTECTED
