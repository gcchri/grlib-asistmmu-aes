`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T+QqrhAAIbpF/3hSreQ/nKYbD+Xd23I1c4G+uToRuzjFUbvevzEWmWcN+pTTemyk
pEQtitXCxNdhJ+GAcSGKz7X7up2uMciTtzOJ0P9FpNiOrjS6lJB4CW1DpsrJ1faQ
dTbE4TLvJZ7XVQjlJP0wM8uZ39HGT6xPTSWXbFA1jxHJ/G2gbLp6LGdlC12KYudL
gD6R9eWqxeRlR+VhJIZLDmFDJ/Fvg8n54ooVwv293fKmtMHqTeav9ySP+1fDoWjY
PLvAVvzI38jp874059/blWFLBSmZ01p5ru4cIGBcJWA9Z2erWACE9p43naC30I+J
06NkDhgTO0eOZDx+v3zTf3LY0CvgRypKAVeOg0FK48l9752G7MucoB3Gqbh6VWvP
7wPINLsgywgLmmzSZV+WthLLc+Bk1VS8ISgz8CyLiqTljDVyngzNxCqu2nL+wAWI
epRGXXDIC49N6t5xsbIWDMDNEivGeeKLXocVxI96fwbqhSUTub6ZUFkXd6aZL4NS
y+XGN1iFauhNB8O0WUvjhIJ9d035SAmDKbjIzltG3KXWVZZqSEKFSAd23dmFMZh2
LJYxH+bsaUIe7Wsw80NHgXLJaTr5IPEhFkn/Tp+yD2bFyDm5sP9tiKzEF/Fb7ovT
eIHqhAmQL7u2uo7nhnepdx/ANzAJCOYHe/8bIzzASLoNNdxB/f9MpsS3vtHgJyER
Kc4TfydEzsbK7tWyBaA6gWCrG15Cy99GQXd1EiZpZjeMQGTa/uHeBrN1F8x9LZRa
QW1At0skjVvceNkFhRm3Ny1dVXmm7+cyhd6qxOg2liaQdXxqEtEWvs9UK5sNG/Ov
nvL8RukUajjHWJJhWcJJuuHwrRiRiS7L8a+T5tMqGOWt4r38D4zo25GpoJkwhfh0
OpSD8lskNJIdG1bGGAUzxx3bWT96O7XTvRQlcev9w9aGTJSQOhaX8C8iB/5+Qaj+
HVBdSg9jo9hnUN+U0E9w+IyUmDovBvo+xTA93xTg3NmlodMZG9ynzjALezS78M30
3kWDsQB9O2/FtNbz9SS3MlQucGEdwCgAqU1SNpUac18PKs9q3Fd51Ln80XYOFF4V
eClsEnrq8IMQvbtgICx5/vMIodvJNBQDVzgUM6U/QdqIGK1e/cyaQG4Qhp+F0MPj
v7z5BEwjEBqrLO1bBfXQY/aKPDH/8+anFhU+pFdbj22qSSUYxVKPE17vRT903AYn
ft3CYR7ljunBgde1Xu5kdYuzFmNOw/a8WFWdyKPmZC9bGQqbXwLJRW/u7ADK0NL4
SqtFPrk9RbKn2TSp8ZACIBPBx9MvCNrlTfuzVcxQ4+soBhSXiw4lvbdCUj1xNKzo
Yt8RkRmjHIaluU1T7d6/dyG4SHFXiU18zgBfJl471eTl7hoiSf0JQLKbO39sy4rj
0ws5n7ZpUtgY1xTtuQNWRPOC7tPRE/qk8xu/Voky8Y1SE70dDQua73HmEPelrrE4
uC3rXeVlxH+ZlQmg0xfp03ETDMbTib7MUzL1GJlQmaKrcaDYndVuiUNig+mnTaGL
6kYjWGB7/S4xLlXYiZGrVW7zNM8f/4b4x4Ofv/KRTXC7jBUI9qw+MRcy9uEZll81
FozyCfRDYy7Oo/JKnsCpT4NXXycUo2v84BQUnkuZM6JdB8fiT9LuoKaYUH3ww5wr
AmcuMOF0lWR+aEXt4/lE4nAyBNrRuPjRrsOwlK/Ozuspu8/hu/z9HgJYyTgBljj7
DvjR/Ah9ND0FY7Up8om/G55qRm8mmG6UnsjR4rX1Th4bWSP+ANg0aoqKD/+VYcxP
xU5d1kA4B726Xb3UyO+79LpWcnRchTEx6kV6z8y375fhRApI58ox9yBOfrkGv0yz
6XbC7By8XdCx2xkLPVRmIUWxlZECvFawG/03O5wQOpODFQlbHYBOC/pqCcGdKbwT
a4hfyXDc2w6XTs2TTnKLmJ5L4Nlp0k3TmHez+nW2vJbYnqFWZv9619Yr5rZxgLMg
xxsr+LXD7EDAdXWzYSbzUUgt0+ZiqpTee5x4S5/leLIoRUH4U/pEAzyQQ+ElA+Qf
CF8oqqJbJoRi1be2ElsZSZA5FeXzix2gw8D40MpFBurC1qgLLMeGkDypmjcB+0BC
gOTsff2ZzMCtcvk+FarE/MahehYb1TuThTlbFL9JES+o97HJiOjtxxZ98T2F6TrN
E994I1XMLyEBoqrfqRXEjTCmefgAQZEd/QElnLFqE6O9QNTLhnAOT50ROIYTm30D
YQ6hqp1wDF/HNOrf4B/LTV12RU60NlumXwHP1qKKIK9KScB5+KePM3Ar6PTvXqls
pPYLTkzQUnA/Tsabyuzsir4NHr2bc5FbZzngi46M+5Msm+iwKf88K8Y/6KKbZJxR
0TGnhkSigRaOhrainyHwsnFHIkHB+ETdndkfIfyo3XCLGqmjqTzPo5SFKL8APT28
b7fP7Nbw2Cyo4SdZnd+F2A==
`protect END_PROTECTED
