`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DPnq82V4MPqDyQtJ7AmrYu7sKGGb/bbVKCMnvxIxBtfvZPrN+0CSl+psC6fhcTf7
QV9Jpjrvn/Sud9aIvBFVHSIzi46kgUKE2Qr63LI0Bx7GDpOeBRU7e1Ur5mGK6irl
D9WmIo8eVxAlLv2FbxRN7Yjxzyiuv9/7VfCrv4hQPqKTndINjtjDIuiq//r4b/WR
uEg/5i/oFSOM2AGyTUiVeNYl2KfRf5ghbJ2AcZ3pmzVupekQzs/nHps8b+fLspR5
0LZjGPLojjR6F7tnv0uIh/3XekIctceLOKZt3252av59PwWlyFLcAV9ZY7hMwvEo
L+nbufN2tmitsUHsgE44C8mDcKOO83QIXeeScSaL848xx8Vwxcl+7LUOJGUyS8Xr
LfPssgHeyCMrd0m5yiz6qraxJJJ2Zc+N9lfIFtXxOTisn0UERY8tVx49Nbv5o1kG
Rra/8MSjaeI+IGD3Uu5u92f1cbYhPq7GLW7vNV0/KVc=
`protect END_PROTECTED
