`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dzBCsz9+cObIMzrgz/hGBhy8eLkj4GhiKPVg0YODFeSZod3lemVxmCMQjOPpRBzm
TRH39SRL9cDQQ1kwYSoNkCKhvRnWURGT1J9/zYjCB6JrVygUXUdRTTwasn6LWIVq
U0wj9L7xPxYSai7nr23W4OpZljOJUAv9AU0y/gWGAIO7mERZ96xis8TtZ9LXXSXg
wx+lXKxQQHU8dHZKSV3qpxLRPbF/4dUsZK55MQi7shyhXGuQ7jHoY5cbucNMqSYS
okXMZCTMFOW6KFchoGyUMhjNxg3qPb1H0YaSw1ARPcHZjNjIXlvYtMWyuhAnntR6
WOuu8tL/yFvIjBDBS/RB3w==
`protect END_PROTECTED
