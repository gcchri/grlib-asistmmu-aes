`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q8iEkkRRhiEFQud8WOPyNN7M1Zt6Cig3ar+SGY42JLB59zumHZnkVsV5sLlWMQaL
PP6TzGuwjNL/P/eroLUupQFsRUMa9spe5cP/3KkJMP010+rwdDNExRdJSGGzjNxK
HQwocrtNJYVoZncOICZYSJ8OhxjVhzTMV9tPstIVJeAxRYqFALmvn7Yc6h0IeLKS
XI6cdUGuZmwW1A5pdntGpoxWAsrZFM8xRsX9Ht50tmdWh8BN1n3i2In8oOnSrzqm
`protect END_PROTECTED
