`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7c9ZSj4GS6GoaUUBl3PylyRDbLElC7KZ/EmxyqdbmdDxJShBWDpppZXe57yB/RtS
jdqp9QeDwfUj0Dm8e4CQMDLxCe70xqCkHMqlOrEi2Z/kHCVF7P4gri+G9oeG3M3x
fN8YIowcuHDTOPu9cKgwp34NzQUKyU3M0cNc/SkREOUF+JGz5ryYeN0ArlxxvhpK
x4FTwy/r1OwBAWmMuma3LhqmWUr9AwDmtISTD716vscfYQ3sVQ/nt+kbNClkO1S6
P13EZkL7e3lVzD9WWMzNHmQKquPpi6nZidhLpf+Y9IJwCJpIsHojR1wSOGWt1pEQ
N70pSw/DGtWIeqfsRdegbxMfze4i6/b6mOMeNPFvuFHB7TIcZl7Drb5iQyafyDix
s7MCC1VCjISo9zo/voLWBih41pf7nPyVYRDtbaTpHIB1rX2aK5HpqDXd+TcP0qTR
XqgFOOuzZYNw3mn9usI0oYIl/091+8J7W8gUWbb529hbAWfl6R7GUD6LB7VFhCEW
qmOPFw3RChdzOX/wPDwdlzozXERQHhWlbB/u/TdYneaOY/KmFGw1GDUbd7YqdoZZ
/zZZoTz+FG2bKW8xInaEYqsDlPlHaggYPXHIoslxNqZzyKIdM8gmxRnDkOdRVYCw
STovCuboYb6VdRDEV+2yw+p92OtCAESkaXs99BbAzjKDf80yfdFItJnEctiQQAXa
tbOGjp24HW4X2F7gBKbSxYi2vD7f2o1nK7VopdQ/KTFsJmddikcyilTvG6fg69Bz
8UHgGc9LSltecv8CVAcXTwhtc1SEK5bpevhn9AwFu+gjV5zC54ocxHTL1G8Kj78w
Au7HItBkUpd159t2T3bi/ErwXChSo8kA4qkUQQBAr6k1d4wJzBU0L8uW/3zM6CnB
q8NAe8ywdxyNeyF389O2yOMkwgAzfeGvTR9N2Ibl0z1yGtJAc2SeXLreMTEoZQgB
A+FoM3Wn+r/ZxUfUiuweTVS84MtirOf4zS1o14m+Fys=
`protect END_PROTECTED
