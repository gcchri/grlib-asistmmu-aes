`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kepcaO0sFUWoBhi+hVUXoiKZf03gSR7h6+cBI+qNZ7FF2raAKGG2qWfgTXRmPSVs
Of/SJTEsOj3ScUTohsMvV00F3mZ0An8GytkxIEZktG0C/uSHTBlBdGnuqiEwPs8H
GuWg4zssXhGer3SP2JbIaXZy+CyVuy1oTAWrYGOhAR5mtQz3Nq8cRL5vVKKyDbTL
1d0yyrSLxnFPXxFJea7QNGAI6BIphAyaQ8qsrB6WYRnTs/mbqJPe96kQ3Pfce8Li
SIh/8YHuRTGbOAGlB4QD9aUwDX/9hKINYd6KQHYVCDPBiywluMNbmH2uHjm42+JC
PLMSBrLYwTsp+E36r/dB/eZ/cXV0HzRda03uxIPuH0Lo251yFYE9W3RyzHzLSfVv
`protect END_PROTECTED
