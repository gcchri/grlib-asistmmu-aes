`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SotPpw6gBbuAcfYrGXcKYoWUg/9Bt61tqEnW6MvwucG7KrMDXUcGg6wb76M9tzzr
SOPdx3io0JwTuJW/H/9xzcokMghdhae7hrR4KI4VRVp7w5E4Ote5XMzpAALEaPP2
rV+fQ0kUWNs4EYE8HP3zLvkgivYht12CuUmEJmCpkSNl5w8yZHnjUJ/Bx19fNEwE
vvPoUGyJnbvhRIiogUDUxXFR3mwMEWVOBhxLavFAjBNCVeqwKVwW6oGaoMO/K8xw
1u0Krm8WAVx3G/HbBg1ILrJpChVn+v76WH479PxuR2t41mgZeZ2n9iouqc4FypI4
wWGJzt+EOeq7TPa7q6WP3IqLyzbOEQPJfQ8HtaxLCsJFNEOIwWXCaap2sVlDGXBR
EgGoMjjrD0LLa3IXBcU9bYf3buJkZ0NCfsKcoiNzuEfCGF3YvRvS/E1Ttl7vSXSZ
Z/4nNPZMxgbsUgcWfGCGW0qbb3LGyJmWsSDET3HM0VnPjKAtKQMIk29+GgWjGmOc
jWNr8ojzXs8RqIYAsHdV5dzTQ2f81J23vpIyAg0uboFtiiBeMVNi0P7jxXKS8Ykr
5fh8YKqSNKYamabm5VZ9Ul0ts7VeplnY534OeDywHJQF1a3nSjZVPlwOUagKUsAc
id/ju9afdpy27hAVWIDYbSz8jpwmo2X/nGtXoUT/BzQcslR7qvF1pF6CX2vJ3M6/
s53yJIH/jFEbzs0DbH5gzcvfJexehp4p5jPVnOfKGtQTauNCLFcqEIKUS3G5q+MS
Vg7IpflfxINy+JtgxNlfQrlWsMRJZ7k/ALlxhPA1+Md8EBAeaGii/BQUkE2Hj/x7
OXOSQr7pcor0Vgfif6L2HIwpHynqaSHRiHOWFE5U73KHcF8sq0rUIWinfs1cEP4+
TuG/yaA3neuJj3Zjtjm3GcOL6uAqaCnOqWzJxsDn7UFCkVOwfQHAd+fcmL1ywQ08
fYhfWIrIb8v2hvb2/lQVqR2ohmHz+puV/48w5E21Ez47P7YrQog52VH+DgRuJK0n
3SRxVAxbyW3rrC7fqhRcmKpQZtzNxWveJPB2WgMKO4NX14ltSOkJl8tA99fVLmHb
86wjlpXjwYGNA5MI3CSjv45IRuG6z5TWKGKIpJ7Ka3pr/0hYlIlFiS9l3AkF8oip
ueFQbuyxfSqx5DYM8ApIpQLGSJseFketwCnVJRNEH4R30hgX3gw4p0v4NiMp+N9R
5ON4NdDn3jaZ6oVYUTujFzbpBLPkHkIFVI4uQzQCArL7kZyclA388R6Le9JoEg1e
tjqHdqWjINngvEFi3smpz9Uuyddds01WtkpsnitjEbhu+BO/ThUgkDO34L1pChI/
6lluKr6XI7FwM+pDLUDxSehtfeZbf2giu/sUvfhSHL9FM2GOX+xVI1Xm7GhhDMIp
GL6n/R7+APcKfG6k92+tf9TvXNVD7AKOVAr/gHfzYSkaZPaEmaVvdvBBHVqnWpnj
q8mEDoIAaaPu4Y8gB2FPt+Cu3cp9qoBtLqfdS+MmsOyA4CA9gvCfDUGcguMK3B1T
Lb91QqZLSYcIBUOgMSUMvAoQsuUSNDtmveQrw6kpYi/92nmWCNDzsNJYKuSMsTmT
56EyFEO56O9SxfZ6RnFIhLWU6f2s5irxD76YdUIuGpyWOie+rPeQZ3Eli9bMCu4/
eih35qVihzIZ+cVZxs+FtQ4BeAeSyyXnHxND/0HA4mjLj3dwYLVu9FlsPM9g1BYZ
f9Wm4OeiGtHOQliW0P9qowDlzpnTgaE9WKYq1pkevZ+VGg0thB+qUtqbawWgfV+P
C3hehXkc+KasCyciRtzjZEfzmGnDxOzm0F6p+xiQ+LVVYGiqV6dgMGi2rzVaShIx
N2gBB8CqZ7X8zUR2HW4zMrbHAHXZmm+ko8zyq7DwpusuDnLVU0Gf4SoiAcpRy2dU
3EHyOBNsLlxUJyde7fk5I4huV+CNK5qRb3SibA25fIXQJQ8JUm5SjufmT32IdHZs
Cg2bLxOPo3gwWKY6bOH6qA==
`protect END_PROTECTED
