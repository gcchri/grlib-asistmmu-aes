`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
INqAxR35+r0ZZX1OEcAJOU7IprreT+R1a82igbGuc8j3BuTVAxRBTTPAp9RpIinF
cpfjtx8lwHiebt9TEhAbdanRvtweBLUfMscvbpLtFDRSUTFnIdvSg7PLv5JHqQ+W
XehVeVAPkowV12K0lFvqSxIv3chO+7K+zSb1zA2c4qgWCs4JFG5V6ITp7+bIBu+N
LwtkbTCiBd4mQ0XXpH5F2ZJJZie/A1SA4C66UkL23OElhKleZJi2Nh59LszXLMGp
xZXxRAuNhm3KJhKlf2UexiwCiipjyIrqWvXkw2EvkyO3d4hjKHRMWWHWKIohCliK
qIVQcy0lmlusZ9bIPhNgwSxNySuk5r/Q2H/hX+O6Lwx1o8+n6CM6TRHIjDzrBJFQ
1ik768YCBpBbbcMQqCzutXFi2jyrcGAC+ZzCy5Qz01/fkkSCa5lqeUab11lrb21a
ycbW+XYS5KtVIJdWBiWQ3NdaG0TVGZ+/YXRPM1SZejI=
`protect END_PROTECTED
