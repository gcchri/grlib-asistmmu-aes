`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rkn6nkDgVQa0aARokK0ucTrFoausy7OcBKPIeNRIbiepmnzyeCDgZe0cjc50DDKX
aTr7AdFOsj5mgTk5n5MMv3PBNz5KvtjXNCpbMJculYMYxd5UIlloLJQHgOmNWs47
yW7CctS20fJeM3y0VBDmSgvbxcVwY8ILXucu/HMeSbd7nSKDPHHSfz72PRGaQCfN
P7zKZzrYEPc+tVigWv3bYwVtH3ywN1PubRgpYVpRQrLzdYxa/lTjRaOPC27Rj0yb
JiLiGj9AEt7Y5UfPvoU7RDPm7xunloliTyIRBSAitC2Jq9YOJrzOBqCy5C5MKYUE
YKz6HIHeLOdk5Oo50QiPkKdXUjiNREvEPWfG5vvIa5s=
`protect END_PROTECTED
