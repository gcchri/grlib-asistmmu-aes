`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8RCCE1DV3yTS68rt4/IVp6/m5IMCSqzDwKZIBzCKvJByrUHg/c8IabtK2BNWoMTO
8+vZNLzp7K6ENsiiCIppgcyEQ8mSUe0W8HQr30m6puKAIDkTpapBhxzGpfM5TvsB
fuOiwzVeIQfyCg9WRUqSCw2EmwNvppqo+1n6Zrmsj6qbSTH8C4zdfW1CTsOke5Ba
N+p7C9GPRG0ZTXLlGhGzUA/H3OTompMIdseCEZNzYsr2Zzny5To52Btg89PCOyMw
WA+ZSRubKw6ezISvLLgycRQCGwBptGNn2EuWxmWij6R3ntHGjIJOE+6m7A4XGQWS
/i4nxCQrVhEUsj4288yP9G4l8bNN7v7bpl3eG+WJ9Hur1dKbTUqQYyQCw5OZE6zH
hXQqIu1XQGTo+Q0lmIuH3gb75eENWhqLcaz/jJztnfs=
`protect END_PROTECTED
