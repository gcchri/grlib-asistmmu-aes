`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wSQL15Z5Ne9kP7acXgY0Yv5BhOBcMy2S46S67Jcny1yNiaykdk7CrNyOMF+zu+6E
nV1hkZzg1Q3sxrUY2ydcGNyPTUG3DtRt3A22PtmMNS2Q1kN/ShJ+DBcpWuChbF6P
bF9ZQxkXrGfNBfLHUt9/Uyvw2FM/zeco/jSUsShBlTPiagINeiqOrWTzglo7wfv/
S5vFf5LK7ssh9KrLX9ELQYqH26Y4QnXlXPkNOdIoKPV5N8QTFtC2X+85Li5JqCFT
Z2MH5tXNOBS8cf/blgNzjlUbOD4sOqKQMRAue4KCZrPTkpPMzdJjGcGTz/XUB7/Q
Er/A3HI6EzO+e6jo70kIRS/LkcbDWp/3+Z1Ea6EBPe4b44LckKg5ZpojvpAB4CEp
q3x7Q74XZej+ORX3supssCtEHT4RW6Hrkvuowe4ZHjBSS6u9W8t3UQX0rVIAU/Qs
f54RtGwodaZFMtn5KGVzbF2fjTcGF5X80oFA4kqIwvX6ZWbdujFRlmNgN1MN+MV9
W0uWLwHLrkhIMV3ebGzRfQT7t0Nj0XyWGJCsXudVHAd0KARX3krWwt9yY5MMWfOo
3fTS67NQTlfZgj+ewKRi0i5wWgcvVXwyPyBST1ooNR0=
`protect END_PROTECTED
