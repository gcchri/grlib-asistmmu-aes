`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UNJreqfr5CdnWKyFqIYf+4wOo5PWbel6pJrLLUdz5Vs1gCAG2Lc+LsCfKfyAonIL
JIjh/54atToo4U2MPA1mEIP+ti9mvIIXDI3EkNl/g5/+SqC+PzQxqOqDRmrzQ9jR
UUBWqwoiJixMKWH5Yywkgu1bFv1BouyV3VihgV0aOgKuzyUH9qAey0g1CRR+vWIB
xLsab/T8uQ4M9MS2Z3+6wSIlkZOATN3WlVblhFJXyE5Y8Rux2CN2t3EQ+dfaF0UD
5LFdb4bcUehPUNZV/TPro9iEdw99EB2s1gA4EtnzQlTZ+UK7Z8QHmJhLA4jBYgpq
msExo/O0e3NqKqXs34QWO9pvQuMtQtsuTtBqWOoYz0o8DK099X2MovoeYSYOTFEo
lsd71hodXJPv4BG/ImDZm34T90xVwWDFxFG4IDDAwh5yd8qL9UyWkqMHDwAp0bkC
AKgjUs36xd0K0HHQIFUP1BnYUhyd2Wb4qXLQX67bOyth2prWypfNWqhuFQewI/VI
PKPl2BXpu1l9esEb9vn+DZeFoiJwyLvy2mVRuuK6epxQqlnGUrOYIIaVRU+EEMhz
Z4OkorTHoRtq9EOiNuuGkQ==
`protect END_PROTECTED
