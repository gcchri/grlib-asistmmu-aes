`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jLYuVjMT/pthRZ4xLAMv3uBVVwflzRIixawreiNt6ftKAb6ge3ugxgv84d9jE/nM
isrpVA7RaFU9G2Zsmcn7Tm0vUhD7p//edPBgTKXa3m/OgTW4d5gylvttp8YVHLeU
fDP824OdbHPIVmYeua6Jwz948C9RSbvz87vgL+cbefw7dNGAwdZEdk35orzMbwHb
KTObmVpTetaNv0uobKRBwjLaH9h67UYxqiAeLSde5qSYRSL9zamAFhTqDniZO95F
J5b3FfVuCmsKDWKt6bZLAcrTLmF76IGKiXFUJdmg3WM=
`protect END_PROTECTED
