`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8brFavoQSvuyOqQx13TOZ4W1WtsmfJ2CXctSWJF51lDJxiez6kYMNlEMbODKNe/6
64od4WI3gAItEvpRytGaZXEKGpVt8qYyIzGu7B5KnAjr/De6w4I0PkIKP5W1HERd
6aYZu2Vnt3eI9WQg7S7usDX+5N0eZ1sCGKm7ojf5GaQFr+60NT9gHzcRIw4AvowY
o09D43llWY6tXM8u2hk0Vl4cWeszg+9uAo2ikP1WuAMVVuqFwvwIeikUhAWe6+kk
3YRBCo10MsYj8GWEys68ogqOd2r55wOn8ht5BszoMH9E4X+I4bH90o2ODM9aW+kk
VEL6q5oZQYGKb39+nSVOFg==
`protect END_PROTECTED
