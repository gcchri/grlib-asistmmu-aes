`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W+T1VxPGpIi8a3w95fWEhpbM0de7MyyJiFhglHiD4MOwVvpPM7PQB0KuiCxQKjI0
sKNGeB59LvHZRtFdy80FItORTl1pJOneco+1zVUugPtqsfIy0PphPzuQ2V92k78v
5bjSmr3wEw6FMIw13PE5lZpN7C2YWPnd5AabmEx7f8B4JUzB++VQf3MPeZkMMX39
aM9kCPYkHcLOgECOPo6wnJLsgTSuqarGG9mGHnVxlkAQfFYobXBhscTz6C7a/hX5
`protect END_PROTECTED
