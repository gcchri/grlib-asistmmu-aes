`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+itytEDTucZdd8f/DsTXEPIg084B6pr2Id6tgUCCPKysPSQB/zifMjf4XmEpZFzl
QuBsudv14zusvNlnas9w/We0/j7HJ5rxxl/I9qPZD8htbGywBUaAhXBF3ZrxfloN
miy6XETiVhVeUUrIsNvM6pofm75cCbuH+hZjfEaGYPeIe6NyUeXyvmpte9LRri8A
j+//PZJZLoSl6tqOyc5dX8z1IcOzkGiaP4ykVoiWBaUKTB7wgqqo1WkcoDwUoNUC
vcfJ+Uz0LdACZbiouuaM0Svn/laT1Qpj39S3HYvPMZucjfaeBy+8bSWEOlQdaBB9
0Ctt+hKwc25AgE6bybQ6YvuZkMON6G+ArNW1D+atxcqaoNMow5reftufJrS1UaeZ
BQjkrDKh4ERrKmotBWvlon0HHdbFX0FqiKUhB1qBNCbNqGelkSpVZfs2UDkovZ5v
IUP0lbk/znO1z1LKwoS9FNg1/wCv/4ziM544JT1MsShafMbGG3JO4xAY72IYo6Y9
+qA1rHPAhNH3BUrfuvjrchbAbim+OcATTs9f4ojwwANsirOYUfEyhao1gfD2Yxpv
ecj7WKFfPkwNcRrJRfervzCi4WDgqLZtN9yh1iq6KRl9IRu+BwZWlWSKLpD6X3Xq
m4yUdldEEeOPCQaUJOaKVpUV++Ouwwp7rtTfZCA97VilhBgptac4I9O+bLIZQE2q
fk5kBj829ZO+uYgdmyEf0qAN58Q/suI0v1+IVPTJigRb4SiAUogCAJFcswTgVRg6
iSPc8XH00j1MAFHN1dlYWw==
`protect END_PROTECTED
