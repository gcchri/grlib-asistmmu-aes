`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ucQ6sJLKSq9l8X0FKmjQgUc7paJv7TZyX67S+5s/Ff1utuFm5UzhIxx4p/XWcFLV
wvoPrWh4jp25Y8CcREwTZ8IKndoqRMVkGxlYmq8igkirT7VCfrJNOrETZgUidV/K
PDbXKQGTwluy1ky5qZdvKo5wig1ifF0/v21koiLUPfZ9Mhhm0gvDFGWAgqoM9QlM
LJtfdtNnHyUOCVPY0Iuwi7vosNiJi7Zz+rj0jWZCAjxCwyhMQ24wZpOwZWTX+wxE
`protect END_PROTECTED
