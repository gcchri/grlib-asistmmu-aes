`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k0N5c5WqTQ7V59QXUV6tHxd5jnDcch1B8eB1Sbhhn/JkPkHhhvSVCNM982lePdMk
Hf28l0xFE6IOFqEBhLr1S/9URS6i993kUEGl+iAMdiJ2ioIa2SEvXNgpjayBV/kr
6rQ07S+RU9SeedS17pjDQI+bfQSC4O5tJvMIVNEQ53k+Dzm9lil+FDRbzMuDK9Ul
Bju3Fmo5wS8a6sTBbtKWsjqyQxcj88c+E3vq2MgsLYmCjBuwPUAuPmJrMeLgdDi7
EX79Gu1W2aeaEiuyj5GCEXUPj5Tq6hOlQeV2FPSzNnpREVtAZt3b5b6TK0WKiV0+
u5/7iNxgFEEATsrrTqd6fFSUN1gPvWG8Q1astOpcgyaZKEDDPCYCKLUKVc0tqWZz
SvdqdKeYwXbeaLyF7sAgRsMxomj/fuHOPnHW6+Jfbtt7x1QxXKHjoIbIwG/V/Ii6
SIWh2gyEeuvbB6ULE4R/MUHFJaI4rYVg7ycS09rGfOw=
`protect END_PROTECTED
