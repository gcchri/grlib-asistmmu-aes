`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lq2RUNYHDi8FSDjetwdQPoaf3aNJPWfC4Zjf9xuILVateREvnd11KIzPaW4BtSRM
k3Z1I5/YldHwhGANM90dENmCEgSLkrEE8RzzQdDBC7LoJ1uhJplWW+M55LYGZf5L
UmaCsSZyfuNjZ5sbqAECJXtvpQeezu63tw1kyqqnR1UvnJHD4XC/19IzNS5qWZda
it837dIuJMQcjffBffP8NbU8QEFaIYhPSwUmjl9/dWKOakrcH7m3/VxvjpXetb9L
1w4FUk+S6iDYZLokLk6wyA==
`protect END_PROTECTED
