`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6OqsJlDHtv4m/sLedXuLIcU72gUw748TYB81+wHLkdg1o2z3CrjhBMBCjSgxt2Vf
9h/vE38h2Nc5donRXVbE1OPfsXpEEgkB5SNg0VQ4BQPZuApEj+j8gt4FFDRySYwA
LtNcHwrDDGBUxDuSVqiukIa6U3BUHxIX7477EzJPpULZE9vYW96uz3WmUxC5eMa7
FlnO+qEhGSk9rBrxHsMz6X+unGF9rh/7Qfw19OTnIE1xLsr68Cw9MyUtyIIcxFMC
O3HuadBJgX1ltUq6a2JwS0XR1dxkrKBOrUka3BvsiWG1d6iW9QNFkMZVEtZ1ha+J
q+1iTNG9vwHI1r8oFi2ICEHvMmx1TKVBmntxkVHBk9MVP8PSQyuYYv3hlurpYmfb
+1tySCI29kskipmA6geDegrMW/UHOULrKjSxzmBzIm0=
`protect END_PROTECTED
