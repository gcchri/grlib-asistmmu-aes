`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SpHEganU9BBr6Rr4rU9mg7lEWvn9PCrwSMc9jMowWm210OVpjWWw4nuJoTeObjOO
uknhnMILoLUEMUAWztzz1L4d4Ss6LBEL9tdWFBxS5uc2rVrIOsfCtdPAx7PIzo+d
fAIyxJx+pUp6qg2I3kw2kn7p0nF8dWx3UrzmAf5asjEmutbaEupx3ipnF0r8NqNQ
Kn6C5C6N/VdPLL3mxqNPNvlZ0Axyh3Yi4olG7/NxkxYa2tgT3gE/jcnPbLc/jZsN
P2cmRVWdgRGCInCxGunoGqaMHmGuGZxopAXJKOn+zPZbYpITLQebOYDGc5jg3zHF
FJknzZDvps0vWOH5gU8Kqds7Is42MIZLrQCDQ3X8Fha8F332f+1UP1DI2suYMwtg
PYYMaWuuIcmQph16EX4lVrjDSwGCfB1aC/Hp+5pOPWkwkIBCKfTvFHKHfNE9JYHt
HbsWikw22yRlwNxUmKp0CHfC4+Q6WuQFaXvJ6UHcLgiswT3GOLhWYkh/Vhvorlmx
+NIKNplGe8o3cqgLjcKdBGHVgai9kZzDK8ZdpH0t7wUdecK8I98VcWp0vs32NEoD
WozHA5rpgbTpqWT4F4FxBafWXR4mDd0rWBX5r2QCd9xoeLlAcOUHk8vFShmEUMAH
eqgJHpRCbghg2W4d7Pt97A8sbwBwG6Um0EXjNuBVSpf5cCE46WnaCPR+AZEm0fZn
JPmBrKtzk8EW7x1V37TlIcrh7wAQWpABPX2TK8eGvTdpk6gMfkckqP2fuML9NFia
KqIm8hppe+xr97Z3wQlwFJrVFs9LkuCw5NCPa2ci4FEVBcNdBd280a1H1Y+9BQch
qdXMHZJjoRj6sKFLkN/j3+8h6ZacxVuiKFBT6Np38Y1Vu4zAYK+I4A65Yu3YPKtK
0iQ4chwqS1i2hxA/MTRDm8Y4vGxsAuw/JfDeLTICvkGVUZJLO4Ue47xYcLeDTM39
/Ra501jlbGIXP1rdsZDlU3swJUVGd9PEVW8ce5+X2nXUDf6OGMbmGPe2i4NA6OqQ
t2GkamlBGN02TlColxyCQJxDg0HE8W0H6uvR4jg1Xi6paIxXjp42i6MscRWtv/+4
wfQOjAA+SImBknB+ZKz3ZeGfgmGVCq00sUepGE+i7nBj8F+kVGZCAYMw0EvC1aJj
3PoKaOchApAYyQ0rkZeis+XM4eV3AhWzsfNo4RNqd8lG/AH7O76na3FezvZfn1/u
za/AXD93CWWEpeAbLM6I55BY+o9biu5efZm7f/tJHKhfIHZberKhqrM7QdputJII
Ihvo0bgNKeS0jgEc/xY9XO3x9ItoloFyTDTy/7VA5y2IVk4ieSEmSGod149qjAqf
T4Y+aPk17lnK0AhU/hzOMi87JpQpKOACbWUJOm0WBBiUnx6SYi6rdARJ0+wOcXKs
XsD0Jn0cnKFXfLAo0dotM+gxzMg9MqJVNX3gjtbwV/hTZFBUuJg8uJj0N0loyB37
nEVn8nZCOMufFjl132Imq/hVgrodJisRcD54r1TvwIeihGrSLwiMuvksp4DpXsJ6
Q+wGfMAit1T4HQcDQFaeflmP9ev/Ju4gva+Fuf9galrI3fqVTNbxCm625cYsPneE
rovPGJI4JAuXocLONjgrgXZUlcoRIRURHkqr+f6V5P2asCTMHkJae2+2W7gMCmga
yw+KyhPD9sPzDRVFWFkXp+WY3DPq1cDV/zmRJBJHjdsFYgWv602urhVZRaDse0I7
U7x4uZS4sFLO30PYSRzwrvpQCKBa2Ap455Mo0L3l1UQTS+dfzKWLbMCvH26lqdg4
JvHhRynRWQBVzOLS2O//RmrlY3oadgIB5TUuLF79+uOU7tgz1FEbsPHFJXSmjnJI
zkMoBaMd2FO0UU5yokCqcBw9nCnKKcxh+LUDz68yCmAPsM5svZVjtdmYNK3wQ+T6
PTva4iDhW2E/fQs7yAgiw8uMoBSzcUpBSVinYWW3Eh7BUUC1vf3CSc14sS4JqROx
v/wjnlHxV6w7A2DCSEx5jCGw0iIUNfoTNwbmbFKXd1mf88Da+esG2bSwIARiynAZ
80+l9uIK8HUDLeo3ynd3Kg==
`protect END_PROTECTED
