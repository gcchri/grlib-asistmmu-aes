`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2EX9j49UIffZERq+CBSJNrsCSAZiTGt7I19LrBI5gUdgoiA4V+I3FyZtgcoZJq9M
xnWZwKBxGdDh+lwzZYSyVKjPMPS07xPKqbVkZlpCRLXN7NEI/j51zSAsHZ1XS81L
XHvmnq/ASVUHeihNtopDzEvxK0z018dI0nyfrEdjlFlgg1NIxlJXAj5pdG1tTYHF
rM6UkXoZpnxZkB7HTh0Nd+VAxb/FSvRpXj0uWc3FwIQlAj8+JokF+538I5z+KsfZ
8oGfZqG5PGBME4ICmVM8QGXYtw4M9FaXWa8/AMbHkINcDf3z13bEeFCxdAu/OIYW
jasXlJ/bL6ZfVPLdTz7IVmH9y6ONzKb9TUXYMJATlRQ0zQfkWx9+aoumK+MiOY9F
kDbTMRTz1SUVyKgFPqUkFk6sQu0ZH0P9z4SfzKqdBfwb/d5Un9xu8BkJZPrdVpln
ZMZexlPECWPZIyX4pQzlElO0OHarGpgb1Mk90yHeTfh0qFy0A5RG9oeMx8fuvlvd
1h7cmtJzhzAk3krKSXEPfDcVToA5H5WxU95E4gL3woIg1MPVT/x4rzUtTIpnny2J
0BEdsHdxvMGhzxpl/pQhwCTVarCiGn2JEt/gwSQ1eh8Qeb5IVcRiWqJxmT9DS2Xf
g0tftfZxrO4eNQjBByluiCXkGKyna+Pitv6ffAwiWhRkIBfWK44Cer/E9jlGIlV1
68XrA9YRsWP9HQJ8ECIXiwNGgP6CZZfsZmR8ItPT31220JYG0boAc32WudYrYhDi
1DDsOViRsF/O7GaROVleHAdM+Q08Jhyzb9xkGcrD1Rue1gEsYI7bRpCM771PITDO
ca+HC52IAAXsvXK6jJZyoW2MJXKwE/koIyJXXDJmHZg6ydOP0MiGzcathQLLfrZ5
fpIc/4d6z1hYUfxUf1IMmKE5VxQNUQpx6XstSzGlJapvM6T7g6OIP56C7qlRz2JE
TDc/hgKXDl63KZFD7E6r0AOoCMeYILVul4BE0H7ysFT2WH81L3KEaBkr3tfQkLhq
gr1NJc+tsuU8lhsHBZWa7C/dyDwdXCT5MKsKehiQ4S/hbufYlHkkRblKBUODyMw2
2PxG+ewjO0s19jjtm2PJwwqBJf3PqOAh7+On7Q45JJFjWcO1hPF2YIisida/fl17
EGcUSzJpYFSO2jHANBrcyVe1R4LaCI0fzGN8qU0/299XnYYT6qyejnRnbNincLXy
6udsgzySpv1MbJ6BzLRf3fKWaLMK961FI094S4+OEBZlPOzsSERTu9zmiGEGWihz
mXuVwyRDXr85ezAjtKx2ckZJiqkrZyWiaayQOcM51K50KXIVhWmr4bEq6aDpoM20
Y6bRDq9YnOs0WGV+eO72k6xAAbrYRpb6NUxLIhg+h/EQ+rJqbRfRMjRggHSK4tAz
UwsrK0BSNBz/ztHIwGoOgYyiLEBbZhLXutf6kwPRANU128B6q/mPK2fAL37gN14O
ZtkGDHgObCLTQqixvtluWMKvf7BHOvlx9UR26XHoCj29SPTw6lKM2tQjSYza8TUa
xIEU9kVuvIbPwBaInUNvMLj9+T7EYZNYeGspbAioPdjx1vq25O4je8uNJEgRlFyv
g3YGMMl7k1gADVCtT5Bk7HUZq++N89EodVpxLzZ4PT74RDy1TkO+xOx/59KvOXlg
fFVIbKRezHqEajHm16qrSZYu14OCO4VuShyfvOY98AS+MKP8ccCyqIWFbcwDUAAu
wOLgYPYWiY668KwOFLM4oIsUQbsLsclJ4ALuQDAb7wZYhnqgNifx2NaIecZa2DqK
F/GkmyV0RGtRSDWWWymffoSgbFu92t4NVOzY+/lfFG9i+8EBaLx1G2thYP2Ptmj0
D62syLlqk/11I1qrC/DGHJrGWns0TPJlFTBfUupKV4ejeIm5H9gU0I0JqlhKp4L0
+lD+TbI7wjbTQGS3FfWap8M3gQYNWTszlnBG8J3RNoERx9bcZwnp2bI1Pkgf23W6
IHUP2U6tStlfOzqVfRgiHnpajqcfG2P5jUkKSuKT/15GgRbnM6LUZrVc7cb8/vwJ
JSpmQx5M7eYPMNuxjJygpldzS930AS6vx46WzmHeKekZGbSAzLG3kIPala35iloW
JqJ5ugMPHPI0UkcHKdSjFbSoIOFUGtTabrd+CIuViPxHUS3gum15zSMKqkYc8ljE
BHe4IHKUqJvvrL2P0s8N8VKA/z0DRlzdXtAJfQtBr7Da9zw5fSEdLL7EuQwbBIVf
H0pQUmAB1eBFk40s3sBXxBAv+jGdQ10qXDltTqo2NmTcehWkn9wVC6Tg2EeqUFJ2
7PfoGhOtf4dCE2nd849UY7+i6FNyC3HuSdAeld8Gq7TKcETZvU1WU2czK/86//Gg
MREJDZTaH+mfoekJ8oVVJ9mDEw1uZq5vcmXwvrvCJPiJmf/wuV1n9g2HFcxTkX04
hZqadAdM0c4pguZK97lx2Vrlny8z1+2xLqj+Xe4bYEH6qk/dumVIz9Pf+QNmAVbO
pKtthxDn1BDOueBIMQqYKp9x2kCnVfTPktx9ILIdbdOHQBg6V9X02EC4kWOXDhSj
e80yCACq9UsEFI0yWEsWKNm+tOGGDklb8pkCyxPNNfQvrYKflH6s9wKtBBEGtanL
7wK5oqSwXDuEVQAV6I0yI7vqOBxRtqba07/d15zx9EAc/WcnJF3nxTxgbFqsMGrf
U9JPv9xg45VO/Tpw5AXlaIsZ8c9V/LIPiVKeYbC8y9y/rqllyYsuLVDhLdCWb8h8
lYc42lQKyEsUxU/HfoseaFni1ThH2wBkQV/UvH55ka3rxSrMCxrQxEsOiygkDA5F
tc6VufUHLj/Hc50KOcSKoGniohqtJzdIVo7QN8cE9W5EMoyT2Gp9XOzVcLB1J69S
1ddZz8cX+XF/POC0c9PCM5ZSTG871wil0dYuaRTKI6xtrzADHzuVXvjbXqQQNsZd
aN0GmE1Hu06GSLf+bFYPkbJG0RHn0ANnSx7jqSOyAx7qqToUyW0jvl0/1DmNiJPj
1mRLPIc3tV43t8DCVxT5qDMFnyt30kSuH+Run8Jp8nNhwch3K/i+sqw8FWY+nOXX
VYPvo8WzUT0TPznLkjA2wSehq1QKVKyY0/6VENiwbQ047AUTcjmuPfnoLQywrSVf
IdVknbWQ9HOX2Tgz4xJC8/F58BxOQBs/YT5xPzs5xEBLH6SBDmdaGYtbqem9Bvtw
th2B/BY+maya40kumgWqNfht1WmpcX+1R4YW9S35hCvGuLKBMqV1LXwdjTBEiKmj
1k3YP4m59Q1I1epulUWrUzH1DFOcyHXD6+78bYN3BXJgCcERCwBaFhUaDl+eND9Y
y0mL73pArQxnE2UKGnAp4cUPmK1GSIk28UyhaU4yW948YBfGOBMQRcZxGe491MZ7
emUnsQkxp+kHgTWUxRfIXTd/LktceFy0OSlcK+gxKnXLQtjtuRfi3udzGnpEos0a
B8OArTRHH+SmM6NsHv0xYVyd5MVstwqScqw6Jwg0y6kyGwxLrhx534JoyW5pNGD3
OeAeRzjeTdPAiU3Y9zgDu4L8julV9j3jB65bOtoiAtIB24q1BeyiVfOfqTsFARZn
xCaTVZXQ9TFEoMlgD0e/drEx/ba7ItYnW+d8ZqsQBf4pmwVttxdiqxAXG/k7Z5kF
r7LyLJqcoeUpqjuG2shWNUhY0U8McLWOMv8BxyHKmyf6ykcM41jAZfSwc0q+7NTY
0nd/n3eJpOMJZIqMYQSLQOEoOsiWqEGc01ZKheuajTh99r58SqTT2zGqr/Ohc8qL
qC8UdiYzKJCZuAcKcs9GqNitsEEqoFVxXCigEfXEFsCqbqUFzjUB3s396zmiPfny
cz2pg2bV5FCQDQ+Dtr9VGA==
`protect END_PROTECTED
