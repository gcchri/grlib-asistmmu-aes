library verilog;
use verilog.vl_types.all;
entity SIP_PHY_CONTROL is
    port(
        AO_TOGGLE       : in     vl_logic_vector(3 downto 0);
        AO_WRLVL_EN     : in     vl_logic_vector(3 downto 0);
        BURST_MODE      : in     vl_logic;
        CLK_RATIO       : in     vl_logic_vector(2 downto 0);
        CMD_OFFSET      : in     vl_logic_vector(5 downto 0);
        CO_DURATION     : in     vl_logic_vector(2 downto 0);
        DATA_CTL_A_N    : in     vl_logic;
        DATA_CTL_B_N    : in     vl_logic;
        DATA_CTL_C_N    : in     vl_logic;
        DATA_CTL_D_N    : in     vl_logic;
        DI_DURATION     : in     vl_logic_vector(2 downto 0);
        DISABLE_SEQ_MATCH: in     vl_logic;
        DO_DURATION     : in     vl_logic_vector(2 downto 0);
        EVENTS_DELAY    : in     vl_logic_vector(5 downto 0);
        FOUR_WINDOW_CLOCKS: in     vl_logic_vector(5 downto 0);
        MULTI_REGION    : in     vl_logic;
        PHY_COUNT_ENABLE: in     vl_logic;
        RD_CMD_OFFSET_0 : in     vl_logic_vector(5 downto 0);
        RD_CMD_OFFSET_1 : in     vl_logic_vector(5 downto 0);
        RD_CMD_OFFSET_2 : in     vl_logic_vector(5 downto 0);
        RD_CMD_OFFSET_3 : in     vl_logic_vector(5 downto 0);
        RD_DURATION_0   : in     vl_logic_vector(5 downto 0);
        RD_DURATION_1   : in     vl_logic_vector(5 downto 0);
        RD_DURATION_2   : in     vl_logic_vector(5 downto 0);
        RD_DURATION_3   : in     vl_logic_vector(5 downto 0);
        SPARE           : in     vl_logic;
        SYNC_MODE       : in     vl_logic;
        WR_CMD_OFFSET_0 : in     vl_logic_vector(5 downto 0);
        WR_CMD_OFFSET_1 : in     vl_logic_vector(5 downto 0);
        WR_CMD_OFFSET_2 : in     vl_logic_vector(5 downto 0);
        WR_CMD_OFFSET_3 : in     vl_logic_vector(5 downto 0);
        WR_DURATION_0   : in     vl_logic_vector(5 downto 0);
        WR_DURATION_1   : in     vl_logic_vector(5 downto 0);
        WR_DURATION_2   : in     vl_logic_vector(5 downto 0);
        WR_DURATION_3   : in     vl_logic_vector(5 downto 0);
        AUXOUTPUT       : out    vl_logic_vector(3 downto 0);
        INBURSTPENDING  : out    vl_logic_vector(3 downto 0);
        INRANKA         : out    vl_logic_vector(1 downto 0);
        INRANKB         : out    vl_logic_vector(1 downto 0);
        INRANKC         : out    vl_logic_vector(1 downto 0);
        INRANKD         : out    vl_logic_vector(1 downto 0);
        OUTBURSTPENDING : out    vl_logic_vector(3 downto 0);
        PCENABLECALIB   : out    vl_logic_vector(1 downto 0);
        PHYCTLALMOSTFULL: out    vl_logic;
        PHYCTLEMPTY     : out    vl_logic;
        PHYCTLFULL      : out    vl_logic;
        PHYCTLREADY     : out    vl_logic;
        TESTOUTPUT      : out    vl_logic_vector(15 downto 0);
        MEMREFCLK       : in     vl_logic;
        PHYCLK          : in     vl_logic;
        PHYCTLMSTREMPTY : in     vl_logic;
        PHYCTLWD        : in     vl_logic_vector(31 downto 0);
        PHYCTLWRENABLE  : in     vl_logic;
        PLLLOCK         : in     vl_logic;
        READCALIBENABLE : in     vl_logic;
        REFDLLLOCK      : in     vl_logic;
        RESET           : in     vl_logic;
        SCANENABLEN     : in     vl_logic;
        SYNCIN          : in     vl_logic;
        TESTINPUT       : in     vl_logic_vector(15 downto 0);
        TESTSELECT      : in     vl_logic_vector(2 downto 0);
        WRITECALIBENABLE: in     vl_logic;
        GSR             : in     vl_logic
    );
end SIP_PHY_CONTROL;
