`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ac6RluTb6YGIiL2FYOWUEtIBslfd2gFEGQWVKysUSVmENv3m0vPHeTCeyeSVxLQ+
0U9tWV7h9m9B9H/6cAoMr3M6hQQ4/0vQVFHGk5JxFLzvV3f0Xvz5VDICKFSPawSn
ZzwC4tJ0mn6J6m0iNaG2SJaQutSuSgiTyWAU4zpmI7Jo0chS8PM2cFIAxo8zU+YR
6RakTkoFKa9xhdjzwbHd+bTWovE5nn+Y8YKWQEAf/5lMrnCxT0OAj0dLz+XKI6mt
qaErsPnQWsQWx2WMVmMoD/7Y0zXeevMeVz/jDfkplHbV+NcXyDNjT7KNWD00hON3
9ePa3l0NtQ7LXRJttLCy7q13FMBXFWqAtFkz9d6jHNUiYnjIT0J0Nbu1KKBTUqPG
wyfhazreFlfY60/0ShT4DnPJ6Zjg5tVjX59RmOfbJv3V2kK98ky76hs0fcTres8r
U9BeniQhqZOBlWYUMXH2K2j5zInQLWuaKfFMQyUOSb/UJvXfgzTrBhj/xlkiK9hO
pL33tytn7vlK2tZRdp38csKf/pqn7/p8HtD6nTrdYAof146Lv7pQUDSwKfKNDXwn
IhDJhKj9lNgh3cMjfHGugS5V+f57ZHx9ST5jqC6f5a9Pj7kkX2XEVd6ASkGnEypm
tk7SWOevEajS0dmgkVYWk6hPO+uHG0jOMb934gQWHLI54uPE6QzF/kMkilPtlBn8
Oz8B49+aUTJ+WIk6bxCTtygF/VnTk5PaogHuIcGSIYCbZ4cXo4tn1Pih9/WT636/
Cu/8weX8IiuYyXoOpNX4z8Gaf9mzjbIAtfz8ZgCz/nHGn9feqYTRupF6Y/JC8OPV
ZHLV4kZQji04f4OLwxVEzgSNbDzIvajgc53QKIWjYu8CGEqrWZdI8bbPl6uHxjpv
Bo5bH6CaOpnZGouYraGFmzf1P3yM76Jt1Vo9P9I9wXmYEl9vWZxWebTeYinPVisI
Vx5+dAWJXpwFk6c9zrHrh0M+/yR6Hzpn00Rilwp2GtW0loWTgQkCyLXtZky4nucS
RSGqIGno7qghHg++f+oy4gs9qIw7FqoP60siY/rvOrnfMo5bUqob+TA58SsQejWw
Uo6iW2y/8H5LHVtcaf5lBg==
`protect END_PROTECTED
