`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OB9MGAhjSHwtVR7u3wu3zir5Zf+XBMPNZQaStia9nhV5UGKKWN3mXFWVO9HtEoSx
K4b4xntID1d8S+hVQeGbtrXmgnt51tdo9W7/kcgEU8Ia4dvlEpcTPXHlXLKdimhq
zmohR1l7Hbb0cQqCdop0RwXhbltzPDBWvsJVEiVMplzTBfdh7VGtm7+vOPm+9sDP
NEOAM5EIbrIDIGSg6QNDlMePiJBEQUFPyFirOLlmpcnMMBbnoUSjlwogoRaZjSgO
U3pwEHXClq0ILJYudVQrxeMGwqDruO22HP/pD7G9zDEOzcfweS8yCOne7j1vlI0g
VwV4Y6F1h08MFjK1F8LwqR2yX6M9uA6zK+PoL3QqA5Yv2GjvH/HlryXHfODRTV0w
SKKDnrODGmJtQ9siSma0sDGjDk3Pi2LO8/aGsW3T7NhaHCdxnfNHSehgU/zHe6AX
PjAlfvmRz1F0mr3rCjf3cZi354qinCiWmjPZOpshs7gzdM7k3xKJhZ/+Qw81i6pt
pIcnOAGz1Z8/zxAXkhd57+RjvRku0KdE9Tz04kkRjpC/gkcObC9wkN17vWtmUawT
eboyzoaGTGpPrbA+fVw5j8S/iPxE0yUSobDfKgdOQ4LtbZ791gd+H2lvMyWox+HP
8Ah9KzBelcNwf90LMvskWs/vzoU4WrNg4iTToFZ9yrZADkDAJ81OuUhoELrBE/aZ
rHYtvozJe6Fcemb+lh0cgmjpyVosbzKheRXE7ZQolOXiIwvzp5fDb6+wRRs0haga
7K//KLCxIf5TqycZ1UmhGqwiv/u/MjwxffYmYgIJ7X3FcChRwJtrp6uNmkHOA1nt
4S/hE+rfcu6pXFcyTVEhgSaevFJEEazn3hwW+uvmZXD+Bk+WYNXf7FV5C7T1xpqn
y/g8brzXN7CLh6Th/jvC4pwSCe7jboFx5G7V4gRemNcVvXXn2ZSUpl9cUkJKZ38a
irlR2yYweKF4fSNxySCo9t3pgegzvY36CsOuoKCQt0YpvwhS5ATvt/0xGzJqG1Zi
DfEjgK2s7s5fsNl3rHWfGDxYw82zVszgmsHrCAd1axc2rtfEC5Z0ouqqSRlFw4T+
DtDkB1WmJ+E20Y+GtUBgt7bkvDwwnQ1iwNb52IU8WG409cAmd6BqJf0VuVvQCR6e
OobXiMGXfQC1nDYK3HuFG401xcdML1hESbdNtHqrawPNFCdVV+wfIFnb+aD6F4qH
9UKjPH51rcyNcSA2rMQwTl13rmkO/kiKPZ1seZYt/PpdJX2hK3p/xhEfLepijEcS
HZT9eeAN7d4dIkK75rF3bEk3Li37ZmBttq5puyavbqBkE5XAz/XBlp5acDn5P5ti
gO8sxpoCgO4Lc+8ta1E3EU5kFGPNLe9W8QermdXEd3q01A1l2sPoW3rdAI9ngYD0
kDaj8+B6nTpn9l+kxxzA1w==
`protect END_PROTECTED
