`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l5XWnlpYqdbwYVrtpLcwgipr2ff6Bl9yBvjkDH/w3dk/DyDCBGNnl48liEXzFCfp
s3E2uFLek9PVC34QOXIgBru9yl2lJGnDtGfbGnt3osG9vaPciC18PnZmoE8aa4P/
iuOPvvWzvsXA8/9QC50xUU1zStl21m1fMmYGUx5pI0WA6/tHa9zU+elAhGZAoZvL
1IDkjxSCDBs74yMPyGzsB34TO893nowaKqeJatrJ33AMIi6esCnp+Me+gLKRZicg
FT1zv4bzWV+2v0jSs9XdgsOk1c1QgtNahjeWzjc1/q8rdJCcS0KMoUPEbnU9dD3X
iQpWRdhvLiqFM3IeScr6N3qxBkeGVGQs9gfdM8swu1j6POwC8F37Wq3iku/6/jmo
8iMEJG0qFIvKl4K10Jvm7c82b3+Z563XWAOBX1yyCAQUeb2QHyzg9Y27QSN8EOxK
4zilvaCOx85kElALpKdO+NuMV17vXatK6v7yE+6Q2KLCRGrSSyg7Y9hTls+3FKht
2kTHo/0B30qLzCVlEsqifD5hhleooRgoRGIFFpSOSsAdy6yQVIHSe6zcnZ9sb0Ma
FQv13g50G7+UhAuYCL61kMgZCM1OZK+SRwoWuKkaTno0DNv2llFHLIiMKh6iTnGP
YtfVG7ddfECQwMHUsMSRQCn7MbzGQhoWKwx8vxAsTK/w2+yf7DFlsz/EauGpSKrP
43xEJmhzfcRJ4nPPr8Cu44hfHMnFTWlB8noHqWJNE2lzoBu37LC+fxuUp3qrq2Vd
CNUAr8XEqtb7C8isvBG11G3QyqG+TpuDxMoGqXlqQ2c=
`protect END_PROTECTED
