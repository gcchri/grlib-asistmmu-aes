`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H0duVCuqSbc1MkfQ1XSbob2hz49fMZBKSpxBxdI4p6vE5DpD90CG+UPrD4glCqNT
wKc0g1c7hb6AuIrTDdBToxpcBEoEo8BXfi/oHtgaiMzbiWJa2S6I1vRx/v6BbzU+
hETsaIijubhyLw/tQpCEAnr/ljLJnqhyYenzVteZmmGRfzQSLhhU3Qm7yQR1TtBN
iU6oCL8kiuPTC74ODW+rLeTjTl6agHLVrPtD9qAm78+CI0xIQEjToXkSwCDaEemu
Ru5s+706EbLfediDKr0a4pS8gIXCp7nhjqvFKOreaZNrvUJdT4jgsPuEkoT8jo31
kQV3D+nnNMLv4BHJqWWXQgW4N3LNSsjU/Vugo/G3lIoux8HOEE66p3gxn6AfnuRH
XAM2/VN1xktKTlklm6rouAzO9CT6n+nb80tgDmGr8f8VJFydrN1xpOHKeUI9Pryh
NZBOD0BM5izX+DuitNYkRHQ0ExFiLhUnPUIu59mNoA6auXckdzdI2dEUqVpwl4yV
Xzur7JgykNohMB69UaSEa3Iwn/b4wADeKOHhD6carGvTQWIHVJYgr3I1GUrMGLQ0
gAL1Qtu2jz8eGXzJRq94OH9n4UAUenv7kxL0cA9rJE0pM1X6WlI8GbSqyYt2bXxD
WUm8F6WritLY7W82JvfLmaZgIQ83qt2N+z53NVSIqbAZmwR4tMDf66SHpuJWi3tn
iizsbGbKzhc3Bfeq3dqpe8Dowjs3/+OiDHMZUdUXAQHdssM3VElKmRcxpAZTfe2n
Fo9o6bUmSDvOpLQJhFulBN+ZYuBTFw3zFD/fOkEjNlY83YdrCpN26/xYjYmLrSiR
rYgJl/FxSiwHc0qlST/siRjhUCStVDPA5P40TCZZM+y/twpu5zjb5zWvfIxsoYEG
36VbajAorq73SVIC/388XMVL1cQ/To+0Ohz6yLUsQL3AgHzVK1kI/lT6JMoaadlX
Jwiniiae2eFhh2fNwfYlJMr32qJBQ7s5E4FjpmW826jwyEw4lAH39qQKyNfC2f9N
uHUDg12YtZ0biz/HKW5atEIU1kCwDMuWza/CP5xfN/rV3ORcYUiSnrPKr7bwXrO1
r3gg+KHm2PdVs32unS3P6/KtA/BOgo4OtYcDPPI3Z/aaaBnZOQWdsAwJEixUOWIj
OMYTPEsOrA+gj41lYUtYCgegSW5MzREJ24OmsLMxQEUq9Xrif72pUZ8vm1osU/Gp
uQwZ9XyosVJfAshi9SJZzhZeBR+M4I7ULrYZWQzb7z2unRcsbTI/o+Mc0Mw57QuE
bqB19/oJlJPvTisxGMDTVCu0/0mOD5QHpUjma2Q5cG7tH8IYPoWgz8Uid4SUyP/C
D+z4vdgTdEPJucd4Fo4jYO7S/xZ+dD5C/NeqGUG52FNyDzQx3SqlU90CKKcLLeXO
C7GAa3XaBEURQwwABZ28M2eo3rNtgPij2zmMnoQ7pqIlpX8UlueA/rd0o/ya1pZR
9/3BNs0Jj+5MjozDmmu1lb6PMFyStTJuSd5Is4dxmpxnGksMayFXIFT7wSMAdisn
yj9QCZSuh7w5Pp2OnBLGm2CiKzkIWoIIcsjip2W95P5xEMPF0Y+yntgVNuVAGRZJ
`protect END_PROTECTED
