`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pPqsM9wqa0sd58d9IEBkYpe9GjaGqITne450x5F34tDhLTD2NZ41sfbeDckiW4+b
ONYhnJ67aRnxq+08fnAesarppq5vd2g4Jnyinao2cvuJIC8u7agYlXRtLbjjDj4Q
UXejkdyiVJde9iGoD/TwqC+my0iClLfSesQHuSblmMe/ZX7Q13iePFKD0tGI5Sap
4UD/16MmMQIdgmMLs4HQmC4rPKsPzBFRQE9aTtph9DieAlw4IufAB0+1Phc6pifI
s7bHDzMqu/OVGC0uSjc+Uj7i4UymmA5Z3muuXRQF+CXGf/05KJKh3iII9pNNwTYa
wBawN4aMnjLMTZ0LJS9Yw6CnxZCh1TauLAy8L9+JNiVwRRSruHRT0+mUwJuyQrWw
nXyUbi0d2+G8frAwa332Vkw7K9S6fc++jaZSdQtVvvjx8Lie+SKZb9+YoRP3JurK
gyZO1a0F/pGlp4p821wO7WmGvTzNs/pHsdhPj6onF0M=
`protect END_PROTECTED
