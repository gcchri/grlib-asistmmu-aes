`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HJXlIbHatyzO9zeqYQ7mClzGbWWyMFU1Boqd8KMpIpdESD4PJaik4OeymE1b7wGW
lJW3RHOUOynlJCtkzntq4W5Ix7TpaLNdcv+AumJ69xGOO2etBn9oL7wzZ1Lkss6W
Lh9iLAiUItFO5VXMua49W5WRyUda2G7DHxynLA4O0A4O9oml9h2FftOz8QuBa+Qp
yD6Froe6ghs+7fnprKsNuxLkQL7bcsM5OoypY+YLZZmcWfdHeNhwPE3rdpeedS9Q
WQejXR4egEveL7+cVK/DiwQbz2sAQEyN4RAc3mDs4kDKy6L4BoPSjmOMKEeMYmYy
Wf+1rzQQcfFO7VTJOvPGDdxG+8j9neU2W8q1HLQOLHje/2BS6wAcsJZTKiQ7jWnH
CyFXlxg9lIiDBxcEo5U37cxHX5zit7a0ak6p2p90fvIhEIyHbLowRulpk/gO+GCj
i/rixkPUU/fxBOYc/GIobrJlBcFbOvw8F/HULP1vANaBTh0LU6XRfPsOgXqnOTaw
lYlnzTJgFSNFHK/j10MDsbVZcA/5z7GvDpN050o2FKyUZISxTXD1fmm4W2a7+Euo
+mIPM3KT2UtuatKbXTECj8/2zqA06KXDCwGh0TVQpFxX9nGHrV1mjQY6x9gHpaPc
w8aQ2FTgkV/g9zQaJgi9yaGrcexdZdGkH9zHWuwTqhAG1aBzR6vqOsyibsY7VhyF
LbesTHitqLBqb2bCZnttT2dVpkwxuwFEWz+VF82APg5KuyMZa2beEDXDsjxBbLOA
gizCZk1OpKIwZO3gO6KE4gi8ilgEWuxuPpDxHUHgorH2Pa7iWQ8ODru5ZUToypA/
Q6pdOXCvlAAeQjxTa48tF+e6qiY4fne2GU86oRY05fCvTcf/tu/2OlDAls4Zijkc
HidOhfXT5aRsafi8jr4vgJJkjkO/SL9koh8onCrj0qlLQmwVagwnGFlv2S7JSk92
AjrhUfM1vGJ1QzUQtfbwDpBb2EIcUV4/sy6POiBK5oBgZNftct/TZ2mdzU8t9Dc2
a81VFM+OrESDxLiX7vzSDQ0994NesI8pvFP3QowmUOMlmMDUE50NguR1koZrn4Ef
`protect END_PROTECTED
