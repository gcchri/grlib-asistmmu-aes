`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WEWomkhJYedOUoaT0Ugy7QADPBuJjexWVG0Gfnnz0pYmcyhM/VvcNeH67AHHPwwz
I6UwdexK2x+Y6RxX/9CK6KWeU7o2MoVqnjjT/Xop0egBT0nj9ssZEryOyTCkmPxv
IHFdLqghVe5rhTrPkmHgd2y+7ysI8YvU1i/2aAwMv9yfuWlmnHRuwPNMihLU4/Z6
DJtkHS7qQl3BHEj7Yzwvw/qldAfsOyprD1jGg9AE5ctvp/mlAemQYP+F/c8CO3Mr
nAbhq5T7uG8l+rcgYg1nzeyJIvf6PAwf5SGy1GA+azA8kWX+la6hsw+eNKsdbcsc
MYZCTCSTR2ud6FyBc/W/6IOXoL7GmpxE3xBCSIdpnkdU/nHK7HgxdH/nm1dL6xvP
O3rFp9ORBx2QIFh2KUFdi5ZPXKxtfIDxo/a/kcHLm67b2DJB6Oo485urQ3RWufxn
DEm88BGoOxpSA5paC5vT93NvZmSJ7CuPB4FzojH3CbQApG6JLLu6iAbxbv7khLoJ
E59rEMRsE/eEYovDFy5lhXWR2FTqAUl4YnmPiFRbMDQRmMrVLU7+SbDE+ZW91A3G
Lu3ARG/XhlBfOO/Gv2HCrMXJTcvf9c0xDJiMfn6pe5vpMyGmZkcq8FSkWi9dB0p5
vp/9dPu0+wtyqeMogAuj2t72njSOYh9SIt8gqljSDfVqf9HBwT/TO69ZECSMOB2t
`protect END_PROTECTED
