`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oS12/+zWgozlpPx26y7I2AGTOX5TNlSVuW1RtGibTMDyl/+NIa1Qlcu9n0YXN83E
VcY7WgcU8HUS2wWykFxchYaL8r3wJ9J9Ub0R8WeuXrQdd2zcOBKZW5Ecc+u/KFIQ
pVxYlaUiXnDc1vdHW04sguwgQwxmEYZ1Nt3E1tjJJTvEIPckK+kKKmkQISTz48OY
4XP/3/x38UkPp5dE5+JXxPnuUHRuTIBN6XkqshlTx3Z4GbN2I+R6949Uyow1hZvm
cPFO6Tl0K6/Cxk1G20OwhVOASzGGI5b5f633tly1cN7F65dWJSiJm3pn/8QPorn5
RGPLWQahjfcBssZZtUsr2g==
`protect END_PROTECTED
