`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
trYWbt3Xz7/rr3ZnWODXdfLJL4NmsShNtZQPuOOCmKSGeKonxRR6q6h2DbH0cten
wJkZ6EqylODk9J2bi7n/xSCUr2adz6EjQCUgAylOot1F3ji7YQqOTxbKNctNEHfc
hUFkjYH/D+1OgfbzxpSC8u1H4bCFhIty8rg4hYf32wIOCOlBLAuYN2OXf8a7tSBz
N3ijkcKCZfTfEs4WLNrYilS53TxFaJtJQNJGwfmOKg0dL+1WfLqym33XWoPTYqYd
5dVcfdDTlyiAr42kdyLAVl82lKvroOfMw7GevSfC+lw7jo0/k/+Fty4UgMVDmB6n
GBgiCIFCF3GMrspUxMjZaXQkrAKRHB84u3MGY4T+Rbo8XKeLmiGPpwRhCeygJny7
PcQs12/n5t7j4YIx5EApFCQ7VoQz0wbNgnBLDIZrdws=
`protect END_PROTECTED
