`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qcmOuBTfhi59D891gY58jNV5yZR5Za9Sov2CsuEmGT5qY6s2P2SHiNw0WokHgES6
mS/eL5+6qBzVUQJzF8R+w+ILhYSyupy2q4nBCf371QFsrHCXJQIxYBNQ9UN6+fWU
rzE5JdQ9KqWyIhAmeSKp7jnzenDviWRn0dGJPip7dG7Sm4y0Nm/M5pYAXUfGuLFd
3GhpJzwXU12izutwCKlX2iXDd43az+6epc1siB0pbNjCQcxlxfLwilgQw7uchyf3
SbtP0r980D+2p3zBSwzlFWUNYSWzW+lhLn2PbAN5LN2FiXc8o8D2W5zK0FgpPFk0
oKoM099A3SteCVeQDz8VUgQZQhYCjXDpcd1PUMuUMjuzcul5IkEEHsNP8Pu0ohO6
P5MskjzXxFuw4KsVJF57RUzJtVUvTYpVwlonu5Nmi6MiGi+uKCXkr+6BotlkhtON
6PrNSKk7L4w6Kpi/waMvgPe0gLfrm32G1ntRK2NDKVg=
`protect END_PROTECTED
