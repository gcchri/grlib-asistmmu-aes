`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I6XMf5ybgKY4Jvxueeo4J7CkGiSyzAEkgQraPnCzshcoBV6cjRlOASAdDVvXxLzv
pC+K7xsOPl3YuLOMursi01VVUJxz+sLhIpKqjO8Fez9t2OIUrgEbeh/C8eKLOPlH
8Ma+EdXgBquADwcWc/OJuEi9juT9WZ66i6hfXvaMW1+pY6S/G3UdCH3wenvc8Vwm
CoizY9IRc5X91EPoa5mPKWxYRY/Gx6M2waNz56bC0YF+gR+t1AGrM0R/AGEezvPf
AcQzMnNRIEp7934NAAPCJJPDHD6h9QSgZ7DA0nBVLIiUI1U2oGr1mXuDZbRXbouC
3dUvv2D0C8cvdG4uqrYbDw==
`protect END_PROTECTED
