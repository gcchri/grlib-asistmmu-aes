`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cqM6LISLOql5cvdNRwsGY0CVHJStbSJma2gfvOFOiLL+2+j1S6e+lvfOq4G0F9oV
AQsbmMvnnrQqOWm9PUxvqPFeXGdcI0tqMduF2sYXmDj6hzcKz5HL6EpRxPumpHTU
KzT5tQMwAZLwVSkkttuYT+DfR4H2ga5xhVuWr6LuQUWK+EJicYDTtFsjGapaSaug
RYhRq/XCPR3ZPoUWjOsJvLwGbItvHAlCQUj+/OLZyzi0Qxswy4n8Hw1KS3j1aC1n
vZ0o5eID+Y9tW9sr1QPvXKI8woHL/8ND8OgeTOOD2PwHZWcdaPEJ9iW883Xi+/gg
DtfS9QSd0vrKj1FdQVbxymNiZX397VtPhYeH2VtS7LPEB335vG43MHrZ6MqW/vct
C5r4inxAHbQ9AcJR4rkvOYNe8REzK75K5R4TgWQbVwKZv2I1ZmQUOY3B9GqHEn5T
dXG5eVvOXvLSpDvNktbMkgZ79omZFv8q4W4JdXXv3pIeM1GCjuaj1ACG6yPcuMDp
ZQ26HOiVIcTkYRunHohuINAYmP3cermPS5460DMIfiprQqmUM1v98T+N6dJBGl4w
Tb4rG/6zYXSaqzaNBeZsYS43ksr/FRQO9elq2TZdcVHrw8TcUA1lt1nQ6ai/kpO1
UDtvj4xlhY+E22ibJGGHsxD8qgYq7aoEepMCqtIlWEo4KHyPISCmrnYjFzBwi9mI
XYI5Uv5h+bbc5FR5QCysnko6G+fa+92lVKMr790N6tbTUmvIIHilviqcJiE0YJiK
0p0Pw003QNLidnnxuvClDfSshZMR3rlgAg4nRBBq+v/0KlPN7pUfq4c1CB8vtxkx
IhtLduy0rpmkBte4/MuYJ/PWlUqCUDWGLyfbaRtPygo=
`protect END_PROTECTED
