`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
umLr3/FGldoBVBFcDhdVwu3sh37z83BiYZhD7dyy+SfcnIgvROUoFLQo+DuRV/MP
LsaIO4kpcyGIPKH71ewW8bnkxXfxTXDxSpOcNHfh60dzwDRbukRpycSBKsvdNdAO
iOowVASMmnyRPVUG10GWyWJYkZk5XxpYqsLrrwUIzkf8ScdW2schfAJd9Y63ShR9
pLpOazAAKhlh+S8BgH72nDkXFqz7Ka5YXHXM/3WIWM3oPdrS1fnskITR6IDSJNfs
Fq59fAG+soqFeNwrrrsdIhiKUBFlNfxgFMAj1Z1J2MTusCsw7m8Gk6RaKYgClqNR
JtWKhuxipSQZRihW1AsPzCtuHl644s2Jg2Y4eUQRzJRYdTnR4i9r6cOXT+/fQNXl
SZHFIyk/CwoC9TKSUjC9qTtB98fpCij5BHzqI0v7hyuMXQFZ+yhKAgivCLuqRGhr
Gs7G4Hb8oXWOrYLgzdfY/IxdDGN07Xf68kiZl5z8ADvRC7Eth0fewqsfvGkwSU6N
ebHTv17135Lun+hyjU+znCHQRFEOZupOjASWGsDE40uvOAiVbxFimVRrFj6BKeL1
EF2jed57i8kbZIt+8uOgEQ12w5bmKfJjHhWJN12P++AEjxQGnqnn2R4vP07LuHsd
`protect END_PROTECTED
