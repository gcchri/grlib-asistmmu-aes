`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3SbjoFaSaDqrRe7roxhPd7P+o7SyLSGI2pzUewMskQ/81e7GHJ56CktSJR8AL9o5
bKbzw2s1z3D2E7kjewZlYv6hqL6+VC0liNTrWBnfCC10cjQqmE1MKILX2tNrB8RM
SFzSj6Gcvmek6itL11Uk5QG7/5MhrishufMXE2QLavzfU4EL6Vu4KYq+gtlcndyP
NoVa1IHm5WeI5Lfzhu/aFOcYN6pKUYMSY734Qm4uxg8V8m/Xtfh6tx62jcSqAUDy
YAtuBabtue1wxHbJe7FyHLfkJYSDd8i4mJ0QogeeZgBGF2Em+u+ABAa1ktI9aazv
/pTwVbhwDgRxy91dFisHSD/9R1JMn7pG5eU+ySks7GvinJMCdK1aNmq7YxxguEwT
VrezfndQxE3wFS/v4VNxpEJ2YIp+7ibLjrXMDKiRAxxPJXvWbkdqNHnIDHxwVkQN
0OoLG5qQF7FIeSpr6N/ravitAk6HANX7PWg9cdK63YQ=
`protect END_PROTECTED
