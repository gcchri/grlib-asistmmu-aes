`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h5Fu3jeOt3JF94qLfO/wgPKcGQD8WEBBJ6FMjheDNdeOPAsAm2qw26x7tIEACXHi
E1825bQGcyVr32+UG8dwYUoMCOQ57OotNzyTOzim786cmK6HZZjEV+dqAU1C8Ane
WtfvBpxDPQPS14bJZdgLb9PmcgtOwDQ22rQB29fSx5vSjZPUVVWHtksHAYCM44BW
2gL/IHDzUJ7RSjZ3VLWVCc5d1mXHWvMJ6plosAZ3W2A3KJl92IaHW3sJAnDCIzFz
tVS+mCsIfhV6CSgrwEBz3z5u5PHe8cloY48nD9AxmL++9yfBKvs/soJR2Q7a3wul
qQ0oM/FYFxi6iM2Y5uYxpg6QzhaTRIyEd2V+w7S8VWVjCKZZHn2dzfaL8lcxVgt+
n0po/IofGOi0iUOzWmczBK1JO7cpL6z9JS30GmXblFXCP9J54VOUbiF7gWOPCn7i
GEuxl8b7xDWLjRk+zO3VqAe2q5rXsXaREKsnQB1wsO6xKNMro+Bza+HIo0UJy+ZD
s4NBYik9v3MB9aLPmoE0SthwFJi/wQKVp4u12zfRtO8lVQ2qaHWJndltTgZY4OKE
AiDNm7MxOXteVY0YWLtSfVJIdS0QMxYZLLA05F5HT25P3f2mJSyiZCPyN1+qHmJz
Ld6vJg9dCzPgroJgxODRVWDItqUfoKYXHPVbK367BdduNI2BORRS4xNdmFSfphtr
OgAq3Rvw/87wHtpDy//ZZrtLtF9vjMQHYK3tG1Bv3X1DuIEHTIonOeDnEzXFx46B
fO6mgVsqwAFqqhIio//Dlcx+kNnpGl1hZw1faRKN1Lp8ghZwY7Uk6z+IycYSX3Wm
x4hVoRYb4Xt3qOqtFk8Kk3x+No13BNIndNQre4OIO4h0eDHsjy7tBHlSsn5kpFEi
WwDzanes41WmcYjFW9FvEWpLdnodv4qsScQpstFLTSqnaSA5MGLPffPfy4JBseRk
HWL2Z5rmQLiKpKWrNLguXmjwqqOtkKTlqBW7ONQy8YY80yhQhYmAU6N7G435aoVd
AdrLevnJ38O9tjNydDlz5f6+N3VUXYKWXHnHIOLVXwSR9l6RZfWYUPoF5ITgegRR
`protect END_PROTECTED
