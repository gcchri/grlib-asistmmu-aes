`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HOfkB+H5K5HwEtV5sk6MGmexOD6KeQDUx/Yf04V8WUOhsz+VU8gJP76rTN2W9BW1
ysF4YqpS/WuQgWxzDmdbqKo/I77BVbVmSWH4qqav0imDF556eGWrcBbrLkbcPX/U
zCORkaHxr5lA1QZJ/T4d0PlGPyVG20vzSwNeq9Urh50EForwJAJTbRN0fNgbG9ig
WXKN6KjqWnveP9L9Wytl0fdBjEhRlGXaxyvsNUxD6RRuReA9Z/P9Q3BoaAKr2fym
khOWSHmPYluETenEMXtjp4ViPcmKCzbmt9nllpuCXdWfrQROJdtp1R6MnsurIrPw
WB/y8xoAOiSHIfr6DXIR/XVyHM4+DdyCUzQlfYh3sQrgo7YznVrAP4uGtmSv4gS1
3WngxmSMjOcXoU/ZFJnRbFe+Ql2CCT8/wQgqy4mIq7laeo0raETi1BhkWJmPR9tx
SjlROuHFB8/vdU8odDbN8Y54Rat6fM+S2bocNsNno1TS1qsa9qV0b4SKCH7WDGV7
QeDid2u6QhtLswgmWjnuckrFAjVISb5DS7EUx9WOlnxbIjFwczf0j73KP90Sn6/z
B4Htt24HKcVMYM3WZjwtRzd4nQi18CRlC8briyBWS/50P+bQDt3vEG1Vw6oNlNPZ
38kJ7e4Seio/KuqGBb4DtaZB1CoAivzcSKJucL2JEUqLjGUqNRgP9KX24+bueLmj
S7eNlQGh5tBv06jaupR5Utqkl6HGoKV8fle8KTqDAcOw62NPqlf9aqPH375HBpWn
EiD8fTTpM0oCgUMh/5MosfovZxh0CU0qhj/nVGUSOunHr+PQWiluXuFxVU0JU1um
5LSnvx23CwZkdl6ciGmsATWDHQjuAQjoPCKdm0vuLHYe2kJ0MRaXD/lIpWfGIf3x
DFSgjtCL73zZ77xTdyoH5U1s0e9V50sRrUNUz6V4wYjcQz4hDC5Ok442uEnkpxJt
16uiASmkhiNmv9Ifr/k7a6bU2okEkLg7xyEuEyrWPRAr5QBVdjP8emDDaD0CwaE+
f/Tobuwtabb6bhQtx/YWkqLCi2deue97fmuvrIB9vHL1HzTgJPuH8x007hCN61Sl
4qLCBAvvLl4rTojhlqaCM4UHWwdC2vL/6vpia77btRV02pv3dKiz9txyEFcenAxu
Q9kbj/tXO2LRECSZt8bwEdn0GXJpg0Q77YrMkkoA7GhkSHxSHRv3yA3NTF31WXC+
`protect END_PROTECTED
