`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
weJosP6U99tRrn7Nb7ZBSnYitXmcekSThLTv3TfHbfv2ntDrclVA2t6nb3ok4+tC
ZoYNlCQ1/VUuKQCRF274gGa8rqZMNAOgV+9Wq1LcXwZ8jwnozWbD1gYK+5m96BQc
M4PVjwpD5GcbAAEE6LNe5z5Mss9BajkU4Zrm5LjorS3syNJha3KppSX/i8AeOtC2
h4V1hINGYeTbwOupvv4P1rVfUImuImyojRDRJz/un4LWJj9HEDH6dn0tO04DepAU
NIBlyQJKl6d/aSk7UXAUZ4CSYIz0SugaEfoQwqud6DaZRkERoosxyUx2HCWog5p+
gAJwPlA1NClU9URdpmI53+FbcYM7OZKHXoYQtTpZO878Eyu4IjzAEbymbQSatIKk
2zFOA6Jx3ET5r1Kosibi3C3cj+CgampVpsnDlsQL6ndG0u7+1KBIjXMFZWJYUSk0
V2WevBI1B54nV9X/N+8HubRxRevkndjitnPZCkCcnw3Fxd7OeU9ig4gAhD4Ivlnn
lEwEAYFNXZZ6Rdox9BHSrHw/0WEu2gjb2uQVzgn4FsfdS9eWozI8lQQjEUwHhrAS
joAWdiyI12c89q8hdISzjDC3XNoD1owxGtKqpMyDeMCdYi7yn1x0Vv+11MU1WTrv
y7AQGpP2KnrQEOmk3va+jFrdW4vxnvsQhmJClYaglGJmamLab9iMLYbyWvoIGlxe
iF76FeXLIOv1GtYImq1Z1Jwu2ybk8LGjTk3cfh0UukEU7MCTHvXVQ20toLE58LRK
vOsgk+jXmRw78nkfssvVm29X48eF+eDc2ImmMVmAa8zwAhYooJ0t96QEY2jSK6nR
qFAcNpx/4Yd2vyBohPXJejXenGyHT7GBrcLYmpd4BEPyeq5VilxyjVhAL8MhavHZ
e3PdIIYR5HO9Fgdo67MZRvav2FDnUUTw2+lhxx71BDqjDFshjMhZbZX5d1vgPslz
L36HRUQOXLaGIwyufQwm1mek0/HfkGS2hRePx7y7IgF2/VEJNWQCyyPndqT+AbVd
qaVO95JxxMsMUxeFQDXZtot+85cHJ96RVOAlad1fJr7ECAbEB8cNHmyBRroogwvo
DfNcq0LIile5z9TefJeuFV99c7fcoDzoXVMwpOh4XVcz7gpyzajoHuxQ7BPBe8HB
LzX30Ut7L5PkHn1MIKLl+/H5oqGDARg0q7WAURP7RUqKCKxr+1AKf6qg7WOf8JV1
CIW8UxLCylCaynYFh0p6H9u+5Wh2ck6dnWQrJMrVZ9Er/0pw6bN/BR57UjBJJ9HS
rhwbIbOg4JF2TmPF8WKFb534wtNsBn1TU9nLYpG751Y1Ya3UXr7bqHhKbxlhcR3X
QoMdpl2KIIBBnHn4nEZix+C4exR7f3MOmcU06oWOsh5y/6aGKLFM+ndZonSxGUAl
gNvRV1jd22q5kW99bRHEYsWw88jUk6jqPUio+O/Da5eAGv7XByOphabqjq3s7+Op
7+glLAfXFsjRIPsev5AJY4hgqPxzZT3hoXrojXTB2AQyMK+UzTJ9O4+1UkEfIXIb
BUP1aERBTGtUNXzCez2RThSai3QXKpKdkO8Xr2e3WbpOnVe04giQGd1JBjZZA6i/
/4rcuVi1xEN+WQDzq9uX8Z0XCtfjhERHXmiHmM48Sy4X2Hw+SULqO/zA0h4P2uzy
N/fgu4j3AHT4GMYaT/VgGPODPto71Ckj/2Bq80kozckkazUdLn6ZuloMpjQvT0D8
ozvyAUJT4kviQ9iTzZDR+nGJPgNqQFX413wHiGhj2ltagG0XRvXFF52o5uGCDJM4
q48mSkSJI1vIeQ1mGYJCUSS2zlVbVLgD0oI7jom6WHfUcd3Qm4F5ClqAoRPLzvvF
WMOztwcsa7c3OsD1vOqCjTj9nOfFJKwThtfNhN1FyGVnCqWMMfEXa+9F7cMqsmzy
r8y2I1DYNbTLvCTqePe7SUz5yGFILR3oXhWd+6hgeE2FxnmtVxbM2BHPdEJZiJ6B
OXByR1M2hCzX7yWnuCTZ24wHMUNpB9B/UYFCoXiSSLXIlGs27nyRQYoj9bRD7T2b
dI3krTDnmSgY9gyNwp3piweCNH6t44CB6/pTVLo5Ckv2tDRkHRUOjM3DS6xf7BuH
IFDRDERdMOX14z90Gc0yPf7U36QJ5RhbvL5ztmSE9n44yOguG5OzBlQyXd1Vk8V/
wATQCXW78r22nJToESb58cmlM4lloyODpxwMDpbnxLMk4lkGvkA5bZNPymbeGPX2
IUDA7kCx8hBbyed6sRlKbh+WKANilwK6eG0l4Ub/Hkwn5TFaVoB0iVG3qJJf339/
JsBei5D14kX0BKIHU5MQKCUYRhvj58GaZtXT3uq/BQlA8swear31ejlAQKQJedGN
+YSYpb1g0AkDWKgjruCqewV17CXv3g9VqrD7jCb1k7PJn0SYdd6+uPD7fcXNSbtU
iWoxXGTFzEVbmn97OTau4yJnbAY+ODV33AAxHEb86ADa+bioC7fpgNshUNd3KWyX
VVwEtKDYkoBmA6XcQvYCqDuRbWbEEoCxui3uYXGoIUqbgqIiPMgrXBdgMQmYoLNy
3NfcYc6NMWF2OJ9gL6sw3gJQrIsoZD9g866TsO5zQtoC5sW9sJkGXBvszJWh8bZV
7jI5gTWCObBbiMt8F76IFy9HO/mKOQhqgmlf7KRwnVimALzc1vVB6JZPiLRbewCP
uiRDCUWZJlAp23M4duGEX47b2crLAJKjMc6hUCvRxqM9CYOdEsk2vrXJPrUHnY6p
FZLgQxnSrg6BoddOVxjKHmDDWcuuINjwHrRJWqC+BooPEDXnnsOO0a0riy8mVoYD
Y6zBBDVbBYqGkhD0tD1q5W2CI6tUyHQY9RdCMooNHsN7xq0hto6IHLFIs7oGuei9
MLgmMrYg++LwyeS0pFK6RxD0a7ErMFI4oAmeR19GK4Dz7XhfSgxBmbR66FvX6bT9
9+tMFyaKQAxIoFhZOCEWejbX3j+m7c8BjqsMeq8i0LT0JlMmxRAPK3FjJyrowHVp
kB9lDDUR7RVPeV+NJsHtSThSlA49BUJNGcdJw0f2DCIIPENxKbSdtP5C1dScp9NH
LqwR6fjHgO4H5bH2xaCKdgsCcfOo+c8BCm3QoeQ7ogwTecZl3PN1m2BaFGmwzDMe
Qm6Lej1PK9tQMj3Q4z6fSTxACY16ciJR0kzxSIJlzk9HW8bQ9H19Qs7+OuqmCuF0
VA1ZeA/i3eSyf2YVfEcxEptrJBOq5+e8lckKFMBBEh2uxTiXAh2nmv1DECrNC++5
BM3AY6O/9RMgNVwyJzFSrZteuX/giXjt9apRaTTtJPxg1JJngmQqaUbj/n7hHbp8
fjt/VOY/mC1LpNieb+MUpTnVFal8wo0p7Iv4LvWiMv9tTU2t5XqTJ8oEe9Ki1FcK
70OKdTaSEUs7fwDTY+S/40v1VgjGlqJhfprjrVOBZrA1GyH7Me+rfQlmt7wSMuPH
PHfBwOjNfCa9oSX7OAcLfdtHGqr+gbGH216VStYomLUnE5WJUcv3H6mpQHcl0zN2
C7pn6kV8ayK9ZFf/cLXsmuw/r5ZjtfPbgGMc5V8tIYDU3PvLUnvRayYAge15oNMj
vQotoH+bXRtANCAxlLC8uyjvWDMYDg/TEhsAalqH1HwV04mqhahKsUtUmcRAAGB7
wz87FO33auWwK59uEykT7h3ntZJNjrg32Zsum41gZERhaBE739TbaCgJIp3r/G7d
5CZzA1QtRIi5g16XL/gI9NLBfFY4b8xcR/G4wJWsqrXQDrGTCk7mnTf0ppWDf0at
oduChp4H6A9ECnn3ioIYVgcS/GjCsby8jCwSHbRpCAeAuGLvViancRd9U3znjNjp
SJFnldj7wjX2DKgxY28oPWWYyc47PMJwFWM86khoBiyBZ3gsj04nwrnlQ9s/mfU1
BAWimHDgCk1I/NS6zUhRjz/pCwsNkI/OjQeYR2XV85ZMlK4DjAShihRWZZuuX48h
Jy1wkfNOqWp/DoZw50REKPfq53h1yKZavqwzfd2Y4sPKCzv2GSXip1Mq0FbraBlK
nZUwkbYfJ1gXlJIaqrLjmvYL2qTXfK9gYSuwtAWrobfsiQsd5csf1VA+N1xRwv9o
/rqTbf4pj6kl5I9Qt2DZF/e9JPlSL+SP+Tv9Sz0CulGyGM/JbwCT8UXpAcWGQ7im
92L+j4PfMa2eHYDMVvQh4/4b53eO12KEsnhOBX00wsLypld7FYLczy/MY94AGHIm
zyNdI8++UN7TPPqgYswnIlos8u3aksqtkAJSSN72hoB4LrD9HU/SZibx9BHhUfn3
cQJDXWUvsOSv0I66LEkUkvPLu/N0hOg5b1uDJZI9/u95SG2dG2h06viTdcf3GBv8
gEA+pkJNXuAAhXy5CWl5Kv0rM1rxzKezMMHXV8zgAs6b/gj5ZMGMHMjB3VZSGyZh
sGCGDScon1G47K1iZBn5IuqLVV5Bmo3EPdRg2tR8apM6wAOf6s4+n1UuHHeg3+eO
3o7V4SGRz6W9/MKurYNukDZhc8wg6DN8AElFeUL4XlgjYaufoQJ+1FAQW9v/HHTh
BQdLzFG70GHokszRL7q4A3Ze/DB/Ak5fuHGT/istw05+zjJq7/edBtT0AXeTwN4e
HBjjbdKppCBD4q+Ui3XDIw1JtOFJAtNKINKnvOaDdGfvvGN+Th3hLdbRfwWm+QQ2
jruOnzfau6v5Qjz2OiXry3jdHUTRwKG7JspTXxHU2Ec89nfosBR1kw8ZxuhwV4Gu
p2rUjgnXXrN2yAVrZ6iQWJJvU9mRNgJkWKtTDDoK+uIfP93pKwe+7xMyACSLp1P/
HsVQloXUesrSacOz6jaINmcswijBcvOGx0bO9rCQXBGpgfekVwhD/JaNo/OjgdoT
rzzL5q4zhgl0mC3J/Vn4SuUtzfVM5Cp9YudY2WXzg98jNQayexUUfGzZr93KnoVO
FfD4Agjx4IK//ZMPJJRCyjdAdbKcbFCBKv914/WmoeLcdeEj01AtgW1bRX/Yx6WF
Ngj/8sjBBbJ0S8TsrNQkA6FfsSKnJzvO0l2mlxnrib0FtyXX8HO+kgEB4ub5ylDG
/mSpgUsOxBboJJUz/0ZmXHO2Coykxwja1DNEgSUtbfODt8WQz9su5yQPoBjReB1Y
2g8RN469BQlNT5FPqFKL7WfUFwqKADDJlrrjN+XzVSmk13wFTd5nbmIBPb/AqigS
arxn9k+yYZvDLF1FmseLagI/qlSlgu03brw7XmEWlO1rIijWBZs6u6Ze2qRNwdHa
ALuEwEA/Q7ufFCruVRDM+q8npMOoIqB4AISE1nUNARo5G07en53a8G0al1xnHmdi
8PtkXrMmN7/2HVLstge4Xak55gM8dpkxcznyKk5KiSAxm0+2Ab6hT/2H4sRRLaC7
3k9xbzfrfiovVpqgeGYtv0/yAzWUZPpJGvOpyAjJbCy59b9Fv5c30jXh3QzMtwzc
td3Jlje9Jzk6/U5ZFQtl1sIeUEGfGhnjkJjNwC/cuUGSIWf7vSTvnG/L52IUJv11
aOC5HoJgMneZSP9H3BdkqkazYCGP/AdxQW36DipEbm0Lzcwb9TbjOdUn5sQPneuP
Rq7lQ7dYfZu1oko/K2zlPpmP9zAySikYUI5tDCBUmxbz7XrZ/RC3+RCw88QllwhI
TYNs4HlPqic/HyQdMJa3kszVMuiEDkmnN6Qr5Vsu8U0lhsUeDVV3xwZZHff2Z53R
Oovyg9EvXGWZCKGkOpGBoV8wILR7wjhvaV5nA9NEE5uS7wyRxyynQZ/EUVR4TEPJ
fojcsiFsobPEiXkuCjCWAQe7PooDK2wLpsn/0L4apQyzl7EIcsdF9cK0nUyhdnX7
zp8WE5bN5qVmntyEFvhPxQRT75pmBm5N6ujds5AFmhMZq8Z2VQtpy6yEIXgwyeJu
ApSRWHtpLjUnR6IhxSch+TMKMhkMmXN/4iIQUImnfqKvb3g9kH87zOTOBEa1OkDp
d5R4gRAzs6ktPDakRxLSSwMimzOn+jduGiqRQBu5nw4Mgji0V3l0qkUNaCwOIMhS
xkPGbefyt6r9lbQLzKKWjw9ImPota4IFys/GTbUOPam9LYjUvsLxDEkwOW8OWq1H
6f9v2UUh9uDXKzGGScy6AQQfdT+qtSGf4osc8/i8he1r1gJLqw1dSHw0mU/hsO0l
qWS7Yr1eMUHliP9LZU+tFHhrFpWnOcLkpUX0e9Ej2HXSIQfdV4M/8ougfnbHbeBY
gwJ9dSvymQRtYISg9FMr9ZYolhkw3qgxlVSA3L38J/sPkoW1qCbBT2gbAqP7QaBw
H6LpK3r84m4T38qEKQcdx8lvwM+TPpXlqJkcJaJ7oxkxvmKgxUrcFBoLdYErBQVW
stFG1Ie9e0A/1Or0xyQS8fmbv+PGWDNzh7gsaqNK/JqcuqiEsH58qCJCXAnYcV1b
53C+oiTZUesmF08GP1PJnHeiKqsbKz3A+9WcTOoE6J31COB0l6/0ugNJRrryVph5
t3cDF7rR6aSnpY80P3UHK8I3lrYmv+xn2G4fauYHpS2NBrT1N96pwAD1sAFLVrSy
WPqT1lnLZiPkfBokksKIscIztPfONVCG+An8FcP8AdiYuVp9TatUHRvbAP4rSBJn
Kcss6aSP8WVNa4a+ifqFfcBV22YAFAtEnG8bYTal6jtCSW8xfwtdrP3mzNWgbXwy
QF5csMtK2xFqmOvW80mMkr992/pDngFYq2iFs5+aSuToTvLNy7BRmNswuxKEffmU
FQUEfBVF/9NP+P6u9w1qZr64mJxPTN1XnWEPiltunMPX0oG6s0KbUs72/z146jjv
cKXI140P1TmOr0jUbccH0VKb38PajvgTcRm2P9iI8kAWPm5C1CC9M2dcRjaXu6hs
BTSYpW2zA/0vFAd/McQhaUrhLUkhlTKZXSezPsHyBuZmz2kvb4hghSUjRLzjzK8Y
3jBq1p5f2Q1tMNzj97cxT+BGl3y+oymxeM3uWmW1aFxFkRf1CH0jw3J5yfl77Irz
RmpbjUSXtx/T0F3Q046k9didpIsxDNuustI43WAv1qii8LFbjLVy2wx+ps8l8smm
NV3I1TvK6QXPRGNmkJoNqc6KZAL4nBzzBjunMlwV/bDEgOAG2VLmW8UrXqxij8e2
8GI+aCzg6OVbxf/l691NabUKSMizDXtFtYLbhiwYC42FrLuSkQ2qKIKXHNXTXpCr
ufWUIcUlcFiYo/8m6JOMoaAtaJ4MOSLxBaqi5NMbihaRl5HKL1fodp/XK4pWZydK
EQNnsdxpPccwGwgLzDTMo7Abt74cuX5CspqqJQ1SUJq7CP8VQXEF6L6Lua51ZLRL
xXjk6thyINwiPUx+CkRKYcecf6VYd9VAPBMH5oKMqh9YeRoZYbeIjA3jtJXtaQgu
ICIXMHcLhJ4kR5EfVsUNFkZyb8yH+F5KVWkZW3VzkF2CLdJn54P018HDLkQjOCJb
EPtysf+LxnJzSWn7EPahuDEhB5Rf0BTNPi5Xjlohf61befQjZc49QoLHi4zSNeIp
AphXjM4AUCz74Kd9xnRrk006FoOnxkN2lfSG/i0U96UTzzPQkhenC8kUztjp4raU
CE53F2FeoFUrUOZ1hmpWil8w4eXpN/6Wtxuv4CX/Z4OMqIBCLJ8eD1576qVjOjp2
rXEbmw1bW7gVpR2ue8ARUxlSJLhxh8dF64AMhH/BI3tFljEfH88NVVqRmF6sRxiQ
Fn/3HGSfJjW2Erwe1OgSB8cmUlqlvqf7BsCBinLlGCuoyL6LMY+0STLGWcM0rLby
H8f0wI7ed5RVxeFsKzSQfGqhWRSl1AQnJEAN/XQei3fHPR6IiIQO+GsHegnhXr13
kvz40XsFVnuZ1efTvjdDOd6tJjLNuFXSa1HIorOFe16EZbVKG7pAN8jAS880xrPw
9N0kWVb4a8ojze+SHh+FnSUnJlDZQVLJuGVSPLBSMFvWKKKoaFPTo1aTEpYZh+uB
gIVGaDtlhF7Eb2143KoEq0OOtX2Bosw5lZHzjGJgn3uTHB7HDSYntXx1+wffUSBZ
WFFj/xzPFFleSBvuJ2RcRxh9EOGT0A6czg8BK7yAPNMEGErpZByxSZAGkraeaOjS
i0bhRnnDoCcEVORBqjmZrLDBWrdhs1bCah88zK4DHletYQ5j2MSVm1z6XeDCnhjJ
zMC1Gt3Br99p4kBWl5qYHUhmSseNIZgAWMMIzaVQ2+U5pSsNb5RFRdLPVUbjGJdr
cQs6Peh5emg6/Px8OsYiYoWgrJHIPm8Md64kM9zkB3m1IWCQ1sOT/9N9Udko+Mp+
/h5kkyPBrqC1ti8eQ/h/iKeDEWhYPWFOl8PEWd4ijnnqqMliwCtzxYFefmX/hY/7
CORw1PFKDT1vrUjhKc7iWxznfOEefKYR5Kr1YzOvkzCdXSJAxutTY8uDmAVBplXs
Luyg4zlm7QmSl1pcCXoMaGcEx5Z5oF9FlekYRtajna/Q9Bw/TZo8zyaS+FkDBUjJ
ZZBr9bAI5N2l0pg3X9xE4iAcEmFBnGdJYcVRMb8fqBzYeyH+lIyv/cl19d177iTJ
+rdkK667KYuBLFeCX52DxMkknMbJaTppOtM2rHhPyLglKzHZr2kSOvpps2Oj3IC/
+iyyGudOZKmovc9QgzorkMU3MdXwbpsvzpDDMYNT9PLUSUM/c57QEjln3/i38qkz
bm5K6bQ+PYYl3VMIfaYGF1MSww826YZczBzumneYc8bXE+srXKPIY0DYlxZtLbrx
D/zv3n2JEmp9OcFLqjzgzCX09QjpA0F8NJEfpnU/HHRl9go1pQeKULggs0Ry+jeX
hEkE/3jSIQNrHcytHtbEnTK1aH8WVwsuVW39u0oBwlJXMVkHxDz6jFv3fyWCBcmY
RML1dUG51P8DZvaengLIQIKl06mvtU8Wvu1keF/nKxZm4oIPRs8WYEOg2ec4KfQU
1FuIdgk3jmN+VBp+NIMj09UqPEMk7XyziOklK7oSRFuJFeuDpXaJ6eP4BYTGqeZ6
DhHX/6tywHjAx0Cdxe2SNKFdWWA9UhyAqGCCBICeZX+0nWA2z1MejPYzEw+caWaF
Br53XJnbjC3nfnU24SLh7pKg+bLyx1QX2ztjfRB5ywfSvAx1jmFq8GdaX4YrrIOP
wJsMDezhWZiGOtfahnPn2gI6w30/uK3kJA+tHiM3kXYTx9bGJjpylhNrExUjAIKW
Q3w4mKwPipvaEpA9KApAXjsA/6pjWohsamduKOCL+VNjDtahatCamS4lYS5rs2wE
7CVyZNM+6/xbViCjkI5ZZ67ZLPJmsIXGuKOJjBI+3keGtexNGNfVaQI9ZujFstb4
4NiqR7qPfqH3aASgttj/Ss2fPWdJwm3yzoOFcacAHXsDIGj5JgdUxNClrpyFnHbi
YyBf/SQl830f3pSrIvegYfuhi6yrMiX/zRBTwOG4kYiPf3d511hjRdxOf2+XrL5Y
n98osj4ZnmRTXAsvTGdR28DviDgfhA+ibNsf1K32FBbLHgGCloYEUmaCemD9anWi
51CaX1DRTSOv8MYdAi0W+oSU72lezlaTCfA9NaoQgycWtIk+HQaXej6kdhe8/ODi
p3Yl9lKVW7plXWl0wkUovs2qtKkZA1IRPHiF/OpAdUEg6yiFYGthnsfg5mx92iEW
nvICYWk0Xcmwlw2L2QK0HKp7cV57AqYKf72l9TxoPBy1ZwpiBNbjl9dX4w0UFsTX
aqshRMhxYvkua2prnkmjxe3xrBx3QOWE7rYh17/cbcik/Ls9+lsOTxnrTq3YEJZg
o2lRLfBCR5tjDDQWhP+v3nloP4bEhDqhHGtctDSSN0TH7YZzO/Boi3BwkDCzUplY
LaavddVXC4YUyqKcMUHhMbXaypzkdocObuYhmQNhlycBc5qrt3heZ2KLaziseB/S
5CMdmbAOnhaRbmQqRJN/r55agIfIlEFbC9P8Lkrutm9YBrJnfAzDG26gbafOMVX7
ux5dRrTar5FK11Q8VO3ObXi5w+31R1wGMtGshpCGy4uCqYydwPHJmFEuCUmA0MDP
0w6TGE1l4slyMb+c4zv91wdpWYJ27Og4tIkH9GH4tjZEkYmFP5FQz4r+CVnkSyx1
xMrzcbgGWfuKovP7U2YBDdREeiP+aer1UVIJdqcM8P2pIwjpyvQ8lZWl2bVZPg+B
/0LTUeQNalGuT+vBp6oHVg9yxDOyTkYyw2Dr8UhMH+WWrh5HSjF4nMn7QfBp4wjD
UrThHd00NYKlf6bm5lt02xWjZ+sqDZDZR29CQZLDo1uUOkCP2XHLCZXLBuLFJwIz
8Uy3M914Jflqd6bFz4+2AkI14HdP1kpDcbbGakS7Uv3tJoZmFMU+hsPvFq2sms5D
Tz523cqfRn8tOjsXrHiBNIfXyDtIYWULDZU7wWIUHI7sx3ZivbCnWAuny0mPA1x1
Mu8rixuiqVmLSBPsHY0QSffJiFmruvHUXMj+x0aIdD5xIXHotkxenuxH0jCn/bt+
EU9hckFhY2XSYzau+xAcFd6gAddBf6segDYoS1h39T5y1YzWeG+ii654L7Q7TY7/
/xklgZXY70C2nWpnNm3ZWcuZkh9jNyVJ6gOLKfol5U94E0FTlD0pcAhbHc9UWVvZ
WdfQZQ+CNydHJwQQDHXmMxAGfKTAvST63QZQZckF3FKz5mCp7tGVDhdo5Kq1k0u/
9SkiTQuOV62mIfp/zXX2KYM5EGf5hxkbGdIHl1pcF68UOZlvOHtz6Oq3sHxZwoqY
UjMuAYJy1MTKX1xyApnPC9gQYYVM8K028IZo5EzJ0J1uHCplABzkB6LZNG34MW8E
vyM0FPe9T+jFubK+Mq+MQO86luw+vQ3u9tshk7jBOXDGq/9o8/Jgy56jBHC18QGw
z1HmyCVYW4thUmSdowGe/Fu1/IXqzrwegO2r0LEOojwlraAMIAihLuQt/Mb+CFF+
IyiegEFjOkJ27SlmxuDrtE+vCQWVva6XH75uYrbkCIv/4ThBYdVaedDZLUhfufz1
CHSGVDWPsiTi4WkQGFYkLXiK4iF36PGG/qOpVbVFJk5S1LS7uvwg2szfpsL+hJg4
nIDKoADbkGiidhBGy+sa2QcFvgnhuo+smmplLsRwkVKBNna+rAhY3yB/c5Hi5ZD1
sUFXQ3Yjgtzk6zRNe25huYKLxx+39CWfo7RYMEl/I6z2+tlUKrP3FgcjguM/61hE
odRYNXh9z9KwQ3fQ6EToxzh/zN/NHwDbT0WKizqo05/u04FMIO20h7alzOi9fTjX
2Ctq81tYSNu1o34JCOAxf2VEbtmbyfmV9ZAG85ZjJdPHF43CxE9m1paLHP4L7g2h
OojwQfw/cinY3jx8zU3v8RE6nlSjnXV2a1cB9Y6avhjADbVSR1yqrd5FbmwmRDPi
ABR24CeRDUIRid+j1qrA7kUPR/9Oj9LGBuMwEA6z6EFCcRhUIukpH8cn3EPvhGmh
oUiigV4tpTITOT2BQ+wqlSp866GcbCoRaWeRHgJz/IQ3O9tsBVUo5Ahq/P3IusvY
bMBZFwkL6TENpoFoTNlbQ29M49jVQ2qCvK+0oEyzdosu4bA5p5LdI9U3wsAiFNqA
mSr1cl0U1HRc6Z/ZNE3iDCd7fdDJE6YIpSGr1kEz7Ga96oFuvY0G/fYajHkW/gQJ
pwKJVGvz4Kp3wWfXk+c5cKS2EhhY1wrb60WN1Hb1OPhvoSR5lrNL22x1cykDsFh1
jZRPcgMIj2eu33BHZb/4VNW1VeaLvuzNVU0ivJREYgoV0s5FNLofsM7jtuwxR5Pb
2gCkLl0rHV4rJa67bSPe+w5mMVXHo3frL7xAz19+zJByhJod4Pj8eb/Lr49GRnCO
cCO4k0mA5M7jnLEnnneWMfHWIBmPFd9tkm0VhvFhmCXIA1xFnQX0bHd4Zz8UneJI
9YMDnUCQTZNfP06P67/+S/5oZ+eRq7H0zmhcYUFmRPDhBoUZa74xtdWWORri3nGG
Eo3WJuiSQs208fcckiqOTgiFJfngAvnmyTiBLtdfir338BU/TAJSr2kmuCbjeufJ
629Q+FWoFMPn7MumTFYh7qOUDWCmY9fwW3TnnT5cGmif9EWbxWbMSxlNFzLYYFbM
6lLpiaG5EKo6ZDs+n2/RjjcugOKtXEApQYT/scZ+oFlo0lcGk+lCE5bBXDbJMjCu
14qKTgQ0WwtPRS/NYfW6EbyOBzv91k0IhwWhnP095LVImkk1YMZIdp1Bo76TdlG5
lxRYRR/G3L8hE/a1BP1WOqPOgRNDxhZ0P76fa8HrqqDrP5Yyt6IWFXR+487U0xin
NaivQYGTqufYNQ/Bant4x7+QvppbtwKIHaVhcthOYlLwjtIBRnUb3RgJLwgRXcv4
Fzl3Otzx2IaNEXhI+6l+YybNuu347DE+L0KCN/wh7sNt50IvKcxqHZYZOP4lx2Wy
ixx6i1s5D8meiO5SJw23h6xz9CLpTtjmxnbFqAD6c3+TQm8bDk/E7y0pQy2DxDZf
LihcPyLK9PpWHSG9Vl0t49iRUSfCBlJZ4YrD40L+1QN6/S8u5Cgpbp2FvVvdWu41
udyVXGcH8QKBrEI3YY1eymwuZm6YzAUlYmjGEjAOZKvouw4qDiHzcJuQmuC5uYWy
/8mEELPeGW+mxu/lGZQKzXn8p6odKkyaa9TjS2cJL8KDmca7fpgf5dMETZ7fHzEa
Ntdtio9g94awbeV+PX5MlkVmO/nhpnvfL3Dfj++EXWtOQclGfLTJnl1uNnVUIqYF
ZB9ZVU8kNkFuJIGqEzUz3KgXd/gdXr+XNLA3fyPVsAmcLxDCVKS708C+g0LIavPs
wP5n2IhJ67GdfuFzsc+wWb0ee6/5uv4m+xXFPdw3/ZGB2+aZ/vrQ+EflBAUcwuTA
G/MwRfl/OY5GU1+1nLWKq/HCuoOb762mqteoFVcRBrOu2x8yUfr/EqXi5P01OZuX
7l4Qh7xHpeDahmjoYeM7Ons2T5XAjKflNQlkJNVV+nWXEzHS2dktyPDDOqU2JQsC
lK6y+CkIQY/gssJO8rACm4J7RxIQkHWWDF+C0L2O9PXfO8t1FE3WkrpwvsObFKwC
LccOScYnx2lyNJiqQxtcAPdRItJhtom7ZC87KeH2uO9A1fTSf9es8Cuttjzf6HuH
+gk2M4cHii+k3nvAOsuy93IvwsQ84cv/o+baXnxiwBoioS83yJDZkk7TKTg9KTdV
h0jMqWxpO7wd8Leih1Bn4Eazppu1kA0/++iF90fYaucn/xglSN/uuIDT1c2LG51S
aZWg+bq5Zkyk8LYsbSNns2N5MAFJcuOUf85PTw/4Xeg/nepKlbW+4EwUJNc6Patg
9f8MTdROQVJPP7wcQ0/YOjc+c1sl7PDtsbmNdRBIKRCd4fGxriLW5SGxifsOW6+C
EZqebq8h1PAQhc2LZ82bQWkOpAgqOweI38X0MQDeT5eBSi37SBQ/A3TYy5yK9YDx
VZva1n+VCQS/QT5pn18+825Kh7HIEbgO6dABChrSYDltrc/hJ+E7l6Gu8rIZowqB
QLVGZcz0f/FZ2Umccjw0BaPe0n9Ez1atbfKCt9svPFiqHw+fJUKiDUL94OhY5A/R
O9ngVJ1ZcHGc+vxxGAQwuiJlfrpq2ff5DEj4VMRdGZ+sOyEXMHRBIPCxiMU4A0wM
aj6+s+YIvRiUgk4kQlR2SavJlR5xlZFsyuSu1XIqZIxwCAbWJjwJ1bzJjSt+uhAE
PpmdkdBKYRh9c6mql35E5wm2ePbS0UmZm/CiFAmDasedhmIfv3U/16f2KQ/wPRlo
G2Msva6fkC0imP2A856uhQ7llIdoPd0vKj+ky/negDDfo5enuWUA9j8S4JsrpGLc
HMOLR7cl4B1aWqndvlXciH+YTlRc/MPSL6OttU3eTYFB8idqICZVoXJl7EBEc0TY
o/z4+mGkKFt5IivrTawnoBApt4WLuSnKG95q5WtRggV/w2LFuw3cnLVcmBLulVKw
DVnUZYS9gG76yA1wxbCIhPz3cMEG7dxxRmIi5nlR6LGUy97o8LiUrHlimG9HOztD
`protect END_PROTECTED
