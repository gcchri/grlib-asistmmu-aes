`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5+eCTgRRFIMkfodWJmhulCVI509tXuFO2fUBilXlM1lk4rGYwcj9p3Vy0BXeJvoa
NG046pf+4FflhwHCXSk2H5JEcXrd+IE8otG2qkkD+OOL9r/q0VwtLocLInUD36g7
jmgXjt0AAyNUeCX/migKpCe4T/ZZyEOdeje6zHh7/DWfUuckotpaVIjSpPFW9dMD
+2ADG5hKBWY+BdbONbEDNuaG/WSfggsRaW3CKe0grv9P3VGLSYKoryJK8kgPXM7P
PPBcKTAm9jzZ95/lEdNaHaBDmfBk/v/hwrsSp9zo6kExDgfB80D13zxrWBL96D9Z
Z52SAJyTWvwrO7dlIL25VLQ7vDBN540dMTp33vTPQWxVsKEkZ7Mn4k6skToGamc3
52cMw57kpfsWsrTRmgGWmQ==
`protect END_PROTECTED
