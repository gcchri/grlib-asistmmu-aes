`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GTtkl8Gxz1TPRx56lLtq5KqIiAWVCQrpYuUi/L6m3hUEdVtRtm97Aj4bu51ivuE4
bKDEDS0W9ayRGhmZRBbhQfsjPQmvJEK5gtNL/7S77CMTFKEI+WQFvQNJU47nVo1X
EUrB3RQh5MrUeH6W+3D98CgJO9bu0A3kI6iWScBaCDmyjE/jqwcJmoOHlosAn97P
ENbPZDjcPPozyOcOMKd02GLKQp22tbag2qxr/7C4no8K4pZIn2139gM6JdiNRT4m
WPg95Z/albdwPLB+BOa94SdOQARtPJYTJ06LQbsgWOo=
`protect END_PROTECTED
