`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5vsePGWqPLwqzz8M5Nt3rOJWl0e6Tu9K+/fMTr1a9st07ynq4O7qG/2+xFxGODzX
+9p6t0oG6i/YD13T9CuYXb/Qqbx76e20erYQNqT6s+fKYq7eRSWnrnFoqpPpUmk8
svu1f7rdPVeSkDKj9oGBpwEA06gv2g273s6+VQHSO5GOP6wYTYXEC5ARVB+3pHCr
MPxvLBLZO02ytwmxkhjk+mDH/jCVBJSu8FKJHDi0OCuk4/PNA7WWpbqivhqfYk57
UHEIuJAixheu3Q2+22Rd5IJsF9YLMxqzv2ukXtlE3B8oxKfPAJG2V+1Xtq2SlAJj
tQWHlOX9+zUzD9spZDb/2sUqWxzXBm1kFF/HtgbYnbcnt1LOMApOuTIWi6k07uQn
EbIHZM0RY8K2Ny0DTWgZjgKYNfQYfoO2zCFxi6U4YRBOkVCgp5z6htw6mvhDVHcj
cqNHAZwfR0E5/YUNiFVzksb560vURuE00u6K7iFxKUY=
`protect END_PROTECTED
