`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RBjxL/fG9376rXUBoZhcRIzTGZZz+ZzmacDRzYpRKkec7ql7bPJMD9n8T07kk6ok
jbNa+26jF5xexkHFOXXO+M/UC3ZgqIqKAKcXKBYgvTm6eN2zYj/QyWd2a63uMCOy
fbiO8taE+mzQh+TfL31DAfIYEFB08t0Klrwd7bKZWkruBT6CjwSZpp2BnuIPstZ9
J0KZovJZXRuqOOo7SSTtimczVA5sPbzVwpB7CXCaj+E5bfWmvWHuh19jxHeCz/uC
Y+Rbg8PIPwRsWJPtY9xTqC99xU7TjBOTWpq93qDpsi8MME+UwAShv4rsky73xmCN
hQii+rNwFJD3Sfo58pnwp6zws9M+QqdkeFA1m1VQlAWRH61mUiRQ+57A9i2tMISI
SLLzn1xxbfo8KPVBy+9lMpmPYEbFKfWH7O4VTE6UBAruU+VRpkxrLbCDmH4cl6T2
6h+DtsDpzLtkt4WCBEhkvgdxl/4pJ0tc2cbjwDls/kIGQ+N3o5pO6ksoKaEWT5sw
9KT3XXQufGBdKd0EG8ADOlE2dGCY/EBiBQVosM7nSyY=
`protect END_PROTECTED
