`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tFI5eS0HAkdwVgd2HHNAg8zaml+VS0eEmRFEMLRrj/4/5ZpcFBWHK08iPg+PDGk0
4J+j5pSWp+IInWsofy0L0DuGYiPKQnNS52zR0DyprJch+igJZIWp6APSMeKIJCqg
m98Hhf/nVi71B2xqW+pAylUpwioHhAZVARZj5UKPlCJYPROIiYUKTGodHQEZyiKi
dsRn8I9PoS8ajH5Z6C86x3JCctRppwQc/uWq2Qx0XkczTc4+Ofm4m5AfB2WQ1Fj5
kTmM61IhEfzVrCIACbBaQ1mW8nqD4SThX9WMbP30WZqjf9NEvV3UZR7pWhKBf8Pw
YdBUMvfyQjQxNnaGCHG0aZwMWCD5JtwT8jAhgS8RK66TF906hb1r5lHwYWca/9WK
fcEM+/2DiKA0UMhOM3RVvs7zcMmkWM/3oVHZ1VnED7PzWZ6Y2TzVvSD1vAiv8RXt
sQ/aBOrT/MvOzZYGMJbVOFjiu52Z1v+D4ldlOdp48ESiR1+nskEHImOcAWoGWSbh
Lvi7flBlCLJXSHCD2f73W2LEi4HjFHJh9WQtBj/BwXaQQF3EN47uSaJqBpMEEy8R
uniLZFGE38d/r1il3lZy8fKX91++/NdRh9XevgdqxzO+N2L4uRoXcryi+oM/tHyd
uMPwQrRaMskefUM/qmeNtgvbxTUgDHi/t7AnnAeXdIkCzeWLtp7TI/zsI2VMj8PL
31Gy1anf+T342HAQVg1NMaEd79IYDb/qsdP5nOVcwmjfdaYXGGwP5nJ7L5Jo44a7
ALBnjC86l7VziTMC6UXm94d4E8PazWAAIVp4npQVQfZjauJ5SlW+Jt0p1T6/7YSf
`protect END_PROTECTED
