`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n4pwpjEEGFEe9gXLNgTutcygzi6uXMBDiLff/OBIK1a3i9gp8SfplT9J0VyvrDow
QU9u1/ZZSuSCmVXUyqPGKDA4x0ciqM6nB0/FxePfmHvX99LJmyudiZ7YFLxJtpfi
1bvfmomGeKPUqWPBQXgnOz4XTusH2cn+/8qjqM42Gd34M9+B3jaMGrYiHo5bGf1j
rLctpGETn0f4AKquaKg+PBXXsgMLEzf913oLFyTmtq8VGyQqnk0EjKrPK2/y3eOb
jowW9aDHQjk8XvMc1CaiqT+v3vjEmxal03yylZE2SXAnc9e7qW6LLd4aJEiY4uDN
FxCnhNB0xUL5BZ/I29UcpJCTkMs00Io+SIKv7JKt+Im+IIB9eBVNkNCeyiAG3s18
AcXO9uXhoXl1/2kQ5MerQgwg7phpmBvCjFEn/YHODsl0AJ4kLoXrcszNnucxm8Rb
/Dy77IJHAQKYrJYWyDbnueStgQ7YZJB5QY0vGKfu8oM=
`protect END_PROTECTED
