`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zt4DKdgkq3EQfMPyFUzN2ccZ/hNxUfjl1Wqx7zv9R3EmIBxU0K85xJI5ZfcS9twh
BGyOuxXaY1jsc2AVVGbzIIvnggcvhzYJ2yiztACEcawo85DKCiqZ2U2tKVTs8Qkt
wd6dmZLJ+dDHOqRLHEt0V/b9Phk+o59oyFd0GMgpWIWtUH7hp4u7grpCTHIPsJVJ
F8IXQigpllz4JCnDAeYj65qI386iZrWVA6G88Nm/5mQf/LaIq5XCGNeWIeOW4HMT
mLphlGeb9k5AAc9pjSniEOsCiM5HlLD9NqziDMsYQ+2bska3P/7k4FcaTID6umZS
hByaBK73LAKUApCjKPYffOAU8iab4TfydvKQIx0DBJM7e6lCQzkZ0ZMRxiK45vb3
YaHl7vv2MXyDNIqSbxzilelnYuci5SLoQf3EP7EzK3UEN800WRAe9VPRWXNWxnu+
52ACe2qnLx9NGYrD155aA4KTu/z3AnHmAhKFnPk5ZsfoVp1Gppec/5dlhB4kzdjR
ZzpjO9FTRWnYg6PmxJC7cKPNhbDsdJjE8Rn+sYsEjlod87/kSty7vneCwywpg2qm
GHIFn/Z8guR7Hnpp4osDTmBP21qEvZ6xhVZR1gso76Rmd/8OSHOtI+xB+eTETxSc
VsHrNNpS4lgT8QEJ9ZJ1mxGGJM7djoekTXmuLEDXzw2OECuHfGsf9PD4PQlienGg
xfDicDZE6U86qak79n60yHRIDl6X3dR4Ldq6VYktv62ac13M0Js1W8+ufMwhyvd4
cqFEfHBcrQjBqgC+LqQm4bTsiMpyiRN97oFNb5llVvlp1VluqyuCdY4LcZ87BUs6
pCtOjC+p7xELEP34xFK8pSSaoeGQHb66zh3ckQj3B/llqPfQ+Mq0CDrLBx/5rgQh
dyHM0ddCGjudHI+qURn61kFnbIOWF0NNwU+RoHvBSBkBe1j34UDx+QjBBfMufgRR
0Fs0j52KThlgkphXVp24jkgBDsPD3RX2BC8FvwNmAnf3zIXMDENBH86PsQpQp433
Ve9VK3lU+G7CxCvYWWJM/DxILUhH4k3KRve+h46Ps8mpyOcf4kNPhRS3KzLCssO8
OyLXwqYLtcvz/jKjOku9TxxFmHK7Nffc4yX97iNVld+FJwsDMsivMHiYVg+5OIwC
RxqIECsyfywgFHzSTqK9El6A8u91maJPvFOYjbAHPQ2PhzzI2iV2BQHQOPildjW0
DrYIgB4yaJ8pucDgx9+txHNEHJbprGBRI0QI5/i46AMUUmtPzL+174u8LDlOFAhX
AYvvYwxmrKkjgB7++LsKZcMQkcoXLavPsq99jLLPmBiEHDP9hFDlsG94VNc3okf2
HpPtmeNvyzDwzky+4Rsfwj+hLBx6vZPBGMK4CHEGQvbTrb4kSTxqQ4OIrSNWuM+a
sGSGwiXA0UCAt6xEUA3t2p0aMVehGO2XEIKhZ7ci+RfX0CZbA+rrolNb5Ct6yLPE
6APxEKJPQThreVIf4lhOts+9XARVbCjGS69O9D78nnUh/GYmvZWuzTrMDZ266ElQ
k/WINPevB5Mie83aNa2tJFMF8aJQwHlWCXvdclNXLake2XONcx5fFuQnkBSLwD/J
XZHsWHyw86uFxM2ILdUqnTkhR099avWfiTIOvEDbiBT+CmnvsAiEFDHEMCkU0oKz
/EM/MAR87k2nm7qu8JIMcXgLq7EO1OM+l9F8GjnAGEEd3HyURAdDRUxluZmr9VO7
TDNo7nf9jX7d5yWNxu47QcObacubVAj8Sg9axlyZheL3DuMQuz6WDZms3TlBcc8j
eUjfsgvPC++UqfBwwXSi5fBRl8R4566OXxEx1i6Mc0ipJnMf0HOghYqwNQXHwbnI
MsmgctZI8Eok8+LsaypMREpQ/n8q1KiBmN0ev9/LYZbPTLdGktyqrp8Y6Ft7UCAY
ntzy9mGcksSSEKSaAsl/rLW32o4CShdbvUshQrIAWn5DSlCVxIH4DHU/fdqRYaGE
KhOwpupR6fNrplcuUjU6c4HYeQmir6TtewBGuHIehQUks7S29OKcG07CclxaUtA3
e67UJ4svgK5lgsSr0IzkAaE8S4iJQDKdZddvCnfbf7BnZErBNyPR69ZL1cbaZDt6
2t+wd0bip6P0VVFphEeDGZljakiLYacXNCIilC5QhKOZoO0zafuky1Wg5LlvvpTW
tcYKKuaXszgnnxUnPMIULha9kQt/NzT5iK3Res/hvaKtZvb/NlWkJkyeUHuV5hZW
ZQj0/W2URZkbkIg3QZX+DzA1u0hLt+A3Cxp/uHL44EiquKLlnT6fWD2yUpylnR/d
`protect END_PROTECTED
