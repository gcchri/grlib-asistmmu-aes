`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YLGeFtPquKojZdnvdHeIfdkN2tWiU6QcMKRFeKmyYqiYpvspEa8LVXhDEV4+x9qf
R8at2zQLrBDSprkyc9BTAmg2jwQF/f1PwoCyb7EsA1bgXCj2sH8j4KHfig1Vr88P
GDIdDFUV/fVubHXGE+CYMbfY3BUQ8IMtxzyv2eTb+nLACnkA2zxynmPHuiC+kJ8x
vZWcvfvZr3sCJ788qMSNPr1BxB3huWkvq8vc5KjY47jmNhS6Pn2GJrgehG79pPY8
TPti1xD39/BHwHJDmJIeBsGU69iq38uQz+bzNIyOTuAl54WVGMaNeAcJz16RW5vt
zwT4Qkp2QA1dpvNrJVRCVw==
`protect END_PROTECTED
