`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LC29b5QDz4fVFfIgSEe7WvqiMUmYA6K0TpOxpgXfJUb/AIR0lI16r+cpUvKOsRd4
b67fNtz5Joh+i1bDB9dzbL/E9S4Lm0KtVMm0zh7Dl4LJuClKlrgmiit2oZuQfa0v
GAKolsGe0j0y3hTnDhudvg9BvR27d5J8bOXZyZqh7yFjc0W1xaWxIhXsy+UbT2m8
YkjPK75Fodvm/KSgGrZeMHkdc8woDnofpAIn+hcHfInhB91Yicomdapth585dg1f
Z3i9l1li0vmLnIk0vteIkL1trxYitrVd3+05cwzrOoXsxexBYij17D2oeUcaoT+u
PSORcEldbQ3e5wEAKhl+uwxGPOyv445h7GWSXQv1tqJah26eINETTYghG8V83pz4
lu8CpzcWocN+PCLFbTrBf9LeY92Fi0IJ1M0t0DHvn7pC2K1A7ICioadlfMdTnl94
bVJc80R9WRSYp5N0XkDOqjWxyxFQ3Im8JASqzyQjMjU6rJ3zurPlVqqw0883pORa
`protect END_PROTECTED
