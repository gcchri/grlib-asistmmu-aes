`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qXJsJfUAomdTIH8z3FhgXz0ppeM/Y0ot2sEEMFGXSs+KlJHKMqNm6x8G6DvVdnhL
R5grHyr2tj3s7Y/uCDdx0qDdGCtNlxvamNbSn6pUUy0O7lsI00d1U7eaIcnJr0H8
AYl1LTsVNsH8V2EcrEjPOx+/jX0UDQbq6hF962p22HzKvq10QQPyAZhJUDrnr7I+
Ef4FInaPmw6qIegCzXtRyRX0xokBTdsqRLelJ9st10B0J+0vlC0DS9L/i600+zCq
m0zeiw+tPcqdLIEPBdQ7rXPusx2m++KHzXZIqTviFZCuQE1QR85r6WgY19obKnOq
hCtx95RoWxYjMlp/q+Fqpo/NaoG98XZqQeh7GUyXpXgEAi8BUDEF4oE/puM1utc6
kEzSelTCF75cohWw7z5/OqZ9eJOfu7asbHlTC+i6vzH6fGdd9wJ/BUsnGenxZdld
szHUkgQ1cLGWUXszN4YTo3lFHygev0EJyi+0B4PzPdfYRv182SJs6Sf8iyRJTniB
0zGLtp0djy9LfudC6oD5haWG6rVCL2tBl9f01WG+2lSw9zU4hob/kCm5O4FWDaud
hSGPQrgveUg9VFOAJ2qk3ascqjfy3FHSbN1mz9tMtyrXlGZfqjYhi0JAwEUS+awb
hhzQJm7233VCMU7MLQhm+l6tzXC14nYSF3hGvvQjtu/d+6mxuTBXNgxMpf0wOetg
IW23ptc403N9f/XHBIpxvxyH3KlcTtxkpG+ScKkqDmW3YGdwnGJq08pGuUywwEc2
yCiXU0eSo2/8J0RlXbr24+zSwvlfOVUIpLmcYVv5HiICC5MfcfZNPASBuIyOnJpO
2W+xliy8DFos13KoboJ7phbolQ3CM8WcVWte/Y1mOq2Qa6S+C8b17bQauQLS98kw
4eoO474h8knafuXqT7LG0vK2/yy3jIeh6N3Ht2DVef5M8DdKGIdUOmqzl1uj0NA3
gSXAFMnrrg3abFw+a6/bfuEiREcdmz0Mj6NMom3ki0ofQisfHUuEd86XKNqG+hMh
h0F8TORdTyVNtV05lvG3qODAoM1m97YqfuAx0mFvMqGQVeRtBMPyCICq/yIXN3mY
p5KLaj1stqb0sf/n+OA3R/31PW5iQEIiP50uLI6eHSjztlPnR1IkSDSRpz3DTXed
UGSoVGWQVEUfXsmDxoXPEPb06wmENz4CN/bmPbi6gy/D6H9ARHQPYq6c/j4jd5CD
4R5rQd9AH+prNTFvOE3sUidEqKv5I/0/WNbQZ4Os7FzP+rGQiBUbnaovqo11NR81
BEUpKHn5nmtsU8zXA4RnsOUHQYRGC1y6pk5kVdeJBwmIG+G2nJCnW3VQ1t2r3d/6
j39p+vGhkfZrHaH9bHuqg55tJ9c0lRafpnM4naTUgdmgPyz61Ct/tCuXRnbIWruJ
wwZTXckKI4Zv/EifCfpsj8agvu5mgUtUcAlBWvkHroajbBw8/IyZ0iOaIMO2yh7S
wijrCHpsf/23DOI+bPgSdM07VmSMhx9JrGNFezB+JCB/5UVjYhx7zgwdAbimpvMT
w553wmCFSr6P9RbcmSTiLcEOoSlGlAUvU8OAeS4xmE9b+l5mXZiE70qxyPPJgDMf
20jToxgQUTzZUR3UbhwR7jkcSAyZL/jwr0XP4XhFdcJPVqalEuRANTUOVW6yhmle
DJcAiZLxaZyTQI+c5opeQ1lZaJGCpxaZTLd7g/O64r3gjNHyRHC8wt3/rCar/0Wl
H+Fh4DR5BlIz3cV7kk/QJwCl5o28aHdMdkFZB5CTHp+Lz3ycBpqQJbU/xhrQFrym
g/E35kndv0oEwB+2aLNVperWeiD2iMjCFub89nqwUvXv8vvoG2Ng/bogC4YYw5lr
ljeh06HY6Kcf5HGYySN1Ij81m2sEp+l2AnTVO7dUrdmS4TUON4mAlhi30bItmd0B
8xc4iqRMUDfRVdTydbVuuUWoKtKAwn/gou2+jb7OLZEfNnG5DBzQ5h5wDwpllvpn
iQX3CV4TysrViIlFJU/lMfy2GngoRtt7I/fRwI6V4GqCG3MSvb9RSnsTCFzYCTIG
cXNq+lO48Zz0oeJy7HlFoAEfeu0YPDG0fYsvBXawXQ/RFa8u+0izJ7ATdbIgMnZU
pDqy2ocINkAxlfJlG1rDU4nTeTkSm7zFbRqCLO+vVZ+iqvluAbr4Eaj6KD7ZtgDS
8HE/TOGtJsA+mt47jD8ucK0TbEsfzAU/m2I7xgLM/uOK2+E3p7CROIfb4SHTuiN4
CAAMDHTPa+BWft+Q9cuDDHtT9eIkXiwPx5Srf3O0wDSOEgByo17rQedibU2cgiKI
sizR3Ns8ZAXyYfFnnVQvxozNeOYgedRMupnHQwNEcoC7t5hlugOnWUqITmKsf1Bo
Aptz5Ecm+j1sOyCXXgiukvXzRL/rZiQF/VcvWoeOuYMKpZIUfZnvXc/Xtux5qrGa
uOgtMCzKEswVHv24B28G2E6y6YN99iL3+UZakvsnZs6t7Zsf7mjgFe8Vw4YDGwYY
op+MSDT6Flebw9GdWBdq7y/37r97dFsytU67CSPp0m1TdD9oCxIGI7dIwQvXJe7W
A7yTspFZde1Npu+sOYT6eZv3dceWe0kzFBewNaPGyMitV+TdBZAY3sx177v5JGo1
cP6kmCUigtSv1udBRg5xrQ2eY7c78yD7iZH91/4SHYWRJAzm/vuZ7eRhGxN35U8q
/UZnQbebSbKs0udyzUbL5SlgrdIYCrQ1D+2se/xTGoGXUMz5VXQDZL6ibLgc6oOb
Mc0LDR4cHno5f+ijGgw4TJRgZGhCoRX0f8cmbfVSsXmaJSVNAK/hpd5Lx9YDBI2O
uMHZyO9Hq7CHG6IiLd/cPGKmxqrqK/FHekMsUYpNcV3t1T6rScX6pbUYHmuG4uqc
E2AiRx5rNFSQmaQhBUM3LHG8BTKiDMy5d7gc3NG4VLRdcitD5QqZefnSGedc6RBV
PRJxJ6NYS4Lv3b4yCj7wTsGhAtbPxaTX7AvNJAK2TOgUm5PEZhAhrHe8EApGWgg2
/iIFk0fdWprHh4u8WcKNV8GD1ODqhuf5UYAoJC/X9W9YxYTlTGcCwreUbCDOCi+y
LJgmhqlTK7HaLV7Sag3zwFbduNAluUbE2Zk36NXea9SdjrdARCEDWuyPDvd5PsQe
X5mHsePL25pXJAwKgyd9/nW1vobjqbfeJjyrZ/ayveB52Y5QEfWgOxYMjreugQ/V
/+I8FhzTdjRr2Q1Gs7endWox2q/n7584zaMPBTCUPPigGO34TD2xT3+ZGuWkhd4G
bY/asZX5iakApABIQMk3PUtmlbw3XnliebTSxNkvwcXhqB+RoO0yAvKxSkn1UFkZ
+wkBysPX9DfDKBVrJ3jPDIF53gooLdoem9FQtI9abdAEaehAP/19l8qMQv5MuxP+
6mQgtYfiu0tVQ/tMQKpIZNW8z7o4rLvsq0FPC6CFBqokBM4YHqm1LHg14qFIPGEt
znHSObuKaIgk+200LJ/1VdwTqrkEKBqqAgwievMjrm0k1gwkbG0SBaauWdkVw87N
KYPs5iD+3I6/60I+4mHUUof4b7IGj9cWTupcM9EFrWcc++4jDj8gwzbUlS0iZXuN
f2G21THL9NzklSHo3VKv84TsSPBsluChS3jQjfJ6K1oan4++KPs0es2GM2jfVuBJ
kcwRvEcruRpfcgM4j+moEKldBo/q50JZR7K0B7aqcEHb5B9faFPdH3qQ1+062n97
A4coYEhcGWOTV3T/VkxuX4hZFqRf20H3uk2dktLprHWEbbOqfarodCLrPLos6Mvr
LDqSHV7FbjESzDI3HLfTbOlGh89XYxmHY76PiLlOgtzhB6vawF87GSdMfT7fILYE
1HCHctNdoAGEsJnu1DqUTJ4LZ0dkpF8+IHNcY9HKtaBJzh0oXxYWq3hh1w7+isT5
3GcKteTLddDAqqd8/wGQLFj4gu4uLY9mizxueNxlgmIlbxnCiIz1XM5HMlC7bucY
db2IxJJUi96qQXqfMQgtTwrAuKB3de01OVQhVXa0JTNdpFNRtMs9UH1PXJli+4JE
pJEyyzTZVw6hIlcHOIVtcZf/QgMOGBlDiLuIhVzuOAaDlcVqPM0tdipD+oIPFA+7
Jthkdfe76Dmn3HHpUTNDq8y0Uaxvd6+9A4PibSFN4A0DJdqfqZqlr8Igq2Q0mxow
fq4YufucQoAtcOF4XUrAjRbb0+8Hi7uUpDa4Ey0m2185f20EI9WT+97yMs+t2N5z
0ifT6mi8Gq8P9Wa02BpLEA2Wafn9EIBkwt/Yq2LHae0uuvYOoaOHvHPuRoLS4RFy
0Kp2gSlcgd2TUZtcOBy0XiUqOP7QdqCZ0SW9owyZpnghYVgIgZVryPZS+2NYZDzW
j9g18Qlmj4kCgIgx/DCvp+6RoiusB3x06DYr200nABRt2yue+3W5cHAX+UoJSwwp
4n0t/6HtirMOt+phUpy8Llc9H8a1F97y8WROpooAkh6HjDsUjnG6u99mohG/gWhe
VxzDPXOalwBF402ej7cIU2eBxrYZOXkNHeNc1fsIpvMiAUMhwtPclmbfyzbDrxw+
OYRPAFNcplH7WSNBz0SKPnycNbbXm9TuxAOEX7gTmvRc3eH0uAeTXwNZsZBtFEzz
SxCtaLUM5uM1gu06STUhf8j3WLcEa8oirScRxAbTilfxJFYmYChKzsAVHZ0/kfA8
KEYEOPo1FMUEZ3nEzI9B85YoZwREj2rkUe+l7xC//Oh+gASDUxuGfFsLnymQg+tR
AUg8qSKExme1irmnlkGJeQWpf+rYHV5OeCH1WBcCUqPBogjfCMhdWM5ypTfSwYpT
npK2B5Gi7jh3mopm7AIK+aL964owGA0rUToL0gbOP9g5hYK13Tkog3fLNg3/H1pX
SBNNBLMy0hc3s6KuXXU7dUgtDzrkFKyd/7exjdkWj3wglMbsncXA7jXM153DcGtK
go7INEUZGvT6P0YiDZJYHvb/PbbUTyPL1IbbWbVLPohJcNLQhFg46dwdvgQl7w22
PygBoGL4wAC3vguk578FLKG/gRvwhD6zfBKwTp9AhbUMTRGLEVz9HnnzidezMQ9U
O0bRkWxWv4tJ8kHPAKCg95Lcy15isWcBp7kX7ae615kMjFGjufS/GN5vQnr8e8dH
m/Gomhxh4Pwt45LruOhafKQDKu3BzTiBBeI83r+562uvTC88NGMjnxUfzUPOKDIT
1G2F8bBDW579P6OcZyIY2/42eX/YI1dN/tXkN4Uh9SwCzqYr7pj9bmk2Uote43hi
EqWYWcfC7uv7FBWDQ5TZjJ8cTBnPQJtJtpDygw/BAJN5Ye13yi3czSQ61MO2koDB
z03l0X/R3x8/M/OlYSceMxVA0gjdCGtmeWGvM/ptm+h021WLsChVORsi86pBoLzX
T8caObsZSoHumwBvRUem6x/8Vqqo901T+l/Bdn/n5rNwawBkIQFqVOyT6ycg6dIa
5mTIbF+DZqnvaKVyblxLnlrNiS9gc8MQ8RyMpaEJ5xFo7QYBj041q4mnrIaminQs
vt/AGuVxXq9pybGKe7oyV9v7NpjfPMtBmQCJ4kvyl6fqagkoUTIMquJ2afRt4M1K
R6NXTaf4A95rqK/DwHyBAEIlAXbkmE9F86PZbJfl2vRpejsCDpQAqiuU8wQWnAMt
x6vd4obc6KGiHwN0Obp5QK3Z694Na+CEZVsT1rOIMW7033JLnIxn/Besj3sNZWVh
6J1jhO7CiUI8CJ58g2fc9zxGaY4lqJaaam13BInlElcGNvxNauwDOdcL4JBsnH6y
VfkMNw2ATtGZOrS1wbVf02kOCvYjwaUGTx9Upa0ow93S4n/zopa0Hin2/Oc1OT89
JnSJq7QeylsWvoJLDa1u+QE12FWYhi0XdPEZt+kAej0qRXP6KPvVGF30R56qUpub
tS3fN9MhlnKL1IoyK31rwQkJc5d5XdZlyaMnfikDhejGvB33AXyX2WLhAS4fxYVc
OAzwgxeB/5Y3y1VtPiAXWwr5Bx9cojmXNGDbHIeJcXpp1JBuo3uucLB87bavNIgi
Eh6vKAV9mSK40PMDkXtsNEaobZuUJCxLkfC5xThOD3hcQCjHEiKRvwqonPGYBi4S
Yhs30guhY3MNw5Rpe+pLQwYCC1b9sXuQKDC5O9ZN7eVHS+9rrokMnSD8G1dkyEJC
sGv0IAe0ts0aumU8HIYZfsIHEe8us0XXBsOZmhH/CdLVuKxJsB6976GYdvzgZh9g
iiBZHAeZ50ZAANiYAPJtL3NlhZM11l7wwGtOBclOvX5lDNdXHb3Tzy6SaluIJTlO
rInJSowoGDaC6evYFE8ouU2EWjWFCJlGgLPhfKy+aXp9Jwnn4pI8ULc48dYJYCEn
F4RzLnI68fAw4QcfPtIhpD/oly/OnWA+uZoi4OU1/Vak7zXq4jMlY0J44bdSTD6t
eHGQd+6MkuuEFXno4zWLSWU8XHgHQyFM2Z6cJeZG36NU8PgeLGoqFypLTT3/dtYT
RpVeaBNrLVckMRyT9IQNgYSTmRBeoqkBF6udSU17iX30evgyHPnvJmy2r0ru/ZkG
+uLJtaAiu7O8vPX+iqXtbjXTh+w0Fo3poWOSaqg3KzbNwBqO3mQSxGGZWINnK3hs
lRy7ypO3nmi3KVY52FgWh8Rtjf+DVKrTcvUce0pWrnQHM5KC+4/2F4OX9J54lGhm
TJHbdjR3HyIfhrBKEh3KzaGE4JOYsNbyvjyTUDOSiiYfJz5yqRDT3kZ71UtBCjLG
UTVwM6JZ9zJjaOXB4gGPZC53fKAIOAmYo1nmsUyn3hX/LOW/bW/sFC7VKLuvdufg
SBD03VZCOvXX90zYlYBvjGuapJM41aammR/vI/l7lCoilLozTCiVnWnDaAhIJy2r
F02AFs3ERvxsWZtjwk9V8GoHhCAw3+Qvg3Grd0khlO5oZMv/8rBNvUx1RQTgsCVP
ejxxUam0ftM4qEGQuNRlzhyatcpy5M0BcALPactQdSWbHS2YAp5bTLvoTFfMVyMz
uYyPjd2fgdBtb/0Ag7T94jv96n4tPQslhgwZ/1e5pV3djCkTga13GcmN3sFhtaju
mvij+p0sg7fRiHHzJmeUth8zJYxdXV8vlDjzz40xBdAc7WpHdVAJdJJUqxl3DJVD
4NiijWEmt43D4Y7kFRzhfq/cK76JLdJF1hDPoImYpY9TaXdR8u+EWxfbFVOjfCX9
gNrXxAk4YqeegbuKUu+3bBJEX+Lvt9Fcf4r8WeYkdwK6jTv1N7lIbGQY/OqKJhip
68YIroR/jZ0SiTD5LunLWs7Zz9Gwkmhg3/uxciFkIGuDxV8VWXoNt7B6l1ng4FoO
4UBKqXkV/Ugc0IhOuHg32T5cC1KqR43qSZWDlRC0M9CKvE64zH9/dwq4rlqT98Jp
yZUUTLQ0fa6nIz1h6eW27xxwcYVznN7LHA2HSIguYiJ+RzxLO/TIpm+z2/UW5bjK
yX7aq+387Di/WaKneTHJhi+yRpkC3Fbahnjyu9jNvjiIOqRxFdlq4Y/AnScNd8oz
8CxFOslJ5PGLYKrwipGCsRmeVZIxwzCWenYHwfmFgfZNnOIY9Or36FvMnRBtcnti
xscFT0SQsjVuz0hBLaVFD1YT++WwTQQdZV3+2hkLcPqqQFZeczuTQ8PVEoi4mMNP
FZjzM1laDNfj0H6ImGtxd8wRVZHjehKCqK85NlGv4LGzc3x1jtvKpu04bwK2LnYK
yRAFkmxb9tud+lWFW+0i+yfXWznHyZty4nQFsUV+wnje6wE1m1PxQMZrgHfOtTkU
qIySHlLbjgGXwEb3m2b6caBWInbCB56F9xe5iz53nK9nMyZpixvjwHkHg2gk5tH1
O1hBkOIg9sieYtDW+XhDSY00vy/6jLkld0HL9FJCiQ5E9e+28VOWFMEEmm9QwsKe
fUbjZdrsM9GktmTJR/GaxAy2r5JZ9fyL/JlTMz4pVarBxIydxl7NWlEiRk7hRVU9
wlbKPNuUBdnxyYGdw89BOrqpd7NPPxQA0ORDng01tzuydJRc2H5IbzxjBr7KoyOD
1fD4+UCwEm6tkkWE2uFmEEsrDZOQtP5rCKQNqGnOonBLbBY0fwfa7SwTXhdlqxcE
vZViBxc+BiAunsWhADHJVGUiXITa9MY3VUHz3QGGkd5rPzUmBHfmlI4zEnJYU+Hz
A9Wv3gx/NuBCFXnIwJ0JM/QbMU3CiedbTemMQ7fIHno2ZnU50CX65bLCWWc+LDnb
WM6A6jCKJOub00uZpQ3jECQkv6XTr4QL4Aw2ZoX63KRGpYabAoiTXlwzDZYL34+R
1y4JIZs+iq3vgng5lXxKAaiko1SWPQihsoPmVI+yAFNeexjm3/Y+L6BLKbqUmjx7
mh4fjxBhkCDMJpGhxPEIgxnUBIuQrd6QJjz2i9lJgxIMfXOvaawlDenOnXya8zWU
SDGAgsft0Hb4Lq/l9AubH4bLCUk/IzmlofQiHoz0lvQB9viRZ/LLIjHW6FHnveb8
9Z/Vbydj31DRlaofXHnotaQiqLtZv4V/GTzbLYHlSYUfX6XrTqcOZoUmf7/jJAfc
77VNLF11IeTstx3hqokyOJC42uT2LJ27d/C30pLnHtr+2DfLIVgaUgSLbpiP9WKQ
zX4O9sOQzv/3xLTXU8qeo0LALphx0tNn+7kfUAiTBzZmAAAbtau49eOot+/he/6S
KgA3KlSVEXghizoIHoxZHunjEKzDzbS8QiX/3YBqRZ4UQqlnv55tQtq1wDHTdiJs
HJIHFyWIKNdBa/dtY9X/7oSbZnTBwsxcxcr5VvHJP4odDZb6rOsiJn4O2aboub8s
xSEZm9BIjKLHkGadQPwGk79608XrDG7N/+YkLK6oIGOD27sz9DKT3I7V/MrPqIpN
43pCEAsK47E9lnc5ryzGL1uJp6+HWvbXRN62jsrmUT6o7ImwGV6sowp1jfVkfYtL
0q7Nl144X+gOVaHK/d26oy4zbdBAGaAoe1PmXlpj9LVIWV0nwXjtHg8UFebGhWL0
HlH8+ma1WJ+ThifJmivI9GxObwtGq8EqsYhhoU9+D0AspzhIZdF0jlCYjhLXIEsY
Z6N9EP2As43IDBuRqFDsDVzRYOoMmg1WmtkVPLoqMuTBK7fGTTEoIWV8u9SLUTwy
ufYsQ551+3ojW+Icsy8v1vppkp5u5ROCS2mljZfTxO1FJg9o7S5P85IrtQyjv4tB
ha/SG/x+IImofEkHLzy0JitIpFaMlOr+YhSEQSpzypFfdKr/6DOb2HEZuh6jHxE0
ZcQaex5y2YIFlgNAZoRyYJBjGqoeYauvoHxLN0kPgEEWo2Je9lU43N6kA1Gbi3B6
ZCzZw27F/QRL9XtQ7VYmDjozsXXb8oGBhqEaJTU0WwRuAa2rZ6Jn+opXRbo+B1Cg
jhocQO35c7Kbq2KAkV2DWOJuSFaqPFriRyXfbJ/Y1YMRX7QbFzSBvsg99s7ETdXi
i8wyGIk9X7fZELY3l9E8+HgVgUc29i3RrXiNy6iPVLWi7XJOPua/Cg61kFtP3PtV
XkihupUFEuM9goDOc+koh5gub58z15qOvgzVKqRQ7hW/M1kyL7DyHK5fDR4VksdY
YKU74sbXeZ2xWDvij9FYCQV8IWcZCyN6qBG057uosrDkrL23t/yZMKI5arQW1tTe
JcO4DjR7IBpQRsDsy4ONvvmNyQjIvvWQz99pTZYRruS2WVs4eAlg/hwCP/AIsImM
hIVAdK+ZVeY903qLlP0xG5+ud6PO1NTLMLQWXoECc+iMispTNTmG3ibvjYJuJdIZ
IImF4VgjJPLU1VelCskRgHc7Q6RPKvhQs8L1+OKcNKSEGAXdN2nYiYy3NxosRrVI
4nOa4dP2b20m8cWXSQTT0Urhfax+qSrJV3nICtN0LD3UiVKkP7y8hlGN2cbMM9zS
qN6FHIAdZKO8cjA8Hffl+NgQy2mgsZveUWOb698UTIRiIJZgmLXUZwDlZLSix5t0
yfSyNsCyskfzaJS7knHPXEVs9RNMPaCqmfIIuKSLYtEp1RoRzY6zH+DJi9+Q0VwD
S1e+JKNeFPYDszKR2SbzRVayUqfTlHUWntIT2r4EMtcsl1kHaojf1ZcI+8taGdaI
9FI04/oYV8l6pEhx98ak4Fdk8HGgxEl5GMhsfOC1POKjYCmeMZkWITQMFAdIP7vn
ZMOTcoEqUiDFDpiUC+CRPui9XiR3EvOT7R5Uk3qmoRsNiBhM37V5nuIDa+hebkGc
Oj+dDe2oZ+BFHy5lUVrVUAEDpcr20Iaj8eb1+VryQ8MWNMSDxjGXZYAcRSz/x/d5
8hZC+vCFpgp0T+PapYkeG2CBENxoxBl66EZqQ7FXMY80HXC45XCaGTDhosx9KeL1
cKpy68vzzHbc0fIeC6FH9kFTPa73XDKPIKWmOwonm3U6r3+OHvYq9wq46+cGuJ5b
hoei0ltwrNeDdnGMVIemf5ii4bSqbs3smVM5y776oJ85TFtohJmTsFw0t0g5suHt
oe5krfMCVpYUTXSfzefcO61d4c+Ua9NrwlQGKuDSH3c+L7Jrnk54v64GGUoZ+9vb
fLscTFx+U8VOmEC8Ekuh+cqLuYHVILRnbpubOJQOtZEyGyVd9KXDrE17SQawxR4G
LkX6ct3ruJAOrlqQNE6um2V95KpmdEdDOWIPtA3CQ6bjXKqqGEugM+O+3HwslSoP
Ph5cU4eFJTrnMXmt9Slsb7uguBJFf28DRN1h2lteffiu8xJbyjZ3Dv5DUu/LLAhn
dnHBCihrYSbS/T3KsBMY6Bp9jLfMXtkDiERdqDRIfQVdtEjMInNhUp+sSCasIoHy
RocQmfeeyanLIc67HkLRfQDvxKSvpOrcM611+ijKRQTd7xJN37npqW4eOjgidQ3B
6rExyHxQrE94YC/mbnxh00zzxgiWCernKEbdX9K/MEVTihduNRbaeWBELfOrCPy9
VQ9pAj1YX8l1XzGe6uaCwdWwsOs86HA9uGtNCcpTZXu36/Jj9I7nuDDpWGqhSrCv
DpjIz6/IxvitxJ7cI4GKJdaoRwOhwvad00RcoRvQzytzVFBVCtpSy4F0jxhGbZ7n
1ZMmp2/3tFfNvLX8QxeSitZuSfsILBJXdR7ApystWgk/LbPs4B9A8UYUco8xd0+2
CHQD5HQ30pnrQM9N6N4kODjl4MW8l3VWodK4oy3Qxr9CjJXMV5gSP8V5Nm50b6ig
sG62CZBdCJYpT4e3Rk4vxHAPnUkiucHfa475DPc4Fjv93wFYNDOifXs6CHpewcqa
AZA4uoa1M4L0haxsqW4f58PAJmVo1ibGiGAeoT1RB2czpq/l9zgWV4EZRzfnVzM0
1rAHFzMLJA6ucHKwGWtGc3rV9k3uQjgukmscO8beyPrE/IAZX96aTCnjwozhVHEE
7Fffgi9hLQwYsY3htp2WcJKekb4LEq1kq7mwh3K4dSOq30bK86HIcJ1wVQRJcId5
o2HcC4+sJF+2D/D/5j3Gy/ke5Iw9SCMSxDCx5o6YrvGpjB+tJomdF58YiL9MPFKg
C0SeJ9pfaofTXNDYOb6NYlTOkGPnnH1k3sV/++BtRckRtBMPhEeqQbj5gdQ7wDNL
pdah2omEArnhWwjHSPpmqV8nD+Z8+D/BIp9/Ka5rxCDwUt7prbRDhtyrbVY+Gt0U
U8cr7GVJgdFUrl00DZ4UAwoJsVeycREZ/xbY6X3jo/xbFVBkNHutdUrHCel7Sjm5
Oy5zs5h2kJsoyL7OYw8gzjiSUXYNzOX+AAe7tPYVRYJ8hzl960kmGKRcp0LuCWqb
kOV4pJ/M3IM0v/YyXLq6e5ty2R46eiI6LzM5kUinv4ag+MQlos5B89vS8PJoiODH
QKqILnLlhIWZCZKT9txRE7aJjMbgZ7ktkcJ+NTJw7zYcpO07AJ00AwmYj8TvYSuh
lhlOThuiB2Zn8Ve0Sx80GVIYiu+ZxglqB4LSzDkbc7oVfFugKnWoMhEZmpA8mexY
JXlRRzxpMYZEe70Xot/eTK7p+EcHEFmitMNVee1EQ5PdGILpKRExng2gB1mMUCk3
4KIJkBrgsMTPZZq20pyCgjOWS1670h9iXybwR84fI/pHj3lW1gmCm9WC+8W6CkNJ
OuGVB2+12YhPc2CBDcFoW6vZWrtqshat7y7qjhoXjYJv3D+atRwtVvPJkjD1/sWP
JmMN4ixjZZF/Z7tLM11Zne8YoVMDa8OO8pd0AmepgbbF1rb6WZKaXUdA42OHvWk0
w+cvX8AD0isQy7vHpMgNarus7RpmID/c2nB+z3OR07vCKa26y0B/iSuu3kNp1ryG
5YLni1nBmygR/yO/cpt7MKxZCjSx1wrgfZh+gA/PWPYwaVtp3hBGZxRvhSlfp2oi
/8qpr/QU5Mal4afPu7CjYCklwVzQ65Dlj5CiF6fRDgjoiJIekZ2yw4t83FB6oX6z
32OtIRDlCqGkFXuwbo5lZcAQ6+iZjNrOUBv1/gmkZ5kWrjYFNKPSV0qHPZi9TjK5
Nc+b3+QNvbgnZ8LS5ypHvWTnLTN1psif+oO4Hezy/J0ONwRcngvsdbcecK4z6dGa
ojIWaCQ8/Pz7v+S3H0l6ava8vxl9HjAJRIM9K26kSYVEmI3JIeBSWOEtUNyRGx+l
sAhkICB+3spHqX3CoePqZ1k42DpsP/bnkLJp8aO9csQCUwuSVSRf9nkyENOmGuTD
/H/wfjy35WGk8mdZSEQnRC1pNfqDIl6WdH9l32h8Z1Z9rXVet1PM5+3apkRq7qmz
uy498oDaDm5WNtkRozLn79TX7OFJmPHxS/hJ+QF6c5gWhMwUl9aE4U/3F/qF+0Nj
JX+g+3BP5o7SDu7bFXqMDeRYSHrXe4S3ZW4gyxZxJenU3zmLU0a/pOo0j2Zhq149
RZWHPcRhRMDgvLTtaZ4AMTsiqsEts5FqyzTvYqHky7uVN9o2O2ywA/MhlzIhhpRy
9YIEI+rQDnZVUUC5W45ycvc098ZK3DEU4hRfp1O1t+dhrqZdEEsRIdngdq9fN/Ma
iGz1F/ml8QPwF/ePvGlykTakMlCi+AO/FqYiG34DiLtBqXPDKw8IfO6RUVeNbE3k
1hSykgTFJ3Gnw34HzHXQeZBvOmo+xjXDYRMGyezpGYWGGTwZc0jmb381NdAOzfpR
Iwfh/FbfJDWUwkZgLeHQ4ot2jhMZw97YfzSgkQnvoU1dkOH/bMVojz+mr1i8IJEU
12N7xM+D9KPu1jZy0j1E77w6ybvoBiXI0s2fmqi2lvEb8DRN1hSV3kUfPUyC1H6u
w0zEAR8+IZT2eOdQzk6JbrXculVgY7GbTVlJbCsKTc8LiXKOByVczXORq1C0DdWd
lncxz4gOUrxNjZ9ltg0BNSI5Dl2ZPtaMtJs9+PnNiKWz8bs2FZALnkKiQA4AWpdw
wu2qtIxHCr/W7rkX/OiFdMiMTkvN+R8uzTXXuylU+vd6sJovJrCaR3qcwO7fGpMJ
5RPqQWX1JohyuMbyao4DidjXru0mC1OpUYaxU981/N4Fc0NKboK8lKY8e8i0vPNT
4CVYOlIvUlFHPpDBWje9OyWpoy2eavGuHgaTBJGgNNodFkz4ggsZg+BAxBYfiynm
i3rdshaBdj6L2zfGvIQtBHjrF4m5oVyDQ6ewLestTRECDQIp/sOVMbNW2ISZoql4
o5tzuWQCCrDX8KjIrwZLtyqbBrGRQfEzTAI6QvtWa3u+RNnrU7NGM7LqtibjGMcs
o5ZyAI/02hx3mpqNUOWsqjSF2K8cfHiFGWNE6a3j7GX0YD0+xF5BN8VeA2zI8crI
mQKMMJNDQ0B3xE+pIGY0nzUHAaxMIb/vB6HoZDnf3q7n+G9kX2fC7vcrXWthbcVP
Q9XZKiYs+5By+Ql8OZWD21MB8TtFoymaFfleSaobMO1Pt7E7RBeK/AynynuMScme
5BDvjW2ThtfA3R3m4Eh7C7QpYheu4EQfPn8i52HfNIXtyR+/OsbxlGAdFbURWvbv
AffopeTPReiIZCJYKREmJyUHYmaj42Na6Ne+EjnL/NFpxmw8HGDCa6gqr6I9dCbF
xb3aUNdSd5wtvNkp1H+bVUcqHO/OS1d+zqlS3gwvyKh8pDJyY3uPOQFbIW9bD4zN
k+G3CN5mqQBpdVsk3a83PnYmtjlrJdsojC34JRN6oSpUDmmxNC5GTrBfvW3bdKMA
P5KeQRdGNPYLUvsF4SDsZRZj+Wl3Z3T3YwGDllySB0CO+gSHqm1RbdNwbxLBvyLJ
WBhc+Qc0BwAocTGMzVUIMB3kVFIXGT31CawusP1loOEiJHSdeMtmC/JZCYQUHEkw
6pc9NzVAm2pEMKuVBbqVBzZ7b9aCzZqEwu8Rwqtv57E4pZ1Np9UsuvlFL6dfejAU
PBci7pIgLtFTP/zdTjaxIwYfea9tUQXdn3G/PJhChdNEjylcCfBS7jCxgtejfusu
2B4P+mdc+iTEAT0sgnJcBWIzmue6FD0WvvW9s6BbR/vewOurDAKa73laFQ6bym6t
sl7ADdjpyCoeTd4fTps6kH4WnrEDwE+70VyP/HorfoxfftdQ5/cdHLhwWXTeZkvb
R2eWijdCBjckeo+aYoifU+h9cFaGFKj4QiGQnKk+0VEyDFT860M5ogIl/RSw7mpH
zwCsebzH06tccXoxYCXQowSTy8uTUEt6PNovMzN2jJkQBQBjp1BGTczkCbCBYfvn
vLwfqW9Bi+dPzZV9wujZvrMkJGTIsArnObl+14cm5R5KlXgTItyYGlP77q+a2Kay
fPEBrXDZFjSaEwGUzHPbDfVXzNYYqPMTXzTiAETZGgBlQ0tiYLbu8OHrHWo7zj41
CvwmBaDZtwdzL5rXSoRxs2GBHxq3xjBv/6zvPcb3Yr4rfJ/6pe/boIgJrii7Cs3W
WOHfmrdsU25W2sT98W/viMQ/yLRIjmsVkKT43gT4fsxW2qdPdh6FA7gGufKnBVI5
sRJVTcgrGXvY5gtX+Y8gaBamJJDiJ1r1bUJTyjsiSn34wwgID4zuRvpvSeSv6PYJ
cwr9hXPJ6cac/stSgtNKpRPsFBTPIMxRkW36gtqUVCJIkPbKp/MgzhXnKPOy+t38
xWr2mwhZaDo8ilwxYuau9VcnYlDrJcBXWoQ8cbw7IdCw/mkDKUsVIBjyR56Wve25
EAN4PpAsZ0c5HMIPq2hsxx7MkN3vGAspjRKxw+Ik21HVzcDPPJ2cH0/2MfVV+Qhu
IXMF3vwrF0N9TobiB4NjT4C24JzTbhBA3nA556UJHHVs5wj6iryDVV6GI1GgTWCz
EbydwlNxJWeLOxjd1mLhNgFXoPDjzakxFoXpyccfmtqHlSzfOB3vwDK2MDWIEs7B
Flb+2u+g19uoHdBEusPPSxWRctzOzso4/2zfp4GsZg1GaGTX4UqKu/g9aIeXAiEF
L0wWjFC09WatzuHicLssTTl8xLOAK/iMgnppZZoga8QBA9WyvWklzb4mL4fz9Gro
EwS0lJIBznolAr+8+cspSmXK2MK1jvEPzO1mPlXsXQIRAnXx53veN8kcbQSS14iW
clzM+LH7iQizhcKlFZU8zsTigLgEhsCOnxdJj2QOk+vXP6Xz49HC/Ofh1rfqKZxc
ENpIfQ41emxorYjqaXDpIVgRACgI0RhVtEjBKt7f1zoljDr5dMI98ArtCm8FppyF
E3y5ecsYn5uyVg7bJhtz9V5Ls4Wx/cNhC/g5L+oWZ5EjgZhJeaHAwlpaGE3qyWZi
//Xfoxivd5kac6FNXJc6AcCdEw8EfaR8hVCdhDzco/dvQLMKCNUgjhYXswgTbiTh
paInvPYevtJc/vtlzzH7CiaKedMTwd8Jwas+SKEzNOlNmQC/U5h6+vuA9bhuyms5
Qs0xIL+ksk10LLQt1GYqODtmw2eu0dukROCa0igmai4w3dAQXNolWj7Q4y4SdGQa
uwwXPGPQ7s5PD0nmz4tnVbUMVZUqwyRa61AT7cMlo/kqZGsd1JhhakVpXmcXNRW+
Hjw6bFzM4LadpG4qpZ+mEkMD3LWlzR3ivRXqmmM52ybLQJidv5g6nDLvGJjzOfRs
rO3ZuTbxpTP4oBo0SJMsWulgQ9UaPczIZZC9+JNN96raNg5waWZT9dAanYJJLX7X
jCVtUpNGVNPu31VOH0tRApBegHg4X6vcsPHbYyNWrzPNqSW9I6roEM8SZJBeECt6
bfrpVUqQXXAhRTNxVshNpXlt+Ss6bO9z4+q33VdJyX/ofjJOyLEaaCJpnf2icnsd
wGcE/XE+uIM1mLc4k+4uqFWONktf8E4tyCySWUwi3bZGN5jZGp9mGTs5rBB4CRk0
LJ7im84jdZaU9o3rQREy+VYKPlyJOwcJJPnWkzEBrilJPiuOIW/9ekBVXrBZwwuv
b0hztlWie+c6WSE6NtPr5OAs9b4jEcjH64dlqlwBgET3Onwu+kuBSHc5oonzvIKI
8t7tl31Xha7H/l3suipyYfK7eIT6ajTXuM6ptLL7w9woqczwNTNF23wtC9k9AVxi
MNM/yZVgXZuVMzp90iTAjjlB/uplhxaJy6mHHFmztYeoAWmL5MgkwNXtPEeELKci
mClnX+CC5RCNbL3/PBkS2LAwZHEeznq6PpyhfXZAXeIw4uS+ngbiO+oVZ+NIFJ2k
mWzk4AS8ThP1MsfdV3zgjGwHzThzhoNCCkvP5bpNCZd7mdnonTFOp5PwTrl59ZEA
0rkKZYFOU7fTwTefsyCaAmdm5WJfkBkczVOReaZzZfxbo0QZXKilddhTIYLD4Jaz
hXqx/XgBp0a6ZoPKlMmyUFU2cp2MKtk79Gy54D5zEmaypTCQNZSjXQpN1ztwkdIw
8Yabu2WJsIyAWdegVrb87/iHsnR3/wbBjQDqwrH12zBqBva/2hbOKyZ/OPqEE5oG
x33OR/KrGOFli6nDOYzT9tNmlU05ngjP0H0kOWnwsOLGxCmlPwZBGzOg6+UdEnW5
lP2KZdW0breJTj/CktHoeZkHaheLIlMLjBa2ie/IQzrYkapKykhRwljodsHME29B
y0pEemdkreCMQTL8E24EKnmduLq+Uwfo8dYDfFjoUHoxKvEFO6k8j22xBqowti87
E4hnB6Xi5wln9Nkb4H+gWSOgbG3RfLTBewD9v0lnhTtYl3ALV2RlMekc+eyBVItG
X3G+4xe9N42yxtlqp5K8HRjfWJqeKFc+m6P+ip37Zi+FsC61QhJAxQLMX534Vwwk
Pedn1Rm1xvHqWjE9K6lWidMaKph4nkpr+VnWJg7aYnH67J4pFsnvZrVtstJsw498
p/b/R0gk0pBCv6O7tVcDLDDWXQwLiTJV9iS+UzVqbfkT7iXuf5igBPIMiYuQW2TC
zN40N+zJsV0qPSUcpjS1XO5SQI8NMQBm0vZCirQRDzDzAl69zvCvGUgSTM6mGwDP
bHSStfw/nOQV+/l+N/oa+CuMByf7cBTKuc4DcSdZP62c5ig4Nc22RcAVUBG+8fT1
REUiPHPvwBMb+pWZ8oZ5W8zxv+RqnInQDe36QvG7JYIGSnieu+eSMZeBs98o9g5M
HQMDGPcBeNzQXKyAOBs4GZrA6HfMv7izsIlJXxTXoGLOrpu6FAcJ5H4/zjeCJLok
KejKgsv3aOrIDTaaU9Wp5AM6KRIkS6+42J0eB1PsmlpUSrOWBI/nfUh11P89VZL7
RV7XsrU+s5sDV12VKC/WlS8fsuZ4xRXoCen+bTieQmsa/0ivBo011ldPFp5ggRxC
5/aFG3tmeZ6nKHl56C9ZHG9HigIMnk4BC5IZ6AITwuRz7YvesXZDjT4CT8dxRcYz
BOp3+aAEMH+EKbHu+uM6aqqiR8FtxA0KrsLZLYpzUst5lF4YsgvQ/I0dC/Pvia2e
L7yQi/4+EXUPTRU5OjYpLXAXss8JrCgy/hPCJagNWTnGxfcfBx+KWoZiMnPDSx1K
1bzygr0bCGCxtIAQBh/N6IJ7oRL7uXpeTe43Oh2ktKs985k47P4mvJ/vPqA3xCXs
JiGv+e17BgIRGNxYQu7gHKLdQ/+eVBJvrdJglzWetV42mPCu3Wss/Dh3FxD1afQN
vO50fS6aYDIZ8FhwSvkcKcv+u2m3A47o8p8YGLZsrJt8bm6A7I+Q2CDiZOWnkkPe
4nORWDBEStWL8ODAaw2fIGiea1pHc1BewCTABgLGqr9TEK107AJx5WW/EFg7WyOj
ifkk8Au8QgkEyUQhFBRsYo0mXOFT4H0VZgvqnubSCQ+ef9eS9z4bVfyfMzh4QnFc
t6yJE4a0GyaR4VKz7j2CIrkqD5xpamHbK9AuhiMw4yMh8OYs0TBr58HVdP2ZGgp5
v7oUkRzP4ZGrTgFvC/u7QIgZ4fTYuTI/ppt/azJR8IToL0XfyI3SXDze4OJJuvb3
tkGo9vpHJj/WZsR98POEOmfzGx+cwN48KeHOrO6QCro7pVOMXBFKKlBKqYk5Ac2n
tRYGpFBT+XtVFRUGwS7COneQA/pgYJxQpN/xM4gJ8ZO3ztj2pDUQDOu8De2kcEjP
dy4PgC/H4Doa2f05OtiJJ8h+wPHQjlmmZq8UlSrNyFvfjD4i+3jcMe9jlmvV4fxO
4uK5aw4KTyKBukA9QRkwrBaTqrIb6vT3nvDA49mHVS5s9h49mzDoU9bSTlE/VjIh
CaUrkC0Yb/M//w1vMyf66YOvxC44kSAZ5i9AaBbBHinD96b079UrGPMuBwsyA/44
UNZ+H+Sjk2EnalfaJVDY5LgyWaKzjOgGTpiuYLCF34ROB0j9L4np7gs5SU/YWGdZ
OeO5c0Izj42iJVmXNEEIhUcOqLJiUvpkK/AEi//FakDBvLAdF92MmkpzCxl0yBOd
9spP25lwu5KP9QIhL8CwRv/q2wFS5dKaAFwge89xQn1zK8FYZTW17AutZiyp9RmU
jGQJlHE58m372xIQ2qlU8tRrHOFVe6+42VLCf3jsv0yEuUX/hihpRYPj3FvylDaQ
Rfl1ixM4YmP24VMq3To8Sg413+DI+Jjrby1q4XGT0BwM6DGRZxiK2Fzo9EPZvuv1
b4Gc+Dur67KOMbYM8hm+0SKKkbZhaw/ynFxxkLn3ymwvFWrmtEQaXsI6DfTplD8q
+VjzEHsC8KRdUzXMSJDZlM1VVzNdpXuh0ubmPEGJGe8I2mDyKb4DvvmEawbgiaEU
k1q349Q7MmBf7uPwQXLpncqjIioFdYRhajbzuW+O/KVhERXNgJK07l/1QZr+Akbr
q7bL70AyAQL6RLiGVEo5O9Wq96n4zIVQHmNcqfgEMmiBUlVnACyw14B5p5IFLDqz
3MGvG+e9+KBxRUINze+fnFhK6OFuh/f5jMLUbgwvc7ivQxlZ/yjhJ53tR21dhL4V
jXJv9pe2NF+aoWEMl5HWAL4RAKJu73hSQbwwz497oaKMIA9cMlObdlmRdoJqt3Ye
Yaqtz+QVf+387+tPtPxv4SpvO6Db5wJlUxoFQVkQ/WthfEl1oButFsX184Ic7qcB
KGtKjH5eX1vNi/4eHCE1PYjXMjBERS3bBBDCekOS2Ul3fLbhUiVGIZUrFKfzdIsK
PkO+cOkpNj8nQUPT/f8IgNUZjjFRKE6kb9MkHUPaR6LvsY3zfP4O8aTx16gxM4Ge
SLkAb0Ocd1w54XweueFEmW56a1GE9liquUeaFPtf03+zKrGsrP00+dwy5dd5RlnW
JS14Ut6IuZNc7SBmzCHtv8Nx3I4RLAAj5tfU/md9ecZZsBueNMLL54KgKv61DZmP
xsbIjB2vcWbv3XToUaMaedpxvGTW1YgZgewkOUfnAw8hztj83AWo+cVKjwRwBDKL
vtkTXLN9whT8QhneI1sXEPEB/n3XqaJEDF1mphcu5b8I6wgqDDQ2xmIiQIAyHgxy
vfsmwjMDaoHBOwIqovbNWH0txflMDTPy/z2SfQQwPTAlMmFkqzaF5E+dfV0C2AuX
4cBi/frv6y1v9Q/FVd4x/+KhPVlYHsPwW5ef8V33v1FbvJ4EgoiMNPnXuiVMLo0q
Hm+kAL0iROGgK5DBiJWSSI4/uUMfN3XEC5jPFGZxZ2XFdq+/EDeb5KE+U2gwpVhQ
Lbj0SNy3Mmyu0e8D1ZIRvOwQyP48SK/wvHt9g+mquFa3gO25ajfoOLLOMZ8hpY72
UcHknoalBRgEHGzyDPa760q80Grih6mYbcJYvkwPQm6wr6647uO7IMtDStJBUxYN
KQHSBBGPj8qzFwfqvSLFYd39KxHb8Lff4Kg+Ox73aJ0ynDjruj9eWt4MUY9+H6+n
NWHRYJDJXSIPOwyn+YLwJGrxB83sFNUQAeW6N3dwt0PslR2RjQx4qq+iGYm94DpY
rFMJDrz0B43GB4K1wCvVf1I++UKwrtjvWOubmpP0aqQmCBfEvxxA4cxuwIi2x9Aw
K1dkiKyKSHgI6RWE+zD5r4mJOvZ0YXu3UDIbdL0LL4I=
`protect END_PROTECTED
