`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jeJ0xldcqCPm/YewmZqeeUu+Clp03ZidTjIL1Y8KHwRnQT1kd6kPPMskMZtCQmYl
7+ja7GpYA3xYZHYaqXXRmvW2zUk68JP0V1kVqRPZSHSdHL5ONfqDsu++c9R4XVbV
ne2lLUNOKYIepw2Jxqi2oN33UjRRNsagCVHxV9UUagA7auV1g9WlvaDD9yzlFM2M
VGgLENwHOnUyDQsA1ylFuDov/hYPXxfOPSTwzvdrKxHFammabuxEytkK1PkMwMNA
TCcqK92o5J59cUVw5e5N3DGBE1RJzqyDHz2jOG0Mwl2D/WRjIvdb37cOkWVWJSvH
eZuzU+/wPMWgH8Jpe6DBP2degOltwlh9/B/FAI/GcUwxEyErmKjLNnsyLxakCywM
gMnBFwpuUAXIWhZPkqOZN9pl7vsRG/pIWfD17ike5xRGNZ5y49ojGzBmDu3HZyhh
LmX2cz1pFpUKCp7/vAMw36ANvt0EH7O8de+SjdSs3sSQ8nCnFlIbLr3QkmO6hJAF
ryN0Ss2DXmlmpJcZYYDwIg==
`protect END_PROTECTED
