`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oXGrEPBDV2cLc7y75VujwZRtDCv9ucXC0g5zgQma27ATPQd1NOt5jlXHo7KDdK1F
yuxxOdWndSK4i/VU560WE7Qy8rLO3wPDCSzxuSS4KccxMSmzcaaDSO+sWn29BVtG
NNTGC2GPQYwEnal3F9ayzOXpPb3quwWd+vfFZzvSM2DvByjje3/F+3ig2MfSyxaV
9LY8RrWJnoDb3CcnLaACxC1N/v3y6vSCeUTNcmTgxI+cjdlBmX6Asrp5iNpnIfe7
HF30UpBwBShgNQzX901NSLoIdKui3xY1pkZ/fMCFn8MPQMSdLRTVa4KFl3J5Bnlu
tZExlztAUttV76aKSOqdB4iHizQmxEV31tBwmPWskMyQN6AtZiCff8w0Z31iB2l5
VUfHHnTbYaY/+mdbpDqmkbriMhJEG4Z8g2f7zCtT9g8=
`protect END_PROTECTED
