`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0qnWSIjtdpry8WUDFWgFrLIYhkrOBZUbM+JUcM35X/Yl5S55EUoK8ETMsLTALGDr
SAOC/2emNO8lmBzhga2BP+X+ZW5uwiHqbwGTJcFy17F/MqAzABlPztVkkk9IPxfE
m+Un1RZUeMdQOlx1YTMTS1bBBW7p3XJQ6+WwczJL1FYIDuW2z+65hJEpjlWfkMKl
f/G97VKX4i3PTH2QvyFwIBhpjc/iBIQ8lu6Qzt1lDfFMVjM0GXbBNEh9JpdC+ZiB
edPpMIBwXspJnZ4wNyQL1bvjdfDBBbnkpxxu5KC8PwF6eci+od2Gtz+qVcCwJB2Z
3RU7+eSb/+YtjrQk1TSqujDctJGKg5RxLXs55e+TW8KVUF9d64mB6ENSalFsn+cD
ww2t1d3IhVVQdTQDY5FVjPda9dyhzeHLq7ciQy19qPVuNtIWud/JGZoytcitGs2p
U7TiUK5/vB0JyuynpD4CqYRzgOqk8R1SeBzAFly5flb0vl658cdB2sJnAiuaLprM
aBI0d5VAxPvP6heY1c4CRtq4kHZZjqk4a942l969x9B+y9KZxsovtPex09V0Ih67
4vOMplbgboWXBn5EqA0QE0HYiTPUEBSdyP4dvCou9ZT3+YO0I/OmTDLovBvraJua
sMXDIeu2MF+6YO63VbiyLhpGma3ABrLedNCemxaRN7saTUknKLRKHX57gztqnLGk
w3auYsWzYlknoDH1K1Qle3PFKmQ2xjBV9KBoSuJRTaA81oPLvXRJllXdW8IMxbsz
EMcjoOFluC51Wwv2amyq2buMOo24Qd9c6emXQV0VjJZ2wFN2VjAr7MCrdwxNk53x
otzrb52P0q7p2WEkfiQJxJF80LfUfTKeVYkL/ccjyRrCicM3ReVyjeCFN1G+sWeq
g0cs8dJ1oJZWzjBUsY/ZXPjFWm+XxTTvDqNieHk47K/Bv5daW5tz+vZRLnAxa0lA
nUVVwjtxGFGCMwY1wXcUwEZVCuMoSqAY1afokxz2OnxLvyQWVrzABqpjQ2NFuKRC
m5RsO/UiAkvHUNek4h+B0zpS0vtKx/v79M4URlYB9TkIsE+CVwVErQmvhppGOz4t
GCcLIvAHl7cfuR+7tYuVmBOOVtia2V+caiqXwHeO+Y8kAt1akpFG7wpS6iPUYtAb
OjJ3vzLdlFi95PdmxqnjbyXk61iFZKJrOep5gXyw9b/pMibuqZc0nnZeNRKK3AUo
5tLuyHYdbeblkoaPoQbsCwVeDz5ZqYdhn67i/Et6tfUGW7Pc7XZ7BdeBpFCiYnoa
gdnjgmiFrSD4OhVMRj1GVaexm5QOLrBCfOEtUotohXA1/cKXCGuzsep2gkjS22G7
+xcYDGJZODS5KM0fp1SsSCjqaj7cI5EmeioQq+moEFGPg4AP0agev1zKFU2r/E2y
26bIeeYRxvP/icY+LUfi60/20tHMcYGBxyweVkaCN6Gpy125ifUmMIgnHJTsjIU2
p1xoNUlH9sEn0eunvR7WFONj3jbZgQU1gfK/7nNiRVVlf76lTssejfBla/riBilh
yaBhHMKog4Yob/OvM8sm73YAt7nTznu5Ezb3nhSb/2o=
`protect END_PROTECTED
