`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Qy5pNAJsLu1GjI6NCZ/atNrmlRhinr/4bKjiv+iZGKFAP0Mx9eYOlAbSoQl+YhK
Sl6oyS0TZVuf7AuoeSNeG27KtKyqhd5bLz7gsvxC1dc6xjw7nyrz5OqCTq9xv6d4
mDX4toySCvREfIctLe7uH+EqPVFyPXMtci9Fp7PuqDdasa+L+Hi7Y4OsaSrg2D4F
EdQWaWzXj5I+f0H0pBEFFjiqTK3bMnw15fBREP8YNCeJeKVuLyiVSv1FCMf7LbWW
XkN7c6vNc/CrdwiTz6nnOXwssH7WdM+2dkZ0Gbbs2WnlF5CSB4jAnDXNOYKnDVyN
I+f0fGREmQMJ+xliLJyi4FNo3LhivWRHvU3X7vKKkp36TAr613wGR89GXAdCRNCS
`protect END_PROTECTED
