`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sYMo/sIuzCgkUcfgW91RriSZvF5zzvtEMnUsVoMHtMDKC2CuiM4QYn2sfVYmuEmm
lybGBMY7brWnKuVba2OK+SJNFGKjJtEfjDm4wPMNB8aVaPm8p5lqCjisEtqwZGbQ
KyAn05PGpiseXse5HxDXyjonf2NjeNy2eTIlQbf/4Gg8QSsdm1CiQakIrkTzFrGj
BMzyy3TUZujCRm4BYjHYrVDZiEEplf0yWv/Rh7LRN/qEXgYhQHa8ROvFiiOYlsFm
Xhjd4XyWg68gJL4PvXdkpmesGW7W4O4Rh/JU6nt3ryPjQsKOuPKMeE6JSH/YtoXv
A5iolanhNCcbX0mpO4a55IXMT0Ak75Y7cotjWWZIasouVrTB2Si2931sbru993LB
pO3o0UcPiid7w9zknOjjd0vmdyST/S36lMZj91QVt3JLYzULkwBrAtXr2wyth36g
f723BSTpdBRDctaNilEQXw05qRoT/q1T/cRBTpuojxtxmxi0ibkaLmdJm2Ay6w4V
UtaEzOn3O2Myj4crN4WAXmvpxYEFCDAS69AjrjSUgtJLMBWXZExCgC4Qqum5fmte
yxoeIUMH3yBQ8pbd5BZHWpElU/Z43lYt77T6c6TJZ9Ycq2Jt/fjN0D7DcgUiGvG7
qjNLATV2LEKlgGA2kQ2MxKCRHef+NtjbObrX3r1lLE4JZEUDoelvlk4stZHL7e1j
7QcNkHh5Q2Ex9LslZE/Op6lEViTuEw71ik/6S/IguccQkAGBIWOW2PRXUWtRh0k7
YLT2O+ClS7vz80cs4IS7EKuEHjQpf+kA5kAAcSMYF+qzeGHcaZh3EE/JZ1bPtliT
Jfqm4Ei5tCNC6huejJr0u4WEeCJRccgsFqoPJ+L7cGhfnlzRINHWfADhuzmeiGkz
BTnJrgA/bCBzF1XnxBJ4VMvsQNRvtA5G0jLMFvUF0n8=
`protect END_PROTECTED
