`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yGPm+BP3Fq1LIR+8iqxRq3EBYnue46fBQveSs4yCrTNvmI1EflvghvQ5V6DPKxfH
pKgXB91KCEDdY8hGfkLWkvRgQqs7kSr0t5+vXI1KTVBV6cxuqm66xslCa5jYjZVu
NEiOsP/VSqlzYxd1y+/VTyX32mZKfu1Myh1lJoGoHXMDSWenYzQffIylK5fb2b6+
V3QiLSJNtXLdmWiFEVYXC4lwun036BiOOtdjo8LQSiVOpXA0HWeb3ublPnFfRFvh
RKa5iIlY0dUCkWdCVFvYJbd7vs3hzNV/heylsOqoYoMpmiqKumzJNqcA4tGU0lHd
I07az3AX2jHLq5UuppoqUdnCeQ/3HsB957Sl0YJiFi2nuF2ahVryJD24nLoictAu
NzwLt7PTxuyXUtdqX6wpeRR0YDVc+Kr78SiKWwGmfE7XI7DvccHqoD4OuSP8sitj
8phoTo004YJnVGldEiO8XGm//kB9+8vAeAC6WkipuprElou9K+ctdgAowcq0fdzc
xfCOvcS1BclLBnqb3DJhPw==
`protect END_PROTECTED
