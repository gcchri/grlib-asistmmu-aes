`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8VuLrSVjr/qisVthKwwU3qXFEE3FkNJ802C1G1uun/z4kClAMfmzF/1/v+NkMSNI
cMHMZkGlAyY2LAN0jOSfNYPMN9RJqW1Cypy3HTcG7wExCEXyDQtjQ8z3ntqNTAds
Khg/qhy4rLWyfCwt4fuvgupYNT2uozjwlflOWDZWkPoxneJ3OEw3CUPx2Yi6slvX
fGm6yzPYg6FPCk2Suz8mfvxpR+J5QM6FdXT90sEkhQLb+nJIirU8sIaZfu7AbWPZ
uhxNfWYfWe2pSN2UktgCQSPW+PK7V6m28oqgxU7El+fQ7lCLKOyCDGHx4/UxqJCq
kPoP+IexP91FymUnZnig49Hyv75JgY5NzrpZkNU7TJxYiiIV+YDQjWF7fFDwDPnE
CxVET4XB479BLoDGEdZuND1/hSQ7PTRuJLekq7iavLzqc0OzH6wDYMetJtSC2AvY
EYDsPY7/zEmZezUxN9yZtGOWI/uJ9B0Ljo6IDPe40U0tfRFnuoi3r/odWfS5QzzC
9DHhgjbWp7QSV4F1LEcupNwf8J3x1wSqey4Q/tW1tg4A06EnvtCt8quqKdWasVVh
l/zOcMF1TZ5Kv2rTh8KD/w==
`protect END_PROTECTED
