`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k7zXawdoJl/h6wb0QRnPZNzJQUNP8sLADqI0ee0IDJIvgNXfjoX9/9EGKfyDAi8d
yWl19JfLk8yH0OP/iQOlpw+A2wrvUor1v9J8nxBLOnVtBPN3dGkUP0GHRwcnEgzh
BKw8YkG5NihoYmKr3F7rEpjkL0QD1P1b55koEOLDJ4g7d3HaMHy0SA/GQ8h7OSri
VuAUh/bHr9oEa6brPiwaK5Yfw2LcoGe65x2TroABkBtIWQfHxCSZMeZmefXsQX0+
r2UvkUfJN6SItkXLWn9GSV4vPenIHsleH5gkKRzCcs7w161sfsJITz7C+1GbTxJ7
O8G3JlFpTVOoxNdvKyx9JPcKO4nDqDlTJ1HWCxTBiu0fOBR+Rcd4Un4YWmLUtc/H
icASQDYd3LVHn10u69epZoUBmx1DjpUnrcMKdyXG1wqyFdNP3hHBoESJ1gFNMP40
8Z9WdGSNgeHl/h4iEIjCFsdrEqB1PxbB8Ve/OkxWrs7r66S89CNl8Ml43l/u/i9X
neOfmraQi+iyMoG5D70PUBKdEOyWdhscXZxOIK7nd5U8j2rFh3Aq6S9GXMqY6KNo
lfL8sZQU2Q2ozYweeyh544pXpWpjwR1KZmOZMWLh3hPy2RCSM/jCqrukA0pVT1du
pn+hPaLBDgWD/E8Dm5VED1aWYeGY0HkS8Mj9e+tyce7d4TZi8wrHhV5iPYXejLwp
IgoMxd8CowBtsFXgtXhqc1rP3VQwh9+MUKW9Q+ZA6m+0/a6Oehwrvxe3nmxqC5TQ
TAw+qPfaM25yHmHuRIP9kIpDJfHDnZ0Ol7M30Q0LI7Y6h+ccEAXPlfOALuqd6PF4
AMvI5pJOrHb0+SNs5VSUKTnx7AdyyC2+L8BswcvS2MRcqOnp3ITuflFYHHSXaOkr
TfpEiGMGajblAkIBtmqA+Nr18pkxTS73OHmhfXSqY9B9rgIudw88KQm1BR/q+rnJ
vvAoB9euixy5HdNVq4IPmEUNsI3H3wij8lOzpAR20e9u4bkqtJ/tMluil6NZsYI/
GOJyTHjKpyBBmhIla8Un4/CBkw6SuUo5JW650xalF9jwhPMRI0gHXyHxtdvBFrTk
kZlejTW2+befVuxSlcC1YN3Y2kJ8S7VMLqlSCm5ta5FRsu/sTNhdrR7PLmpNqHBJ
IPo5D/HL89n79+l9S/QKNQFw2vWpr7sCDvbEPKaNypVcgwF3CHkaVP/RLslLRBVr
y/GDAgQw+mPNNhPqZ6CuaOh1hulhvTIp9LBYzwHPlFiSfLyLRA74oBlgrt5H/gY2
/jznnCj00PVTipi1L6KS7HdcThXAkifR3pMJWSN9y2Gq1QcEDfTVsC5eDmDCidQb
fcBEnr3kfP1ofLfjl2CY5xjSc9w2+1BbCr9K4qs3AqlHiuvJ1wz7ojVNL2Axpw1J
d0p3HOT0OZ5z2BH0KWuEw6bWUGigxQyqQdtxoWSGTPJSE/VT7Is6jOLPM/ZcFHwh
+K2eMChravGFCbxwq0QIx0oWwvG7X6us0ReD2TLfT2kB+ua3a+rG4Oq7qw7W71sV
JG+U4nKGIY1LphLUUjNWXPWE58A4EpJXk0eSORDi9VjDOOgLHDoCDCFdquuanD5W
83Q/NtJYDPjmHkWB37H/7CEJFCPXZV3mWiIp++ECiJmSvxV0RFhPKkkky/DtoESn
gbvA5KLH6Ji4oNsXHjujc4F4IEsvYYsZj8eN3g8x9QjDWwVc6zzgYO9o1SL6zmdy
q9CAkQyrVfIb0LpfQpZeyfA1Ru73G4ldSg17mbO9LjFn3eCTKdNeOShrp9RWN3tH
wuoJjWXN29JMOcP2zSFEzUuemvqrVzwnXZw+cNtZFLpMxgyk/HZHK+WelZu0Wtk8
BJyoGHrltrsJEf3V7jWg02RRDifw8ZCj9XwC3IiN8CyfVbup9munF8a+N0nx/hao
E3Be/IbbRIg8+vQx76jR8L0/DGdwdRLYl79iBcMWm9A2+Bu1TWFc3b7dpNsjmQx8
lkZUHJ6sWHK4G5yYI0qhOKaXEH8nx9xO1BaiBpdqHXSv2wURONb+dFRlR+tEjugO
qvDEpLt5IN63Jb9zfdiH23rqilJ5jFrUHjXp8l9CBBProxtMX5bTzegtxfyoKlu1
BhWs/qgRzqghySHBQFtbQTmHTZiizv5BlAqXU/LwuWTuKSt5+kj/CaOMiXHLDDEx
d+3ei/1/H4PLOQ1gXLIz5DqglwZtsUAZjMhQeFVNA77MN3WotHKcYqgGHrInd69a
FarTY/zWn8muLVFe5Sw/P4vKrkafI7eDixrWTiebAhkyFxwsDPnK3ix/YPpbN51j
knJQ9v4bveuHjPE/NORci0BlPcH/Aik+b8rkMEsnhpwL+1+g+ujSrIV51aEPyOO8
Fuw/XnzORATd/8qeNzTdFR/UC9zLgkISHRQVwev6sLNW4KoQd5JbJKBVQ20l8ANq
ezdyZIf7YiHCjALkFHfdJpRK21xdVihBCRHnBoIjMMza7kxOFQ5OwyhTgQ9LDGA2
uzJeqJ1wMwnPI8ykz+BVJ29s504LGp2Nvj9ZKdT8CSXcC9VaRpKa7RnivMnLivFa
RWdZx7FErlKeMBQZZfP/vhv4OA2smArunMSj55QKMZjH4hKFKskoAhyu+cA/EzYy
Xetzpt1nZjT11zP2yxd34cQ5VV78nD1nSi0ZQEeZoKIdviFji/w3VPNIc9/wbmRb
ALuPFmeKMQeK+ndZFScCvxVNSaH+N3qcnR4xM8NoF8ecka4770UzYaUv8ROnloaN
AUPhHqpaeXwJ7HMLKY6iefm+QVhVK2SSGRnboMrWcMyT/CUzddLa0jL9grLsqS8U
51+huUe9lTXWcndJVkVsmkVeWCu8uylUBZgG01zX1mOIoIfp7zmEH1giSFvf8ZL3
NbLsa2zGtq0AvvhPzmYzqNffI6xtKZJUceJVayF2lZPmZinxfifzXB3ANXhlHUcz
SeayUdJqOSsdTADPuvegMP77ulTqD/6mQ9RpM5BJDIolhytzVwS46V1p8HZdV5PZ
d7svq/xnIiNm+RsFATj8hteSMzvquvxw9f73mc2v9h2PRVqmjMulZ1QxQkUj5rJI
Nkl9RkzmqnI9LtNCOWwI0+4aNk1DgFrs3izJRN4eOgfhvpidJ9MjGBG2i1xiXsgp
1+9uYhHZCgxa3vRjV/3wt5nyb7AgFlzseMj0VA2EZFpxzp+99d7hpeYF5QXEgC4M
xkEmWvnKg25REgQn8lozl68/rIoP9llcZhivscyVfYm91IsC/EXLVL8j9pV2K08B
/q9pSSjiBS/Yv8WXpkaz4/Vlx277xGAkBQT5WGC0ZA3hEDWrj7B6MgPF9C8x7736
nSZUsNr9AskvKtx4wvzVueZ2cTEC3gEtlU+qKSuigoTjSaQVP091DIkFk/8Ai+sP
59tOFYteR1q5UFmOYonM7m6JNKTtuJNt4ApIf1y7aydhJ7FPB87oxseHj5lx/X02
zcHBYOzrZqYAJ1OmOpLCfTE3lOxekzZR7KENpmum0CfPwUg04ofB3lvs+3UZUvAk
hhtumPNr5pb+DjYQHvyCI1sHAIjHHZvBfbgETivcQ6qu9GY8jHpLd2sQo5NYRmP+
0xZQW1P2YhsZGaQYQtJ93s1FB0mk/DmtkkT5B0c9UcPsn8C5SqfndvoCH79vlW5d
+1PhxNEvlTVGR9azillMB0oY2wzJGLn840zx+5hLNvY36CQwIhe4jfX8O7JX9MlX
HAQAwsjWKNAPRets8dyODhZUgweNtvX+ykwLyyFdebKq+u48TDTzJUx346/pFzPN
kRoTlZeosdI/v/FhW85XkttnRgg5Go+s2ds0daibEMt4AkVXISZjbbZWIWSqsYNC
RoduQTEsTIdLqFJ7g4BsSxNMZiVYPOEfcA+3R30qaEMLR3zQc6ZS9fgs9zx3DT9R
6s3Qlb+JIzGj+yTaYMdX8gVfDpgaokfdCRlZChBOYrtiP+T7ActqfC7TaRJGoTkm
lSod+fG7aMof7az1CaK7BkSa8PZ1hGbdi02ci2RfPp/2uRczyDBPInzAjZG/nevF
lq7n8imhIRGRE2A3jhmWd8gfJqAvhUQ6jgj/QiMRjQhhTB14VL2neZgUatzFQsZd
0r2qh/KisN1pvAXlRDRuOBOWi5pUaIXa9nNjFS7sT/sC57A0KhneNnEjuinGKN7V
jK2fsDwMh18VoES9o5zDd/uQJEBIrdqhOIBsDdxxYxY+ieQVSKePEDc1B7yjtmxR
cwVaL9Ag1wlsr0phcXqGUml45i+IoAyNtTPkqDdma9Gua2HeTDLfOCfquCTwj1eA
lqb/DcdCx9GWN61Ff6MU9SnsY7AR8Dvt6694aEOijKj+6C6rUfzD3/piEzDYzElq
mVDCJd2qltY1guV8yhvE3YvwoTpOFuDHlfZGIOGfgRKa/pkVe4Z+LmyVuDOLG9y5
cgGKPNG20PapyXf38yOw4zQ/MKm27IH5oK8LM2YcH/UZAxLXwCdqv7HYWphp1J8v
shqtGuI+3g7qmSlnGBislnWcS8G1XZXjj3Mc7zzplWs=
`protect END_PROTECTED
