`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eNV4QPinrYfuTna9y93vllJ2ZE5uzaSr9Mjb3d2e7Te+gmakQyCRExUMwAAZAApv
W1IF8ScUUlFFB+6njmtCfYAFPhWRvUdDnH1Xx6zVrEAZvPrEgNeq14J0MdrFul9/
eFi3HPWG92XO759JtvXRdjVO65tOpckutgRXv7uBTHt4oitMLaDbw0THbnnDjwJR
IugyHXRrv9euzaigkTa2Bmu5+m/9+9ymlMNoAF6+egIq+wjuc4Ny27Uj/pr1sZxq
ci+3plKAg+1jLqZS3TA8AphNh68RXaO34YZtmLNpF0kF5Av0f89RSZGHFKDeatyj
Bi3lHRnt7Cem8fb/Wbfv3BCL+NQ5y9VbSDcJQvWy8qbxbm3dTCAARQZHaFhMhv6t
3y5ueO/rlhyijgSdpKf2tNrZxUVVIozGcLg1PNDCpiaa4rNnZWRs2Ys3JGAABsxK
`protect END_PROTECTED
