`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EwhZr4wUBOiyUW/X5CkMWHE7HSGwDD7PaQ3oztZDDhgiAdkXO99dDUeXIidudLmp
D/ShqGphJuZOpKG3yaTVZL/xRvHPsd8dpK4bHMRhFuBSyrtMQ5jNeHzYs+QDYCvp
pwS2TqWpoPf0Dry3OP7Kpu7Fc6Tn/SjEVxvsHFr2QSp+LKfGNIX76B5RUMQsTOtN
R8uHrlHHGMdoWdqouBfa1Wsz8kS4jT1tZMduKDBzgWper28FhuMHdpeCTysAnNUa
t4DQH0N8LmxFdKYi51jhhev76CZqyS7LRIa3yts1jgVoUeP2pQz4PZrawW7YeYrM
5GSei7aznTyXqFa6JShWk9bXg9MzVhrWebVpeLsyujTfBb/7VIEMzVrss+01V4i3
KYZ4HH5s2Uu6EEA+rQDWo8v7M3PqY6akMGl6q5TQgJNl+M+33CaWDhT5sL42qODM
`protect END_PROTECTED
