`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hwGbljJJhe5MY4z8y465NchHTV/6NDARQfZXOep7ovK/qaDbQcCz/2SyF7CB+7Kn
K95smEbPUSkqGkHPylEA9LQsyY+PTFt7NKVFdzx5NPb85cgp9X1QrSkTKFPjPqn5
C+vu31HU3nXiRIDU8Y9JcdVIIwNtpVYVmWUv/WTtRuZ7e8VxLL6WnJyL5OwJa9ts
UKJTEaI2Tn56FbsiryWZ8S2PhoBLyyhC6k0pIHs6DCTI2zbzZTzPcnBJZpDXFACq
7oY0BoGimpSodCxrusHR7HDWQu3SYl8wA8CpsXPtPhnGSjvmX+s0baKxCffLCgCj
lhCVp3CF3Nry6Y9HwwesVYHjuRYrKkhZ6rA1ZAlT8C4IMl7/iYsYQxNuNZVK2EX5
06Ofncn1N/vjP3DdIkc/ZTFeX7MZExRE0AGb9npJiU38Rc8OANQ5WLqnmr5k8K8y
AYvFXJnspE9Y1RrjwqA/NXeP35aMjJ9HfbfFRs2DgekscCtAWshtxIkE4KpheDic
WOEyeMUjdDyH2yWbO9KxtaKpOguEyvoUGx6VzcVujoRJ6D72Ze0pap0RJfTOfqPQ
wP9giL6ILgnrOAGVTKkboYzzuOzZcpzcgUx0SKvpVJ1PZld7LNam2sO1daGgkc/i
DkBI6KWYqyfTdDenVmhAA2n4nth0l+kU3PZrPFoocIcIAlTnp1zU+yhVqphMBO9W
K/4XqyifU4s5Vy7iS8R1BPNmj4NqpNKQqSPpGG0rnWFxVMUv79nmdR4BnKk6k5b+
qX8hcp2mXjA4BFsVEitIg8FEm09Zp7gx7ZYajRCSZvUZFT7+WOnRtlPoUTT+8p4G
qNqbrLMq7EA0WaPwqjQfZHo/GMaGXeNTYLEKzZZ6XNRpxILAV9bKiOJRS5XEcPmL
w7ZfffdVPxnzukAdoU0/Wr+cjg3CQfOBF+HahFM7FkyIrc68XPcXrbwNNOb4ztSr
J8vzIEojp8/HgrUYT2Ek85QhVDrD2zg2PPtZD0t8IroAtuQRCZSunC8Cb+VIY1x+
V0Dt0UzfSKKpC6mYX9bb0L5JYYJvx3qaZ/xCLW+8YW2/yi7ex2ADIbWTiUPg8oBJ
VMtSNUyNPA0I5XZHOfe10+FQyPxRUr2gbUROyRw71Z4=
`protect END_PROTECTED
