`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CFkeut3DbaF6faTB0OfNHpJcuoVClE7HkZzDf5tPLLkynuZvU/5m/XETlk72rWoY
zmSMPa4TtG2ipNaLJDkNHjiS2BwaXI4Z6pNBd9A6zBTvjd3nHja0E9jqQ7vgfcFf
aRxCF8R1U7IHzRCPjUT85Q6XSK6WGxbfsd23Jmdq7BF0unh7HyVd0ujalWu01JI5
ZmeLXL/EB8fs6cOl2HIHGuD0ARJiWDdb3wVWbIJTff0Os9MgPsu/29I5Y3CBWUUT
ryn2LKvJrWDUjoXBSRhIvA==
`protect END_PROTECTED
