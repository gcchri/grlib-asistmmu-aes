`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6fe4Zyhtrj35i9vd4ASWKFaLzg/J44htNHCw6zyP30gPovC1QvMBvqRGWSMP8FvD
68DnlV+UJJETqk4NtaimwGZxyggIHsxS5FpF8xp8PITsvXdgyaoIXLHO4uPN5jEi
1WvXKNr8v/aJxVdpn8EcKZ9ZV7UwuOf+CNXRgUBWmAsHdK2o6Me+m/ljn/HXstGL
E4WitQ2ODewhJYM9uIZSfQ1jBK6quHYJ6ufol5dxZZVLEc2XZsMrUVWu15G/FPzg
m1iDfuxrzY9iMs+LgUMBnlVnPCyD1FA1JhV8316xjdnQGmRVPDBBlZPrIe7KFE3A
gIY7f8iF6XGOXlH5trp+snU6cUfZT9+bI5cA0x1wM+o4WbXzxs6vMHVA0LyskJts
LwbhmR5CUFn1NkTc2e2CWgbAsfkCDzlGUpKVPjZhkQmRvC6h1C0ZNCGqn4xmzLpS
uHWRfg1nHB58y04R9ud8B5nmQPOhqqj7x3YxX2WE94lapDd3SNzYRHeiBFK/iUcQ
`protect END_PROTECTED
