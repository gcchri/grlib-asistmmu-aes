`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YNSSBG2qUfVMH/XsS/5YRzu70swE/jD33N6L2cQLvOtO+amyXAxSvEsDIDwRn3kf
DzkIw9UUvSYY3pqwStlLQuWHs8RrsivH9NA0lchSC1/8tf5zHAWV4tEb2rzxknqM
/M3k2WIS/a+OS9NQt5IWNSEbaBe+p0/kD/zWVGBhKxD7JA51Y6EpMQLUesM+Fl6j
8MX2KUlgrhnPp2FP4J4BE8Pmt4bD9Q6UQwT4+Kgv7iVmiwIWoXAlkdo3jkPgWF5s
3Tj2X2uhtIysHpDkcq4yFEht2Z7i/78WO71X+/rW+jpGZluQhbVINSWzrGCL5u/x
aQHFX62z+vLoYCH8WduXQw==
`protect END_PROTECTED
