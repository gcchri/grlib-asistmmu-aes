`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eo9Z/iIdAg/C0pnKiDQjthLOfvcBmvLfLetf7iCdeV5lLJ344MbyLgyAsskQRzmN
Sq9UCu1vnC80t49JrNImHL9YfmscdPU5uvD8t3lRAv7PY2fq+Rk57rCvC4UKMz3Q
64blLf5+wTObvgKselhV/aSm25aFYyLqNT2lc6lE6NVAJYfL9PlVeQeC7t0E3Buo
fsYv0s5rnUftA/SYR6o8/Ze0s3p1qtvSitw0TzHrRObjZqXk6nPatRaxPujY4Q4B
gsGEL7IZ0KndFLMfu/XBG5+b4nVA7HtoTUtzvQcEXoO7JxK3qpyjte1o+mQHQnqL
YNil6AX/XYSUR4kGrg0U3Zjh+V6AVFKyCRvVE9V6OOo443+yqlZ/ykbcXaXQAfeX
PDSwzQk3y/Mb5H/azjrlWQ==
`protect END_PROTECTED
