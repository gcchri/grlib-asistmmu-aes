`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Uh0tekpdKRtaIXSunsJippFyxMhVG5B8QfHFIjxIOJgvsQsACmv+AU/soelyRHM
XQg4zsPlDG5tTLFn8NJbfFWtJR5vz27+nt2svb+YfA66tQV5/D3pn4HbAoNiqcv0
lpmUSLhS02HH4iez9ULwel+URYvKUzL3ldeNmdge/dJSnfxwrP1sfmBOCYAnaWvm
QxIAd3C2dbBfexpvg+QIjZw5He+25eMFwbVJtVN7Hazo45dYCzU+vBAlmF8JTn3x
pAI8E7ZZS2y09QckVDHTpxjnFC+v7VaigLJXKXtmLAXS1P5OM2HAc+1uWq0/giUo
YJEwUcumfJvc3vqHVXrT/dbPjZ27+pF66/YbFkLz/5BcJS6Zovv2beGzbETFPyoD
pdzPtB0vNhkyRpbkfKndcoh/ygOK5ApACmb4heigAGvQ1vHH3rlzPNQCTxVTz/Xl
I4Pr76LzM0o4VkrFlNOAGwStrIo17pDbEHEfK2Tg2DPC5PSDLP0zC90APseZn2ga
p41l0IwlO+aX03R1IEPR3x2hTVBC1ZatUknoxYhREsCAEaJ+ctGISDwCkfzZg/HU
JiJaYcW+yIvFWyO/Izqriy4vnvBCgEVuz1UqggNLkGKMEv7rRRBMG6wvCapdw9pA
E14hCd/qP116jDx2dVfevvl4vKfhaP6PpJuMpvtGcBqlLpZr/SIRMxo06olYfvpR
HR/ThvhVI3TNyoZeUAAvDzTd4TbuwyJmh+55iznnGD7brFBVE1uR0Kw0ze+DKGaN
mHSTYW1lgm841x/8eRINP+b6bCl5E22sBLoPZwZyYzX2PxPHNCJGF3ftYipFBQMx
DijoIJGXFUFPTa6wV/OHTvp0CMPw7XOaWZw1tAQbVP8EcWEQPvumG1++w+Zmliyj
AMxl7K15PkbTHoYv7Q1FIY16eDzpXGHyz2kN9MQcSnmqzbxlaUaiujvfQprTi3Vn
0C3yKcWjvhrGSLsiP12TuonF5dbm8nJWVBc7Lb3umHzOyZiF7NcXsCdRSWRcgu3h
vVV+GzJ4ic6uqhjIcbxaPWnUt1y4l801e6MwOhGb3xNvZsY+EBshunX4Tu2+n6M/
qOYMZ6cvHdp3l5+q6tXzCRNk1www9Ya6mvGGHUzkgOJS+/9/6ZOUMJKf18vrohb0
wtKofpJrgIqB4tPCnbtVvvLX3MyOBG16zQHMMMOsRePjEif7AOSPA/XopVfnnO0S
j1tRGswIg2PD/spSm/hG/ag1T6/PcBO+5HvOFO+2UjNOFGxE6iqUgMLwjsyKSCVC
nMgNdKJqLd855COvhNLI/EGNL/HseJ1TVH2B0m+0C7hTOiPeGP1+C1mcrlwJ8WgY
1LZqROSHVNRqNCRrdRIJlaRvqBwYW01o2dUJwp2fiJx0OIwf0ZdcCCYkGKcMpjjK
WrfKxWEOMq1EwIs3Nk13z4bGQXnDDB07qtjfPbJOVkOHaxclmuYrbKhL11kfF0dN
hwiVoXCxYzMnmjC4XlosTHVC36X7DoPke0fEbhdhorBAFW40TId/iEvreyDgd79t
mD02ehXsNipYb2gRRNLnzE/gcIPi48GZ1K0d46HwAYW/etewUxYu7aLL4yxvCYgN
3lEAI2qL+GBSSNbzlm8QA1ZvW1xL5KOdCEltSh228VlDFnkUDAZ/+V64ko+SGpXq
KCQ1O4nFsws/Acuu+zu/y/ZU1C5/fJuBKkOF5SaP6dOakDwYDKoTu86sJweimtNn
rPJrirE8k6FXZ2mIt4arpyQIz6STso0bikI3DiFCKy9M2uwfSdVsA4e71Ivbdys2
dQR8v3WxqUadMfvyB0/y/mg8ZXM2CEajRiiPMVEglVahIm/9O1+6ZKwcGJxdXCK4
7vR7VLKyqTTUgt2gn7pCfBmYzeLYprwUYR3iKFy2IsHlFF/yoHoQpuBTe+GK9nq+
fkvqZ60VSgH5ofx05Vsf4zJWtFmV+9HhQ1Tt4wRdieUkQZgDtuVrgrej7HKmQMna
7eOJTabv7oj2dVQtCq4u5YHDgLlC6EoRaK3tHUGXQPkwuHpjhkcR/iH5DEIA1OAc
/fAfubx5Z+1vRqsPty92+QVw0zY658jKRqussls97SVQNTSmn/gXSSCpVMR9CQeR
rUXWTPl0EKa/0DRxTbWWW6aLx7D3529Zfan5bwkWZnEUfB3JzV/xcQPxPmgaVude
3cAAc6gVlyTNbRaN4v2x0my6XVPj8K2fo9xvZ2JvgutHt8TEEgOCNBvQ1W5ozeHb
hYRAu61+Xpz4nB9eqItuPsnAfLl8ulVX/zP85pUUSaMcI/izUWZNsMujp32kj98N
eHhmEpA3tU3Uy8DgESLKz+8LT3xc/OuC3pvSfDQ32veA0sre+oQ3pduqn+cktsMh
ne0/xLUwypOFkDoF5A0j6meSRQzPKO4Ih7scqMF5SO/idqiuWHo8rH7QKUxC92hh
7sSE+7VzDOb/7ZVFnzTzMoNRBhEdEXGrFznKhZlFzPwSk7HRNjKHV+aLon8tNqIa
DBF0zO+pKhy6DD+0WhD+aQNYfuuqa5cFrCafF8Upz7juuSyqo2DGXfAsCQQqIXo7
AA7xDeZ8UVMa8b0RteHDB7DGouxmFKMxr53V5t/QJsyLjKmU4bh+Hjsq8DgiIy4Y
/Xu8irxuE+RNbjJcvI5zbyhGQhOLELOMYNN/is9PYwUjII8ZQQs+VvCDkBKJSqvj
cciQLBtpP3nP7J5qsjceb7lxbVdw5tZfAOZfNWakIOpbvLraIJylovTJV12HjmNq
OAioRdyRp/Qxk+qqPkB47WmvA9iGr+RlUC1Rym2cajsp2EL/F8vc5n6tIaiIxXZU
dASDh2Imf2j/mrmSQc8F7IQeM5oFpOvIo6By+aveZ4Ey9vedN6IQMWBITLE8G7do
qAFMMhKQiwVvY+vltWlhiNAlRhmwQkLVME57hy0zfSeBSPu3jY5etc4XIKJP1OXy
llgVpy/qyoGhvJBvcNObc3QIvvFqGlPCZyL1oBOmUYLnXQ8C5xPURn20CdTU2W3V
u7GD2zMrxH+qcg/V0v5VACEEkDFB8/otN8ZVl+eUTdFLIhD6VKete/QAITiCYYsE
cr74e57bqLuL5MUrO0PGT5BAe0EhKeSGsLPpnzPvs3AFX3Grgb5DenghLsp0IfNh
OVsH3iPvT4AzFDBD0AaYA08sDh+G0kSDOKBOahdYdh1QVdMIcsYTmOO1B+F/ImsC
YBy2qfZ4FMQatodz6GVWaHowpzFhCHM56aFZOT1bW0qTrxiElruAs0v8owSZLvCb
cO3NILx2RAEjJRyJ2wBhd1EeLHXWYWKewCJZEnzvPmzFItEW2h/WHAdZ5R8lz4kP
NN2Qp2qF5jBlCyT2E1OP/8h3tVGzyDu4iMH7yZJM1ODWF7MY7Axrkz9Tjao1e0k/
rz7Q4RpRMOT2C72wemRYtqkP4oJhHtQOr3JLRlW7RvfntH4vyQX6+3dfR2TkmX1F
SUWLKNxsG05w8YxK8pTtCe/PFKZv/w8vgv1b2KVcxCkt4GQ0tD3ubrqbR5hYD+k4
oNA9U+2GwtDB5fp7Vf+HNSU87c2+ASee5CkytsQcM+SUVQdQH1UCVFAj5TdE10v6
UNeNob14GNV6p9PLNDxlxBkAGEUJ/uZUu3UMWHuiDM6U9mqcBDN0XTvZ+p/mPxjo
qCvpDKT398Xop43hcc5UCMD7jvzzDCImztORTJ1jMGV/VjsbbIlxpRWBI/XE/T5p
r+U/ezjxLJ8YxWt9lKoiFq0vHMHYO+VPjLXd0ENRTl0/ZtWVaCXyBE5yeT/9dxID
bm1bNyVlcQOW+EMNX5wBkwNLDd08bhGH7jmyHaNjzVZNAHE/2+MD37d+p3gdZ7Al
nUV+IYKCv9UpS7pZkGQAXfScHYR4U/TC+jZFi0vFFE3AYvsVecxuvPZE6HtJX771
WJ9TgMvnOzRzIFOPo13U8AlChhsNJl9WpFRi7pUUxh7Ty7ooZTt+QG/dnCj41VO1
f2CUV+rGn/lXMsMAnqk/CAcbQaORdLor5rWu4V7fGKhqvv7q6EcDC12yq8ykILmB
g6A1j8mQQDSi513taXZW6h6PldibDyKeE96m1simJAFnuV+XkdhREjtIjpwlAqZR
OOpLSoC2Tw1wn7l7LHSDU8otmAU/0gBe0iagadQNTXKH4YLg3D33ERZ0/SARozur
QWF08fddq00KqE2so5+vNqrUadnOBA0BDIiTjZFw+snipjevU99cA4xQBZ4skLl6
L2Mga9Eqo7VQVifB5tpcLCXRzS5DECmPu+Erwn30t83dPZ99hoYkfe3NvsqwmxNX
ijjzgvnQXXny9X1K3KbhrLiY8qywWp4Nynt8DUkKXUMYG8Eg7f0DP+b23zwg0Dmd
8Ma9NwmUEyuP6KBXwZzKvMCCdBc6MrF2JRsXHoNfQ8F/7n0gH585LGKELKqGgVeb
q+pTirMd3J17EO/llGiR0Rjuko/MqwH0jmP3vOgi2jqTl8o3K8SqF2o2HtLJhGL8
5rSc8Hqg/7lNirPW1pJSaWLI1bPweIwKFbpmtMqYXJ+zHIrcFA+xapjA9nL3gtzr
wgPshDGi/nYjr8yQWSUTFac2wJv9RNsEDapRkH1iYs93JYXUXRqtHvFgF6MNV+U0
QegdwFTqyOUTqLdPhTYU0Uup0+prvsEzA++uV2SlVB8wzCr3Dtj2Sq10NRd7zFVJ
LJy6QouU26wK743qGYumjzgxL4iuy5kRTKNe8OnujRE/DyYaNTIwjuk3AZbee36e
ITZED5MtD8C4wTfvXnhoSrETw9lk5f01RJie5j8bTn9KjYuO4JxQrQCU1wCtnCli
6tK3AzYdyzj+fU/PK2FGCeWxW0XVgB/Vvss1D449IAd05/c5T+YVb49bi+KmSFT8
i4Ya2Nnto9r3ZpLCeODsTv+60bHw+o5mYcI4h8/iF3DrpVB2vOO4kvzS9Nm8tmv6
f4Cf+ZPcGgK9ha19Z5jvIxfIgbIDJ5VaBdBIma92UtTNqc0K0bRdHyk6rPe/phFn
sCXMjg+iyCff8ZOgYCFw1LKnwTQC/E6e8M1HuxAmnaKKqM3T0s8z6Jxb5EcPD5Rq
MkZSD1OBxfAlCeTd4w6Qlu6lbQy6IqBx4hr2y78m9iTgys8qj7nADHxj6S/0+t6/
9yyaSTJxDhjYYjBkkcojJZw0OdXuYfoPWyt4uCD2VkMal1StUMf7X5qjYXh571WV
FYk1YGNS/kMqisXrbyeKzTsVgmHRMF8nLsZHX/qW+k7EBIS+0jhsBXOxWWGNQJmb
5hdkqHpdrp+OJe+9cSFSXRChRIcoJhfbE+B4y08hPqezAdLB9nyk+5CajYZtWf4V
qwqeP3MBFETJ6+owyC9vqEN4Ej9f/reV+dQIS3zjAwpToyC91SOvirYv/Cn98rkS
wSteFbxt1OF7szup2zZpaXqzVM5oQXgy1A0lmfNol8Jl6jd4qhH+gj6XXRl15It6
aH1MmBLZp2Mn594RGbffA1OnA9ivHfM3jpPAqEa3zTlROIX8JlQGxfBeTtWz2TNG
Hlig0K7Wkq0nhrWH5mHPW3bj/7gzfisvVWVRWgK9Sd3gj6uUNdZ25saIsvWvbVe5
9FTtrbAjfyaXzLWhiYSXKPMgxjjnWHXZ5TU9EJxtrq7qIpiNs0HfX29022jdYNJr
6oEq6t/71wL5rB+kFUGWFD9Vd2y75VRws1twm0LYMJvTZiXnTWi1wPvk9yN97+Wz
VJp7jYZ5vPl34QUlqM5GCxLs7Lijg687xBDGuUR97Xh2W8lv+Ki8DVIZmgyrbdSe
7HTTC/V1cNP2PRCfHRbnVCJ51Ng2n6TI2feYkbZnFDOhDAWsS3txkzl7L7Fkh1c3
swV559IuSpZ9UA0TeiclzddOb/+l1W8/KqPhRBT58ElsgCec0IgDTZolxq9R/LT4
4TsAKzLJtF09E0T4UKTp7mjRKNHDQCYOgseoJX+YD9gAAt3OtdREqEvq9+dARI64
9e1twhgiRmi2s4C0eueTWE0ZnYoKtd7Ivudtu37z4Czp0+z+JmKCqsekGXaXE+zI
I1+TWR+khajjNcneM62nyISKZ0Dxj4ylIal5SoXbNtLgzAqDHZc3yNOtlXjtNNsf
raEfaBZ7/nto+gtj0bvTjS/O2MZQFycb6Zi27XFSmLR6b6+wSE+77hUECW81/aTb
/cce+1tSxWjKlUae9lnNYVwZBMLORX3AXgBn9QJyIG9OAfUxyLb9liAzUCYtkKnF
IYM9K/sFblWwIFDEze5UHBXLcH3J3qbG+wUp6zZJBnkvYETz7MVglkxk369Zh6Cs
nYerjhBVvc2GG91Pkly2/zsF3vULFYmlWL6pgrvo+vyIO1hCy9m8el7U+CY1KtKU
cDMsAPMmBZHfr6iaUVbEq9JFy2Fa+jgPGU9BttbqholCVh3eYC0sbjJcm7A52lMV
y5ss5q+cxU1WZ+YKM915JLxwO5qZLkFUl+5bYtDRmt6BQpdTYM0T7+GVNp6ziGwO
mAw2ofN0ALf+gNbfmTugxekwsBKJ+ajadfjZCTM454LTqmHXmR0VLECQCH48ohu6
xCtto+kfBO7X3nX+pJoTguTEa/kOHGFfYGNuAjZC7Y+a/j+EE3yCzBagB79dq/+u
SwNe8/aI5W99QGl1EeONvbMSCwHol0RaYllxu7bkL8g6wGMzYq0pRI0S+iWaP3ed
opvQYY85AY6Gc2HZiuy71djx9h2liUhs8MzgkmkvSIvLVsLNhoS4tJXGiAfXRmab
2/VDAfcs+aIPYiyuYwFA2gDsfTg7S9AOKMNGv43SROKcFaOjtcZgkYssGaQ4mJ+W
hrY7oq9QkeHLkVAeCqDkGjapPBxFoeVVUT9urWJtgqeULkK+LfKlNpPybGYTMABO
PhNqL1p5RFGNmm8YGtQkOjY2tNZmFrSsUWyLMf3poFmIWOY3/psGzg60Dd13VsmL
KhMO5rTZDKpJJmuvQR/nrUzmjSaAK6t5HYXVgtjRvTBqnD5dT5Itbs0F7TbAaTRH
pRdkaI1TNeYuJ1vSeb60bU/Gb6URtZg0tsM//WnWubTah99FfY9ql6zDBweHX7bO
1XQYvVmd6vemN9IQUqY0miskwS3i+MU+Ra9WbzjxqHwfmSj+omEYjxLaERgK/90n
xlhx1CqQPLISKhwOJfUfYReDeXaBJYIWTJOPsbHau17e8tcX/LhR8sm9KwmSgWMs
+KAyL0DhOGd6AaVcpTp1pJHB+5p4up2JyRX0jakI/+nde625bTe9650Hz+Y5mOKn
uzlpypBbYvAGpj85m8fArqL1uzfBxFJSHQInLXgNy8oX0L61G2ooPB3swSjI1ijS
z0gFYaotlSq1D+TN+id8hxd1EXTQbO76YIACFfk/6yH8QlnuypSniACmZEIFcTwb
swHwO7NeuRq2oNXSutiOwjRGUSHIEJLJ4AzG7CE1eGqP9Fe+GO1NpUlhKhM7SaB7
Z0RI7sJFYNKlzRPpTVVfKX6A6F2dTo0HDs2JbFn198xxr3vfZ6CX+qJQQy09lLls
gT+TTOlDjj+eRUK95qsQCviO9Tm4KGL7EzaB7tqiSNMV5iP6xqOI1AFopFnSSlrt
2dR4IrJRMfuKxhCV45fj6KXQa3srf+QtVi/XFEZOFDQ608qR0/11Ejr5tXj6Rt21
36P3Tgy4rqm0OmIc0xwhut6w0Exlc2M9GIijBn9EBjNY5esWUGkcUMEw+gkG2oA2
04eK2pwZ8MvTunAQkm1xDoNpjXU3jHldxiqtIlwQSMsn3CoIqTfLO9ZQHh3McU8B
Rch+yCPqRTvmeH5mPxzlEuVGVxwQ2Dl+k0WQCvzAChwMydfqDz9J0tDm/mJUVwgt
jtE0iyaNTfq+kpeCiGcsy/ri50oY3XTkK9KbSWdUBMRwHt+1sTyp2PkPMHdji0w7
AdSe+JQbu36ltk9ZByS0cIS17tJ4ScXpyk3bF9KTgdWYwT4oXH4T0KqeDfSYlodC
FYhEWDvjNfx6Gko0J9YvPwXryl8ifFwuxUVRcWinuiME0vLW0Yu6cWphIC1IMT5z
Pbcok9Myr0S+YIAeEATKe7+6FQ8h6cJkOK68nnIOSYVoC0yhwMQjo14kHjUSCIPc
fDAizxFeppJdpiDHRyktXlfR3i8Y+7qQ5w00m3EYRq1nOolWxnOm1GIveBXjSOUh
hVWCx6TPFr6Y23otA1Uvln+nS07LapXb3/ioUVW63ckjSl2X7pZlTEOj/VWO/Pw4
MzKP1ZdkZUzslXnUukRV7zxgq0QpW2vW/mw5UMbGuaeL8kiaOESVR8fZw1NZbY+q
aHdREJKnOxQi3TC2YbdRBJTXqXjPXHBMfMcMnNDVTuw25XLnXXNb57H5kMcAutOQ
zEMW2hTbQzmHPH0mRqDxEwrViQhazL0MAzOeeAbiZhWtZRl5/wGxeisM/KBuW6OO
LPr0btHb2Og6dZ0J0fXpPxfCnFuiuQ3+QB8Usy+7RqkIjxRfnuyQ7h9AUSHP/nn+
csUL2gVtvCuMq6VLWB815wtkO2OJDcm/Xm1c3sMpAjQC7ev3BBOKjlfKtdApvBxA
cXnAk8FcgrFbcC89ZTQ6tWzGMMNtuespoCcyKlzkMgpxvteDbSK37yBt5FzV/xfp
45vTL543ZKm6WzbAT6j39iZFxmCWx9C504EBhANsjJQo8WQr9wONVB7mX1J7ABbo
FoqwLYvqnzl2DY0m1WsduSNiiu5034YhiNdRnR5D9xIPUDfZoZQ3bgfflF15SgOE
slfFDxt6ZzK2mMzZhNwEHc9YcTO8ghI042fUp7HgFHJ2SgkNYZhMCF8pxsQkjFtR
tFbiI8fstCegyc59+QttsClHQsPtj7XT22CY36fwHnB2qNZLi8bSr8hfPstu7dNI
OlhAp0iS1OieCL0QVj99G5DD/EJgBZOrNNk+3nt7HOjmsxDzqmdzrGS8vs3fhcXq
CxleOlGJQw+hAIZdP9QBye+a12UqnEKXQ/26fJhNngMS3TfItADFRcZc+p0zV1Kg
lZ4P6Ief/sx4DawdBRXUVlpFaC6f+3qAccrET2C+EjbHFN5VsahlWMCmsuDnEnbG
IXkfyPu2WjXsJotB6qdcg97gAJf0KcZ78jPJCO/LdSYjHiw4Xz+WESbDKRcpF8Yp
XeMnCxTuy/DwgFmhQOhNWiwaa0z/PI66jVUkckl2eKcUdSIjzWYU7nOcCsnJLQnC
TUU+OJh/Fke9RXcV+fH6u23/qhJUHfwoMDzpIFSZfza2aWWWmNbY/lRbfyHpPKgB
cEeDQL+J29NdVY+eDrREDM9KHtEhoItOUcSXEWN23WbKxQ/ufKijpOkO0BOIH2y+
3XdS4pWw1IqjTZzfjN4DyvtRthXoM/emK6rZYD0ZHvU0SYeUhCZ68xA1VU4NReJx
Nb44qiMEuxSSoXfl+Ece0eUd2W39xlQjo75t5DgfTtsTk31CmW3c8ZUWqU5BwQhf
/dQ2kfmx385DdXNI3xApgGnBZmo03YNNkyfsuwv6JSF8giUR/n6rmm3wa41YWV0W
lOBlihO+o32tA6fabl2+TMLBiWrIR1ZiWWIQzgndiAyLJznjAMXwQzmZbrVmE4nb
ws/1/YY6M63+GI3L5XEl+iKnTehGxbhaKThJdMtc2CSlKCr3R8i9EI8kATSfQPkl
8arl9j03yb1LyH4Xpa1cLDqgghCcF791nzU90tviRcAsR9SR4/UbmnbjMiIBiKXx
7l7Oum9MG+7u0653+QjK9lg/ErpyxaE38sEWB52tqAq9s5Zo988o+aT2iiDfAQcE
nqag968Zq2NM7bZzAAsL9ji2fnnJcIBo74pRuwH1QhX+0hAOJq0pVlGKxbAB95p8
jFgTloMaW0PWE8lfj1o2Digiha6wNWWBgbvJVBzgmZYSqSZy3oxlWXOSVT6aDJmf
Q6tSrnDPiwD5H1oPzNWH++70f3CskgI3Eo9kgT8ruKN1kc/CPHQzA0JDwLAcFRNq
zRH7xzjqS9bE2P4wHxYePVNpuxxYBhe5kAtAkJXxOT1qLGw5BeNybfpEXVkJqAJ8
6S1ZWTePyq+ahmeFcowIeuVBCFqI9tJrZT/vf6SwJgC2SqA8NKmJ3rESqQ+fxZf7
nzfkWbrwYbuUv4cdcG29MFrBTdNhRulPGHCSfA25v1YeBZycjrnSK0c0GnaVrZ9l
jJFBkkjyet0RtYYc7MroJCZWmj27A7tZ0FLGOnWi4sCpa1OBov5v1PBc+UbTIHKy
eAMgOiE6md/JwKxQR30XOpyokGQYSKVsaf7a1Jx9BSHUIEo5ccw4HC6IhhoKsPWN
2WX7P82K4u6ozuVxZE4FyiFhvOd5sGMwysy8qkVTTSRyLeqy9gron01X0UVkyqTZ
w1EB3xPGILbW4N75rSvGpSSBaV3tYW/QJdkbKJ64wv8lblRLeLOLmNKZDocqhc+o
vXYSIi7tAIr+5+Wa8EMbUuRciNyPjxaRhnEtOInFme7qRyZ1WV1bWPWtf8IjWFuP
+XeetvCdRx9UYHiyGLAtrNBwtPTQl9tivHbMSrj2k8gq9p2gt7YPWpPoFAN/vUVG
+BcJRfLZ12eiI1ISfTryqBEDq9Gc1qFgfoI86r7Tq1ie50pwVR09NcYTMnEm75M7
CfQXtY6TjDDmBcsCvmiouwsoaTDf7BxtyrRupesUDvo9N/VcYWpDRvLDB4f2GNu4
Tl27yoAHtFoglhJlHaGWX29tgVzUBVpVpHE2ESM7+DniBsk5zr4Iju4hq58hECsq
zKWSOf1NmzxCmcO9EbqRtqHdWdWaZdMhY7o1lsnRkjFNUEquroxd3sisKsbzU4H0
TOGQj6SqdJVXC8F3mEi66plvcVLQfOIJxnzuzJx3CvOQIofeFpr5VLv9CS//Rk1b
La3ETvqSoUZ/4NK5vQTRDzod8QyPNtV9P7TfCL9EmV8DtR6IfcmnAfRfXaeuWX4U
UeI29N/kxvhEIOdgHdlASjswxg1fQrei8CFwbhVHBYef69kDLcCsEoKLXXdusVcM
w9xGTtZCkfOWgzke3xWgwR3If5c1h0FNZVFnbNUnMHHtQOLfZJ46KKiNwmiZTqQQ
2coYP3icMecY0kdYZ2A+Hf6oK3lFprrZyNGIH+hzDuKuUblxDdTRn6LPLyCTY+dj
3xF0veIOpa0emo/fBNHc/eAy4zho+ldPwbwK1nx6wNq4j5NV4WPnNOatQwPLWAWC
OOhGOMXoFR4+YPen/h5IV5i/moEYeEJ2QzJDX5SdGFPBWbz3ZpbswQmJInrbpta/
uxBlkuk1BQQeqsaTilfksd6IhJS4KbbIErnEeA9UX0MTWiqD7Lb6FimXkRFlGmvL
wRMYd62cH54qwWhT7dethbtBoYEb2CUoK6pafS+7hPcHAAOqDYthhVaXB7k3y3+D
aseG0XMzC9QBMhW6hYdgdbEXBDlbwzWI7BiTxlWBmzQgiC8ZClYaWsQmObJEmp8D
v2Cip0XIB3hC0bPm0KdWhR2v/KmXR4thVgGKB1wXSh3dpRUBIy9K1K46UaDojFdR
lwgC2p9sibYE5zUS9809aREzfFjuoT039h8ybNMf2ZXoUf49MlSXeWt9gGzD1ZlC
5wtgezzTyilWX9mmTExANkaFPVBlKr3Caj3LrQsSCFetFkvh+YypblRBRcc6CVeM
T0eDXfa8SfX2RwIyy7nboWKieYud8XZhSFT8EfcxrI2wdp8p5BRFkx7WFL6okN+N
Q/HRosFuJEDwttXGnQlKA+BSpaT6eiK+fPDJ78yDeIN+EWrj/eE593p/UU40Gd83
6oYil2aaQd3pRSQszAf3e5Ptxm8JitDGAmbbQ1Zul75uYDokHxJKNDC5Clmi4Ojk
djgj8VsbWS8BQjnBumPzXHADoEQCNLM9wlTTdIMS1Cau5I88cajJVVa/N/P5xl5c
KIpOsBcittCELnw3E0hL72z0KFJ1cVInMZa//+8+L2k64IqOFj+O/1T4mMpmZ0xp
OgE4YhSh4vP4lOSd4BhQxZGwvuWGSswDjE4RbnUvlTGvLN88GXF+D2fbFEzuHEpB
/J7YeKLTgIPUhISpBl6VR0UxcbeBtGtOcXaNwxw5Urmh7YomTKmH5OyhaIoBAjhW
RcpxSPBaBXfCl5/gIoilIoEO8BnTHcjdkc1kdZQpR3D97/bKfbUTL/E5/+A849gN
ZGUAi9oclwbV7ju03p/pWavzuY1mi6SDm14aqzvbQBTeRY1joE2WDbHQrMn2S/ru
czGgTLp2F8sgl2ohHpoxeO3Ge+3cSkN05HWZY4CYg5INMeAoTvPfAejTynPGwVDJ
22ONN/hpXGxtHxZfrd/yW2vgMQjg/1wTX98RTpvl3Lpw/TSHHjiRqko0vg6Hub9C
LYSXFwMp2KxacMIxHCRTvLSWzIRP7TS9feAG914Cokr9r8goy03yk4Mifw22W54f
AfVaGtADVvVR/84Uly3msMEZiIjmmwWAZQ/pYwTTacB0M5WvOyGAspNNthc90Im7
bj8LmyDa4JhkFT5pv42Mq0XNyUckIBKN+d/lnEGY/Beh4Sr4izTs5yR7cINhQYWK
AXiIf34FBMKjUNPZ3Knn3rAkOdOhpfPhqXlIcQmyypqMq/CE296Drr75FwIR0b01
KVz0QZRKpRAHUbuHDqXiL103145lPUYiymxK9D3D+UoD7s146JwetYhm6Ncwr1i+
VK82wlZAkz9xx9yMERlK8aYCbC5UqQ3JtljF1iI2sY8isgpQ9lVSMhoVpLKP+/bW
ftMBYDs16jI7iVHJcSXoc+mF9vlrSGiD8xn6Wka9eyvf2o21jjhf+Yv8hM88SjY6
z1+LqYtuKCj0QroR9GHHAp5OZMI0nVLa4eZ9VVyfOxVtSp5R4LqM7TG/Hd9TiZYf
NVMHPeRuBzWCy1A7x00YX7a3bptkt9qm3x33LryHXdllXvczclphzAW5Qr38sXGN
192eU3Ov8A+E64XH5gLW711bEVzwSkbEsIZutu/EdaDv1cFAbDnO+1cNJFKuccQ+
XH1V+/+ayd6A+nMSL+2tovJTVzZx4fQknoHFalctY1bEvQ+dxXziBTK6pyeheveU
OiXI0hylqRfHBUz54TxY58NizkqG1n4ncqRbZZBhxZKXTiFuVYrtiaXzxVIhgRzf
IN998vYfLMWjS7PLapIgLq4J80PGMN36O0BRjx7kVe1t7au3qHCRHn+/SzcO5ZBM
lKJn+HmeweP5et0ZvoylhVJFD1ep2mxVAVLqO7+pvYwWhkmd9HYkqcfQpnwJwudp
oygfZlHkUEM5VC3QFHQ/w4uVJBHpr/6PwXsWQZC8bqqzltZhbR1xXKqi2RQCNp6B
bNtFJVD+tFZavHajm3p03TqeVCzSpXcWxL3Ig1M0h6LjMjOHHvG2bkOvODquiuJc
bWYdaxY3hq06T5rlCh97froadQjPiPKd1t0/KGSTqYIbj1/ctUGISFz0MQExcrXF
DcUZkB4zCrPv6Y71OCRnbN3InNuHLY93rKNpUSEh86WKC+1lxb7rISgnXjTGZYBP
uDo+wjUkf9h6LSl6O7Hvn2X6Xu5cIqecMj9uvxeVegtIeqPZ5WmuH5kaXVVorXte
FAFeLl1ZcgOpox5KanPsbOVzUhYBmnKLQSoQkVoQFWYwtUY8QfGlSFxMYWtN3Ryv
Y4XSgYuc4bxgscSXxrYxudBCueKZhE1TyPlrmy5G9ORQ7LlxgZecavKV6iFxilEH
8DQ9YedyqsPLPXpH15w5dDCsVfLrafKgozYbwzUEjnSRYz5k/gK89fhcC1zjy9vL
6J/q16C86uetEKOwIQn/pnqxmp7yANh//VhzBmIV6TigaGOp/O1zaok/u2ONufkQ
W9Cthbs7MoJzSHhXuBTMD6MUCdAplaoYorTYoy0lWOVANZg6aBNzwO/PtXQ21R2w
jjyyBLedf1PEpt6hFvuynyyW46e6zX2/nxJnu4jTRq62DntpupbpRekkVl1wD7k+
MCkOBUcoVmXQRZqJpJm0RDUHq5Pmhg795f2evTeDoWVrf89/ZS7p9iafIRhGxHSr
uTXTdsDzvcmL2kGuHLDjjaX2bVC8cx4Fg2PgPuzkP+aTyO6pi/R3LDCKTE8lvQP3
ig/xlovG3+yYJSRZsQqOi4PcRnAlyZl2aEqNr4p8UdRxQGXhYVK3Qp6rgpsfb/aV
SKQYXAIL8xR7wuix66DCMVZ9Jaoe5NEWz7Fx7QAOFq57FsT6uQW9kFqqresJQQYh
8iyiYkGz+LP9sMyrvh1bFSnp4qv5rFLWqzD7Jr3tlbEGKmv9xEL+cvZQogfeqNzs
DC/z9ZWn493BXGfL71OYWs3QxOwEn/l5B8Gyk+QuYY96Qln/N+dCgcnbk3xqnfwk
1krRBnmwjjIxcDvpB3ur2JR9PZM6nVONjCZkPMV+LeWNXH7mQSPUbI4M4TAI40xH
aIMX+rd9GCWdCkiaZ6NKDItyhttEvblM7H71MAxE5RrdfS9UALhJ3ZoyH6pJ1xKk
+cEUmQ23iAGbaZitpQTPLsqNY0E1nQDofOD8rELY1KmUCtBOawGySTWTYnQRtfqx
AUwY9TN2UnOfbn7CtvNsAoGPMMXL6qrxSVcqdmNrYf/1e9oDvfmjT4ElEOS6T1cS
rpmtpmp+OWWrpyiaOY9YTBM1TkKu45J6Z0+39zYRDTUj/yva2t60tFOlGvtkvaFn
//OMa//2sNoLI6DGLzVBnzUqiXGIAshfhzb0P600NXS5RNaf3B4oFxYegePigAZZ
+mF1qDXp0LdJbam6gTUh9xISN5ZHTmjQlOZzxr6v3w80MIh5bfwxWZZuZRIMmKwe
HyNSD81pJFN2W1Cxv/2NM36H0suUxGI94HEv+aCjeBOOfHeRumcmNoCv8nSnPTj/
/6mPCAxA8NNM2s3nmObGfUZMvFB1/j02Gp9G2O+DJSQ+QAEUKt7iWYWi2w0BJqzZ
/sR2TYS0WSChlIyGXdm4w4j5Ze7WBCB7drbXVmwAyxN3As4EdSUKTFmT9nUoBztr
RFf9nWNGfj3MSO33FMgDr7tAjLnO2l45O3jv6Fal2vNOEV7O64pf/5UF5jJ1aFRH
B0c7T9rcmO7Hhuqpi75WRwakVipjNxP3hC9pN9AWAOL+8OG3y68Ocr2dXwYtn46I
AF8ZVFDRiEQGWoYSaJnXK3jxGFGOaDZXKqYbxdaaogykkQdOuOh951AL/DrAyss8
dYV33KKff+RWsU8rVHK/FuqHcwnHq0ddyal74IVHFsyptADEDy9yKzLl+DlyDlle
QaHxszRnreMBDxaSWUqVErqk79nRhmAqZ1eGfXN4UMTmAsvwUcK+lsaCOSc0OscF
7WZcIy4b/pV9KEbUlJ8JNvxC+/vceWFYDvEUdaFP6cuvpsyLoUiCTE5ffxhOSrYJ
900ZSW/Iu0OAE7FEVmvVGsj7EPszoIdXbPqeeXzgF3bNOTDCkdVafV09b8JpZIaC
DKcF6h3p9Ya7zZ8Jsfmgak7hiyxV3rOP91OxHkzr45iqP+mvulX8P2atFY3xDCB5
/prFzzF2obabHaKg4cNO6IrXeP/WsmAeWoUrpqFDmJJifFzs9JeWp2obv76/2oFs
6r75CBsP2pL+7CnYDGyfKoqkvcS52NVYxODzz8RJ/BH2ZQBZ38BlupBPWIyYQO01
PP+jgzrIw1DCF5R5Uioc9dPwo7X0sN2sYx829DrLrQxyERWFuYSpm5OB5QHevZVj
QKLja1xW+z3ubYGjSItQOCBQduahAjVzVBREYflLP46EHbd/bfaU4xhI2O4TF/m5
l+vHMAVIvXSWxd7aaufxSwCqaxOg0sKLTBxXyw+oQP2nsnrdzPfcw8gsDV5Vm6Cc
Rf0QPcZ4o/05ahn/1A6Ff4r3ySnFWewpGaNiUZVPxBSGQ/C6AIImlQFZtmOyvwVa
t7Txiah2aMKG5jEek9Tx8FsUIDnW/t8hK8Syrizu6Onroaz+2tlGgQHg77PqDNT7
oRZ/ci6gPGZQNELSmV+h+m5cPjhMu4od0DuVcVdMHLFxbJgIzTofM/kd20rSL2A5
psajBy7ak3Y2XYHokf0KR+APR55qyTvDisobmh3pZ/YW1Q0E2lpjat/0V0RR7io+
VWaDzWd9oMxGnV6oV43/y5IRzUtF21s0furSx/L9HtJ2GflgGIXT2XuNKRAJKsQx
85ey0Vw0D6/Zifd/HErXFt9AZz8O8xYDbSKICuwVhg0dfeip/XvdHirzsFu+wYyA
ysVH9+0cMIhs6Hk/JsGUREVtEuHk9ql3JpWbTj8nnuuWySLbYi/NXnh9LlZv6WOo
tygIkCU2pvV9sy/BPy459tV8irbU1YtidwTG7FY04OAb8yg6NYlst2ypfP1S+rOn
fNj5uuaGmAgBygvm5uxRnaOHVlohAQRshaIquHcDwMV5LOgKMBXN+yDqgGf3qtu8
HctmIKmaIGPrmbXFOZIlBM4tBFruAGWl3fjqobvb5Or/NSYnS56GSHRtdeZPD3Qv
ulbhrdl1qdvsR4qDAbGwjcUG8rGtLogDqHal/UrHENqVDp1rAZZqT7KP56bb25xJ
wOyQXOMmFG9i8vPaKVHQ6ZHv+SkaxcXqmjcfIhIl2DlmxUTLLI17T7TEXIZrOkR3
n/hAcma1jimSaNuHypePeIT9knV1s2CeCEUuPp2y0AKrtK9kLWUbBMcPlDVpDyE5
puzvJEwDNINQd6WGp06O46LDtDvlVov/gwZ9ntTfCQvG0ep7itwzx1b8i0ur2R+x
YdtHu6sD5JdslNL5ln6Yk0X88SEKTiG4V+47jvQOrX5Dj/qQxK4+Dct/LxGYzj8k
rTZ8MUodeW/yXhpcAKsgEYSKlrL0uegy72TY7e/Nxz9ErOYiakP/UVwgvPasJchs
XvEotFLQ6WcOWKzN60jpsrdJTz6Ey53PnrgDN1zccPJ35GvyKrmrEG1auKY9NTiA
jolQu01WmK/uA3M5I4oYOxov/vmLgJgr2GVhzeTMPH1gGobc66W6LUkPcGhTSL55
4rRl6Ef5AS6NAets61Vl0rECVEnAIR3n4atfrqLbR0+kMVminbDQ2R0MLqstbC9+
pOOynQWVs5p369IZdZNo3RGhuij1bZLfOCJ6+riYk4Q95Pdyxp0haZYKD5Z2HB5m
qxc/XTKKETb/Rva+U2EHXYKy1x9NwcUuQgvVePoEPi15/g3rVBe7Xhtk/T1O6hvd
rBua6xoyJdBxmdVN4tgfdCY5tS/QkbkC05GJmy1L3QvXX4kB2d5LHXNtLpHNz5n4
LMqPTeMuvmVhaoJgkU8SgfSeBRkHIKqpaNoaRyjz06UnS8ao1ulNQG8c/OKaJYbL
aZfM8FdjnNo5B6fANNMlDKeOSQOSajj0Z7SnK1lqAreUp0NIE7GShY33x6fZ6nnm
T6UNL+KzmXr3w5OTedP7H82pWUM85+mudZlPc2XaUc/NvZks6LxesmcBS/30JF27
ibmvuuLnNWt3Oex1SSAQs5YLeCcKYHDCfUzaKhMbXWKZdANoUWL9QKNCbHDorczb
IPYFWmCc1ADaRt6LEWXQgDhOPsVpBGKvU7NH8EDJREwyO3+AcomYeCtiM85NkPO0
NBJMgXGJHjlnKPiuUNuKUyHfoFv4SW1gKjb0k9x5U+x2UqlzXMHqa/l7RN9AX5vR
sFZEH+hM2Iuan8YOFSmnU2fbFqbfor+GT8BRUFJctMYEhNeAZHKjOenT5hWR1IdQ
t5tj2xmJvzk8v3aLrWgu0ysJJ+qnwhrNtXjEXnmzgZRfUr29h5e1fra/e+iwE9CO
IRMZX5VCoYRyPSC1uMXwTHMyCOmDlPYfNBh9wE8IUxRRRjtcalZiZ4R+syLclFM6
FV64NGUZd57EpiY5Aw6yvIB2/1eZypiQJP9ebi6HLXwa1Xg8imhyAiFZ/xo4RV/N
7OxmZXmImnqu77qCKOIxH2nfihYkISRUeOiN3oPseyQM+wthwAqEeCwXnKxlVLlj
biSOH/EhAa12fX5akVtbsdM3sqtDlkXHZtiMy8HrtYiq0FTeUHCer+NLoYZhwkmg
6gYvZwq/L6r4XeJ2/OzYC+jC+kZIS7X54O+WeHOe6NrI35OXcZs9YAIUYI99V6Yr
OIEjXUqQIPfDEZkyK3v6p6ZTx0AV3sRnBiuhsAPYUGIRhCTgcfkAonZjHJ+FqIkp
qk00QwsxIEMMQR6JrVUU3CP8w76WfV5rCmaEhQli38JIrXOaCAhh1oWxpYnZx1cb
9oOX6fWhLq5kxoZ4HoqW9qzlcgojVNuxhc7ax/QXSvYwj0txiEfxDvWkBx6sQe4q
wIVzFbcqh2U1i+7z+O60aCc7YltrHBkCFTo6DTxtmzGDXj9x9Fgf/C4tIBy1ehr9
rJlf7a4Rw6VmteLUMjzWmI6FRomNiG7L/hnizlDcKx2OAL0KxBZU9jRQgUSz6tN3
WnCGBJsLMjFD+odQfvuQrd2I1xMKChbeo8dcsLDaG9BV6tDVY+8lZRGhD1sdWhrz
ZzcxdOc31yaFPJU/ZFdqondF/gFqPgnGlJnwBB6g3eq6VPBXpf9jMU4rUvntHk4x
trSfq4M1V3AWBzGaPKdXBPpDM8SnGCYc5Rd9qkVJMcG+YtmC5yrwaRSN74oYRsit
Lr/HihEfAi2ltp1MCwdongeOZhCs7oaWCQOyMe3GXAoBoBxFXc8f2CiH97j3f1Gq
uUXVNj3OnGnBxAmLFrPYnpvpZSRWsKL3hCpB56Qc8d01fNxRDTlDNy7HsoOkYKa3
vSxB5NM9/WLY8I1ppc0DZ+Ec27t/+mY3Lydbh63WUBORcAeL/bpBWr3LMtoTDbOu
1U8RxfiHy57hX/WuZzjaNlbC+Uzeh7hoJaxKlLbRE5P96K6nmtIT8zqWqD/rn46p
dzLk9ESAMFAVuZxBWw2AD/USkF4H4QOP0RBd7UBFysoYF4IhbLJPYpq9sJEAcKaP
i4WCLtFjM5qW/ClfDmWeQGE/S6tgbAl0niR+LfNtymKjNZPU/iyPqhP1yXHVtf+9
M25vfdfX6wp3tJ67aBG6TX93OauSqSrO8VZCWllLx/A2d1ViGhtwHLFVb3rGJuWf
VqJIDnWzOP0pjxbGwIz3xpeQk3ehKISgzoHnx38TPeHqD3C9ozdrihFrWNKN9BtT
RsitXbP63ONfrqbDZJ315gs45V8FgUVUs99jGnVy2+wacgimnp/JVBcXQGZFWY8R
IAZKZJD0qAk6ybe883pefMgMDxh/JSOA96JfzGEPHK+EqSjfMR6E+usijEvXsKhX
owc03nN/xLFW5DN+JE9oqR2UWYHCnBpQsdk3Rgsq1c4xYLvvQBRGyhr2ldiBtr8T
b4bAcZ2r8MFYlEMYWJVlsJ/SE0QYI8D3+aBSU4cZKpEcb54L5GpJHXyqbbmRnl9j
9xT/yM3E7+2ZZ4sdy7Tl1k8kF8fVRCJap0f1BpQvjZhw3FcfaC+9F5LTHSD8hrWQ
dcFeyJLd8b3EHb1WBeM/qNIsDeQqC9FsVCF3NnWIb9N5juafQae1Srrsi+5EnwXz
QppkUK5Uft/NAthG3Mo/ubn5OnqjIIMjCCNcl0LYHpvWvDkNNhr5zKIH+HnAcWt+
NR0+WSWT4SwB6xrJxQ51CroEj2hWrb3o4REW8MWPtbUcG2vhoX8H0aBBLBaGORd4
KURiQNm4HLT7AN9LK3gq5oXhantqy+A3TXkNfLeM+vVLRHSs4viY6LVuTycTCKEw
5Au99erRZlTMIyuYeDleFrQLiEzw+vEDyKvtChV5Lo2dnQsDvTpweCvns4u292G2
4BijCOS8JM+npQurRgtWYEZn/wNN4KJ9IvBMzjfnqmJ2+/phRJdd0/NOoh92WX8E
3eUvm0B+nsYYBTsMdYe1H/Ky7wfHrpGfdTi5uMwKX6bm1XvHqbZIOCnY42vFdOeq
TYLnqRC7RiMzfjaOo/WmYugP9LvILlRjbzwy3LvLEbVYuYdxJe13b0h7JkSVvP2r
nxobY6q1P7hFHnmjYHg7CbVwbSL7ccvtlGYXk7nrEC/nIx3jmAluL9k3sImZD9nG
DaVASrN04VNki50whR63XxrGl83E9nQpwoZNn+Eyx34VKp4Lt99WnN1m3JX1dm/U
bffD2EKl3ofc2AslFB6W6CjeSrfIadYnFitppVoJx5eGXUD7aDK2HulKHhP1wZpz
M5RQaNTVWxJ4Ei763PGpbZOUdUd/gBOZIEQ1sMAs+DLgunKdV9KslaZHIdPptEsa
q4tQUg8SGzHnSn4+nOWzBfPbLndE3/kp87vfOGOq8TItZPk/q/pXBahL1td0D9QY
aZjDuDc0N2PrXUXSa65i+qT9MmEYSTUpmstWFHJAbWZWIkC66dclVyjv3ItlsjNH
IKlG8+DCZfju4nAqMR1J8bABriawooIiaiqPDtLbgpaC7cJARx4G+C2Sxdw5Rooo
ukPKrnIRBlToW5TWk8K+bFtyFfvfrJ4cHqMb79bBxZioo1sgqa/UFJpDVEhioPaI
/Y0j+f1Skg4EC4IjlXdkyp8lAo6UNVwPv+99RVNAmyVi9J2NzuEbqn6C9OchnMa3
LJ1138Pu2RQZngrV9Qwcf1sPt/FW1n8zPGOx8jKcupeI9k1E2Hq27TusR629rpsd
PM+SRv0/hRgdhvjK9VodSXb+X+YQ7Tsu1InRKbtvC81FVFykvIlwFfJqcYD7vqcG
OxwCR1NTKCkZk9HivtkgP5hqaMfeSgxJuwxiEF6D4kQ0V8nNV2IJ+2jgneOgB+Kj
liJhg6Hc+jZyM3MPWF2bWbeZcPzePbR+oiz4N4e4sf4BAwWL0vf5Tm8dWvPVkSVp
e0s6njqpZjVUa3BFlleSjt6dOBGzQoRHWB6j0zVbHpxa532H7iyJZk9h2JkeZfdF
NQoKxWP5clpNIxFExpFrDKKrX/a1mElQeXl1/rGm0GvbQIW95ZD35IK5O1Ilf2vA
IRfJ1wUXkFK91a9UEjFNhWPrMqhcnlhqhTz/lw6cQFdVD1XqKCJ9QUmrSMzWZqR5
4pDgnbaAExy+JCdAciDicdUjoS128WLTsswdNw5Iabu34aS7dQ4JkfmrpnQcwvJh
khbn781sq499gkplDnQsWMOw+F+VOqFtltI/YiydYtjAJYlczlO2PrOBgTQuogiW
JsS3cc6yCw2wERHkKHNJDp+LRM1/rPcaYZRpol3kOy0QBcR4e0bTj2BATgPY17eB
ZxnBMj4bVyC0npHS5hbNsoeegINbnf3xXJQjGZ+MzvRTTKZ4voMIBQGK/0nfBja4
SBHSFQ59ueUTVj3I96o48XiDDB9lQdEzndSwmyhf9XO8+U+mAklIylG4You4GeBi
ru67VaWTkc6mc3LODz8UYm9AMfnFK795U9dugVjMD7QohQhbJQdw1l5g0m5q/G/2
0PK53s9wqk/hjKVS3KjkexUoYIwlYdGDJtHsxMETkOj9teMc7fU40uLdAbF64Gk8
nOX3vZrMw8+AJ+pEYQnrbdKC9AFSCP6IObpT5QYCJTzkEDYHAu3ZTJpJc0xhqFSE
jRQGtPg2xUQXnvjTH7mdqXTMe2xC5wlllnD1wjeuTtKDnAjvSIvJ8i27FLNp+TAu
T0gIm/IqrR42p4BWwbqFngb2sA1IdSMupMzpZQ/X1ID5YvoBzZo3c93G1I4bWpk8
PZFrkRS1SO6pgmUid0u9UIh/Odbg/aVfIVFXDo4C4HUoBi58bdYp1gYYUur2S6uH
l45lBkeI0qVsJpI6bGPiziuDAR0n9ydvRoN5lztXGdZ3dqxEq9m8KTIGWndQaA/V
u6eo4/iDWaYYiAx4m1poRPdk0uDdaU2eHPsMXwJ0o9eRznKNs5PPPGCJaEuM3iid
p3DRo2PbJ1kvCvaj2U+3/laHJfitJ2VXFCEvHJa70RP99SawBnxuVMLfALIrZExi
wT8V1/c6xt165lPGEwzBEjWRYOPYr4R7lBM6Y2klpcSpiddK6mR0TbCKazC3Q4qB
XTorhJEkGEAZla7RU8qyIBJmJBsu7TWwR4J3ECDH54Aq+2AICKbakZ6aFFmjEAVV
aMqju1zIPrDWlu/uESVvaAr7KjpxsXbvrteUSQWNzo3Hs03K3CM6KUNvxCG7G3GJ
woU/Zap2cmJQdsVTZTeSb/Fnb2i3XI0pWPEIFVzO1loPU3QUgT3nWKSRonWrGNdm
jtuWfwlbb/f8+J8dQl2xeDivRCw2y95ZbbsBZp5h/6Y+Yjg5jPbvVsFpvEEn3u+u
5hMJiQ0R2uwe9ZSSUcmaKqIugbU0rSpPaR2ArV8bS29jYPpgh/zN/yjXi9iXPQOg
6kuv3GPw57ue6NB4qETyr23JhJuyChIE78xfpeiVZ3AL1EI5ggLxLe23GFiw1JBP
EI+Hdl8xzaAksW30u0nDcdw0Sgy9DCSocRtm3PtUZthSO5146tceq+U4IJGa32mH
t7tpp6CgGl2eCSbjVqPO7a9TKJZvHVfXG4toSEo51V3zaIdBoMbb3H/tKemh79cb
l2gXwFaNGh5KCvkFINTM20hg5gL0QQKmvDr8GPLPjxvKiJszSm2Jvv1rrWY/nNLv
eEnacT9GACJhH2/y7fJlS0FOWBxByr3tNuy9JmU2nbDHi7lCEOHFf2GefseRvpnw
GsHMKLnjeZBx7NSBpZp7nqRJguGCZ7/SpH/HKkIdkiCTC4BrvjYAKVxBlcddjTaC
/0ZNbZDK2d/+tABMj7q84jzdS86zXOBZImKEWDJZ+BnsfoCVOR0hzI200+R1rlLR
KKzkpRVCTUSQ6XvqZWUx7vPWRp0H1kOmaDbaSK/B3XptB+ZwfchTYNKbvm5ZREtq
8wZq0itJpn5Qui2PVxK26T0T24p7DM18QofevtuhpHjCPk7C3EFhD7kKDv9Z5BLd
gi/1JHQ54H755T2EMwcOA9WNnWnUz0UvJtjLl1cA+AyTkoHG2CUx6P1nLZWMnSbm
aK2yyxKpkWtawYl5Fcr10krLizM3rThO/vRtcjV9Hz6O4c47l37SBM8EAcovgeiQ
Tid1D6oRQWNRldtMAmoQ1GvZeBeHOF8opxPpUUPcGdtbGUqfcUzUu/kLwW4xx2z0
un2sfOxpoGF179QlT1vG2xD/eGvmDwoLXjgs28Z7GI039DJcKbywgYOIw4zDt/G6
bibsRtKzXUK+Wx/2RxM4kLFfcvo2HRPP47k7rtnTFcUU7i6YNHTOHW1YRdYbHtn2
27lRpsM/C2cRiqz6++q/j1F/2AQMbOMWKzXOKcP6BhQn99bwMhCyQ1WkUY2fZBOA
kO0j3Im+JVEd6YCXbKaGmwfLuzA40uS3pfXA7zxG6tgau7sx2pMKKN290KrywSln
LjMm19aozJPtyQBdWjbM8LywtIviEtNBaXPR99qxjHILTQZplBdEMiJm0WigI/ol
SIjj7NX3B6Rd4pICOxcTdg9Ec2/gYY8sQt88ytQDRWumb7PeVeqJMMCfXIaVhlti
k9Meu4JbbFLImwqw9hNfNqvdmKa1jPMJQYdR5Gp/t3S0Vyw2AviYVYvAjo0dFnCJ
fbjAI/RYugbAaVnLY/MB//UU7wcxnwXWjzEXIzW6/Mgvjch5sDsDZHt59zN6aDnc
bb7LQ0Vlp9WzN168osdVdzGK9g2P8qu/rqHwQs1bNbWM4MK7KOBsqtwDcCEW0S9X
VkmFGTbOeltLD+KbyNyBqjJ7FfEFn6+FbTZ8yiMCgiwrVONyqzXb5Myfskk9kjex
iqVErf0xg2M2ndlz5xr630wIIPNg2lAYf1Qha0Zp1FeR8BKcBTKQyS+huU41pRg9
sQJ6r1hZt5WCoiwj6pSoccltHgwRjb6K4ePiuqmwhCAU/So9BCyeT6idYI+71+yS
NkVIgv0Lpn8/CTwrE+sOsvE6w7bLg6bsWVBwKQTEfVl/wU9kcYX0bOsTvdF9NMro
rNfHSGkvppHDxCqtVw+aXDnOzXocFkRxdFoZsOKoOhTxO3Kk3DeAh145aeB2ouXj
gSYBEQ5uySshq6OqIPX92at7l9oOPvKELeprW82I6yS6GBwu4vX0lBrNox1k59lX
CbJLjDcsvoxZ95uTawSWZcElW5lzQvaOibAU8jNKhbuzH5+oAn0fncZX2nK+n8Bk
m7YsVbDk/kKnvCb6pqg4XghlrKI2WGDjA/VzKIe832UgBpJXxuaI2R9yzE+bKkcC
oXaa0iNjVfZIE3dvBUwcXkWQHWLQd7e1GD6CrnwE0qNCPrVRht/EptfZ4rG/4J9P
Jkn5wJLNdpUpyDKFtp5wvL6SUMYl8j8GBhrJUY5VJQOf49wLj3LgrKCVZw8erctT
mFxHx1azi3/ADKPvxbHyFnISo+YeAqbp3rY4Yr7jiY1fgmt8NrCOXTzFDyt5a4Go
GXBqoHANDcRzfet5rcfilBXVqKGREJZrEOvP/Ynk27DwzVe90ugNU4k1PJSkyfTM
CaQG1Lqdt2cpPBGC72PMq9lJ7Jrm/WLAZtk2xJzkcUbVJyBDwUF89RWrwZWOu865
xAUYbG9adeQj6adw01GvKaJryUBJEmLGp/r6dxk+Zh1h4PQtKRj54b47EPxqo1D1
UR5y3nQVDDkiEOz77CZaWoAum9XXYRuJnVN6dZES7gg8JrB9tEGfmT+53/aIS7zv
19sa0VIKK1FwhEx/PKpOP1JR2QkkB4BByxi6/2+hyE92faJ6XTlgOyBwl80arr5V
+9G1Q0s9mcy5BrQzqH3AQw7Jn9Y97+2/NRIsuJ7Enpm1C4JCv5DvjKjPD8QQx4D+
1TsYebOlcT+urSMl1UEt7UqmgY7yMFOXxXwp986fNnJUUIuum5jt7I8WrQx5AG/o
408dxtvowhgl3B8h6Nn1gR7h2kYioihSei8UJpDscBSJpJq65iaoiylgmKW5gNrl
/DYPq7jahtS0i92faUZB0j2+30+y26ltmkfigY72zrHNHaPZFfozYukaogRjO0j0
mUU+OUU9X96hIq9Xhww78zTqK63klY4defEV3Ir5MwWncnFaxevBxULpRQ4V0WVO
ryUw2UdpzInqIvO8zrjgbYAOWfm5yelx8nR1m8xCiWkYA9WHBkDYOSxagTHOfcb4
ROZldXPzmaDQRR1nZ10TMYuhb1iuy8WU68npAR2o/Qp8r7cEN57r14s8MJeljwbR
t0Bjck/iCDZ6T+CdzMX1RsTWDQriU95mQoy9F0QDRb5cNA+yf88+XAsX7WXE53Na
9V345R2jMwiolrH/DNC3k54Zk2VbFurXikwvymgkMeay4mjlkKAJeRLwz1MFDiXw
JkeGYSzrAbJDREuRFiuNo1AF9VQUReFi3/U/ZoyulbECvuPQNnfCQeuxRg0yypn6
a/V8MJO02+YlnnL9LGgrOOOElrLbJU0U/7admpj4Y+hWu5pyv4yqSqgEuDlueO9K
3HrarSSwiW9+uKBSB3cgOxKClw//fEsF/ri5VNfgWOUSHQwIVqhvRrs17GeMHaes
mfpKpI/YA9MVUUQkea+vFpH47BN9xmjQOPyiepVZIL5dH8NJN9vXoSku0kFIac/b
sD9I2Lr0wUW9KA9+6WoqnqhTV5UE5f9sSYvyZ0ornKlkiwcXxEcgBptYV6W64e8y
Hl+ZBnVx9NLpQudEx+URVTV554FrGSi97c3+qUIsQypb+S6TPCJYQ6UQErGokAoG
KqlETLhzdn4sQ/Tw586v+pkBegUBxvLa817unmlCpPrOW6cVJwB2CMXxPU+6sL9L
gVFaFFLxAeU1Y8U6j4uRDhLCMStnJ9LL98ZN/NnlsfXM2UADl4DX68eF3wOGUpT/
i16sI1tOs91Wt6NqbWHbB4x0FkIeRnsVsaMov1LW85uiFau9qPjb2U21QFZYEb+w
2MSVlMyq+strSmCdXW7bJMVfps7c7rTiFv1cNeUBtRKFosFWS2VijSPy6GUOUO4m
q2bKwhf7T5BFDKdCQ6I9QvwVmF/aORxrsplvdg+J8xGoXLLbcO1BgIbW/XsqYhxV
hYDdNwTdThoFPs6W6FekiiioRxT6N9HecFcM1MAloY+uwYa7C7IjGrBdTQVUgeM1
Wpd+5867Ayc+jcfso+R8SH1B6L7OzkuO0VgVhbmZl32EfG7YfB0/z9vKhxceRyQi
sHLl/kdoZk5Z5wPZfaxSTITYPKxsK7lJC4VLlOO7o450e29hZyP56hBCkjbrlcrY
uVlluaqmMrt1jk3Mo+wYaR2Qr1qZ4j9XUE51MXbHxCfveEyVvoBB4eyjSadl9Kgq
Mvxt/H0cYgTCHl5w0rc9hG9UzIxUtGM6ClFCbZ8Gsa0E0DjYaEZyB6XBSkyAwIvF
7WHJ/3BAAhYJT6STUH3owj5x/AosiZkRHmXToYQD+452mVzAEBPqW/hC75UtBUX2
UFfn5AXWZfbRUKI+d3+QjkQxxa7MNuDqankohymBiANbrc0uVB2oDwXE2XSSazpx
llRXqARMwmEe+VE0kapmYiNmwevA0pb6g2SjyQMDeIT3qXf0PKJBrO4dENqAwU20
gGx5ztEMHjpQFGYRN4zva24dJXx72xKLhx0+oDcfbnot0GQnV6qskGbF65j8PukA
hZa7hwrKEENJDloXTCAkmdynjzNqQ8/RH+2ZYyqw0L4yJbBplARnyinXgd6oCR1S
Zu8RSqhoJIoYfcsl5+MbTVunQNN1iuPEgeSr/eUSlmVB3gjKOp7LBQAdIvBhIJLB
8+pQ4ThDOAu9ruPcd8ZWeD9mLAcEwlZAGJ/VytlnTtdDolq30JtepwaUiQlUxiJ0
QxUQ3VAMW00W09FMf8C9N6hOrU6fz5Z/Gg7jqn/5gxIDAwxdBWviKXzxrGbEX9gX
u0tGMCdG/4ZZl6HUDBR+0iUfYLNaWEjQShFLxh4iiRP2yb3jX0T1DeDEJxQI7LfD
F0oniAFSbvzWkJ8zgxCGtrH399sKh/m6pyusaaQBhIto0059gXkGI3oVtXmqZa51
8+1ZdKYz7Xr4BzVKN/QTAbmOzLEwvsqg7W8FPHSgAgZ4T6FXmhWIpt7sJnPaoyJN
s/yY3Orb1CVkTuWUighik1sl3AdLbvXyBPOvfgSNGvXuemsquQESLfZbcq/KdHDc
cTCGAvE7JIkug2C13xZkMHmzphT+kea/1U6TRFBRkxyX1QyUP8DVshn+h/Z6fbI+
Uq1Z0r8abKNBGLFFc+LOcViJTsmAAPE6mPdb9TQxcb53wM+1mvGv7lXMSx3Ca/A6
psqlFuYUb3Gn72l80igvIJxoMEX31tz3Gtd6QQOV+1JOG56MJLiBE0VkMKPsNHLl
xQ8i1QvKuobQaXE9nS8n0Ux1T2lHC4ERiRfgjb2D4JkTz6pXU/0aF8Fa8NOXs6do
QlBfF1blG3x/SZIWP0V6emDgBX1khHo1ywQXkSd9JIiqVpE/cEmWJkIkvy0YZt5d
PJ0S7fTHdYbOdT7j3xXsNYqkSRIP+5X4JL3DdBm5afDvaw1ApaqRNz8N79lV1oVu
AYWJo5F2Nhan3gve6wkkCPs20D5szGKMDR9wGmVjNC64ovF8OfoNcSd8EgM46IpT
mv6+vdvLaV/LxMk1yGuBj+G7OmV0sT9bDAoemusTyV4qSyZ9tD5Is3EAYXllBfyD
9nUaMi8XwSQlSsCRqcpG6NH8PbbBoITmTMVdsWOXXlVD92ZzinOWH2xburX/80cz
SVtE5D4XiYwrTkGjd0jbR0FqsaLrDt54PGhZS1qX2u+yQGWmPq5HjeDY0LDq+II7
jWN6IWT0HJnOIOCZKqdEuNFwNch0ArHxsY0mmKWFyE5SbzWy6zp8ycVLwJokL+/a
D2Sg0i4Mcwy5pmo1xLVUY8YYTdwezxCkIC99aQ3hy9KPmfzed/g5GF6QvqbgnAdi
VSNC5+6FOZ2KxKXdOsuJGxW0+nSGauaP0nfoC4Y5PtJ3xm/wFdZenj8kVu0RCKmY
ef+22P5nAF3s1bzCxg6I867Yyi+crTsy69mLfv3nk+G0C26jrr3QcT1p7IMcarLm
q+sqMJ3XMbySy/is2kUWoh4qO+b/RTsaA4CGy78NmHAhd3k1iRfky47lDYKu5hUu
bE8QfuvMuvUqY44krPJhnt/XTqmL+MA8wjP+lEniL2NIgYJKBL8SLtn9Xhsoj6YL
3nt04GvmpgktS7wkL0Vt8NmxTZ15i46M3F1leLyU8vi52YRYuTfvzdIzKHl+m5wF
Gf7ymVwCw4xDxHqYaBBpYAqZZph27bf90CigpTCO1ioEOps0oUKHwPTQnvclCZIa
J54SJa1p/1/WO/7po2DjWB1AEM1MhdxMdlWGms5BM5gWi5N9a9SREtu6d0MLisSl
Xm6ueNXYBbYBNfph1xNCP9uZ2sVcdZpj+HjZCXHoEuyFW7cllHRnP4cFOjHzEgp/
A9ZsHwkJTsRYy6hi4LOGRqnP+2ACD2TeW++1jTGctgF82SDzkk1EvakWDSHA562W
QEK5XxaHK45c5OQBvJ82Bvel0Cm/lbY4J3Eu8U6pqA9Qi/eZHLwgzACHV9fZ+Rul
P6MeTJQVtcn76CNIGZor5nP0X65FKmopo4I2iQzdGYZi667bVeiLVbQAK0sX9CRv
H38QYC66/YaJir1dJbZ42FlUXFix6MAcO5/jCCzKOqgT/1GVV86DNqj8USR7W/Qf
PJclGmYYotFe9CR+/M8TlE95lcVx/yGa31kn0IclaAq/Z9J74ajH+X+UluhgWqwi
sfQdK+GVFEfADWAVAyYHyqEiRU6oqYLQImhume5/21f+qr2rR0Hk1sgzaeOmZXBO
uwnYroOeSR+k4sD//LwcmXLXqD8MZu6zPCOsX/QCXmMy64oh70okh3KOjUWY48A9
qW6PCBGe+eM2AMgXy9MgNX/LsbYhvkOc8xF53+OvPLtS0sS10gXigQRf+Ih4dEx6
oVetlNkLLamZG01bL7qrKK/m0SgeXK6+zQyEqaGE6J21nn9oJ8kOJ/Sj4LlKDk/u
XtioZsWsa2NVy9MIFvLIkoGmryf4SBM7MEa5qNRyaWklFtAzRtuunpEqCy7WqVhC
40mdiM3Td3e3lJANl4D2fx8ql96p/82rF6BZmeWd0kiv7JEGC7QZ0J0y13ohhsGs
DP17dN/d4pRxZOszqKtnN0CtR4gI3lSUpDDW9KwTMaZbVJrwP6+XKbuHHvkawVc0
ex39488IZeJnuekcG8NAFrlxUdNVIiTzBVkaBN4jjQpHGE84ykVjs//stmV5+ALu
1EEExbknNXeqe6AFVJZB1lbOJneW+iFdGiFLCMepb3Q2CyBidCDE3Q3B++KpwZsy
qUrgjCI8tFmFMfVi/sJ8NHxi7OU35aQHhaW34MmQt5ewdCahjA+0opjEinow+EFd
Q2v3t7mf0nclqCE7uecBWsYMkjjV6G9sXGXVHFDyg6d+fqqumudqtlFFmfpczufO
svc23pw3ODQgCMBT84D7rjKHI9XWQN3PomFPb31aBDODgXxV2Aq1LMrDaPE12WQq
Oe7M5o+XavjQnzWRIUc2fQSXbEWmxe7DR0TOn1pndOGBTQtXgQhaT5IrFOGGuiYl
NhAfRewRcRpby3sboeT+VSgfS1NZFj19M2tEqnpIi6sTKjeVanpJI3JxwbFXX7Ek
IVvgNZmIt/kDPszePSY+RkhwIRVNlKhxTMEaUdQMJLe65OUbowOLMm0b9tm6/6V8
t5VgymXo27quMp7YoySRvq4Ozeh5Pdunc6K1s78BgrJeUHpS7c43q/S8bcihp8nH
RagEPVlIEmw9+he2AbCMMgjjk5R4AI7bhrmdU0Yhat2I41dpZMTnctBCJkRX78au
lr8KylTPl1nsH4/pMx/6t6KKU4unY9gjlJo8IC3MrqQqNIr4J7TC3X2C7HnNVDyS
VlNyoKTKyhPHzDymI0glZIIzcxBWnULnFzzkrX7GQaBxEfM7tE4XdiwsnMjPrGql
4z/8DYg668OGPZDYHvyqN6ASpmPZ8nQvSqzZq4+MuQJrIZi/5HWUd38RCkHDpCtr
9kuA6DYhIzWgK9caoo66KyNu4JZ4+TkCrBYeh2lsNaqkFus9VtzC5hAi2YExC1oh
7ouE2UQzKpxwNPI+rQbIaakTIQjGKiKkNE8jzqD166j2Rzy32kxllZq6KCP70fGm
airPOjYl3LU0hRlcyGhXO1bzkD2GV0NvXwby/wNAeHcgrekB1Ua16VJ0b3ZRNGfr
mjuPptspfUlr01TzgTv0TBmN/sLiXTD/LtKmQlKD9Oxz+OGq1VpQJl5EAB3h6xrm
MzEdSg3f06tNmYLIXrTiv4rWILI6otnENOpLKvm3BQlxlKSWbOmk0vXUQEVn4xfq
JDfdw0u7Yo8A+wLjm5V2MrFNg3586TnV4HpS/52H3mFgqRPvQ+7BgsXlhLBHzV70
bdgzqBSD1v/VoJ3BqyZFiquexySa10nNzJgrCvJ9dqLCygyOW43k4viV0JFYQQOr
IY4O3IlkIyhcIKkc009ALHRPkiGsAOf7jZ0PDhE1P4uJKDLE+fOPFF4uN2R7hh7s
vOKpFqy0kXFbA8YAs4tLkFwzung6NqSkN1zhp++bj9SJ3R8/vQDfrqAxXqrO/wHz
eabQzjmMBP+j3gbz/uzRcoy5RoDOv+8Z+Y0ScXwMfecLDzvFaQNywhDETDSjMnjN
s871I0mIlfdrtCUWlxjfZAzw8++NUxiy60MG4Kg9c6x5Yxv6UvRB0yLyUOl+Cklj
azVZxH0pVrbK23iBru6gJEMLOrktuCGcAouHh/vBZWY4fiNk72tX1G8/GtIbbhhs
8BkitVWWO9Jvq0rDQC3eBIcUdbriO1H0w4OlO4Z2G4USbLQCUfqtyvXZXW3aIamV
akB7tW0a3BcFACgKhDNQ9NfoJAoPD5xZC0y7ecf9sECtOY7CwJLv0gipSKcJARxL
IDo1oofsGCgT4oc/abgKCYO/doakRpmkOKdFF4Vu7oUlGDyCWwRWhOI1USvNuqKD
N1qIgGCUvrPuMx1WkDjgt4MO0rLo+CVdSksSKdCnrL09Yh3gl+zwnQmnMSiVD+8e
U2ItA+9tzgfcjuD3ENJwHo94ioHcyjNNTB/AEi6diu0aMYoV2252t++gwx3VEecX
xGQ5jB/97h3qErvYdATK3XYwGCkYH+Szmvw09+NJspKxCNK6gKD/1v3rYSLKmWzP
Yks4sI6KzRK6NTWGr6RKNwNCKq254N6zC3fm9uvDiYD3qTNOevGX8qxEvnl/uNca
f2dHUI/PROVpllULikDHpdqZ658g6oxxpRYW7si5M8yLQWD2lliszovWcTjJcLyd
sIzNpi1+esZz9slz8JZhUOCYkZ+Zy5pccHXpMwR5/cb80TXQt/6P1FZ+FWGyM+cx
HaAlA4Jn7CAvKpbt/3IiLpfWukc6445EioMkMPNs7wl0LelY5kxz376O8NxA4CJ1
djRl4PQqaNy62CiwdZ/7Q9Q9PDkvxEptNKD881CnxYj405iieaFceZXSUweI5FrX
/vZ8yksfw5op17Gfjqrh8Ir5YKNQYhPEvyjJ6258N9hfK+OXAA0idSo2K+iYGNJG
b34ABj2ze8ue/zCAaxuItBIWNNi5HX3rs1CIJFlF7mzPd/JNF7Q/YXPQ45Cfx3E9
ttktdozvzfX8JwqkI2lTNALQorkMltC7Fo3WMGVfw/1mqllsS6esGTQPF+hkaftX
bRYEg0JL+nO8fXIk77bTGnw+JlHyaDfQkXKrqn2vdtOajpEq6zv7Sg1VrJlzxJk7
HuLoxlYL6iLqFW2mh52qKp0W4dLrCPsJbd9rUAKWhQsD36Aq/6Fo690unTx/2LWw
CIF/wR+nYgtjeGCv7TrP5XEWAJIJDQFbiyBl9gaTI9Aj7a4cwhUwMiYv0utwnxK7
1sbhhojZ49IKTDxhQzi7xVZour9gDp91IAp3gOaXv+eeQumbjEI1NS6Dba/lZIS5
9vQfeYOujtKfOSosTP09qCa22PxpjokeqxXKT6yzcJb6FLr8enn68hRq4+UR3nXZ
8uojJA+lbaHbTKN5irLRbcGsU2svxuXcIpkJUY83gG7kQh+/LE1u3qP7ZMzZPbvt
ocCQG6Tu4s+P3/gHl0fPEBD2lcQoeYRd78lp5QeOe/Y8+gwXq7Iwn3MVsUIkpQZG
7bAmdfizgO9KNYU/3jVltloCAhVzuFlnrEKubY1hlsMjh6spiZflwDtZbx2JE967
ne64itrFy/ENqBd9zJk8HtUZ4+PA18AP58Yz0RkuihNSmc0VyjuQO8L541jXKylp
J5TSfNiOhuF2LZWW22/v8mwmNnzrDGFBmJgy8DBXuIRDCiwluGvnGL7sfJDaKMJe
XTsoPLD9mpdzMRzWn0O2q9PZKWxfDsrWUAbChOGbJ1UIjUNkh5Axll1HWXhbafO9
JtiP7g3Br9uQ+4VfXUC9mPVkq01gzFL50zVfI9WdkQ39cSpuW62xwUKU+hSDZKsY
EDkjGK6RLgF7AbFky1zGh2FGUAL8/uslqr3lw+jpvlWcFIQhk8eohBKyVYnyw+dO
7L3CevWvjDa+uWX1BRchuHrPF7iRSYLmaVwQ2eeD/MdhOBV341Tm/xeTLL/X5HHW
c7+V05fKKwIZJ4qTSEDgxSXb/k1aR5PHpp0kqVXcg8MX81RDbdHNznQytktTDNIQ
PYVOyXcjvUJFg58DRq6xgTypxaszUmUyOapMhnZGdLWCad1QlehzwT1avs/5LkES
J6XK5i1uWP4svC06TQxdLVnzaiNnyyd3xsg6NnsR0jgUKkpQYf1v+vasd0evw8/F
iKmxhgdfO/kJ+9HSSpCtFWaIGUV+kWKz01N8x2r1s/ou6gCVqKBS3qMHlrZ1gIZD
riVsTYB6FaPPdEE+RJYbyx81p+jdztOMzR8mUeaY3A6abGzeO/xKcz23wtsy0n8C
ivLRoc/25NwifwwjWeqM6jiYZYEE/F1irTNlfdJ8dGWeDPCHC2+xl0Qr8nzF+DHb
lcOySaeKbD+4+ZgLcVXCun1A3QtX8vzJMo+SIKfcukhkxP1BBP0x4R54zZFzinsF
cDXW4aP+WDSDE/ONviJhEuq4zVQ65h65MPW+1jDQhUzLz+mMuXxYVbHBJ4/RUBeq
p5AbNXoT+1qSEMO5T26xl2WLxItMOoL87ncQTIvGU98lVID7hYqbR67HGhg2tiFU
Y2cGEnwyKCEnad4eILRMRmamC9/YwearEc9qb7VPCBI1KZUirn9nPGQ3iDtZtXpP
qrtDn1QHAHx2WkCSSaPwqA==
`protect END_PROTECTED
