`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8eV9Uvm8L7uhuRKvo2f/mac/AJwx6GFsPpSM8cMpY1jDbC8VaPZDGtG2c/bHjAyb
a5Dw2sx/VQ8pCxbqY0gil6ewHpqLkNrwfxCjRJ7YeZb6ZYm5ek17PYVxoQyZRPZk
Zk+bv6KUDfHYZWW2gQIcDGMqa4H9zrDggHZRK65dcnipgVmEGtcRnTBkhxnGvibf
bCIwC9EG3N4eRqedg1DFstijPJ/i96anrxo/vsGBqRUUBP7njG6Csa7iBHU7se/Q
ZesXrE36XeFNpOl4p0nshoU8txYXBKiuw0IPDftNfE3JJROzuGS+LhxDYnYx8rr/
4N3UGT2IiyiBZdiCVIjNmRZXPRIA2gI2NY63GBOI2wUOeqh1pqQsJeGRY8FeQeoi
4I0FovBi+Q18Dxanth1DMbCsst7kQWNUCbgEQuZ72Q04aGLc8HRPz27rIEnAS4po
`protect END_PROTECTED
