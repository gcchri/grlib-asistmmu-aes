`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GVIci5rBGQbyeICNfllEKRxC+htyqis+qzdcj1SvrewgaRxANAxfYiDZDCSGWoEU
9OkYuPDMiMrHMabKXFZf7qN1P61VAXdqPwZAxc22qu68oocal+SzKM/ViOCXJirk
ok11GYmYtbGZc+K8slvefGoFzz0S0EzZgGIsC/zuFJ1YG1PPrxgCfo6ggp3YP7K4
i7KX1tCHekDMdb8S+nohYC9w2y4ivBrmxHvZOXFEjdqlbh9XcsYvYbO+MaDLMhl3
mjiC+hyEyUw7IJJn3TgVnD7mpmSW/3EWiLZuY57pxuGbtYhYRpFEieuddFMEkItz
1kJLRJ+XmMi5GuKF0oMmv1+dLoAzAr5R/fR0gp2zayxoRg3EPqo5KyE2B5lf8GP3
5DiUPA5U14XU4tDgI+mrrrtDw1kqf48C0++voq0l41T0oFzVWAevvZljSMVV0Ohg
t9Xnn+Dfv9VWIYt6RnBt46a3+JnDO193GDxcGmpJppsnpW2ioUmw1cvrAXiYfeJ2
/SNX0LvMS+m5t8OxKrD+IdH2DqYLoghcSTTUcfThFtZPVf5hepBIIJMNvGUv20Ee
0kFM9FcxoZsTjDhr6tobHA==
`protect END_PROTECTED
