`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vdq6c1qfszRCdLICJRpwyoEonEDMDOmikQBOpVPLey75dwu2S0XBg7lwdej2ji9/
CTUnhgt6JOq6AITmmYHm+t4qZc4rePN093BZJ1Od2VCQo482qX+B9vLaQbN4bQOy
NLbjBTcjFZCyRQanhVRqVqnD4Yz+nl/dODCrbHtxkiH+1+m5Dym8QJaBcSW8sOht
7mJVnrifiGs1TSzjLefRrmycGmhwFfXiI+LH3a/+mif9Uf45IW2UrW7PgmiFdarY
IIWvlRX5YRzBgUdTmgxK67bZXBdtDJI/del3HY2CfcoyEh/OQhbh8e699XphR6Vs
dugQWPN3M4Lu5CJ9e9PLDnJptUpWVMJzy2fJYdKnz1n2O4zUD86+3tLU2gSdVj2U
/IWvCl9wkBpcJ7SPWf9xqL610XYKn672PjquEgfYQ2T50kULRPuLQq8qReqKCyp0
xGEWvZro8IvrOBcAjebmHWwKZ0ytphCwG6p26CsxY0K7/YyQcW1g2JllPXkaYZ3j
cbOvGcHEtYlFVwe8mpvtDQ==
`protect END_PROTECTED
