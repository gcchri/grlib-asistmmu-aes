`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PfAB3XzCqDsZm43DpoxOOGRs4w6dbHrC+ZqoPPA25ppWGELA0maPAST81jYnilAs
S9dK6uLMf2iFi/N5PJGP6y/qPq7s0JN2eg5BdhAWC4XabXwSEGPdmmQ+PYEMjUyD
fQNhnF9xWokcBr5foFcbNecEqda4j2iFwkGNzzximr3QLMcboNnpEKo6EcVOaM5p
30/SwDmWg+SonHLpVRu7G/+WSVAeqez6Wu1js8eNAIoAo1ufSwiyui/bti/PbCz5
4MNvDS6+6Qa0RdbZf4Mz8cwzanOLfAyDwC0k0Z/4x/M=
`protect END_PROTECTED
