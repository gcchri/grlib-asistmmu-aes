`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dOFh0i22fXpA764fcRr57yAQzElEU+aPbipg0kcdIvw2EW/ToN3Wx6GEjZ9KpYGo
f8I6rBh3LQ91EnrIJnCnhTyNJ8IEOw2vQdtb9gtLhA/NDy5vMgTu3v+EQVZW/lzs
OfvBhGI70iL+tQ75RNDsiy3BJvR/faDcRa50Rv9DL+8yjapSlMMpvJScRt4GsMT7
rrDoxPtJSkyJwcLsEnQU7TJCb91NQJsKLveCy+sw6kOoGxogkxmal/wZAdJab/PJ
oyfuRML8WHlkfKavSUGp7DMMG2Brwu9HSJig6ga5DvFQtb8OlRSYVQtDXi8mwjoS
Alk/r1T1WrZCPPLw754edZy4UN8fhv7f1VaRo5fvfj51yKrx1jkYIlB9BUn1Xw+9
0EaYiUrO3cLWyy5sgcQx+9LHs30iILIaVw5O70ycZOw4HVMOnBr8lBBKEo2Fe9eF
YSsZt0hehkmXZdsVyBRvM0O7uQoopMygwHq9RyxeEvWs1cQOuMljtrIjwOj/unCX
oarW+qrs/+b4nE6gtqvdViBE5gRL8Dke8wpo7io2iZxegqspH9Wim/Z7EKCKWMB8
TZ1OY6nM5N+PmXbR1+ayPrv+XQc6l88c2IXmIE4NzAV1fApyPkr0HP03omFGRoPb
H6AT/rR/FxmXcBMtIrKTElhuoB66KlN5HCHkLMPadX1e+fVS4+O+IBCytrAKv292
j21lC822Fjjpwh/2ryUanQ==
`protect END_PROTECTED
