`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yknkt9YEggVIMt8mY7pb2iNtJV0ZpMpRBLUzIKPEaBrzCk9mGhCXV8GC3RoU3FJK
vmXUwqBPcFMA5sCFPJU9bBiaC4Nq3bkO9JLJyS07c18ptmBUMzPoZBVudWy7pfbf
o33qVAYFJ82KIQxvbnVZP3anHiYwPsd3D2TFPi7gyASCWQLUCgmKuZwzEjTLWSeb
rki4f+8KDDls97049y4ig8Vn/DELv9UsTFi4Up2GmHZcf5eqtT9A8Hd8o7yFvxgd
5OVI53qw0plvxbQA9m5AWe5rZt3ZSggcuBtsGzU4yab1+qX3Ebea/ixVhQ/G9Z+e
8zpLi/pw5GJmb+NJCu7FwrFmHf0h1pADPArVryuK9cdUQycIM/S1I4/3piaK59Nn
CFah068B9+LIPmLXnemc98SX1e29iBtFD4rwpb/Avmt8rAtaVmFkEreWwP4n/Xwa
kJzO8AkvDQsbNQ0nTt3o6S7hEiUjZume2r3GAm4gsvvwIdUpWlmUVhmFxwgJHMCq
`protect END_PROTECTED
