`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vy2Qtz+rAN28lmX3vnwVN4PRMdoft17q2qOm6DadKxc5kFeIUadhmvUJuun4Vsjh
7szQMeJlCMC9Haq7AI85ARid4LkyTpRAYxMEfJ4Op/LJGbngeEJ9gS75Qzfkznt5
24zBvAKLylo8SqivG7HjYY7lXb7IBqw5xVJaBMZYYY+jfKOtT/yJS30BEXNy1qUt
Xae8vlTSMEJLabyW4FEpMoVwD5DtOiAjjFXneJd05gfhfnWP3aXknUMuOH7y4iTG
Vk8BXuWqCXfIjIWOCYgFheF4V5e34MjbZRL8QoQeBs5uJMEoR5rrcteIfoJz94Fm
8RHq76HCqUb564svVG+pS2g3hFFm8/YbnJyMnuYTGIukBy/rsoujeWBWmAucbfvR
TGxVJ0yQFwFaya6Fnm6yXsqOYWSD1aRJ0fYyhGqmjPE=
`protect END_PROTECTED
