`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s+HO/per6YgOHbX+yl/c7WC1UGtL46vCelYSDR/oQV5osdQ5ZIjrkNofoHLqiFd2
iVSospGEpoZR26AfD1HzQq9+qPjR9gFAwHkEHz4jNT+zV42kAu/9OKxSdwLO/Im6
W79n/uCzP94IWMm8njIUONgtu3misB2qBo3/eedC0BIjiLGlz53Egr+pxG3wEi2K
HFbMJaWN/7IMsVCXyMF7IG8ka+VIy1dckFM08Mpjzt0rOuDSZ0WzuoKWyjb+6vC5
9rBDuZUviuFDpuM4OX7oIw0iPCszsC4Dtyf9qZpEQZ3Ch3p27UseF2LGcVYxq7O7
tQ+InupknXVq6cLQaAGG1k+rbIsNitd7DmJAMOblblFYKrVFyij/CF62iNRYhQDt
ET1rZUvhQ2hWIY2Fl4QuKRZvMkDyNu8OObRaQTgiK9mp2hSlsNXkaZBC/qXRAWpX
QUJePCgI/9OhGOpShjXf39VXyO8AyWai582mseU++YlBoc/WBTu3FSIXxuzoZCOq
EqlD48lzmNYFmDNdBIe0lL+bz0o/4IeauBm8SRnREBkHLs7RfzEkvBfNzSIOv0lF
fgcFufWrO1FnNHh0e2WvpE3qf/1daepNAsToSDjOMAKePCoqQmFwWMzv/PEyUDB/
+NFztye3TyerglMc5APdtvrSFtTlQbFFSYA5TsthvxXJqz5d3VaMTQX0UqOvgUPz
qiYiYMduj+EcPsi6qfS0w8PHj6PChSIrH8Ow/ijAUvHozHMU+fL6wdFlDvfffI0K
eaZWybzbT9AIKGJPDoBIxP/Z0k1Zk6GjlryTV0htQxoM6ApbHyivjidZTF7NcdEY
L7EJI7wtvchPSpwUxwG/43Qkz8qRZQj/UnUiRb3zUdcaHj9+VLpWoQFts97qRR9b
4yMHMKVAge4KueJc/42sIdcwXIAPRATDlMEUnSPFAeijuq08MQi1PcI/ZDbqxavO
zbtTOUWFR6Kp8dMLzhJIqynLkLrcMs14BL8t8wTywRxQ5wgBVqNJiSSDR6Vehuw/
P3B6DJCNov1QJKFh6lafB9xF37G8HQsE3lYeRQkSlAH+xGTv3+R89FfQn2saaAiO
xTuscp4GGSFAE999+DoaI9+DajlcMmKKbo3IMrEdRNIzhSodFHXFLBZmAG/giR/3
773Vj1MS0Qtwyla90VTHgz3zrM8m5dKW2nxNB4B05hyQ3zAH9SHzCb+7LZfcw7/k
YLD8OO1wb6S4wrFbjGOgkvFGSnjsy+KgQB7Ln1+U+Fo/XDth/hekHCc0YnYKMZFI
VYAeiHWRu5RwmDEUMCiSPI3irNd5N/9GgyAtgVKI7twK9m0SXuCGPYVmoAxlifZ/
5x6pA6Rj8oF/A3DW3aLQvumq4aGf0ryoq7gexk6yFy1Zsxs/R4n5ef6sbI+tsmeP
`protect END_PROTECTED
