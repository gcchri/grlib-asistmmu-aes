`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m02wIYSFbn0O6tmRvA4PFtEdR+bW3q8PWONMOe/TZ9UQ54T8VWx0SW/8k2t+S4RS
xujUu4Yl5aSC6bNzVdNc8kkL5bB+JLpiS182QQLKeO1uQTB/dNYv2Z9cpL8wCzk0
Pjg0/Im/VjdKbUS8i3KtlLLcEjwjLeKpE+1hKQj1GmWfFKoC+rUHywR2fvAiA+hh
dFYxku1ktbOmebdM3JC+87UwaITHlr4L/G/LxLOyQyXSCnruzqhcH/FOhTWplILF
1KZrZUhJ048wPOARc8jFOeqfSWNUMcQAnEVe5/4tVgpUAW6LHiCzyBX37JfQWwKo
dUFljbrv7Kdl7Dubkfhobd9MT9wi3R+3/qvmm3pseMpxODoKCTygVhY7sEO5x34N
ZPoWm5UwNv8dsl2U/uTduw==
`protect END_PROTECTED
