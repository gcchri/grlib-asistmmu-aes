`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rAiKGTPb68QSWVF8YMworeufu3Qw5xzc23gIbmTeYR7A2pPDXCvzXJdLkBZzY2cQ
VEABB09Lq+Gctc1H1sEIdIWAfrtidB4kBTQSaGoLayxo9AgU22zEsxTcP0meHCoO
duML7wtgR4LV5rOx60n/5+Vp6yF87VXVgu3L+URRYpGCb6DBoNC3EhVZIPbunB3c
RqQEA1022hkrH1PzASGTDhfJpEs8w/OKnwNa6QgHBrpRND6XpxbvyOiHL6km5TrD
C84ml+9B4wvPnghiqwoJhfBV4Wgcb/HsHjY4rUjtU4hYj14RjTeUIsl8AOF+Y7LK
RI4+/XQFfWq8+81ieBwYvA9P54IMLZoItyF80PqQi5EjjTdIO7yQdtuXS+pudj1o
9RaPnfo0JVjGRe9QekYnvAIFt+4AVJch5pPmAr+mDXV2RBug5F/fGgnlr2p3xEEa
`protect END_PROTECTED
