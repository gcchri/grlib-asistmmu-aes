`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CxBc87k7f/F2tiMuToN+cxtAON6xnPgViGXF5AhnH3oTCluh/fAeiOOudA8MX4Uw
0n1z8rnf07trFDaduuOA8Uy7QW3WSz1jb/6jK+hfJNP9Orfx13G2gquL/sbzZpUy
r0M6dYStg6VDorH79P/pWeSFoUiJg1hu1v7056H5NtW0Yxtteru4qh8x1r9JMcJM
pEPxoZXWu7RsZ7P+8rFMY/ELlBgBwt+tI0k3vR6KDPZ/lCzrTe+xh54tmCHJJtZN
gdtbI0A0XaeGanpA+CBqe2ZAbMx2chhbpsJuGuIXKGCebctEaxB1wi1g5f8Yt98T
G17xmIkXzsyAtr43YBNhFbj4Q8UA20HnY1zlR8ExRSylbCYq+VYNX9dR0mG7Mp1h
VwZgiv2mEPvp6t/Nj1NZA+vMU48yYy+2Z7PXn6+pSsQ=
`protect END_PROTECTED
