`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BI5XCLoe+sz1wmzBxcxnXsAXa9qMLhOb5Ad6WVPeOQqvDvJxvgL1kZmlERFl9YLo
tx21KjuHHPdtqNDsC8DmNJwHlYF/bu6E1hHQcUM5y2BngwYW+zmu7gLo70qGnxw/
pnPomqtesRbjUxlRuSBGaz3Xwe9DqyY2V85DPJoiCBJ9d0mHGrDlksIMaLkzHN96
D3cO3B9XorlX8qvKNua3cTIglYBkonrC1pkVtEilWkwNEGUQX/zn4IW2oZBIqjSH
F1RP0IFqq4dLQOm5JXtOVtwBmzHQJk0GRmIkCyei0pJPBu64GVO2f1dXPvdXIELf
RzUw07cUpP6VY3lVRzl/ACDDHvyp8qZl4mNCaHM/2dWnN2v1y59vjz+WazgZ7yBd
rwe5YwVz97DjHr9qugd3ES6rCAUPJeXK8kbKMSO7fpo7Q+tcLXkTqHgSiyUZK27H
aM6uHft2AkX6MHiNkMWv9BFcBxCFtYZ0edHo6ODuSBYbWaYwfzP0/hX2ZM42dMEN
4vmbkehqR/Zolq6yW8/wjf9BzxSmLHscI0xchA3cgFQjBJQrRC8Zh9HbQkVvWb4u
RxW8onIwMUu5Nfk+7w3CDswZjUVJuN1hhX7DyldMKkFqhOPpXMHD3C/wcdLGR6Pl
8FnfgQy9rMwxkj9YI9laf2jRBzhDZsCieUvElHB1IxZMnWUrfTR5YW72kaNlyZjY
JpMbuuHthCNVbqX8a5TmOEDMBI0YhRPWWjm5T6DIvZGaIJpkLgnZ8kjpFpPhQ8AW
DvZJOBbXLFYO8ll8JGHnPlPTPqj2gYysHOEm/o+pHMqL16EkwQ6LXXHVxD2RyXKQ
MTvKAzaZz3PgGY/qVNBUgQqJDrz4KYMt8eSDCU0F/BMpyRp5NCeJXybS3MQqKl1U
hgeL5y0NVN5m+kURcgIIIjF3AVZL9W+6rZO/f+9AB39OhnHdyIpK3Y5MUOYDfB2K
qGa9aUNx+2xETltRcnNDjt6I0htVAWyIJR28gAhKzbWC+xuLzYZzxJsShsNZ7Ch8
pdavwhCD9PSOY8EfGJKaqWv8LTjZeJezojMWVr4C85c=
`protect END_PROTECTED
