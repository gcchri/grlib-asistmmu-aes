`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MFJx6paxFkspX+HPGGDGOrcJMV9simB2ofs/j81pyGeXsowTS9Md/16+pOMz82Hu
DiOkyWNu3Tg4TxMG+KyCq3DMu0V4wCnpt/OilV4buu2TXC8d8qFRdRSm5sY6PrVw
uK0oDAORySlpHU5llvC2imNlsbDxKPC0fuIyGrC/NF8nu/Svs09hS4kBJ9hMhqHR
j3246Ow44M34n8XZUeZkf3H0Ehc3yA+lQmV4lo7W2dQbvAQbwWFwiqCBaZrWv9/F
VhPwrjqF5k7PQdAohA3LE/OyLnKTN++un4cULWmwaEyNMe2q0myDvfULCZ5OJ+vO
Y8QrRKzf3MCn8EaECN3+woIFeXiNRy4R/+MyA8xiF0t/6vL35UzAdHRVaI0svaxE
JHg3dT4Ah8COnRBqqmKeldOe3kNDn10l/iMBJo8l8OE=
`protect END_PROTECTED
