`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VfGrjKnKfU+k29tT6m9gvwdEsmOCW0MXYE0strXoIstaw7UJ/srtT+8O9vdVyS4F
8uijkYdon9LbgZK2VMySupJ6kw9EmnxlEULqapTl+YBL6tmqUnu42sWLoOdR2non
2QApdT/nA+M38uh304a9xbxXb2mJIZk/tT0uALqpOkX9+NVypJvNm9yy5YGpyHGP
xI4dyyJVmP06uvbepCpS+7YLGdPJ7q0BMWEuM2LD4pwyyrudf6InKYk5B9SR1Yr5
OAKnLEucVCRMtTzmbaQZim1VvDYLWoconH40UCca8/CD3cevihJw/ZCKGFLDjODT
PnuPU0IxlgLSTA8YWUj4XvnF4prZ3OVAQlSf14p6+eN7wz2w06quQ5SQRvpBoG05
Wpzy3eSCHesg4EHNeTSOfGQ02w45spribS5jMbh7KWdBCNlIgnDTaEC2MsPpq9bW
isE5zgDakg3QIel/vykogKWz7HuzN3U0vxNibbadDihjkQqcKk3eYo5fEel+0foL
UShBiZ+v+rYveFogD1p1/cwwhrPcCVgEqNMhjED1jCQpoNY1MevxmAyes/ay2jys
kwNpUq3dVKqIHdkMPD2zmemCxOOICuUwKAWRsvIcCa+70JL8olBAsbNksRzrgXVk
b2n5JddI4QQJBpOCkXZgDzcm54vbO0d6KOgsri9k+zmNS9NFJbQAqX/JSbsL+VvT
cgvwglznmo1TiXCjYhpMZ0b3QaBq607XwprrzAKc87U=
`protect END_PROTECTED
