`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FKTr/rdni665L6O6jtigWnCKL1/oWCF+mZV5GYE2HLBTMhqjBKhejUZGATvaLYUr
6Fa9WwMafLHqSpiJnJV1p0gHU1HAhbKm9AU2KdgiU5fUluRFg7MP9bpd8qy+vopY
2tUeW2iubgsEBnlmw0sRIud2aiPGSOy3B9IkIwp0pIEpId7KiXSaz90JDNWwHW6q
xgfkUZCs4hQuKEhuGIXoGkHtJs4M653cIiymu3O+yYM1htXGHBMAxVN4hPIg0BuS
rljxiHqLXpLyK37O0YNFDA==
`protect END_PROTECTED
