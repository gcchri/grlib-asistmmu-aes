`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
84ln+l+7aKU5jzHymcJIdgCZHTVcYhK8/fH4yt9yF9V8rLB7nUZkk3WBGSDRgFaw
GfVvPkPp4uoUgozIZDvzvZRz/XhsObUlzO6TJunNvqnHJLzMobRUTr7/VoctB4m/
fNP9mIBAQS+tZ3MwOpglqJFoMy48rAQClie2+gO8NlGLwag23t098LrMgkrOI98y
w0Rdd7ml9Ht9RKrwKoMDzfdvVFVBZ5HWirWMZANN25Drf0M1+sC5BryzO3eH7cRo
iYvXt9/HT9V5t9YEBBUxIfnzCGzv5TDl/CTyha2bDuybN/iepumWvSY/zo8Ihyxc
Y8ln/c+XaIArFo9ymqeNQKZmTQlTKdk8ZE4CMwl21DmuAabnL8yslEkeUlZKgF7j
pQOH2GfRnhqV+JkugHY+UufFXC4ffgAcLIdtRnCF1z+ZT4e1dWRffOW5/3STZ6U8
h77KB1KwiMKWpt1DI7USsioUBrhg3lqhn1oAd0nb4AmZ7ySgqmae/RYGZ3vUkOG2
ed9HGLTGTx3M2QyT6FzkXJ3chBUVk2IXnackARbB+4g3gvv7eG+QqtpP0wJ1n3HZ
zfUbq5iA4HlpZQJJIUHdqrz1e1DRWmkZy9yOUc3l7XYx1PsuXzWV1sQW8VIPmbAy
QLzNm6cCZq5hJKDupJvuvdA6ujKFpLsOkYO1gg8WxVgNZqLPrLsr9cj3w7ZSWZFV
H1fHQUCO+FwxZxiMQoK8OXpjz7gzNqe0qrp3Fq1RayXguRElriwUMFyWHpH1HFec
zUlb1sPHbufir6ia6xypIDMgHI7ts5lFVUUt9RRXNstbKNpQy8jaxGxwl++q45WD
5kD+unX5w6FZtsEASVuNqQ==
`protect END_PROTECTED
