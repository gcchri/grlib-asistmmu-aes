`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
luwj4oGUfcqs+FfThvCULlPUTqANZNr4V4FtfAfUc9tuuXK3c+tnrp6y6one58sb
7OflUTps8zPTfIy9BjeLzwv3o2hOXlyVlkk4Y7UJyywoyt9Tt6glyN5DPs7xN8oy
DBnybOfSadZEiIYNDo9ZMUSb+OisOVjiwxRNcc5icLpSJM8YNE75bdomqoGLW424
l6y079FeUt5FYtsIm8XsKewjanlofEodPZ8cOX7x6Nj/GkI+0I6KdPxc3scUnlc1
7FgaYcICCTaRDyVFmHeOhRxUEKg4EMA0nB1vI6G5svF/GlP3PHTXZQeoLKnarW3r
R014jFEj/EqVHfYa9EORjirsOAim2G86MLix8eoJ8hgGA42JM6V+QpDDgQo/rpDw
eqBfPoEgc5oMk5CPVH4ul87fdKsE2G5rxTAIwb6tv6hvN703hr3MqH5tZ0OjuXlp
Zspe41NL0Fk6lq5/bslVjOx6gQ1mXTNhS7aZEVAfqgALp12Ocxc0yA9Tyk0+jMyX
R6e6dE5M6NImu2g6LXGS/iOeOsRAAF24BKYBkDI5IDso0h+K5w/6DHRP4orMAJHn
QozYlrF/cqbcr6jSi6jcD0Qv3iBAg8fAGfemtEDK9vQEOXakfZmWpY+U4PD35UHT
`protect END_PROTECTED
