`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0agTZTc3n5Eup6uldU/WQwmaiT8JBpAuh6M52LKS6sx2FaAbJnxzbmB/ryXt9jOj
w0DUhLyaun3ePzMl0jQveJ7fMQZmS9O+Zj89d1qgffEuncMMVuRa4N7QlCjHENnA
/SDw8lGF3vX7Rv2E19wYddIWN70qQqu2o5XkoR8vN9XHxmieDI//UJ21MtbJeoLh
9ftM99bWFTSUgeu8vrbly3otIg6XfLxqsgv3QRrS3fNvZeGvmYT1l94bi+Oi8H39
wMyFoST17A/pO+DGQiUc/hGvQBnh+emc+ZhN2/TKyr/50867+fznE6f63BiUQTfT
6rJE+zgzFMSqtvmDog8C+bAvpkijFzVNKzLpGmK0cpm9h+Z1O6I6XMynGIDXCci/
U343cvwvc2AhD98qLTrVYZGQPXC/b9ncOdYC4giXCUhWCKs5Npvr19pq+4TxkSgP
EoJlYcgtz3XloVCRTikCG5EUW6AaXeriqr1x1a4ksFo=
`protect END_PROTECTED
