`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SUqr8xHVCxoqUaQctpW0ZP7SFCvVtGdN9AzRbkgp3kndW/xoDDPOhvnRsB7BqNNL
yVGzhXzZTxWFS2PQdZfrC16JERF6m1iC0Q57+ZKNf/P3/L5FFEUL4kyARdzt7KaF
YqoLRzLFGS8h2s8bEnPiHy32v3zOGgWHSLWqgUCymVIvb6xhAToBNhWO47jGNZ7G
xWeg9XmFye3A6QQ8MulhOKVKP4LyAwtgwQOmTetnNr+N6V+i/0rX8vBn0hyC/gx0
/owvlYbM3+00QcdeOXaYlDOPG3vOTOnrNnoIEdODmCwLEdMV5IorolMrAMb/7YCo
ORDX730Fe3LekjKX9n0KtPINd1tS23MBULXZbl6OQxVdQcOULzrLtSP3aFFJSN20
Sj75BzNDacQ5R4t0oOCCJGwH8knjJaSYZqD+OIjcCgPrWdLF0zuk92qsxQkWzAjE
6SuiiL0CA8tTfHmIgJP8CpnHFBQ/pEMo38VFruK9Rim9K6lcHTWP4bqcnqn3xDCA
ICyLQZzMYEtU/gU9kQybEY5tU4uuNRczx40sKLhINn4fmpXZkNnQrAyDJld0E7o7
YuFlr0BuIAlDSfZFycKiIi9ZtvqjeRHRhsZxMynceRrEhqAaKx6R5SFwSwrPD59P
TcYvae5lOyNw673U5O2wVehYEsr5BereXCQaM4RjPoURbFeSNam6FVsokYrqDyZu
93+I8nMnE2xDM0YxRLOJ1dlOOOYTGZLRSF4XBdn3aMQ01/9Xv1syAS8vmjsNCbcq
`protect END_PROTECTED
