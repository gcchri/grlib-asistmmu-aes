`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qRp8HLy4ELIq/TsHYtMPOGiDjK4pLSzw1QVeTY9bTZFli5Ql/MwmvYj2OvChNa3t
g5hMV0OO3GwRMknDd/9JJOacnYQr2W6tiZ4MpKpTK52ic4JuXc+6f07Dl/Z7/z+R
4dzsj47P51AXMTxYoDatDmzXMMnSwMjNLBzqAzvTd4Zehkbn0WnKso6CH5mVXCgI
apdCZVwiIwW0xSmc8HqRNAhylogJeYTdPFN6rbYZ4Fd4tT7bYx92Eo5rhwpbIpWc
m+mNiXYMVMvyj8rdn1A2QhEiEQBpDysGBgP4AfUWESpZu6269COd4OFRk/PHZxRr
vtPvI1UEJ//pwj9J0Shm6uV1Z3XkyLKyG/7aMTB/G7CT0/MBrqDm9IwWVxmY7/7n
3kfEERox9q5lSOK8xpRFJzY/hDMFOGvF4Xwpjlge4tLpWGSWA42Xsf8OsFSlYxq9
HHJTKOfNM7izTGzWAMwQRg==
`protect END_PROTECTED
