`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TNA0GigCfe2uYUvTRJi0sk5GjxfQREuacsslBu9YoPD+mLNzQHI6OZZ69tF24l3C
OykBmckkh6avrWPQ91UMl11SrA5juEsMuC52dktm2zJRid/ZHGIALlCqHoWHB63k
PNnYhOpkO/hb3Qbu9rPm1yJBEP7O8YqUpGD9+1/RdxsSOEC8//di1YdKPjvCjUvJ
Mm8ndLVC/Qf4ZIDNsuH7EM5fTYuhATeM2UqsE/F3tTRXvVjR1Y92DuunDwASSpi0
nEL5Rb9Pir1oMqWSPmGSG9NBG7Uo7APeiqPPVx0932wXVmiRj+OxfTs5XNIQfRHa
`protect END_PROTECTED
