`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SNgwavStcG/q8jFK/gG0tl7WUjRf5pqJS5Kh+ac2GB4ZXD114EIvNg+mUM9EfusG
l7D1uISqXoIwJww90Cax0KTHysmdG5MXKfZuz4N/Ms+1jSW4aUBkGGWHSN5kiRnT
Xj3hJVR6tKE1HZJ/qL77Gi/9ARV6gkUISFEo4t8nV064ShxJBkoiFYyoUA/cwE5N
K7rszqF9MarfYFdz6LSVmVk+eVDXlv594sh/KAwP3TszhPP/TVCrOS3iQ0x8zhaz
ZDQJ9Yyae9WrKHCmLayWZmFAm515CXDX5DZfuFozflAJBKNk1nv4lnPL4yNUMyCQ
+suuqGbsXM4ZL0k5WWG40Q==
`protect END_PROTECTED
