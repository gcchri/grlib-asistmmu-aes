`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pCVpv64sYl2S7/VDvfMwUxETSA2UoLQaVLFeS9La5N3RRcoUgwd6LXPLlGkRHP3Z
v2qHOh4oZnYzg+0cXMau5NWlGGvGKYjwEuxJGkUEVOcramRHyJb/NdQu3ZxMCd07
V20K4yl0pzb+7/A5Gmj1nMjVlwRKwcvcA/OHpHYNtqk6O+XWi0hAPeMUFMtEL2zj
u/LB2bKInipl55fZOlkLx/U7ma+GXsj/F/GEEtYCNrFFpyTMjVOljpYzP8J81I3k
+lZZAY4jGLFv/v9Tr/84CzpTiUIOtNQbb/4+lRg743dwEWCl1mTW2BcOXShdwi9a
9nRUJS7y6LPxUh1z/NqVcXCwfSdQc6NQfXMr7bqRj5pbpbPqVp5I+nVmBnQCA2L8
Nf3u/MeZ+1Yk7E0/4Opb+hLqXKSrco2RoQazeVbFSDrVuIsX1EkwNWvkiSWb00SH
M0ZwIT9ajox8L152WfEYjqW3hnx3IRV2v+XBehJHEFg4G9SfvEMHoY12fb3mCX/A
lseDjncrOrBZqUYl8NwikQZQLTUMsTWkibM1xs0kdrlKx/DpubEaluMahJib6iCa
MPFJsKwAURYujGUXvs7+6+FZ57M02dcbuKFmK0VPvkbRsXSBY8zQqGHvl3kxl9In
CyYd8jcIt6UWt3kj5XcIZA==
`protect END_PROTECTED
