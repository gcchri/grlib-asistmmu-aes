`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6I1Y64EecVONzTA94jQbauaN6QB/MvVy5uD4IQrUGYs86mhf21by3VlxUTVrdcnd
2ihaTP04F+5rTMYIOWA+LTmPD0iAx93BLFhIPJIVOpFs5mFfz1KNBgZyM0dcgUVY
ve9WYHWZnZn7uxW+u8rV2fyYPH/iv74XuZraxDj9moCHKBioFkIebsPE9yXuNRzs
PgKg2YH/FZqAJpwjXUyGAWIdC/uGd1oFv21I7EjintdskKeuLXbaE5OxgT/uBK6J
5qugjUez1oxpD6sgpBSjojmzisa4QYwBSdhMVVS8DdUMYhJnOoSnbUDDbUE+szre
X7oLZddsJan9/v+3fuf9JNHYQ/WLoBGwesE1SJXL+PCTPL2bNrPHpU/PNQcMefTh
XZvahiuiY00VQbvaQmIYXI3qJ0lCC8Nb6KYZPZQsZh4YJsjGBPRGmAKCKryIeu+N
N+/lePZhExXQeoJyIP0NAkeWIGB82yw6tA70KBsZjHg2s6Pwu+vWlfIDfPnwngHo
GcG9z056tt8qG2EXB4BhH0kgB65D92DgaKruk9EvMwo=
`protect END_PROTECTED
