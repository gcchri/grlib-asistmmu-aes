`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y4Z6w2jyutqjdIeFcKNuJP7o6N4/CvGs0+YUOivuAmm3rmkz6dR5IJxUDXUWQkfy
W+bO324JkEPDTYHPdTTzdjVZApM31FQ4yk4PES74q09co7F05DEcNx0jWB5TF1hz
YLk4iB8OgGtAd9+GEgZIuFFDybUlKKTdv7mEpbAVjq2GqGIVGYYOIa9fGybv5Lm1
y7+aTSRt231FcRclDbDhD3vY+yz67rsL/UNH9hUikhhLmLU3FFjYdaIUjdwwo+5B
YLoshYxR08038cJCL7PZ1p/LxME2/2/ByJJjNzfsPGRje5CnMFFMz/TuVR2v6dwm
Gf3MUibwSIqtQPtQKndiKngUvqVCPpBrI6QGfAz1A8ybiDXmuOIhpCfY1w9/jHM6
wYoXgIFO0JVKDqx2SuGtGlwAz1DZr7PmKgBWEcX/MCw=
`protect END_PROTECTED
