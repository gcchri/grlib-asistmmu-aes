`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mgBFvmH4d54sWGVpnMslZ7gcYPCTMur6Okz5zK+k9dHwTrjI0XdSoTM05Ti0WSl1
8uTEGbqGQeH4WqB6j3nDeqoWeCODbAucEp62g1X/OVGUhIy/mzeS7TghVgeYhRqD
UKo1og7iVtyTLeoSXJ6NMV01cP4Mlk8YjoF/xpshFNeAbQtin9Y3Q+sKBeejYCXv
Hd7VG7wqey4pJDBtjkz2JHUde+Xek9rlnb9yi8E1nCW4Pq4mOj5tKUxtIKdza+xe
5NcwcKIYyQCM2hMiWd63jwKDS43kbwIarsLcKIH7d0F3lV8nBdcT3FWP2m76kdMG
zNKnr+cBlPnih8y+KHYPKLBjVy6fGegwVTy1FgM9JGpwUaZ6Y38BiezyE19USrTQ
yAW0dnjpGG4LafPftxz7QIFRgUJIpkzkKOTBow1WxWVSZAaGZPhi/GyoFwc1IqqL
85VdtDw8K1gALEfUIrR/IGYBOhBhSpSQdrBoZHXKO2QasxlzFjBSqFVuw2mZPI8N
`protect END_PROTECTED
