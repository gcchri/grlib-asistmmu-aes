`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UC9GhXtgpfxCQG4BykK1aTqygEAGFt4RfuumKKQdmUoxQILvZ7SUFRtwUsn4peIA
ETh6VgmChYh8+CXe/2LUkt1RFgOtRAgusNNzi9BYB+sRgr9JlzYKfPx3GCpxVaQ3
09CJ4rGCT8Js39SYcElvAJ0vvh+fOg9ZlLrAtIxExjTGiJxvAk0+r8zovCJ+gAPQ
9VQVkzm83WxVSqb9WFlvOQ3x0Eo03vwvuJRyBouhcM5iqKTnMZffaYTNEvY3aK8T
9zA6bs5CuYSjzxxYRRHXdb+GMPkyK6BgSnvHPhkkveIHa88VmY4ry2f1qZIZxdSb
`protect END_PROTECTED
