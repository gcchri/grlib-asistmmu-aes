`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L6TLRO1JSPtit/PKk7+FI7EVHr8gbC7s8+jbhEG00EAmcSHlKZTZG/KUfqtNolqX
EzqZC8e2rEfvZfVP2q6hklSOIF7kYeqoFXLGfIbBlvU8NB1ssWZVtKhs0AOlHwSx
0UNBL7qcrpD7+xt7QnA1LkW+ryyukrafUIwi+q3rfqw4NFCZ4oKm++QP9Gl/rjfX
xBza91sXoUtqxPYS5ZerAMtdf9CcOB7rcXCEqFrGc/QqFLIKhz8a52ZyvBKUTbvh
4wIQ7k1Qep3Copj7JvSapbhiS5MKHnawtOBfH9j8qv7PfVw9T1Dg+Gok6aEuRqM8
BQjwl0UtOTWC64H4cF00OQ==
`protect END_PROTECTED
