`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Moyjn5WxAFa7F31FwkNX+XDMdZQ6kUYSZACrm6+AMepTxPSEcy1PqiEWWOCqmwwh
8X/iGLw7IN8ULjYZJahKMhoaejssMsT9bhWBWBTuHhfuG1UvyfM0NexSx/uZ+Xlv
E/nH6dC0P40AAcItiKFBKN1gN4ftw7THZc5nrWQ8MPADim9lUp5PouK3dYhT8P45
0Pkc3dag7e7y04c8B/EkcPYw3JiHlURTLS9umSwXzbb1XrXnKyLZWEIJ+FO3jvpw
Z/e49UOQlbs5YgT0lyYKcCEi0ZFNbS9U+fm4Ga3K8jmDgkUG9IGh4+ArjXQQQcbZ
YVglPjzAeZuhvSsROtcUdU8IWIgUL1O+4Zj5qL42RJ606I/QlnAdZFYuu3B7XaFF
Al7p9FiRLirGI0oH6VKlbpVGNbQjQyuMc3huH6fnn8Zk1eWUTxkBeYlMbByQFng+
0Z5Xa7c37wIulYDJRKcf4q5g3F9QPMYhFB9SSmumRBOZzQQiYUaHDbqg/6GjT1PE
4CR8bp4Xr6316/V1lSuc2cRmSBwz04gWKFDpoojm/A0UqDDkxGZdw1NRveLoIRC1
kes13+oGQPZASDMIIXxfTrbfK/AaW/+hjZlFcYuejc3avzAfffMiFBfYRsDMl//9
xwZbHXXq7iBIC7VkwenwznbRNqhrYlmULsatE+fLZPpg92zxp7qJLf7RFZAJPKyU
9sTiAq5yiGB+SV6u0HiL5S6bC9BZn+VNRJbe4zOQIN5DpeVuC7aP5E6dTnD10inX
hENOKAoS1XanPRhcpX02qrswo+8Vm4QmzXnfJSD2DCRfsJ0TbcYUp7mlsftMuAvA
SMTwoN0NvRxx4lOJwUwo3zxx4YeoEATdlcVdzN/XMottbxhwFWzQ2fG3P7mfRHTr
+UxtYPjK9G4OfJJZOOYxEM/9FlpPrQpUAhijzu09fmpL5lAnEUuBWp/3ekCtMVG8
+0Gio6Rfpp3DnRSEimUpJ2KwxKIvYXYKDlMNG5b3nITBOW0FxPP1X5uyEN9Yung7
333ItpYAQOdl07TGwBitstYSG1iKFIU9+aZdG3X4iGsb6LqTb8QCkp/G6LrjRUHN
78fiFqgBYRW9f+EDQBwZz/ubOMyR6oPtiTGuGFbQW0za1kLkKwKdSLFgHjZfRrMI
yqYCYXISgeuIKPeUAOAAV1/tmvqvmLHdKF0zaNpBAQB/kjWYnnlrG+LFYb3ob30u
4brW+ctu8HI4+5FtN/pWSRzWeS/6/dhWmKFAN4+OSYiA6YWddzGFfdAwac1ckq9s
6npRC/g/2HXitw7J3iFNXl1L+Ix5IPi8xPdrcK8bUR5d164RhZBYmvF0v/PYC9XA
UxScMWXDmjF1Azm2W9M1kEBkAElP80rOj4hdL8alC7zl25WpRbm9hkqap8WMfyFX
beqMGoQ7QaCUx8jl20/R6OEpGJ+RRj0obBHARdCds0F48uV7O6IEk8EtqQQ1k7kG
Y3Y5vCqBUPFIXWXUzJ3eDJ6xDqoeteuVRmQrQo3imoUYHbD/lJ+s7D4D8Dc9RxUx
VL8dE+LWDsopg+r9Sq7B+mBb/ZsnIGR01nIW1dvpIqIYhzRdJO8Spe5I1ig6ZSml
FYVPmShzS6N7oU7/DijvQ/08S/oe2shgoNAASXZkRmTOow2JpLFu99BTk4Wm4pCq
NO1eKI0w8Jp4/tOr9HNsbP0mWgQa6u1dnRdK+wCiAairWpqLIHg8URnZdJhZ6GwJ
W3cAQT9L4p+WPUNnXvRl9EnDAObVtnZ0j8dhBZnFZo0NquJeYrqVULY+MCtw4O/F
s3TDJkuotPllEjZHfvAZVK3FAffCHyAi0gBdwsgCa+tbeSTyAwAUoBZ15yTdvBs0
9LWm1RoIa8OtrnR5eNEyA2KAgrO8k20eV+FaQhGq0QDPOrHV23nYxHjFHbm7UjCh
FYzgEMjWcnVH1X6T1ZG2ddX6+voQS/+6hmFEYwA7iTDR0s9Tkrn5FsKr3xUuPoDc
U6II/ZB7vjkvS5/3umEzluAS6VlOB3nfnFubuSmhWgX3DX6CcsyaaIjK9RjYGOTM
7eLl4CGHSnbQobLYzb5lzXtMrEswWEvXLKzVk2lANnp/L6nlNk3sirXy1R0njuA/
p59/01Ahcx0Bx7L0c1xu7AbRPBOrxYdM7bd06as/S6KOnDYQcMQRzcCzrHvBGA8x
tB98J1Q0VOcEZajIuR3NPYDix2dCsVTtoktsG0JHYyystFw6jRQd9hqzLnHdpUb8
SoQQq8gTv66J90/LBjMaIlJsjbyYaS8FUq/NFq87lGParf6U7OtlydeIMYdUPZzA
7OvoZvrb+Ze4uo6e+qWIsvYTqieBM2A5SM7OeXRD0LKjdTXgtkIbJaJPKk1YVuRO
9NyytELBiriEroZEX31d3mi9/XZsfJRmK0qHRK8WcZr7FwkoP2I4FtqwyNamPe2i
7bHIVaZIH7R7RL76uSNTFks121RjoHuQ0NN5cdcQEEOxemBXp2/Vk/jo4XpPlmAo
7bl9EP0maOhStdGIyDCTnNDcTuBj7w+PVYtEqqK+vfLju/bDHjbUJNvxr8sVRn0m
EawX+VBI1MSfP9Rbm20Fuscx36eqhCpFj7cTGsM/4tRKhBwENMja+wHmyRWaXWL3
JbeNRYTFDjRXOlM24Psnh85GvD5fsCz7G2uflXHV/+d/8E612BmX3bbpKz/2BdxD
Vtqe2WQzn5cvhiE9XdENUIvJTAvaN4045nA6Aav2v5hJs7A4XNZxgrmhdSwLT5C7
j1qNZStvjkDC6I0R0xM2suAYLpua+pxdDRpZ98Jov6FPWewQau2tqPaTg5ttAzf3
DokUFcKGF4Rx7ysHxS2drp1JLqtlKlzYBOoCvsmW0laU3HQ3TjneTRK6MY9MQrl7
0zBGDm6No3rtgKb1YYpVDfBMuOdg2yTixbjJeqXW2waOTEpbA6Q0PG9vwK8t3EBQ
XwHukVk1fkV/QCsBtV0b/6GvR4PpgeJvwTUOqD+I4HBeqdlk4EA+DxELmPwa/dQr
RU37P33rrpN2nmz2ot0Va7GdWwrbuWbxzjrcwavjiFn+UdeUIz8yXjVNW3VJZoiC
1eszmVkKMv8L0Uwd+f9MOc9+klerpUjU9TBHpsArlbGcySmnWLw0ZE76luajADHO
gHb49XgPnLjSc3HfjcWl3DRwfL4K67CgxtfzsdneYktXMJAL1pxtBhbzTKcX7BwJ
JoXUr+w6JRdL7XJ79DmR0FbivkCf8Bpc7Gj/2hI3bkuS7d+ej/lfaqE37L/WjQOk
SJk60nmijZmEHzJXX6OIywYvXuH6LyV0P7o+10MN6O6alk0DWZaxUG9vEucHy4op
L5YJBXIW219wX9ShiiRGTLG/UfJkhnLn2RJj1f75qYY7+WOXGzj+wQj94AJLgbc5
IoFzBMAGJKuuTilBzFPuUXZrrN4I+WlA4cmbCjYybUfyjwTXrVzAcFnCnj6M4ksi
c/DEUn37htDRFhCXkdAQINtBNCRjNnBk0xrxnlxZE1yohTmPutlFAwQWpukYxLWk
d8MatqFoeb+hWTRBAmkp2YPhkk3HgUrCf7HBMRQq7T8D9AYknCFjRiPx02IUTXRp
TszIap0hBrvB/GuC0fDkR7OxG0Pni26vD9W8gBswnyZ3TALKdmnP2rIplicDcOTf
M5U/LCqx0ziwpSHmfR42mYMqdnjtUfEGRWB59aXGDEgjMHNky4d9Qlk1eytvmZdv
9A0YIQClhLymsontNPFmVyalHaBI9lMxxrfRrt1JAPla6iriBbtc6baVtnxyBHni
NQhgKOhFG936U4/HCzLGTJLZxv0MyMaIb4nKrdphwZLUDzKYTyt8EdKkaOZTKMUN
pq2h5kvpvm+hWFjNpEUQfqpxO2lVnxH5wXhHVHCWJejo44BKdokeaxJi4kjUWGEL
a3S1rdhBwXUzspMc2SoAY95J/xM4MqfE1hnIc1fpNTWJd0tN1S7LEGd5K75vu5rq
n1oXjdKl1aWfLvk1yACeZ/JYlCnD7HAIITjRCQx14ryBbVFRg22iOnYcij8Q7enl
F4zoj6vNAllm9DgIz4fciR2HXnSRxFOXN0funQWu+Q/EK+ebQ79F606NHJ80PEdA
H5Wg13mhPCDaPDH2K6mJLR07RMA/IN/UNcX667TNggGpv6zXkDHyDNNi1nMIGrGb
3Ys1aFrDzrAWw03ARDJU9z6KaK+tBWl81YOves9ktyBAZj6M0FFSPwX+LvHgB4Hj
6WB9Kj2tBoFWHSnmrfBTigldTe5KJU0UGsn8Vq/gGoUqVvMAzHEcao58qIuUHb7z
GCAZYci4Rh+XLGBLB6mF+V54SougoKxjYKS4B50IfROyylsT/4gfLLKLicxq6THb
Zx1fCIRsu7R/qKtwyAfYoSuk9BFrE+3WDEw5tODomd5X9u6tlJNo6UJtiQEqwa9R
/AZokvRDe1H8gZYkBEz2ZrZajcdyM+HwmFHVyzfdmc7/P1v7AAhSfozebnijNnOq
8BFkQztXOG7cHZ8bbVG9vKgVOTI+3VT8NWiAhzeIVFyWKqi4ad9BY9WBV+oJGxqH
P9abjujp9S8JH5KdXWfn9gaclYsq/xJgmj/DZTnKigqvfNQrBJy7VoFC2dShbPk9
PUOMf7aSwaLD14gP1H9u+FaA0ISK+T1pYMmlNue5W5a7z19mD/pgwnpL3isx9fmZ
a247vss1P0+fLavuxgvkIUoK/1l4sXqdx0G88fmifKeabQj699l81otPxwdKxZkk
kFZJr0L9Yj14Sr6YZ0u+8Q==
`protect END_PROTECTED
