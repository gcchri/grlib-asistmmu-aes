`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fqPpA3BIVftQTwlFpxcMf81vQNcYql/zpxxbzlgELcgVu4eSNbcf/oWZCxxTNQiA
8a16B5b9XSS74B5hcoQMKJTeyBVJ1GrxRp2WUjJeD8i9FyfEoG6Dud6ay8/itp/+
DiyfvgNaXDS6cahp8E4/WL8DhOe5VpCOE96JCcGPKYg4vtTq9tn53pWz8RY/BIcE
UpGKZjfG8q76QCn+VIGsMsJungmsH0i/VcVlNmc8YEWkRk/LfsoJMWq3sioqDBpd
Em0+ZzaMpBUHugbJQdk+xtbGlDYGR82nRPmludVLAhNgqNZsXiAjc5q4OnQOJn2m
3YKKKphzSiIjOIJZ7nDpnNl/li71IS4Y5ZQjbJeJwJjxvf2i3UL9dFdvHOV5DoSA
bts+8F5cY/GMLpQefYQCNA==
`protect END_PROTECTED
