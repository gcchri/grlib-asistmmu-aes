`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OTvCXT9ByH1+ZU+/2gwc80zLf8HBXfd9ZP70trGiqaILeVFPUHot90grPFOdsNmX
M4GZ0sXCEbwZx+TCtfkFgqzU3YpboGceuAKCXBZFVsWi5UUD1YlZaiLCRaTw6weD
XAhrNpeD5eNhlOHpFZgzdfaYjVfUME/rmamGYyJfF8mex4VtWAenZft93i9Bw3FZ
tvBM4uaQIPiAUaBxU5CtQUqohT9IsmhpiJccjnZeZEL3uWj0UiHAsRSr0JMkQITh
GXLh2/5pJm9yHx3zHapwVdeW21Mf/BShWYr+3DzkAtYOSrCLHwJwDvjsFiix92rp
xrRxY5d6yY0hclZpN3kXzi4/xcmfR/4jnLX1mqTAD4HecldlPuk7gxLR+7hCoFZ8
ndHK71pc20rrBGKFhxOelwKBFm0d5gnUbbZTbOfeCo4gYadP6y5ntJqMGe+4XANU
DpL2l+c6ZChmKn3d0FrUhYJThIkkG+LFzjM8Rfe829Y=
`protect END_PROTECTED
