`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M8xaH3kiIOXdEEzUffXb1+H16SaCFyIswUp4uvYoR7CTICpcJyr0SynuqzH9joVD
owInqKHCA7A+F/sW8sW2wWqmAgs3JISsLtr1YSf7g7JLDH/pezrAAftgF3ml1ljD
IjviSVb0aX48w2c/THyKBuQOoEWqRqYhsa+40H/SM9gf5v1DpVxbWOTBOEsRVGdz
9fPIsqLZV0ud9ysrnCgXhoRWoIvJPB1Z+jo7GfOyn8kB2P8Q3O6ViMFhr/wF/d5w
NRwg6Emwf/pieLWKcM83wVlgpqfaYW/fSfQeUVw2+8RhN056pmHGJ/G+wptBbMG3
3hG2NuEY5O/rczgRzI3CC9yAoa6BH03TDE5YMHMjpHI220I7t/hLtkYKKyZFZNl8
aNKGxm/oynOdbsCWKWGcBa70GXSD9uV3Yzymq7kUguWqOYiV5gCbvzcsjBQ5bQBU
8fbDgC9oiaJQKOcAi+qmQnu4HbxnkdMVCFbd/Lepd2YRXMEHXWIYAm1nIIm6cU+8
nReFTG7lds+Fuhr4sP8hpMUeMCr2xwkS1AnuFnZ1Ts/oF9+ihL82IJp/ARcRglSi
5zbNSUW10KGtmp5Xnbc7aiv7LKCuHvRh3DYoKgpamOUDQo4IQcXm/YH7z1+s3JSS
KzXBEhq1MrvR9919Wr+8kguykBOPlC2cGWEgFyZ+ZkUifdzucrGjM0e5w0ZVYvYw
UrJ6++WWA1NX98OZnnOZzcl5HmMavfM54+EI/8B3jBuykBYlZzcjENx3PbcNlQBR
ndVazneIDihKazGjn0dgnVVN/RMBssnVkKVMpXdz93rsDO89JvETOqJLY6DFuU/S
Oss1MLgRmTRXb3hGiRp64g7nuw0/NEjXZbhynGaNGm24uE+J5dmb5Ij0l4LdKFlo
+4rVWQWLVw6T6gaSyPbeZJ1VNhQ4VHOIynssz8f+tvtT5vSNS4tE9r3JTZFwJB07
QiJ1oieMMQVv6luatPd2mZ5Yqxm5PD3bMkis8fxZUSYyOXW37ITYa97dTENqwxsY
y/vcn/qbCwZsqIQKxdVB6+YsHEeXAU9FYcl1ASCjfgE4NMzeUNGOkvnw6wTohfJ7
LAR5rXTV3tTxjf9cs2b7kBLAtHRUyDQ8aj+s+MBPwQ0YE7HMArrGB8WeDt4xUbba
p1bWABwX2VJy3/SsfRTHoFPrbRG1/5mzByHKsFWoE5XQkWPKeBNy9KHHBqnnkX/M
9TUTInPxfM9+lzsD3HASUe1jcO+zy9rRUe833b05dUBYL5yg5Kt64sWySHfZGG7G
EUWckU4TeexzzzPkY5nyUqGUQeMYLn2Dap/5s98h820H74ln1YhlfUBh9ErJUwhB
MEM6lWM4yCOiCLF+5tvfKCCQ0tBknwddzykrp8Gw+1ZGEnMYVHx/60QElmHYNXUs
9i2ApubFZWrZ3xJj3tffyPGhQPEQ3/wNTviBoA7arQFXHyH3tqRTPJic6CzCtOu+
Qpft4dsMgyxMzFQ3Bf0zoqAYNc4XhqFF+sswAkWCYGwes/I4FzKaPA83CA/VMJVQ
racouhmRzZLCnZTut8O+2VQb8oVTaPdjrYa7+tjeTHS5l9E+suRPm+GBwIuaVO8k
zsePcXxM5PIcQhh0kM2jAq60UTQUEAx7T7P9eG995xyLGSiehZJStQ0dq/+PiiEX
`protect END_PROTECTED
