`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nDz0edncOfWX9n+PWqyp7kPtbwAwvW6BKulUD7gpWAJmkDhq7ZN4fnXX378eCEZ8
1dZEUyTmCC/2gAr8uB9Fp82aNYNT78j2LmuxE+xaXTYfIeQxcTyt79NYlMaDr1KN
gAaaYNfQYHUWwViCUFgWSY4ldOBiQjsd6Tdt3hhb0vwxOEf9+iOAifj+oZfaAQto
atfBSeBCuD/ylk+X5WXlkUUEUju3wblAN+etuk2TlCcWUTDaVdbaxtw85MMPZw9L
Oaks9NvMc10RVbTNM0nTo6vwGVCi54krMtg2kdLz6WeKyMOQ6EhVGEuxPWxPDv+v
qvRDIejS22DtMqryPgGSS/YFCbOb/84qCZjgo1WFE00EMFMt0Tv2RSAwaKUjb/Vq
7mQ4/3EnMYDzYtbiEokNZSsU+04W+ljAJ5zdN9fvVDlBbQ44klxqEkoq2KJAhvKD
S0KSLxdeOj6t+Rdfqt/UQY7q/tZWmn1pxp1ZGnQZ+dYzpPK0FAjPak5+/uA6EKIo
asHYVg0pcHdEjqlxVbbsj3eer3g1U/T9Oh9/tLJJjIo=
`protect END_PROTECTED
