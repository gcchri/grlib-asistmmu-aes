`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RGCqIDSssQ04MPXy53B4F8ALHJSzQ0LIHJ74/RI29WnctzsVotfAU0luonFjUJGv
dhwphkjrwoAV3/Aq0C8KLR8WAQXqIqFtxeTwJW3005PQ3HzWxQCDruEs7IL7ZAqu
BBFUjKEdqM7dZw7k84JPQfSZCJmU6w/yq2yYjv/Cj/bKVb9ZckdEjNYzRr3NqEMz
3lXyVSZux7peBLtziNYxC9Tjor3j5cWsYBtAJXmE1dgek4HxvF3kf0Ub/9HhPe27
0xDJhKP9ZPgZC83OK3dY7BDmK7BHJYgswsLgBxWcTCXMEfHS+oFg/uXFXstr1L56
uX/MavmppaJ8eJY1Z3a1+baiwsAyx+QQnSYBRX6EP3teTpk3R4rX7wzPO9NyLnOM
fH9LqJLhxL91N8wiGI0trYDJsaHEXge1fIOc4QcFPNgRGXGvkcf9qdNa8DyP3wwK
C1iWxB+elP2rz569E0/no/lEejjLGxTvCN04H8LVnBE=
`protect END_PROTECTED
