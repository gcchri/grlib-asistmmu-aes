`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yLAfmAUwI7OUrLn9chhaHDaslM1dqkdUuocIocJI70T5N7hG7I0CfLh4D983NxMK
7hbjx8kOHXH9l2pSQ4xIIFJHP+VaQDd9JHyKcYWG0B68awP7I6KuCve8fS+Dt/WB
S6Svb1xFUHrPsnc4k9OJZRBQC1CdeG7GQrKd70g+3gfeX96nV9r6Sj/aPPrN67BX
zYbKkGKLCtnU+9D/R+YuYkBaEbN3bU8HR2OVam42kfGmu8ZLCwixSgUDhJrg0y58
Ai4NnL46fcPmAYXxZT5qOdNTZ1EClJ9gj1rJO5wfCYYT9lF7kmndiptIMRWiT8ah
coBO9m/F7uFXe6VC/+fAbJiD4YH5rltEn/QD7d3V6WRYfk+kL9D7umE0XhUyE0Kd
I50RocJfrup/oTtU5X8ksVKnH/ukA9LeuSOGQrUOzq65tnP9h+Us9lGdSCf2NWzK
lW47ZPieRgt/sCz4+HW4RqlUBW9iw+ce5UMnfrEl9lHhhwR54UJvMNk9xwNFttCh
eWDtxNiwQGEYbb0zgqu7Q6k+6j7lbIl2ohBwh3kanldB2fU9WvAxv0cYyodNB8wi
Zwjo4VV8nn12hV38T+YF+Q==
`protect END_PROTECTED
