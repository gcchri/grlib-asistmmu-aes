`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F0h8w67bF7RgBqcz/uSa3YMBt8TJ2inXPJOAOAV3aWDEMrWLYtHoJuQS80BjL7xS
FUEyPwQEnd5d7C2/ZhZEG3m3fHv5EL51ldy48xEMH4+QOg2lg0OuVnfo2OJBS+P+
152D9CM69hXOW26RXol0FKf+X7r1iFpFA/nVXvvxhcoVC1fZz+SO13gZltYLUW42
3IpTBbhK2qYNzpJMNxMtlec2Pj/nPkPaAk89b3s5QRs45ck8l23/4X9/XT+r7Fe1
+DfZB+GnQvoZUicOzu6NS6VdJBZQtchEFpvqbFvXnFSuSyLdGXVEq7jO5EeUv04p
iWr35Bd3kdsHkJi2AOowcs3t56ry9rPGWBQ7C3jTiq2xwTywuzcBHqkEUjo/YV/n
z7qX1ruRoOOHcjzwGQbPLhnDugHj2inx0nVjBCbqaCd8NGt2qpv/PkJLbVrEEEsP
0tI3Mcur1yb/Wld3xELm7lDCaJqehdu+qKpJRc7T5vvd4DPcSozYBumEywoU/ORv
hTQ0y5MoCr8F/8/KPeKISa6sHzcYfYLdOwKtEG59aeg0uo6ejAfvh4RylY+cScdY
VAibG8fowf6M12ilFF9vVQaBjyrfF2pGqxyauHmVd7w=
`protect END_PROTECTED
