`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OF2oH8egAJewrxVaxiZ5CuwBqTwAVyxip1vOUXt5r+OBi2GOBpCSZdwsy06CH5VD
yiL8BCAJb3+MGXKV2BeZbfyO0ms9q+xI8JNKPXKBd9igYQ+dTXcr8VwTk5qd1FWq
LCQN+nBcyBaKg7xPL6Crml7BSyHSiUyX/dYBWvvd6/x1vuNF8jz13BfyGDjlR3p1
yvpa/TOzLIN0erc8bYyyYfzQwjygCBoirfBMvWejssHqDoomFZw0smAkl7hj75wh
n3OEp9/N1DeyZPoOoNVM5+IcGdCFYI8c9eMlahVT39j4erMepzkJeGGLSFTYBOAR
KgOeWojfeB266tqBEM+ihKJoXAc/uA/OnwMLLy8un4AVhlnuJA8JNwFZxfzfqj+R
EeU+mfnz+ggKSNfo0k0dYmPuuGMGR+ZcP+UvN2ou7ogk+26bZPdw9Or0JvSg/Zp/
aJF1DW9yi9r22TU/cpsGilMeiiL4R3haVqQXTZmca65vCX++IJ/jYVf692FSP3ol
+yebfW/bO0UOqiKBibEBh9WFfjeqfAtz7HEnvukhih1UlFnUY1tm943I0vXWJ/gX
I57JoG5gW4JoNlFB3+uPxGU4IqLEzZzm6tJGfZme4qLt2QJJNjcRLwM2vXxg8CdV
509hNPhuKdkTly2164A2VQ==
`protect END_PROTECTED
