`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EY1JtfaKUmbAug1OWmZSy/N1rE95IBEm0stwiC6PJblzaXjvYqGtdLNaaCxFbCwb
Mmw2QIz7xLv3zthqZ4vxr1Ys4YFBpsusCtyWeyrEdVaXJm6R9qn26k0EVLLF/crq
0SKIEIOdQ/YjB0IenJ+3+WSckN52/Z27tmlIopSsTWFo7bMREbVTSTlVrCxAcUeO
w6Az9SIYAHGBbhE0NPA6EtFYWhubMKZHM/01lY6BYY+PkU1EAi5KYCBmd7zCl0v2
Wrg5xOqULMbAa2oxTE8gOmN50u9Cq7j6bdi2dvWEc0Ip/Hb53wmnYjK3+TtLdsNc
ttxShl2u9BQEL0Op2E+TesignB3qpf0KTPhVLSp6SpkIB3ifNg3/yegRvQtbQ1gg
`protect END_PROTECTED
