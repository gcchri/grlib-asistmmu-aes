`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0dkQh3qkW/u3EBu5L1KvyNVqOQGJVr8YQD88hwQcTKcuoZGu/w5oYRvxyeUdFu3V
zQWzPl05FFEV2Tem1cslTaDDWPrri8a/f84pgIaSqhk/mL/T6NLLjuvUiWxFoes9
s/rEQTZH/66vgDxG8lAHEpUm5VoCIqoQZ3mLhIWh24XhebcVV1otcb/yzTa8XXuJ
tZeUbhYeUW5nQCgU0zDKthbMvx1FfJv2ktBxGHwH/6sJAUGCvCHcrb45vr/GORHI
IIstaFApCutYZ8NWMf9i5LHQbtLwA+p8CV29p7kuFl14dNFDxGQIa9BLCb7U09Vq
Th0YKejWs2WXX1KST1DikcKy09aDrEHLGwLblOPzcRLzfRsQghI225fOi1kv5Xy/
JGssEcmwIdGS5+Xy2IeN1eOaZ67+BSHKTk6HUrtP2bdSU0caEMHfmZCbCVmBzNgP
FwT7IlJ0qq096NOFDTBk748P7GMoCnBatlCklAKcpxjO+REdagJJGP3EQ+r8ARYp
s9EvaQ1KnXZ2bgxxQUH/+GfvhLkUZfc28ARu6vtSBCRBipborJEQEqVLLhNLbW86
Z1ng2fbTE3OiqmOXi2QJ+nZLcAJitEkliczuD+k7PfWJlFWGWVSJ+e8hKLCe0KWD
kSRGPWInMIGiBZWOqRXQ+o828fphlUcqcukJrfkHWUqBLiEy2/KsOe03ONjjBZfq
d482O1JjrMak4G0HfOP4qYvQF676/BBY0j5/KEN6BxVmXN4/4CPhSkr6DDG2TPx/
kmTvmbcnCEpHX2rLjIHh/V7Forl8mo1a7flCrhh6NGogYcdpGfwrse7sQnEOEGoy
Z3yoscVctyBNnz/Mm7L1r93KOmqlitAeCxLXHxsf6cietRVXcUz/UbHYTUJMEtlU
wlprQ3E/bdUmcmVR0oaZlDBPXqspAcCH6KKMPcnvdEGfvgMuHEucY8sJqoC9pvh5
IzoR4wpby7FGoxdgR7LaNzWYHva6xQvj25C0lfbDWCxRBDabJ5k5Xv2Mf1XWdY1P
41WSXR7RiPZzg+YytpyqzqYhIMYcCnh4oCbFB4vDCqBecsl6ee6MOFRR9A8+0J3x
KI6J6jysb/0Pef0Lc7YDFxQlLPwodmDTCoXufWEs9hH55yF3nQsB/jvbPni8Z/jn
poLewBKl3IXb4rvR9gOlJfxVPFjrhBo6K5434ivQb2/LK/p9CmNBAVz6IqO8bRjK
vZhIaOp0+Mr0pb9jOCB0Cr/NYgplJYtbuS87UPvB+PgMNKQeImCzYCXYgInvdizC
UJFznYPyb5YxWw2jfOGW8QDH8189F/0ZVjgHuixwlRD9+FiVqnQnh41lZhg9sGBX
7X6FZ0W2ha8WzKSv0TEiWDsWoKWGuykqA5gAZ+hSz4E=
`protect END_PROTECTED
