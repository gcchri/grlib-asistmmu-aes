`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RLADd4EsMiKNp4PNl74iQ4mcPQ6Jt5bK1WJGpgz6qaS/DToNLOa0jt2xPyDcSakH
kP6mV7bxbaU/iPzkHG+v9ulFhxZGHNhVBG8qWxC34oS/Pt7bOkRzvN2H+EZGbf2/
5Achuq1Z8M1ZVoYS368Tqvpurl819NsVauTOgbZ/niJEzcFQORO+42nCNns8mmWw
2cuKXnjw3mwA9iLPXd7RgrXtm8R2t4OllLR0kaBxLA10XeOcD1/CNbLX0PFsIhVp
RClAPGCN64dmsYly2OLrMjDYlpSUn0r82dlU0jT7GmmWw6A6QCfWkNiDeS9c9G/D
TF3xDvr21hKZ/k9yOAe9NIpht+CX1XgNrprtaX92+QTfdCTljxNvrm0/vmHpqvjf
ou+ZDaMSy4qNKhu02rLRWQ==
`protect END_PROTECTED
