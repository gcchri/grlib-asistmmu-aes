`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
idWvohRgmk4aMo+gYQ29mU0wpFkCrHUxRoJwj4UVYrqjvp+76XLLXpUsB2JE71g0
DxfXZasvKPoOPEF+FDFRsTSPIt+0W8KbSGNPCDoBn7bZBUgVKT5dYsBjBbqyS08s
9hMOOsUdnvaoQGRiGVrDnwoK6cug92Mx7JtNYq8doqLdpZq7nIjb9KQhQg9gf8CA
yFrOIR6IA31NrrvZpXBwXVUGlA0oCrSdQ3qHZFWxki2zw3ysIZebir+vJ2Z0akrw
w8G1gFQ7DOiJ3u4AwRmzstF1udPBcoJjCXHLzZzjGwo=
`protect END_PROTECTED
