`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rWLDu9B0YZc0VCxbN2DRA3k0Jfx6IcIkSW/s7PCPyHm4n/Cad5ogmqcU2Be0TUgW
i8oWOC87I8bPC6gIJ+tS/G+Qf9Wzr9BgdZ9QUwrQnxLScFrH9JS+aI5DYmgHl/i3
QBUgxipvEHT80f7cWCtZKaJfH2+joNv41k0GWvOTZRIxfmbsuefL3xPFclO0fW3e
HdQEqY1pOmsBWG5EcNgJPP/hNjlkhcNB0A98Rh1gs0aFuSsBBBKy4YEy3Dk6FzJT
P6JV9Kt4yWymgZ1aL9UFgh5mUUFucEwEVRPP+WcQAmpf6Ql1UBxI5zaaPKpkO+1v
ZjWW/gOtgpyLSCOUhdH0h3YrUEpmr8NI24DCfiZoUeO4ERZbjHG9tFmq+uK+oDE8
8ll8DEBS4CPnPmvdLohAKDNMSHYf2GncNVJzV0hjKJ0=
`protect END_PROTECTED
