`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GQPMbszYbByjOz6oz2POuht6KWnRzQsQZMz5S+aqKtKWad89uaRN+DN/JRrCZf80
L2dXtvPQd8yUgkMB5I0/Dnm4RHTJSmNHCAzSJCmcSpLPpTeAbhAV0GwXj++tV2F/
kC23pENiiPMW1KmycB3Y8eb6S6LGnWyRiIzJx1tb8kJjQQeise6Cfa2egU2/6P7x
O1FeqFAfP98/65mGIX2z76r6Jumky6dW29vHhX1+DNA/XQ+FtOt54c06U55K8Rha
1aEEeskLaP8S0rPyaRoFAWraZuAVLPjpVDpobG69f8PGeQNePWDa1RPqTcG5GfIH
LNS6zrajewHVlXjClcbgbKufNZNbzpOm58jQ2hFwsfKXGDkqxJyzHDuzGYHnYC1L
yvfl9QWuc/KrewufeGEaMSX84Gy3tUXtkNmcTu1ho3OTLdr9ju2dQyJHpb+qbwNk
5bpJeufMPJ51H64fSRZMGp6b8WYWCI33CwGG7tS+1YyIKWpRhrCh8lMOA29fNY71
gbgq6rDnQE+X8vuAKAI0c5ikkD/FloKTMm//yOH/wYePBxGzMcMiwDd3EK2u6JY9
36LHidbKH0QmmjraqkNp8h+wOIo9oivPzGn5bBj8A7iMUMobvMzbXKuNbtgB/0iP
ZjlOZtOxuQDkt1FhDjkPVIB6qKx6VGmuCfdztSVRGLfrQ1cwMD/KJ3syIP3G/cb5
j/4wFAuNxjSss/UkZtb2fHcJaVvFjuJoIAJwODV4xt+9uEkya8aMEZFtjftPtHLj
wf5fVqNfKf/X+qa+E/ITR1w8KteCR/b2i2R+ZBEN4IQQgxbD79FE/2Q4PaNi0GUw
e5Z4qOz4BSdqyh7xfwLPnVCqseFrO9TqdslfQ1lWkENegDGlQIQs8v9MyZTWUXHD
nKgDBfAAf1V+C6YXy5eLic+Q1AHo0+0QHqun+mHoJzqXfMRjEhWFRHlhUsMTlGLt
7G+Q6hAAqZGbB7kmOhgpe8NlCAacAuYdSaUnTwCtspyjLmh2uwcPOg2czEF+iVzB
jGxx755OiJNbdVoIdiBXUz9D50ed1nqoiowhj3X7aUEvOdZXo717z5iRnisbCi6X
V0fHYEGmUWpPjDBP9MgprbGzctO2O8nBHWU9A4H8SFWwI3TohiAqa5JkWp8rcf5x
OYSMaCEupk2XqM7WbO8kgE44jUTiWt4ktvOg9w1gezBZF63Ob7WzLZ2l9XgJNr/C
5HZqSG8OpaNdnqcheH2TGUFndLKmmXZQH0OzeZU5Nq8Dw54l/tqGJAps+e2jHYP9
O5WETI1vtSmwUfJH6Y0kZmFd/O9RSjPdYnayT0uTHSYwmI/VdPr+SLNAD/w0QeM3
ajEHwjctKfIXVJ49f4FUxvm+zlZrePrx/XXjocQArcfUWySenQwhJVgYBZf37JJz
rP/uY1eaMVWtV4E3JEj2QoTC8npfWufB0vN+gBN6EcGqWAkE7Ueo7Ac6+dC11gF/
mpbpC7EsZBMUWPGeFzeRDA9/WmeEHRYy8W9u77bNe30grMCsOtQ9a/nfmVxkxYBB
r/2fcyKqPhxZLQRZ58nOro82JhwsVNVSx+f/X/HiZnphzeECi9y1CgGd6y3Lx1cD
cztLWjKdcneYw58oR30CFArWfSvlUz+QLpLgFnAr+1dHC9Y4Sdj+TrmgQa/0YQFX
DV7yzsKYp7gxeYsfIElWWfh3zabFFLuU08imc5kcTSMA5dfSwWwZPzclb5LZOh/H
2auJ3JEnaJkoX8pVvI0tz5flg4h2qeYxMPCgnTFQ9MJtKcU4Zd/yFo9zcISSMxW/
ZTxFdKcdAYlGCSnmTyzgthCItCHjFSPVl6q37mpkNnbrzl/BvLbvpILIsQZsAbgz
C9iV9QmaleLUbYLp5YdlYQ7KHGAvxofd9W1Nzb+aGlmwz3/6s4z9BtVPiwccwoNU
qTJrGFhr5rSlczG9v7hmBCncwi35ZHJDpY50Vr5iPih5SNhxJ1k0kf0J4cWGsGG2
kWseh4HQXp5SnKMK8WzDa9fYxkL7aSvegF3RVrV/MOegaRsszbhEalKmH/D5fZ4M
aIvQn3WBUuYJwpwg+TPzjg45ppQZ1dSNheRlmzHOVNZcuAD6Sum6G/Ef+mhWBgdy
Ok+yhTACZDFV0VmA+cb3kjpssa0IX3YVi27RY37AsNXA42mwfafDfVXcvbpZhx/M
CVS7Rgxh3rokdufJBVFHnICeIxzVCM2DRq6WhO+wAwQAQEPHV/c8gI0mII9Ff/4Q
wQwlkrL+A+iCezDnnMUXH3Dtcm9JZK2raUeqfqklU/KJ7Md2uQtWH9iQY4W6M0dW
/tCrhCmHDjKZ67Zfcy3cnGa2wpx+kj3ST+qIh68B3gKkqW7BhmGe53WGdJ3cHXfC
9ZeSuJAKDrARKsZgKuH2aEX5iUoDW6VIv0dLeSleYmKYuy8Giwa+RICflcRqrO/G
mYmpw7RTh0bZav2nvbAglH5M38/3x2miXw0ZgwsCvfDkXQPP+CQJJbu5Hbe+nBdM
ah8wTpwfODQgz3u4UVdTP26Y1g/eER62qZwwIhRj9JAYeHMesBpI2aDOwXvvp4ZB
kid56rQuFHpZqbpy7eRghrTgck+j/uf+fNrw9zSgnuTwwtbkAgnb4yCGVH9dvgJL
IgtOu2M8nGphx6Fvze+74yxbms+fh/Gxbha0YKjWhSJj+SWL79RDUU/fvCp0OgyG
SulYJBBicy7AH91jNbrfqEQtqsrL5qZbViTy0RKFBG89hAaTS8H3HqHZRXPer+Ds
YGQGlcJDq3xsoh4Mji0Rs6iwPSPvBb6aHkqBytBzvt0ykToFsxBmDyuoKcodT9Gq
eH5BOdyPyMA9A3CeuS9aXj1cKMspP0yO4AOBIKSjqOKrMpb0f0AqrL27LbvO4MFx
kjy+MfshAKkjr4+VmqjTxb+Ioe8ij03uijdNeu+HHL5GgegB99tCZH5lknjDKoOo
EMoNcKVD1qBqpkpzgIJuIvPKJmShgRIVIjC7zLckrfdG+mWmw0mTw50u9dQyE+Tc
GpvDeiz+atp6cFTHz1LfbmIzacedCxeH8ruYqf9cwd26CZCCEQquqLN8EOQmb46O
oK6FZNxE7EosqyHbnGcoPpWRcJwJ7a3MEjAnFUH84VNQL9ZAuxUtkWTzl4nwepdn
WIG3gcgToi287VTd4+bAbskXKxS9cmyjAyE6p1d0g6AikIX7Xbcn5bLcdK1O4XyM
ojfKzUCkoksWcJ7td4fKsDFF5rLRBOW37qhDzsuWQWpK5DSw8VAWzrINcp79DTWw
V1Xb9V/NxqfBfdLdyd2KJga7SLlqgZlSqYxpj/tYyeMBJVyUI14oAVcMWFWXxwgx
R7k1oJse90hOa547VvGcnOoyRt43GRE8kvrgfr/qQDkChPgTN5R2aK1jP7BeT7Mc
Ee2NeEOPFilVjr+WrVjXpPYfLQporhAEas9nPWHhZyK7Wq/8fWYeGMhRMvhrpxsd
EPqeABu0gCra1cdqOysZ8P3u0emCtTJ5p293eFdZgYEhtMveaqBJ/U8zejyUKgLw
IWH287IHfdXpCcxJtX0j+DxkyTbljJVSoxe1uy9kSlqWrGDKCAkgAvmUVUWO0qT5
EHpgNxA9OKsrkwvW7dtiuq20UnD3zF1iTOjNiLS30/Xpdip78vbXlJD/qDt+CItX
vZg7ZwknLiH+fRhNdpEdJO0jm0QBzzUYym+VZi+T5qQgTfIeoCb08AUv74fzpJYR
pGf4MRLBgL/2V4vRKJBE1BiGrwEtuM0BlFgRildUMMuVBPkiy6HZ0G3OF/2RbPdp
xn6T2K6LlvyH2d0JBfrNIvMeCPOigfYWhSR+5KpZSQ5ggKizC5nLFOH1I49lPbiO
dgO2qjNTuAAzEq2GYUqpZggS0kKMPim7MJV0NGz5mqODjanJdj7BfemnMzSndoxJ
9xEXDrF3yEKps/5DU27oJgPuWuK0bHC7U9AUY+r4XBqTeAr3ZglW2cyyLUZq6Ppy
KkJJ+LPCSh5G/VGzdBXnD/RkUaYbI2qZJ13YPjhtCQPUdEX4xl/Sk9h/5bkW4Cn8
A+H5pTVPpHJ0RnEEet4M0mSglMcC2GkV46xj+vovuZk/fv23rrgSx9My0cDdp4yK
mjYjuePlNv+94l2Y+U8PlKUSUkLNEqjpbcsq25du+tnzOS5VibE23unDItDzDB9r
xy2BLuuzV1j+dLln79wNB+a1AZ3kWyMVhkyugvf+Mu1R9B4+DONHOWzDIrFgrOvJ
CmwZXVf/o9hqsqZR9IIzL5se6j31IVdXCSrsICl/Y/jW5kHZf1nmYC8ug7mbDTY4
LcU0JVR6ssYFQ43+E8F8UVE8ALSMFdFWrbIuXiRiUbrrDH/ZpRXreRF81v2tYPdW
dG9zW7YTZgL/V8xeBTxM2cuJG3NB41/2LTPHtMKgjIQNByCJqgH24kbUB0vwkKEI
hxhkLuf+N96e4aWq4CHI2OBSq6p+wuJiMXZBmvaPfttz3WOun+GTbEhY4SM33CVz
zy1Ev5xfs4S24RyQ2wWyp7jKz11tQJA+X8nzeSD4pZgyjMEcPOZGQaphh1OpAHHI
Z+uIpb5rNU8uiHhBt0I/vJ9YfXvB7zteRdNMSpBtj4HrHLL6SSrECz5zl8mdxWz6
zQ1JfCR7kRy9nGSwYLVBdGxNQte+1cPtbAWmuHCg+PYW1/U8kpoUGWRu5apueppU
vXYHjfyJ1L+Xn6JKt4cfiBI28/ntavpB50cpxvUqPfuFRw/6etGINNvqmVmx2l1g
yVgRskvaHeBqjZaqiYouq/leAZMMeat0m4ikbsIVN6BJNtb/CNd7vVHtNokWLVgr
l+fQdBBClA/yXI9Oi5/1yWjmgWCepy0RZU7+J4mF5QCBh4SE5528AB8eZwGbRu1r
CYgTz/DfaL0lvzQFL4S4wmrjfYDt6SEhr9pIE5/VsFIp1rcCa0OOvlVqIXpWpq3g
KImP7CBQYgVNQ19qV24S+PzBJb2oW26KglDyf1FJdrVCv7g2lZMp72e4MQr8Efl9
6uYAkr8V7Ju9OxSOfLmLr6nVb6Oa3YLtoJTbAC+kHUR184WSXtbvTljXTHhAyHIg
OECVcPa8Dl8AE/F7hyA63glbz6Z0gqJxodnXTawJzMcBZRGBU5p4d7qKo53kWGQx
cNXHfj2zE2qi+s/3TdEZSpCP/EiSwgacRh4t9bE814NUS8RqslEIGUxUH9Zy/DzR
wu+rD2KdJfB9+cL26EMcHgEAzCe3Ij9NStOPIoMVsBXz0vO2BKqUbbX2msK/U1eF
B+h5kBY0gJZtcXpBFllsGHpvggsguBZW1xx6ZL101vFubNdADcqEYA4N1aTQeGyI
7smd3TdRCHlMT9JGn3QNaygix4XecgAuI0AttkWjccxXmyW8vbc63intWT9XRKB4
9bDKApobQDz5X7HxtOx3wAcTO8nhi6dj7yzCop45Ym7AVcyTQ7O5L46OFbPskpsj
yRmAbwhkyz1GuqcO1A1KNbAUNhv6TXQXNQuCLq1ycVbeQOdh4IoTOJX1+qhFrC5T
v2fYzG6cR1tiVnMaFeiGoiW+o6WDJ+uYVVDxsH8OyVqEO/zyb1YTCouOdOezyKHu
JnRx2C2ouLROUBwIb6z8QoxS3yoTQcZ3vWY4fzqBbgyho9GBEdT7TqIfQOda1HkW
czRrRvAK2U0/+31cQNPQbb8AmGZWuViIEQ2p9Rv5nNjwF+e6gL0Gf/XxnDkDVApH
7DrXwcGyaK9vhlNNBfUhemvkKrKZvNXO7Z/MwNdu2GBJGNqs47bAneGmF7dSd0C1
ZkmczIlTrcfwi7o2eXxzjteIE8Tkuiqh5ta8V/Be6ukjMS5fTvy6q7C/f9ls3wyN
V9YIMEAQ9PCmFOZmz1exWubBxovijOND9/lG6C7XYRayYKwuaWrQbzRi+GX5+qd7
bRwwyMQDklc/t8Vx0SyMivjdL0GW1Iwk+EwthbYWsYrMh5f+aaME/kegMYUpL/B6
W6hGfDBRlZ36QzYYQ5vrNZwVnZ1o/BODxOJyl0wNmS0syVK4wCvGXAQFfQIPkj1/
yqidhm2k+4WEX2NHW9itxHTj5v+aFSv8WAhAMxJuIk4pz4jHkjr/YvFD/oqt6cb/
yqibJ/3gpweOKXuIT5zt5T31eiy021fPXO1Xsfgs6NcMbNHweNch42EUQ4ZlwYJX
HjlC3tAMqcXIbU0o2+WdRzqeyn91VhKOYniUCHRE1GETuYcuUdSU1Tw67rXPM2wp
wJsOC6hg+4GLZfxeWbeoDwA1FVmoVmbtqnIi2ixsiG60pXEB17bWN16qX+ZNdQrm
2GJaTQHxsjJ3/s9Sn697/1kiUgcokPGHCFeU/wtGSIlEUiAxN6+E/X0/eiWMF0uj
ERwaDTKn8UIJ1BlVbCLKYlbUAC/24wnGovhMkhgcQJQs+LzcGMmQ8Mn5eytWCYim
ROhCLp+7QLlV4PrgT21Pc7sEMizsP10WJNSNdA+kPTRGAOb6yd7KM9msixX94trX
RM9r/eYbm+Toizop79XdIqT16YpGXsypUmIGvoNosuPs+IdFR6IP+LUp4KzbWzzQ
nN2ZgJtHPOurytorz8G4imbggSiqb4sl1nRbdP9F7+QWFRqxZcj0K3FrOPckk1NN
LFplSYDT6+1JiL9wqNPOFu4t2pB3Te/G7Aw1qPd74VkbV0SmOywji/Vcyg9tkCnd
fs1TOIFojMkVo1rF3lsrtYQlZ2WYx8wahbuGvikgm2zGJp/ubPYJXd1uGsaqG078
LT4UgZooTGbr/Eywbo/Rv2i6VzODbOYP1cj5DK9uD7ZJ35gCenS07y2XirYCMeMn
yckGf4qnDGN0wqkRHYpQx7WpuB1qwXB116AMMlEUWIrwOTt45LnUYieEtP4gC6ew
CZ6zV50oWeAV+S9nmK32EkbeFPQAdLnk1pO9jqKQtzva2bDONBN5Tn3m+UPIvMW/
cUTGnaUUY1Wj/PqEbbNeEZ8vyL0nKXYHJtdvHJjppSyuI8TeH7kVOdrzlrYw4SNg
KbJf1asDj6FGShEuwhI44XWYtf0b8dbRzllU+B1ddHeCT1J8rWOQ/MHNLJHGCL4W
5zIgA4ABUXKABHH0+pjKfa63qQPlu9xPi8CxwuhmF9i0m9jmnIxOl386FKA8w7lj
FMdBYkC0CfVema6f7Efr3Gcxjx63pxQBQvfJZ7ztuSONZbxz6HWFLbq42NvSRuzI
lTxaaiLZmm1cDiaZ4u31BNO1C/R2ivckGicT6h3FyKfd7JifHPV4M5ayCZJo1BsO
SfUX7xknIn3QGRVJztaweSu466wt3dfWuOmH452O/FFsfAA9EwEhB2NA4QkamZrh
fZcBAv0PHkcDILFIQ3pm61fUOyMVC04W69t9youGeIrDb3sEproUP8+qyXDoaN9A
+yJ2dQ1re8vpINYoeXlcjL4PaH9CYoiA4sErwQ4IKl6fFSXUO7YsW/9RbhA/Sqrb
l1lfIoSGDH6TFNFh9ZzQ0jlYHMk/XZ8Q599neebgVuyESegUS0bocu4/ngJPHz1W
ZU67DF1rjq15KEFdTZDwIJXL30Qqqk8mVE93ejipxf//YalRKBcz2lAF6LnusP0z
mJDLMhjntNd1zezSHggrWSlBX+J1o0VJ4mHNX5+IGkVC0kdXXrKSgc/0HOi2N6tJ
JEVE1GDKNfIg/utgr0kUTI53Vh7rTwhX8azuUMVIceg8B86T011A0DEA7zki2iIC
b4fARXV4EiVJaxrDWapWE1f9FCGyEkYAkH91mIZhHRJ+1ZfNMZTwViapJ52BQZtm
hWalgSUwMo63Tg7ynv/w2KJNlK5mZ8UaJwW4c5XK/J3pXfyWZmx/uK3Ch4c9qexv
ULxq9Lf1z1PBOVdMl1p1TBSVct6ZPstoTvTTfhDfyBZpLPrY+jiEvp8KXaarlrI2
hwhHxUdphMQKIlu5dDFfn6FpHTB8gAkvvdXSVuXMT/5pHgFG80wtH4Dm6zzo/i9p
7E5cklL6IgpdiZbQj+GHwF20p82vD9wCwF5XAtpJVCZaFTosiT+VfWP4+8+q9kLJ
LA8nj2fXJk4lpbKEdgpqX9J0t61DgK6sZcho0Rw0Xpgj169WMqce929bCRmuWpCc
QBQOvAhzPYqJI2s0FlcwSmT3Ds1mjLy2j5BBtGP+HPwkqvjC5hd6zasknTSgqLIp
bwrI8dn6no9FIDT1VdrziUo5vUnSnZ6EHAWcE9aFixHGQDtrFvN3OGH2GQJHdvlb
So8dMtWnqNDJQfNyApp2q/H7NajhDtEIuf3Is9MLJyvheAN6KclhBvVIEDV7XlX5
1mfjuj4VogKebBXmopZWPlrb9MNzmMnrQLDBnN6yEjzSN7/L1XkVTDZDa/oyany3
+qTN80QPrz+AqyErs/VOqw4J6a2cNKVJ4YeXuQqhjTk0S/8H37h/vfMYU/n0N9hA
zSyyUFv5CYwOm+KT3FtNTcHsoym8z6sxGsB5u3Ci7qO5vMGvGfw/Y7++DAq/LiWw
08oafaZr/cO3MjC/Mx6d8H/NBm6WCE3GvwC9VhF0IR/IiGz92zsZGqsznoyJMF3u
rPqCkFZrBUSva27Tmk236nsFduEMyCgAERnm1Rebmf5fRZ9mvtJRFiJkMMrElkMB
8UlZRyFG+YlJ/vVnpbsoFZaPbz3X7m7crq3A2SfryevaB5I72XmR4umaCNLZgmIq
12bc3D4ElSKqcVlQ0stCypOHFNpwSSCsd0lip2eFqSX2YURZiVeabheaSj37sOgI
Rtnrmn4yRH82YcF6vMnn9LT7jumVmIEMJcNSjmJXtJ45wI0N/Qi2DqhK99RbZk+i
4p70zYhX+V2JNmT3GAHSF51n7UzJL82YE+jvo5LkBcxrpXtrBbq/vu0mKI5VDIPX
6ddIf7zSIcQTMr5WZXKtv0HMsoYp+o7p5Dh0HSVfRWtThE8JGByUu8+9ng4Po5iG
AKyvKARcoC3BCpo0HijUNuh3po6E2n03z6LgNSVPH3N55ZkLSFveYfb93DDhVa7P
f5y5WyxVoY1UqnyxUR40FY0RExGQ8800WUe5JIgbGyos2UvMmAAxr3m1twPi5KQZ
1V8u4NtRvPrs5piizHJyDQTEM98Umyir+Ljo8YQyIX5+UhI92728jhmxH9chdPak
+udbHHGzkrc/WxfDwtqdUNTgQy9PVYYqc+2eFcAtzFi+ZoX3xIuwgBbaerc21EVh
MN2gwBXIbnitoE0gZsaTn3DHXDLoa6ba2STrFfBWsd+Mq//CNZXggkr2kYfZZp9w
f9D8Q3quVB6t/dx2IVjtb4TvCjTmbUtRrAadEmFL4z+aGTBfYl1mIGQYL9AQUbuU
2mz/e0hRqQGtUk5dyogOPghkNbSbxykBeyc3RJvZXZMYXWIuy5pEjS9sR2wve2QA
fP6t6H4q0Zv/rtWu7Nl9fwDofwwelPLb1luMZ4kyka4U1TLrdUq8xwF4i9QwNlQS
Wwrj9sNN/nwOarA5intawHOy1tpd3TIz59twDB8GAitns3MhfJq1BpfuPC2q8NJT
Ey7ro/K37FNLzLe9JRdk+g==
`protect END_PROTECTED
