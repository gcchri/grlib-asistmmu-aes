`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7NV0h/KHmUDCp3Sn7f+CI/gKu+yNUpEaBNXcJMJx43R/t3eUleXE1C2jfaxal4Dx
y4ebVtbXnZVYo2GLEMxSvfBZ4HHcdoBIizfT3/limpSyueT/sRRSh9Bs+Cw7ZK5l
XlygHjaOGYQ9KCF9emzaT9DqSjsjRNC9r7gUHwrKjQJJ3K1mfjuJPP9JUz+hCIIw
KDXa7wSftmhP6WgAyQUtVLeafC1IFvx4i3IkQyK5XfS/4mq+Kn1fquPl2adsiqRE
eyALxgvR4Co7kGc71reVvRLLH5YAlcWzhkFpfWyhn16S7ZbMshwSfOk1MyfUgFAo
b0XmT5kSKOgL5JAms7UJbGuDUtENSUbWHFDBwhtNQToUqGeKiXWeWzNSN9893Vtc
k1nrnOZT+15MPKthYxIO73AUMqs+mXW9heQ9maJqUawgCAqy981dHX2PLQaWY81z
stODgfvHr093IXaORp6kt0IsnDAYcH9+Ng9ZJ0PxJ8Zllz8nL098ydcCcdAB6d9L
NdqiCyc/W6o2XyJeXKaCLuuwrQeKd/fr/XK9+YrCcLw4xKElcmVFwhx+S8mhWxqg
evsLdN0tFLQY5wGGmzBlkmkSjWWp7D3kDEbhMHRtlMXUMmm83KMjHWCI7kRAfagI
jkP5Zs2vSpD+4GK6iC7h5iqZtXpdYGHMewSA7ywdqeGhKP9IV+/XVjRRgajm2+3x
dxiLJ1sbxBuP5PtDLkvz0OI5/zdYhAbqOL+uKrjI++9WOP2BCz6PQ6zMHFv59Z6j
75x+O3Aqu6YVqf3dqTZzMeBQF3k+VN5vawu7wvHu5XnQWNU0r81ZMaVxrRjAlpUt
l6n50Wy/4mt6MlqAKpNghrwWhoArnh5BMaLwuO95iyOwJvLYZe6A5KhSxL/M8Yau
pfOuHCuELrnRpw+J4kFViKIvAlh2ehhcgHcWug1RrQhZS0M7bGpYD+fzH0tWx/XG
2XMcRNAFlgCoMDffnuN9Idke+ct/G3gZJ4vBUazMAFEAysy7GgjXIKXiRqinaBIi
QDpTSY+1ZWeQmkjkGo5JMQlspkMToAh6cidZyB/J0LFJXv+qJFZ8XqOqHOlPf/kw
74OJsbyKNFXoS4FZygcsVb9anRkDLJPGZ+4eFM5G5ebsHxlwXBGeQ4zpvvBNUsee
ywoGvmG9ww+xAyaPkpEsdKivWvbXxh6R+XdXxn0NVakgNZ3oNtRb6TmNIvJU+8pk
l8Zhc+02oV2sR3vRXH0WY5vLK288zvqTrKFgHnaCgjiv4lAEExZ4pL7OdZJXqhnu
EFIg6Hawp7NT/ylwmhkL/bGckZcqcFMo9omNWYODhS8bh/UE3WHX+/AaOW6zZiqs
1qBuoMA2X2z529la6T8LfbT3u5dTe+RRJZWsneDfvwvcmhIivGSUQPnW3k+C01Og
JYfM4sc7dZ6mPbcvijb0l98jk6Vl2vZGtwCpPYibGQTRVPceyDyPU45DMpysmLGE
l+hlWpSemYieCsiDMJ+ftUQoTOK+GBV+XSZmEmcN/PvcktKg28k2EaFNONDRxLM+
in9gq0m5rVsB5ImUsnpiXdcpVnENAbLGYik5i5RhDDZiYU74w9E2GwEvDU4ArGIF
oL9KsWUmhPlhKo5SqlO1sN2Ee0ARjhX1+xHZnLw+nrQR0AdkqReaM8Czrsss5yMj
1ZMGszHRT0S1YmX7jWB2kWlD76EnbIGoM3htghOLhYXB/U482ir7otsQotKGuSIz
jiPhp6+kG4qBtlsP1p9WUX0fC+jO1IjckaBn0JYggKKVWVgnp4nJVuM3CIhPoL6O
FOz0GA09ClOdc7Ht1lL+iXgWsxBP/TwbQ7FZdwJsPbzoFQvB2mOWVbCImnc3PlE/
SCvYU6nHsg01RqwcBMH4t+zpwpQMRpyXGGobOWbE0aOVT9D9elz8+UWvBFxXVBQW
/KjxRIRMsHcBVhabPyChdMVlFskF/T3F7/iwWnC3ycQFr+PTgTwq7baYpMu+n+7c
lA6m+RGy2iyxNfCtQPguJDqKaWVCfbBNgRV4/zV0twtwx1br+rPpjBih6DxV+nYL
xtQXH4uR8s1sl7nUbqVA1A==
`protect END_PROTECTED
