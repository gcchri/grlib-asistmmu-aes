`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LxN0Q3ic+B85DtZpDiGqecCdAHp5RJ6JwSHlpKqmN2uj0WzIYH02Vf7uMkmwtsr/
iBFOjJrAa5pKbWyt507VItoUfM4JzANCvXfMpHFfUDfKgf63nsTiZV5I638S+Esj
WmFE7fKn1yWjgnd5vb4mvPB+Dni9Ss4bXyYjSCdZ+JDXntYwQzm13HxwwCzQjYjn
I0rHLJydLjXDHo4Lhg2Fscq930OdI9GwXykaUFTQY6/xvbX62LJphYJwLZ6/lOM9
JY9StqBOPFJarYYGuQZdRx2Wer453ArwoOgQlzgTvU1lLwrKKCbuk+LzsMVY5Lk4
afiW5X4T8xyhUgJLHVjIAZXEAYAZD4RQ+4ahWUmi8/QJHBvTFUn84wxoE6Qk8rxM
5jhfymBMMsHqO77Gpb2O7w==
`protect END_PROTECTED
