`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
imKNNlxQNhRwPjXR5H1BpiUPjv3DDCngiH6MRiU1ctMvq4yYLQGAnaaq+0ebiGOu
Qj1cHq/lwaROO7mjNQv99sedHh1zALqXr6a4sDuLHMWmfzjdIYu6G3CiXbzfS1kM
x6GHwd+5T/t38CHD77rpsS/Wmyk1Do60u+Msd5R+LH2iNAV8L2MH7cbQN/ejIBWx
40kW1hMuUf3uW1uXwp6Fh7bfELRFbLzvxdGVTqDr/HCvtlCAtm1/owsN8F7Tis15
rJZRi4gUrwrKOshawnifivJdT2QwPCTJMyuBOydEkrSa6kboTHj5iEhyQceQCT//
TRiVJxTouLKS16PGQ2MbYHUhDyQS3dY0Ov3WclLwsmXqmRToN0yoJb5nRrfCJDGD
N6SiT5xqGPj8QTpAINGYb1gQgibSJDtO/ZagBbqzbnwm+hBjjyikSSwhkHoX4m7S
7ytyKAxjSov4LAhQiBap5O9JdT1zLFQxhv1CbZVfwRdKbEd4CwKt8Xwx8jJNPZaO
Ea/0Sb73uMbOYTZ5hmtRF/zgoJ4Vuztmo08Gh8DFCf8TL961gOZdVuJjG947s7dZ
1qdAA54hwY8yyqJQ9kYbZMba+vwPDnvnzjD7iNK0r+tzXN5s78JNF06wtri1/Ipb
VV4/olU7F9eigL4CZz4jJg==
`protect END_PROTECTED
