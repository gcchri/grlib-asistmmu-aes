`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rnBjQoMiRzc6/0Jb5PuNI7cJU0RvHH0VALjfextTscpyqYkLX1expFkE2ytdxm0O
srcuUsaSRJ3TiB65SJ1y1iGi9BqD3KBD1lo836L7u1MFQF1b7l3PV7Ze0Pc5PmeT
bKQjk5Dtd1bpVN6OuTvF5eogIiavhTePzAkUt8U63aZLBkle4s3vrhdjp7xCfbtR
RT1rG54pRgocIHgeB5Drz6taq4OzPKNOgIJEFBu7hukSN0IZzGODmws7rv5znBwg
aeSXCuOjz2hlnCGbJ2JUX82KD3DN69bL7WScEc9bs5Ew0ggK2KYv+y/px+Z5FmmR
q8BqkrJuxIBZ2id+jBUpOce1oJsgtFRci8dArU1iCFM9K6e/cDton7fkD7aIrUZl
8WZBDZJ39SurB6XafgYAKGJnNOqDT0JbvNQtO5QowzmuIiGn9e7e3k6x/9yQj8sF
fQsdx3HpdZAZCewOqoUCq62uYi9uTP3ITS/My1MD6grNMrtVLN9zGK93NFL2GKNc
f32kEf9dlkReV8kKgMyiY6I7JBrAVMLQk2RWzWK16Zq1aR7Jqxlzl6V5jFIU7vM2
6ycNRzM69hWdADv/a+bSPWhytkbWUxdWUioAaw3lUZt0O4mz9hrBVZekuo7FUTYD
Sb6W5MjlNxTvBOBXVgGHUrF9D643d9SvjS3T/uUDKrsSJfWPILZgdpLmhHdkf3e6
Lhojq8H5sI3OuINebVjPHuixeTK88qccEIE1vUn/GkBYOLiv0y8G7cOfb9ADhMur
hsQkinL/6+UNVvMoFltn4Kd5ZZg37Cf6xNWg4y+lmdvrGyUB0cu21HE+Evq9YgrL
pDMeCegPKepPHCQuacU60OTULr5AIYz7X8oF/LGwe/SYtbedkK4HMuVGjfvsQwsj
rMtbXOoGm/tI4rrq+34u3B7uNQEW9PejvenjnMXnH+uUotiX0D+PrVbhQnRZLx95
`protect END_PROTECTED
