`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JAoly+o2kxZ+P2iR/zaZZ2PlQLw/LCcU7bU1aDa7b/Ok/AlxtMf2veAG2+/dUl9B
trIhBS05TgX18p5I6y4bRvAEjoQpU1AJIO9QdkDv/WV50DyMEKTcyrvWHmBEuee2
oHOtx0e/u6D4vw0ilDaSVgHX/nyANkoriaoIXOrsmq71wRPJPoxyZLFd3E7NLMZG
ciezfkFdQro7IX3KJLotVlM8+cQ0znFfilfQk03a8mgBanRhVeyF+ddCBkEQ0Zfu
O5yYddCkAlk5jYC09Vfy9esXfaOUSIWtLTuNAG6OQghUuy3UiHqAoGQqQ0Fwy90a
AbhRjcLC95m24QwFyqorN++6274FpTQPWMBD4kZhaxIhuvrQeng63C7FIK16xx0u
xPywPBdUfSrBhgzugQ1JAuObn8ugzyIGQos9eKXE7qd4VvbnmeH6Sc8HWdiYF0vr
ZEgBSuABSbiNlapEaokkgCVmnKbvNKsshEVoKGyfya2u7oySm0r3Gdl1Vj6yW3aT
NtL8C1vERx4fxVCWnNhloy2liFntQZJZkHu42e6MDNEEqL2p3etPHGDL+a/pVcUW
Mbgqqg5vOto1Hn/72QYNRrVRCwyB67XA4VrDUvWLhdqurz+VLVPZEsjPwkkZxwL5
I7ny2sQeuziO64EsnNU+oH7M3BYsZTClw9ZHY9ngHaSxEZBwV8OoCsCrb8eQR84k
KmKzCBW6D8d1p2aWoNWQ/5xZM/16slEhRgSEmXOb7lc2aTxNpcdZCmEpRN0bzaHg
A0neNDItVM9Pyeuh+tWwjj4cTnImB72Yb/kXQHtdHvxz0aNAkuRs3yVyIO6aS5Ix
bV8o7p4U4gCCGcU+O9lBdk1jaZXQuIxwFEWcJnaCile/rmyDw+ji52shyem+9pDJ
g4v+Yd1CPIg/T+n5vvZi74l8F68lJjU9EGmsOg2kf4rJcfHVnBThtLLMZdsThodX
gSZZ8IBqY+ev2MphqfOvMQ/cjS/57rkTSEDwkbKCjdsIdv/l/6QrVDEOoYD8ORbb
k2LmriaeXr3xNP0o33cpB2jnmaeRRo2K/jgNexj5PvzTErosuPoBd5c86CGpGn0K
k3AfwYtiXp39AGreCvKEh76doihUuBAnQMBFWBntV6UAnvg+RA7IWeC7Jo62HFxd
0AG1VNTu+BgOHoIh9rGSgS9rqgsKdDqp7dqUnOuz0BBaLckxbr70arSMOVf4hyxR
mKgAWX5pMZOQa77aqXqFdE5dRuFLsNXRmE59fQ4iy3aOUp3TB7MfNc2DMpBiPe7v
2kFeMN1gZ8TYlX+AHwiCpfNDPrvwIhuQtc3T0DQDXpdtk6EKyvl4/3/HIaPDN+5R
N9fhCLDV2QFzDqyjR9u3c0gkrjca65AbvrjUZXyHGLWvrCXNzuxqcawHqYJ7El72
p/J8TYl9j4i7HTFrpzlnz7hSYbWBKCAf3u+Sk6uU7dXXylSvldO134scPT+hgaHT
WVr04wq0PfVAGH+fhfjYE1/dh+4PFeM4jW+RKIgpLjTQpyVbM16Nx6yQ6UnsNLXy
+VQN3WEIYXhvw4bBXUEcrOCtsmo9ej/GTwtBef3BMp03Fk7xHdIRiGkF/fUBbbI8
Ez+SKQy7p0gvnZCXxQfe790V/tvoiolK+CZku4l0kvT2mMK8PH3jKDzDCu/4xp/C
qB6TzqfbfOWsdkL6JjdN9G6o01KxjKjZlcoaqZMqW9Z4MYwVGzVqCJM/pUBgIbBF
WMpGhVCpGtHc6lr8fj7Xx7YguiF0qH740l18sWqqXnWIebzefjrfpIVPfPmKMANv
GkRTMz2vDp2MBniPPqZav+E3Uf6H7xItPFkhtmCyoV8sCarGG5UADz8+ttrT1dY2
+5HtJd3vh+Nep3vKpI5jAMYyFlWRnGZL4CtxhWB6vDeLPeI6IhR1nlxjDxr3FziQ
Xu6LoFrZia7V6aVyX1iY/jWpkxRl+TAc/pVWGwFD9FXPlWB9qCO94eGl9LjmfjKv
GZ2i7n5NSJY9iLL2qlB5twQMhaIFIov+HgDPkDh81kmlCHyFEn1nrk3dQpTcJ+5v
NnbltNGH89YRrwiR1Y0fqejoEkCH3Gb8vjDpSVHi2HGJ7V2a4+sQP0oFfXBwdi/8
3j8WRQJxWUn5fcQv9aZquxth6b7F+AOBk35HTRSJQjUnTW7RtRtIUT6sDvfqDVfh
itt9PrDkT8foAn74qTYXS1yxCEh5Ef05IDKsXZoY9is+2LPIJb7NCrtxHJZgUfUV
1fLZXo/R5w73rIt76/piDgWsXG+UEE+FDqqqn90rU+4j7j2qTBaROSBYdKWjrtqB
1bz6mMPODX/e+Q4lhFXlRsYG3qNugVTVnZiW4/rbm4l54hYuUNL2dk8iHJwnKoOy
/Vk5xSWbZbu+VR/0eC5AdX3o0aP8YG6reYo4XqGSRrEggdWgvJm29+3SaKYJ0/Nf
3+gJGfRCsMBTOURP4t4i0Yh78bsflMTVsfZqVZIFEfTPo2zHABiWw/il/oO+UvMi
TOp8Wq+QT5FJCZH8mNVDsQvzFZmAsaAEkm+mnacSPaqwNLcBTl1anDkal5+DDkP3
zerYzCc1uuhbn5e7IiHpdHnw6RI09514N/VcpQ0eR129vdYG6NRhF6Ocg8uzjrV+
w+YPEKNiTQNY/5EcNMPLC+rt7oXn2GcHfTjqMkiO+6hkFmHd2+LAsvSoKBQzCcGq
vo0vViNOzS5zvQ8Vk4qpqtXfFJYNehgBHdlQYWj6RVtvdeEFtoBxHgSb4p6IVw0U
nigeUy5n1HqQaxP3FNP9FNdQ7fmnZE6jhb/6IYXYtoNHjsYO7YBM48zHBuf4cRxB
fzMUmHl8dpU02F8JAaF7lGtRZinhqMYvwyHKkeajjYBWikU/Uck7ToCSSxYqGvcE
0/RYJV01ryrhUO1f63MMpgG1tpDPPsgEL9w/2JK30tj809VWJ2OV90bswZa1s5Ll
HwvpP3vf2CYCo31j3/WLKhdfqWhd9viBIO3mm2MWDz/c2SGwY1UQvsCFvwoWzxYk
nLWvjdeYemvy80BuKLzxSICKerQSpKrq3GYzJNbLvlX1LvHGK4kmfY4nKtS/hXCZ
8tRNcTIhuB4U7XrXt8hkph//WiDXM7HY8zKiBolnAoF5f9/acA3U/ewp/bE8tdf/
eiTk5leYIruIozXY4qP1CRvpVKoGWDd1tvM7JSjpz1qC/5KMSIl/9j9jtW8UdbEh
VlMRbkyb5yXIFMpFF50ymx78oKc5/OBzeegpCTIND8Yf4Kyew1gVWF7c0aWu6qzK
xznIgIOzu3+I0oGU/om5AL1N4huZvE7uLNNw0GBND1emwuPGtiPMebGy3id0t2L7
4bqRoJLVhdtO+jfOVOFPcw2jGIUqQlw+4Q7Oyy95dERBIN3fAmThFh/fkM0rVnyT
eUUeyIpDsKVgfVrmlaNDvNoANNlD2ZqjXQmpsZsSUnauujEz3AoMk1tu+cuIYHCI
saRphg3WHijWpkbmodiFn4nR9hqv716pWaRz5lYfBEV/VFd+gK0NxqdAIOdGGm5c
H2jMDIaV+zsatxbv7rV+U8rbSW0yOpf7KypJPJw078OyH/xJvRzG+ufho2hih8VV
Hq42kJkoBzWMiPIzJ0v+vp24+9oITnGEhNVIUohR0vX0VRrFtyj/HZmmJZ1bM2is
xJl6PMA0Bi4KliJ4z4b9wuzhf3zp6tsCWZxCGyZ84KUrXNwfYcNQWcYW4S5rSzeP
vzw0TAfyRywnVFPZ+kHpHPQnbvAh5JdZAuIlldFaMWE3gB+CO4BFzz7OADWyE7kQ
AAkazJ5nDfBUH2xcBdZvCBh9HnfFLCCQBPeWh1WBUJuSaNsAbK+whrQgr4ezfMDl
Rli+4c/w+CGQXKz5krw58k89dKUPXNMXznVykhf0dIuYCGWCxHhOtDJkXWKxILec
++/3qA2Cmrt0KksiIWpike+bNLgr2w5AYsTeuvCNgwLDHnS1hpY2gZidzLgKF55+
8ilsGhWkTRz1zLYkcNdbFzeFwzU6YnsWELDSDz0RODS7eEeJJc15OTT+g2vDW7Yy
8JoU3SGXZdL2WljusKs3BW1/zYXMaTI7rTa0DqWD64eaexIOTEf0nEZecgj7nBlX
BZZiLwi9j53f1IjRDhEujSyUUk6LzlmqJ8ZxBTHqJQWwxntIQKcB2eVfgXIRo2ks
Ui2CDejmzMcldUySoyQ93upox5ZKgNarVvIT7mbcmh9G+ea3ytdrMp+BGOg/PeRx
ZqzQSiuJ/mkX7g56bCnYXi6Po0msbvPja+GKnaIbZwptAxD0jCYzfLXO9kzHby7t
jeoSxodNHRohd0srK0LCGqmFYpfn472Zn90l8oTzBNKej8JKD2DesvRfmk10FOvZ
Bu8O0d5VbUFREpZN8Prsh6Wg9QpavhYzcr7QFUE8oOAB3y6/gPSgvw9AeHoCfLvu
g90q3q9d34vU7Vxv9hFIcxBW/hzQnIQvzHALhlfJL6xllplc8bSwfzzkZ0SVogsd
+uHSBAu5zC8Qrd8QMg0tBlBM4VCXNgX9/yXA2KKkCJ4Sh1z9GRZ91ivxB4Utszt3
JCqBH9tYhIo4FODDk3OoWEn89ISyY+0v517y2w7yGxJW6P/HQqo428uxd6ETMG7E
XErUhtUMc1EW7V+/PY+K2Ub330EpzS4Tt48gbZtrFDfoxBfZHEI4wVkztpTPv8t7
x8g4bUnMBw10sl4b2z5L+0t+WNWOHmJJi1v6IH1cjmEKhxDC2gWbDCXvCZmoVhvl
wzjyKXPbntK7drp1oE0w8IyWdqTDOvWrV9ZEANrjlZNWPA/y7yJmsv35mvO+u97H
xOzhOyfeEm/PuXdJd8bkuDdzDfg9u51BaoRRglo3FCKK1mBdljTpOE+iQYoFnhER
stmLJRH7wRpoGwUod4y9O4wQqcXHvy1YJc9yJPtdtYLgYOZMw97LzKJpqDSL7P/N
CBRVYasAlT+crVDcjosEnygpx/gxQpj2Qw1MAnsNdALn8AY123maD507LI9FIEcH
bb6aVivmfBE/tiNNE3cPv99xmRdwynJkxchKWawiQK/KGVJrQJqDVVzgjEktplzW
NoIerkD1JafEI1W8cDcRQg0y3JGMpK+vSlLjJHrmXp+FElcxhSM85mWuW0UAb3xt
5hne1MiIYy7RxCq9ALLyE7u8ozs6C7oh11pLEb6ThHoIayNssd0cy2PGv5T1RZBW
wKONkL5En/VZmGFvRshjsfQmj6UZZOvrxGdlx7AKRjMAm3xSDpmLNwLAXugT3bLp
nLr6xy9GJHMzM5OpVXJ4o8Ad6FAWPTJPkpKrlGIvtMPip69+PPV/0pcNTS7ZCOQD
icsEOpkNcvO6Zzl9VqBLRioGRolEqiCVsWA6eQzhpmnz24D/Aa2QQz/o0XUlCA5u
Yo1B8h3mlipdhETrqR+ZQN9oqlWXJMRxYALzvPrj5se0+RY5GwzBOxQ1EMH31h/a
FAJSzTnBBY8zklKjrKyI1Ua6K1woJGmZI6g6ywRqusp5smxcIfdZpYukv3vCCEZJ
BtLTbZxjO/w62/64XljzZSkuKsxGKpZzWc1CiVRRaJwlIrTSbLL5AwQJ9ibZEIdT
3mjy26gRT6o/+g2j3wIRdIFYgq7RoUXsFr+KLudjF1xKqBQoY17nZTwqaqsFMNdV
YL2p/NrZAqViZ9S0P+NITLWHgrqUjuqMuRWMNqbyjcL6RDUMcljIYOkfRd7jFpA5
0Cn32wXd7QE7Me+v/QJZbW5mKXh01J4w6B8ZF9EqhZdw6F4kCMAo2NjhQMx46mww
ifSnypbgui29w3VNu0GxeN859Ctjj7bKTTNXTz+2gvdj4Grg1Xz02emdVLxn0BD+
SwVM/7aEw9mLiTCcLW7q7vxvtSeNjkIed5iCzF4v9/1XGtQ+UbR3HtlBHGiC5pBj
fl5T9j5Gn3kVbtlNP+IbZ43bEvHwGDuwwEXX08o4H8Naa0whMqVpD4L9NmSXJk9l
K6fd6S4WUDThwehOXT6Xq2pIMeSAXt2dZVE68RzELOELXBLNUx+HKHxmJPIGooHd
NU3HSFlUfpeP5mCI5sCBg3/NeuU4aX1lWsaiqdpvHV10HAm/VKlMuVUGzkMqrvSd
D4S/fEibNTKXVrWYQWjjMLOtnhJaN8ix/w/0wouEg5ynW8PN4fe9Nuv1SqOJhfWa
dNcpmm7FNBVbpSwwZIxV5yBUL3ijtRaCtWs9F5Eo5PY58xrz4A9aMvkFDEhFbTyX
klasK7jZC02Xtyg0HRDN6hIaKEbl89bEgvTTzvTnkx+ikBKITqYXM9yLV+Vj8Jn5
rBF3mAGRF43M4Q3rZbo8PyPm7syh6epC8jzHf/Cr3m/bfYQEA7JRA8YdTJ7RntF0
cjE8v03nFuThVfcrWTi2miWkFnOf+GhgYQJPY53oGfRGhILVlNfBcCVugQDeTir3
JjCs69UdhM/N7SqSWFY0wd4AGCwLtACk6MQW3GVmc4M56AYVJ+chrD4OU+Hd4BHi
dhFSCjGbTqAsvWwp2lfkPYnlZebojoTDCdH+46vkMdHMSKLI/pg/uiEBcYMoLfXy
zBrHNruiUokSI1+ncNe3cd1WWC8Gd5XhwHMpBJ7DnJfhst+ToEimYsl7Y75NrEkA
w3uX9SU0uNvXOzWd1pznJtNWwJ4icrcylJ7+Y0hiLK8Qf7mEa8NHMqc+9QIGf69o
XscNdbk2PVlBgKSyfMZIJDJ3FS3v71mI/NVnQPXURwi0js8It7tGZ0ftvPKcXn4M
QOygRqEmpnJZWgAPUJKQFknK1VTE0UokEXlfdhdo3sChEQ/gzlnJ1jFn6chGvUIn
xvxiSLhS6bKNttog7j1W80IFSGw9wvSpPzbC/uZNbQQZHkwPDd06eeieFzRFQEtD
oqAXiRgY04BC2iSS9sAk2mOHgypBubRuy3+iHIKBixwXK8Hdpnl/XIREJ0QIjVNl
NXuxO5jJuyN/uKQIet4VuS3lZIXdSmnwXFq9ugv8wRWrMn/j9yDsDvfzVC712k60
BWf7ezj1Nd27uVJqPOxAR+lQYrRAg8zq4UsnLbTAzfxO2UjCbHGpD50GbQGG0zJn
T1uBJWNjYArgdas0SM3jsfBQSXlubA6wcXBz8Lz3+I/K+Z1vcl5CAOI6WtNE/OQ+
TG5ZPW5ypOZzKuibtFjANc25mJqSVvZg19OVRkY4ZO2Yb22ai3kUJs4NYeqqq36r
ibL6rQZxyZVBH5vx1BpN0/v6sJbX5XELD2iNDz1RPKVEPPFdUrScFOkFNJq5NJYz
SyDnUYDr6Na5u3xvi/9rDuMVNBR40ubCMwGt7DrKuu1HueKw3ubgG29tMp7i8JPE
ufwazL26wklTlmEESzJE9ljI/MsofS4EqAfHukT0F1roVeR7bb+tOXpx7v5+I5II
YobPhN9OlXTyc0JHd/emuLYx/wUBv37QFj0LJ1vUNfkR4ik1V8zJOAF6AEP4dPVM
suKexgsXhRR966GJnRgfvVgT8DZHx0rwCgA5jM/OOm5+3drmZ+SR0H0PCqS05cxF
YIUcxLwRKFIHDjq+3OaRADalCAPphh9fHRN4qnRKN6bO/dkmzuCJqddfoqm1OXqL
TpOC/pnj7uLSIDs/019ulpGcSvuPf0XsVs5C9jcPGjfaxzbGL6Jv9JwO4R5IRrAc
DZMu8aEgtP6B3V9IYacFk/3p5QMzBebt8wIT/o/OVeLpzsfdG3J6Vjp4UYRYfGBM
ZnGMZO1EcLfkaTr229KjT7xERZbKfbrBqCllQOymMtINR/hYtu49mNxfieFObo7M
H4eD/Z8A0Fbjt+6ZsHrQCLCQMCaizYCMseu1kGyi5+3BKiJxzM0KdFt+QcNbQpE+
jxX9stauwnGMEcGeYyz8iUSXWb6trgSoDZ/y72H5f9EOhJqmqx0xCnE0dCKqEnJ/
SVHeKMNYh54sxiqkHpHyPzDjyg7wBSzIr18rgEaNVtfahxY1yrjeWR9zppbhD/m2
a29odxpoR1UFCRqxIG97jhrA+2xfEG+KhhpDkCEDc3Yuq5XnpqWdDSz3xCjI6xuo
CJbwHNoBe+/86ZU/XrNuILthvqeUKKyS0LimSuHVGn3BMxhNjYVICe5V4CuWpR9E
V80wOU//krsot52s1yu85LKBuMwxKICfSvoATxkbVsm9bas9LXfjSafncjaBINHZ
lYtsfQ3CrDXPT9dniVQgqOWAsKwjebtcauO523ytX5G8pwAVOsbPd+pTGEwDEL7k
wLtEy1dwUyue9T3v3atCvyQkOU2eqKottfINPWT29qsTo2chJ3Bi9bo+lIZB3QFo
FTP4h2dNwYyxnYKJXd04VQvatvz6epbUBzg51j7epPkPOQWzxDGMd1VuHR0nitHS
3MUMfclGfj8oyMsiLQmprEfz0r4i7CmLPoNnidLFBjurqm+dPvDo1xKlFyWQ3Uyu
kyDV6vWIv6w6OyldXz6niBmLE4Iny/dqFFhUgdDua4jmSvhaqn6Jp4fnSrqJwtM2
Ktgha913SX+vc3KuNBZlO01CHnqmBCiOk/oxOAdZPPSImUEZkj7IjoHGQ8BDDxdN
uwwUEB2DX/1Mvhn1hR3SvmkZyLWw9Dtghzj0K+PsgNbzzWW0TP7iRTA4QPvX0/Pm
YXffGWnNH7ArokDpIpkchQgDsNx+a1mzKHLB1BswiNHtxilSiDwzgclTp+Bqt4M2
1rDDKRJwIt63rRf2Ay7jVhm1WHo84P5zgqJ+lLI5gAEIiu2LmBm129H0VAstxEo7
HD/u/eRck27pnIwtNh153ofP5+0ukr3tL3okPe0Ppaz1LfZElWQBA3Yba9mLHE7r
opmPCl3fqo4T3vSgzG0GwSHQ4JGjPQI1b+kE4yEFEyXxNfImVAEN/2/KFJldjzj0
TIxbORb1Nx44gb78ZpDyMGRwZk0cp5q/HAFrw8IUuE6hXueXBU3obSPR1Zoe3CyM
Y0mn/Yv4pRLVKiCEpML0/sl8dlE2k76Y+PAK9YUOFMiu0HlPe7Tz9MG0uZc5zATC
q0rN50VXzeop7KnQWBqfhXsXKm4/Kk0QeUCL2RjywjHFOLmsLLIoG08z+9ZvCR7H
VRNinANDRAs0SI8x1Nl2k4iYRn4QsjgoQsnqDmp9UvXwoJKw0WF/qhwwfktUWVAp
dVgnNbO1pVQujrZo5C/ORWkFfcpfE/PJ7aI1oOdu5VzGwnBAxBWBbQzJFzu5JEJe
Q8vt1BIhEyff4tQ37mSTx8hIoHNh2mRXLdil2vcFIDP2DEboRgjH/yiuILw05WPU
QLE+5kjtyxYNiB/XkRhLV1/Si1N4a0o6JWtoTGEdVDN8Mu+atqket8OfKdLjpEEu
O02i16if42MtaLxR0pa12lirA6oH8nreteMDWJNdKhZgGz9fqnyHFURX5nn1hzck
Zv8c0NvXtC58ZMhPGWxsdikPuel8fY1Dwc0m8Xd5KKUJWU43hiCVC7D/J51SWQII
QGWupadFK+5GdwPuZExC8lF5/2rSH+EIYR/wmvQO6jYN3CJn7rXJNR4kUy0Ek0S9
Ec6xHMUjyIE5UiGsnDpD/uqdWauE8xcCoajE5C0voKaU7MUZvQarJgExPBJeUdJ5
Ux5xFwhDIw62Jbbf4nAxj41o9MP7ROUTtLGPNIL/ctwTy34YYtRFrVAtw/FPb8yO
fEvJ94AVdHiBtfh4Dmj5JVkpsdtDOZslFLOfR4fKb6JnwBXV//nqGr98l+dQsasz
A53t8KyM9HQBLwLfuBuBK2vgSyUwPeQoy6/1VN3TJp7y113FxlBVPLrneal4At9n
Epy1D5oCceQ0bZht7JuWwXR8U9g941n20yFk/5sdE71JGx90v9rxB1xoG38rtfPm
Sk+So3uJFhwRzpG3iA8TA32P1fXRzFuFIp3ufW3lgWw7wsoql5vr2uw0c2ySBYSW
ZyzHBP/PZFO4il+7+6mUez4cePsCv1YnR6P/TDGgomRBv8n2BOSB/PiQbCPUsgr5
HTseflSa49N8o2FZgxQB9PB6GZiLHD0nLAbqLr4UABqlOXRy/8IANRcKNNu5E5MW
IsWnEZji9pUARp9hQ7dJi8yzrRoz5xPEUegZWuzYWunPL/Rjb2uj4ApqXBLLr2q6
DX0XRsI+u+1X2IQtX/H6aFrlfxIiHrdoy96j6eHxCwhp777ljKIoG0ugWLhaKQkR
8CkXbX5w4sk2tz4vUX+x3z/wx4fDwkKUe8xZVrCiJHRxSosoUCqh84Tnbgro6FCi
nnQTwFy3r1qROJlEZ2WpLLn5rOcxLfRxHlBRIVb/x8a2RJzcEEPKbrLYim9QZ28A
/+iOZP3bCM+N5IaLjsEdAOfXNOR4CmMFpIbgUKjdhHtpTVG7RTSVncBGyUalBfD0
0gxbpp5aA9ZiXzicdFw1SJE+7aiTRzjdbBkH6aXctFE4wBgNYrajZsvWLcqHJsY2
IC03JCJQ+EE2ElVuCRWZ2Eobuq9klHsqE8uUIBosNAvcEA9L6hFmb1on1YblIFLZ
sj8y5Mvz592jxjVTTjzUTTrMr+tYcKpSzg5Dj5ll8wSKxe5rrCIPMT/yDB840ai8
9Sf2Ufsf6ejWy22BINEfnPpch1tgTBzLfJZTJa9OYI+CYV334vcATMtsAJ/ns5ky
qSWGQSzWH5pox2kt+QOJOOX/GoX3/A3gViH8gBP+THGWIcwlbVtocBUxIzF8Wogx
N+CiB8Z+tH2gMsRsaNUxZTioqpR/16VUPDvhaa4U/d4tsg20Pp9RZszjOXluMqDr
Jrkah5BpxgkmvJJZZT+cdFmIM93+4vEgwC7QYdCVyqy68lLi0rGi9gIUHJBfj7oq
eGG5JjCEYIOm7rkfVpTFyQQBD1Ppnhf6X+p71xi7LIIAxwQoJj0cgyYVydvD+xSD
QDjrBFP8Brn9jgqs4vZGrtLoHpoHzX7al8r83kDNY0nHo36S4jJd1UGboDw/QRv2
OFmdOCGuOaIw2GcPiWppXfMaz85IX2Fw5/69HYuTqqBYTi+szWgpJVxWOvejvQCP
rCGmMqlK3myHsYv3ACRcvVCiSkv64rIuCzNA7yVWF49yvitijBv/YXNVy9Az0yiS
4EDlp2bdnZLju2TR+o0sgNnQtwtwbkqC96X9SEQsIuIfrDzvgIhTS5BCvG+yW4/k
Lu1F+xy6xu9mrzWJWCnomn2P1bxTXjVUDH4ImCkzBwEonwMnRzQRMX0ZhFfWjtcZ
7dbo1/lALCeXUII3aDxOicHjZJP4PjOChftIYU2ZokYJYUb8AF3oyOA3AkeC6By0
hAiA31uX1lrolhaMk13TMrFxdj0Hqh9Y560Itto0PXGTINYVzleDG0qxhr2CBepM
RY3lUt6TA0Wx6AGYiGB9enIk0L5T5VGLwDQcuuUALsrhm1jPMti9l4G7b/kyAwKD
RtS0JGJIFJOt6ezBNhXKjrklGduoJUTe4A+JmTqQNeSRRDfVDSpv2+Ddp8T8vaZ4
oIn1bl9qms5Uu71SyNqbIQsJAhhOlW/zk+x/IVw2snzZFSfzxanWxwxO+MjiIZC9
4lRswE6Da1dsxVMeD40gzjI0Kv+sb8fAJ5CyXcJhrccza1FRvAD5YNNsOZ8ObOdS
6BUOWbVh8gRCeSPJ3/knm0tEFrgcd0tjAn6ticsz8rSauPWzTi8pqTWn/7X0dUxC
1S18qHZtWaFK8fega62R8V7XXu1hchIMiK/MWcXcWI3I6SoyJ/HGFLtzjOk4xkYZ
waHllSuuKYJlsmEXXyxAZOH+9YlDw8YNIr9sJpKLq6AbqbF78rRSwn5L6HESD9bH
KwdQ+OgFmCtranouSLnh+VRht1N7yXuNp9tv/2y3r4sG+3rTDL61Tin5ph63Onw5
ttVEfM8YwOPxzBhOFErX3/JYc7/CRyTDO6i19X0aerj8/i302quj6i6oL2T9ArlD
ORPal+SYwkWdVZD/oEJuay5bd2EI+GdDJxctHXnMAKwKcC1ek0+7WENjkr1qsh93
xXhv23eA0Q4CsSPmyLZ3W+T6WNDN9KRLVcPU8gdIRXXkLInoGopTqxMMfsLG0+Hw
CS/T+h984lRrAL2UeFLjbiEp6sGA4SZikXz/nPinP6OAIbkVX6OHrH7jPRT6gp9U
fdmBVPh5Rp8C+kr+AMPK+EghtAgngQmHprpdFOa2gyK5uD+SY+6mYW1YNfFx4jDJ
F79Hb2/t2BwAaCOK2xB7yOJY30/4HFCzTSalP5fAFTyApuVFgUWzAFqbAOCI/f0a
lTVVrujxL+0gMZb9X/5lTuPUUZdbpg9kQ72SQG051pI3EmSLzWmqrBYiY8Ukqe8S
EVbNDnaTTjUwJl0qOSMnJFNL2AwIK/bNH8mTqkMfZPOZR0o1CpkD093Q0tXXlfy8
198v0jOtVPNEXaXMI2NIIfz1SErJEkCOSjL3qOz8Di/pKTPDelLkmzpsnpq39yZS
JWgfedzcoSdNlgwEbucraKZ/C+GnzzeaV624CCQlB46h8FPpoSDer4W7n9wqsF2K
kirRbNuhuKg5tnDzCcKQeFIkZJIXHh5lIH+H+SHl0rCSIm2uZYn5YxDbjqA5Cug+
3BGl1ZV5nTib4pHts0ULKQST7ORCtqPT1ArMG1N2A/Krb7jJM0mQdOo7L2brpD6R
ktamM9Dx4T8ZAlQHaTNyjqOzpphfG1Ij9HbuNBgourQmczW6qKONYC2KS7F+Bg9e
LyRCracGcNr14pnhSiuceNrYtlPSjLI7leKkXKas3lsK0OflmzONTc5O4kTwjfGb
3/uxlE8+p/eVywEBEBSknYBTqfnYhvyELLkSRZX6gxhYnUu9V0BriPIZlcqS+6zN
n1CzxSNI09wX5Om1/OtIxWanheOATKgIQoQBTTZpqx05505ZOmcA1XaMHuleD5Pk
3BW1ohlCVe6TYI+mXL37JLisv8rb7C1moSu8tlN0cgpF7G4HZgtf7Kgro1lVE0r8
LkxTSeM/USLJUUkxrSK6qME1NHPKdmMkobxhu2PI1Buh4b+cHduD055IX6JruwUC
fq5mChyvzHb1v57hNU9Kodt1CgIWMWDH9etqVYFPpp7XIrPVUXnDTZR279+gP9U3
9VeipHXu+h6Ri1PmR87hkYqjo090HwkucZDrgX/tWK69sIxu/25p/OEevxiz/m+n
GWyWC7Kc9kaEwr6TEkfH87mvsZVfZJ/zV8ePIMBLKPqQOHbNkqoy5me8ufv5WX9k
VW++09BrJOzYIrvbKdCbhQzbayJA7CFLq4R6gAeejKHrMnh+13346sOSIbPgV+qC
k4pXUf4npdpuIkxR4l5MCOEAYPDkXTHFmV2Hwa4xDLK+YMkhl+D5jh5+pGcx3/CO
YD1cBZ83eT/5Rshy5XNLvE4TG+IkmP3m6qfXX3WMPmZcJzXnSMdmk9ODWCXxYzT0
IUko8Lf/4EHUs9WfQiaKjEqmIZX+lelg0w7x/yjimlho5A0cFEdu5p31J6u4KlE8
Wsj3rZoJG7ZPXLHgD2HH/DYUe982cghG/KFBQSK/N5gofzLRoUrvaV4bzyzqL8z9
O7qPdvzgNy2euzcoN5WfYFc6xI17A86TaV1I1OnHM5sZngXH4H8zcJ0bnPuW6kPW
MSFO7Fcw1rVgZDc51Ef98pakQA7M5qr2yrzJ6qdTdMoY8uK263ulkfmG8Og4BLBt
lkO/Ez2uoeo7KyKnBLpKPYmoCRo8fhodsgGAQaETPOqSRf3gICd5dEH/P8Wec3Do
iIy5MwT8/CIAw6s/cSOb0uz62k87X5c/g6exX2UlExU8NtiO4khtwx1siyRRNE6c
qltJWCTMnhKBq5kyQXqBP0aetzBSZvYrDuB/GdOZMcsNTzNM3Dm9sclKPxH0+4pM
VkEojaMEaCQjbQ0gDYwPFMsyb/74d8i4TaIiu5tu6p0kOuUH94It/CXP8FxmgBNc
Lmh1cWeiCtbKFM4l4fG8rBs60BCy4GJXaixVjtwW4ebU1ZtHg1IhsDkTGHMYLjhL
7/mXoVuSLXvPGNfqd+VYOsp/W3WUnnFlz+QWk3h+FCY6KHJBsmkZj3habZkSJigU
3mn1bGNE6TwOqWT49+9FiVPmjVZ2oyr6HFDROLouWXUr9FTEFuxMAOJsO7X1pfqO
7/XdMt/iVCM19nhBFxtkRHAvYiaXmrXJyfl2cGhkXRQaKkT0WHHkUDesyjxhnGgz
2pK0RCIFxp0U64ULaILj1RQGgdf9rDE6wNwVTFOANE1t+sTpppe1iwjCiwL6L03g
pp4Uk1m3wk8i8sAG/2LSYHrLs3cF/oDm89UGw/8WOjnVjnwxTelbnU/cYHSoROfN
9u99vNvGZxk5U4rvjWfcRV1cXR/bmBiuXRmyMR2W08q0i+MAk7WPQDFZRmVw+ade
cFi1SGn4JSPOk9NVqtLRSdNpPbU3h/gCagN1K9mPpI1nQADq5S8oirSTkTcovS9H
Dwk4zIVbKIeLbslAtjiJVnxe1yihgcOGsBHW9tte0SiCebCsaA3/rrCIXyd9f80k
rYjTJB+rBsMcoKtsXOXdBe1Qr/oRj9UlV+2mO59c/ACKwaec4sxWs4gFbeAR/Mn7
cTddU9DO1oyXCql8gcARmLwslolWYyG3fQUYZEbIHqu3GChGu+2uKsLClR6WhsN/
Iot9xmwic3jVPL/gpy3W6qHU0HlEcv1SXo7je9s+lVsg+4NM6FEqDYghUK4NpVLR
CT2ZCKSx/cF7qtsWyMSXWcOspqKEFOuRXX9WXOf42aPPLk2VJuefnyQXD++F25cJ
Y7bju/J4hgNZarLkhSWmq4fKQwM2bP2/2gyX4Qy2CXdz3NCMX2uxxSb4d2K7hBCA
amyJX8Y7IZk9nxqdynpMiKoSjMKOTEg9yOzqPRoHS6O0yp1cAgiWct8ar88QxI8Y
hyQZnCDKTxkYwyUVHDNqzO/pA4/ZO1Au5OLVZsU+k/JLZE6fxIqyafU5Yn3EY3tD
q9dNDTSQZVhuy43V/PX58m+e2/fpdyfcgxaCfWEIIU5NnsbGBuDBDThgNcy+/gLs
5i23TlBxNtM2PP8eusMjNFsg4FziW6bSWy7HXZFfPA5i4Jsm85zN+6LrtVis7cFS
rQKzqakt6AQS5LH5gqgcZk/NX9a8+z49nJD+4ydFQ2Kcx/DPo2+bm/jkTKqjyais
jn2isD0kXjtTlQJxSHkg9wXDHlJZ27ULdPtucGTlG2K2rBVNQmiCn3L9Pj3nXZur
s1H1LHBDyZCxTmUVdwi5Se3EvMR6CaUI61rVcKX39I5QxNclTc4QktUQ1KAuI9kV
R/I1C6WofNhVVs3pAJn7iuAFkXw6DKq8GxQkDs9rEjYqL9N3A4hLneSUIJlWx9hd
ANAdwWdRjlRrzFfFLyRnJFaJ9dBr7xM5kSSXEypiaAMgJWbBJN0gUWczIAFXz+VN
fhF07vY6oTMnkwDXCyG1ALiz53sGFGYoTGJiVMsxoJOndgLX7yPtrrUinS+N34NV
areTI4BxeQ+1ex5BF5wIjgIsrrqSmmQZPczUz11JqHYsYzi/RJeDpiWbd+uK4mE6
i6+NVhqFH5sGJKwsB7KFlnAnr6ibP3PVe+9o5ZLFn/hYG4a+CB+27OVoM3wBKTI2
EQ8HJitf45wypyesX4Wf/uGO5eb5bzhoPBqZXPVE2omyazOBZJlZa4atcHbKBnyq
2FTx5t5wY0kE0lBzpFD5URKs27btFpXYZsWX3gu9DJoR3HugBTz16k5VhrXgmTAa
WnV1pvPfEtCn0p4LEevJuX9tL13+RVbPIy+YTzq0FI0qsbbaK6imESDd4k9HCs4K
V+5WSpnSdjl6wwtWfx9djaPfXT31FDH4tpvhVk6p44WwM0QF3/aAv5Vv4KNhE0eV
a2KNCM1PsDC5YFF2TRK5WKMFVfCvFyhS/IbFzo7PPn75awiEzc+Tf+IKXWF20VBv
bvTpD6sAYH8r2rTO/7WWZyplvjAGpY/0NkcHeGTQljkH7yDJGBl4mJsbVwk6Cvuh
p41EhamZV7IE3cQawrfovoMGp/v8KdAQFGrJj2kCcSPx2im+HZiZIwBx9U0pgYc2
b6Mcdixp+dd6WPeoclkuTVt+j2TDB2HZxeUGzy1L7hdpBD9AMoeiCtodUm0QDrfL
uF4kXagHyhuoMK0uAnfa2hQQExin/z7DAyXtcrKiuAK0aKjWetufJSQY7sWv9qkY
5R+Ha5dPevs7PV5jpUtnQ8zc9Aj/o+PA+5+DbEP3eK6k4URFDwFj8QtUTB28Iic2
J6HFnyfK83Kkgswd7MRNM7i6kY4i58jGBNVvTHUsjd73G2b0W4wvy9wtnBr2Xh/G
BUTGHS2zRA8APLevSG3xcIPKam0wA5+ZhiN/+vKN7D6BlmCIMfO3RzAWCiB7/ZOq
tZX0up0+LlZVlSAUR4SdsXWprdk3BFMquic4RnzUCJJMwKePlH7ZyuCl9bSa7V2E
ne+OVnXtQJjTkBl45NdJk90OikucdTbfJw+kkqWFnpjiuO0lnyj5QvQSKBDf/Od9
4jom6f2CK/T7A0BU/Nx+9Vw0sYtdVX22UYWrkxbNGMCH7iZauVuSXeQBz801RMLn
U/ABG0/sKM7Dp49EMUCOQ6CEDWPMF4xKgQ0ef39OPK6Z03VTA7UcyysNbvBWcxWu
yM1acxNzlipPzoskeeYbTW7UBl7UoHufbMaFUQxbJ7uuMJRzaLTd+WkoSxTmeOM0
HdWsH//+GIw8WsjuUt/r7vYe/tUy0HVC76UzhLXZK1QJx5GaxS0Qux5z21PvXHsm
Hmhd3s41AKorsDBRvWV5GVttHNG5ErWxIQ2W1JIQGIsSXU8ApTaGcyXD0jctWQr4
/YlLBBz+TJjCTy1ghog9AaahfZMPl0nPabYe+CLPnVwZVfaEMzbd6gHS6lsz8U7F
tq3aSNtcaclD2gmxMwUJQDSQLEqneSuV7zWVK4rqtJq8DBrO95Q0m3L6LCqYVjj3
sKM0/uUBM6EdWI6UnM5DOKEsFqT7e7yBFfsPLAjAF+k8dFsnP6P5N2ennwZFO7MM
sytQOYf9a59KH0icVpem0AW4167jZucsGBrZaPq1ljiHjB8TKojekIvOw61jfFdF
vIo2ucRT28IQYjfk2oZU/niisEI9b66eEOKvNZRWASf0sU/ACq1I5uUS1eVTcyXa
Cgo6eogRfyCIUJ8xpK3LTLGjmf0cvIziaK2y4rXByBMTDuRHaykPgxdB7JW5DY0I
civbLmNHi18j4FWghOQKjSxg8GerVtah9PS0feoYwxYM0T9FNBq1zXhagAM/mecs
li6clYmKNBrl7BFDIoDccU/mXUUZTuOc4HEbfM7EQveSzUD8ZwUPV9pIczB4VVmw
vD4TnYqW9Yo6eNFARi0V0/K6FJqv6DAUPUIY2wl1khlsDzTeFhT/do64Ok2c+TAP
wGKEue0PhLkj1W78gojFuBwhu34muWbcRXymskaKOl5Q84QCL4IDpU5CxE6fvtsH
ZCJj0/QqByT7g7OUnQFtmmt0ykQpKjEbZfP0L25BwA97D1dJtWwg+VVm1dKS+pE2
l6AETNCrN8ETWgSznkwrdDHsbTVVjaeVnTSJVrernAz93lhZ2WaS239XMaFTTTbb
TyoVVjlUc6qJujMIkxAUbYeJgGAGpnaURuX81Et4798R8+TbI52QrY3Imsu64h26
ujIllDgciX0bWaWuQJn406+0lkECO5V85DdV2Q9xp+yxJ0HEHCGPEQ16KNtGsjNO
jSZb08JH5AZcUKhGnlL0CBi692Hnb5lcBy3XPpqpX6B2mO5VWGkz6qHQyNYc5SpI
KVSBjtaVD2pjqwA3OHVG+apxoctxsgLxskaULae3/hujtxKMzeCLHi4FBv9FvKyl
moSzeeztx7awRCQPQatm15FdrmXa1Q+MzCCMHXXv5odpgs1AMJ+F65vmbHy0kb9+
yFkjmo5MDPDeh4LGbK1fE52L0pWRhoL9FkYTGcnK+t0mf2xVsYWHUHMRMHCIRpvG
lOZUkpj1b8zqUDYOsJSF+jE71YEhgNRViwfJqow2ZZlPiUEUT4yR4YaxYeilbCsJ
g2HynLDLFqfDcEGNvXZ6eNK/NHIhVDcNL9IgRMTsS7IMeRCNDzb/algZ85Q6f1wg
Q3MnKf0Rr0YjUHO/TGHXv1KcOrR9Zd6SN/G3x45CNPnUXrhkXLmoMOMLrb6rEhqc
Rnkz+PL8G6/58ASxrT+XCdzqNYxgka23mDEotZtSVrd6MCMxFEMTjYAoPsjwX9Y+
eMWlEgtdxx+HuFXEEkQ1kmDLE/7F+F+4laAiIveRk+mRCwG5+cLUhBPIpBH+G32I
B+ryRGn0r4vl8hDeO3+gM486MNBnSPjxYQ8poQsujVW2nc8TrhDxs3rED7GGsE1P
wrngAc5CVOLu1s201fgpYJJLizJwvpGKKj4uR79bbjENDaVmMHKAVKvWxt6xmWRa
EWQoxC34aZ4NWvrjJqalhmv+w0EJBddpFZiYfyFTVTRLFJejykJMR4lr+UKV9qIP
3TuzT5UVIaWmg/MSmhI9hZr9azcMy54k2wlFamFStgj8dUN2tHhznQj0X2JN4Gem
gFmKFU1080OJezLn3RZcfq4aA95hdjJ4Z9qoCUSLa5bFXFwrSIAmySoDbZMXnR2J
49EEc6yJ0SDggPDECGwrm/MESD0rhiOOA6vG7OglHQoCD8oXE+ruBszntHZloEXN
cDT8LAdB7lWVMFJpC8JbQgWwEVKuFbKcMisuUBIRx5mbkdMVwu7ulLbyXnYHxway
CeutmhmyV/sN70f3ytovanAWF5JMw7I2ge7qjXqLY7BvlDXUbO9FQcN15NBoQqAu
oPmcxCGYWXgzULozoj5ZBXKhdyRqfs87zydDEdNlJcjPPTwQ9oOC685AyAiPudUM
emLJ/pl+87mxoxFAlABpMhnUyRV/vje9owCxt4LhDwlNUqV0k8nNwUPZuQjAE/8p
WaNs2AItysh6TCj9FTxOV1Wx4w1YuyQVYPMOl0/7GKUrc2UL3j8JYVOWBQswmS9u
P9AIjfsxPcD2LaRm+80DP/El5RLVO7qUmTJM+RKwOO9VO4qGZR826ZEQUc7GP5AN
y01EoqbGE6Kto017l5kFinEAuxltKhgs8+cXKp8h6J/YSeuf+JFIjyN4XeXwF8Ac
tIrAYwofI9IbgCRTtfGeQxNbQkQDQ2GfarIXSsup8qMhAD7FqPRTqBzzF/A3AuUY
wRbf0zpaoUC9n67Qpo/x7WoW5t4rIOuPzIoZLH09c6HJGgBYxbBo4Z43IZhnPKIS
oGwDvvoZBF44CiFiAuy6SyxU1lUWRGuxEKMXQopzLfL60d9avYO39aIIAJpNnPSQ
qkkWJ4Sli2d0GOq6sX9d1aWe2yBq3vteWSkaAGiqLTap4sjLdQoRur574HDLU/Ar
l05LnXEOYt0p9bne1noj7Xh3gqPNnXIQCMCPLN2bWSFulhxXhYNX3tQiaE/Ie2A5
2BYzOY2WkLW2Uo/to4enHVKSrh4C8FRi8kkUFGZYOBJVudNat9+WOcSnjpnsLToa
eT7mUideEhTIFu0/fzY/pimUCr2pIWdrgQhS6ia9CPSn8dffmocvo74jHH12VuOv
YigReN/oX8uNj+QgMXUEAoO5+hetOotMQ9AAy77b8Vn4dE6bhKqqCKke6l2tI8J6
+n6zIF2iTlLpZG7TQz+AP9d9Qpm60Hq/0khZNFeh+mjb1AZOWK7W8rjkrzGygqvQ
yPHnJ5GHWv93NV7usjm2oC2mvCK1WVaNwoXdPOc+cZTdR8CFtNErNokLs3+4QJpP
eI/Uaa+3KQfrPFUQT1/5Uar33j6Fsn/l40rNIyE0KcGqrGNb2jmsWh3mFsWjv6O7
oJwzr1GNDTCYEo1QzNsyhJS5BQhwurTYMgkQQnFX4YGhJNdshLBtPPiuvAdzgSn1
jko5XqCkZpJI17U+VMtDHPxMs7DPpx6/1i53YxAyKnlcFUfSpyc5O+ggzJsOIzm7
9hO207L3e860YtJ+Ec9MnIcAtPgQqm4DvtpCoiZCQg6lVbshJV2jmF9aUXZxXVU4
r0/ewiuqJkp64O4w+YOwBqsMDEoSuF9FmL6sD1kDDC4WZzTl2Rhdv6qjfSvoIPx7
m5qu5ytvjVSAC2pHNUsSgFI7aqw7s9vljGiqAsvHZKj1AWCto7B+9eyi+Y/KJyyH
ucLhlZHKsPvBCKMjMEn2GyTDDtftwep7/rWx3+luVu47WyPesdEZWggYAl4opDCA
CsqAssB47cIpO2N6oQqEyld8bRQ7uBeFLLqZushe2bucPQj+fh7eRRmaAizpVVw3
SCFijO+bHU/7Upi+bPHJPxL0fNWJ3hVBbaTkao5Hceu5d9C/30qHXgps6oQI+Ul4
HwXGaor1H1SqalLPM07mvIkjBIiT35g0FAgqZ1Pfdi3aRPpF95k+43y4HolxcMYY
4xsagv2wC5/Z7iwtcJZQ2YzLPVY8ND4yiVme2RjkKoJfl1gzQeJsqipCpmPQWIXx
VtDkxZhJqKCzQVdy5E1gmTrD33VhsXl7PzvOaL1j2qx0DdoVGbjIQjoNd01Imcn+
O30ucp6WmDVWJmlfrKCuvdX/qBdAPJjemFjFSNcSCC2tgwpLFVSn7eipcxOGP/k8
UiD1Dd+Msedx7tI5flKOmoVYX6etxNeoiiLJFBx+BJCryTL5lWC5qFNPBwIMwg77
5lM9EYSLQ6oyBq1ybkM+iozYcPVaI0V223ist+lc+ZAKA9O17/BKiXP4QNYIUPWJ
+TfNtlU5YRSq3OilaWo/7oNN0qU6Mu1gVvdMwrqJlkgQebWqJuYCKWjaf+8LJvGa
/esGGbAft9bwMRubNIO2cwXSCwTs3OlacAdyuVkFcm/6+OCqLJtwpV1A5sCfIP6l
M5HEgDmfmlN62Gx2k5m1hSsfiri5BzQyD2htRjZmC/Udo/LemoeaO065IKN05Glo
WEUYZZNiR/Xeo88K4EUJYK16PabjOOjijEWa5Gw52ebHLx0OBL9DSdBHlOHvMVLi
77GqSoLWETMzwsCmzD90wJsFLRyrWBtnoAhTYApiLYIWOUXDJDzX1IQozpiW7UQf
5qiTWS88Gc0rqhx0gY8Mq4/zhlLKlqefCNEYi4gLDgVrNyZT3R9Kj2x2UEIA+8F6
o668mHup7fXFkDOI/+4rtbNkW/MlTPYAN3Q68r+5nkR3AIQ8le1dIYJmsBpG+wBY
uJh5/lgnYPCycWNxysQbwDVOMt5eqyHE0LKd/lLaykOx2T/opV8OGnchTcSxe8+x
rO+g3NSJzp0cgsr3GlKV/2YNyLcMtFG8VZmtE5fT2hulu+Lb2NXhp9LmKYhi0Abo
EbOJlpWxDlKm5Bydc6rHWqI3svkYwB+Z6fjIc7j9WlqI9zg6KFh+6vuAFtgfwtsB
jVyWaqhi+VyikFJkjvQm19DYZe2rnqg33WRDw0UWV6L9SPvprtnDc8FJ2WsyhZwB
6DLY5+umNvI4YVJeKe1QQrhCx6TWq0Bz8pmkBzU0ENWI6kLgB8WP2w7CQjObsbFO
RNSTSQ77L2VNnGyZbO8h6E7xY3sRQSa6TIxtYpjQIJGyfeK41rQz9MkAW7qW47wa
Rm4z31Ht6JMhiB0jbTJ/iBByhBioRzLCxy3BhXsX1vSpHdl41DWIxMwNo6BROHWQ
2xDUfwECIu7x8FcaPPRfgPIn+YnzkWaI7T9cLy9bGUbS3qTkVlzssLCPKKq+pscc
X6wYtV4fQRUvVap0iFAxCLP6n+Z/uPRZlpgHCo8zL7wUyuxSQGHqCr4VPVMuCeh3
TlFE7iyml4ch17tiDU+pG7/NonYrdg1l8Lkz48xedVozXy3kD0KIn0Ibe1LeECr/
7SLB3OmEVvLAYXFf5dBSeN9xJ01T+hAfX+wOsI19GGSl9HpMNuq+1/u2VDUX9BWH
MGW6dr3JFSGJNILQtTrqgoe9UdjEuVoZFEhZQ/L7PRMx0bRcZ/Er5bGB/AcGpjeP
NoWbhVtFR2yj8KMrlhqiKICC/wPyJgTimFCxIq7fx332l8aNPFTp/GietugGZqVr
gyVlyfeIsKhJoU4vv8gJvHIfXiQ3unU3BzuyycifDbuZNqJvGH9d8Zvuie8/aNOa
2kDHuQjHoY+8FhZLv45vBpRemMpkwzwnbx3hKDqBSu4M6DGDHu6mpyID/HfG5xK6
ulHc381Mib5SEse1Yk1jOmyZdfOT6ncDGsyrsWbYdcnaaphERPwzsm1JcV1kclAD
fI5Egqr04SD8nvu5jYyUHLEVYOiCJdlqsHZA34h/9+JFuXnKxSvLMOK8dXPKX4XG
grAK6FdhzBuR2zZM7/O5GN1gVAu+rxfySaY9UWRH9BwJ4X1D/RRh/9G2rrpnFrSB
raG1T/bV7gI1pTbmYTVZUP7I74MdjkMSbbSSIE8ykRyRzes9HVtGf62YQo5xoMKc
lIUn2KrOzhRK84L7WXNtdk81BtlnI3vJ1r7TsV+3rOQKkXcHGrhRT/bN+1xF5I8q
Uuq6Tx6iPRykJe7bQEr8QS/VwmHeMzOVT5crJELLVWxCWYZb5DIdDKVpDG7ys+zK
kBVyFfErDbDEaBRhy0B8xQl/rA+cLkQKCcIDJEAbHz5QbcP8eMLNdaAWuDAJAv6s
runcNYZLb4I3XswCvTo/9ozgD8v24GDp5uy3nJHyZcfQJAHEb33KHWfTGAS1cMIZ
75D+k1p7xdhs5WTkg1qWrj3j/PMWdYCf2KQNEMoM3POV8o56WB68UG4WFUy1FXxU
CpUiWy7ug3x7JX/pASsgtQGEARPK2hnqYpt2s1jtmggns0WD7eNqHyrmNW0G1XWk
hUcoQ7b5xTUvgW0eH70sIxqoyZBRDkxPybqA3Ecb/AKD7nfrWblVI0bfXtVRWVmD
EtNPSSl4stbiOIg3L3hjwr17xcc8sTi94ovkqoeba+G+RFbkAbYeSjzmq3zm533J
39HYe7jeOEFD7/xyoqqwLRaF7hgi4Rs5rVPn4AlihTScxx6WzqaBr7tGFbD1V7qg
JoBlvOVSGYw5NurYDBCFZI6RRMXVv3aq9X4ziwcoc/U5zNB8iS2XcGhvQHvMT8He
yQTVj3mZDPf5oQbvOm897Z7FwaQewinCbsVMdH5i4jK36aE6Y99bZX++y/bs3g6I
8zOE9eShArUAnpnP29li+8oWNsVD5o89l0UsDOSMkDdI1N3wFOqb6aeFpMGRsv0c
5ot40dnH83RrQ8/N8dPNAbzJeZ8NNVwgR7u+fC5oz8uc5Bu/DnzwyDXjnQrIfMDk
XibR+Rj1zZHem1yrQ0M3EmDTrm3H/qh08ibUNBblY2BNvSn7z9GTKBY6sHmfYuDH
Q0Fhq875oLZr25jcz3yluKyqU3OHIUgFTI0HcrlRfV4SJJAXeAtW1OojxQ2vC1+1
gfA4c7WivbfMWNH6+QvBv6U99gO+UiH3ulB9AJyl6QqlVo7+He699pQjI2GCZB3k
opJ4BbXyegZZjoY9LA3Ksjxw9hJZEb16dI3zFHsUFzyRU/QonPRaHu8QGuy/ED6U
IZ3sIHmiWBKfI6BLned4+i+3RpvZOKa2YCV+ZregUOZYFO8i9P/aod2UmmQtFYN5
gPnVO/CfwZmVpJ7zTUmzi1uidDt0PHKuS97yW0QABNMx9WQQMMneUhbFTyimYf43
0IZETZ1mDEfrx/nQLyX5HZFaHSNQ/wHlplty8foAJwT5lvrnsM37An0mUsOzzLFf
XLzCEtE2zmPx0KzHCNu8L8EtM6eYBdz9Wn6URTRIv/Xn9tG17Bij/827STt65qhb
Hyg/r5QBBFsziCJ850QQ9a6y21bqnfF9EaDKaN6ap7eo419RO2YOtwqcNpXzQGtb
T5e4Dc7+jMXg8JeR1a3wEKg1vNKdWf5cMZeaqZWjHOo71B2Ycop90UxW5LspL1Rs
l/FFIufX6q48juCcaUv4Kx0Kg2pmTL5S7nHqAmXbhe9sI6CS5VKB+N61c6na0CVG
7cWzU3L3xqfdfJtLdYfO0QFSkwncwpGMIPO0EpBWHGCIBRNxyVHg8MC0c0XZtWu5
mHSKFhWEn3RUYN4NOv5t4D8nodpS+kAxH8wS9PxR7vsO2JwEV959qtMqjC9qAmBD
jtQbyobyJUDbojJo2X372pF6gf/5Yf2cI57LW4vYFwted/xpZdiWyh1951VE9iR6
8wMWPhOSQjuQdzB2yEitfOYlOXDgq89UOcTsq1Baa6fMS9rPBbsKte6UExEiXuqG
KO6jtLZEBlh95osu9si96LbSkUwugulwvLxwI3fNzMTBUVrq+OZQquQI+HO+OQoT
iz5GigQn2NSHmXtwn1JoruVruCWxnfTmwZU73x4peQaGHaW4C3Xid+RE+b6JaEz8
PvXuL3ZL1YDwkaIK5rWf8G8g2+RaUXjo4XcoQ8nu+JepGABcpEUJSYDVx/J6YNfR
cud1LIQ6EMJLhd0GFiNrarTU9YZSYuEKWOdPtxJTDruR7T/iOlx1VQMjxRzzRHKx
X8s79qsyzdqESSU9a/T3YpYquWXJPDhJnlbTGAUqFh4N4tFxTw2SyDwc/JAlTWok
SpnDp6gxkdVc4/eMzu3G16LgBcTaY7e3pbyG5mHOpC98TBIWgjFOLdJpxV3H1x9i
f/cVd5vSI+lRVHfO1bFFIy88G89g4XCiop1CfybJvUxXMfTOLg3D1vmph5XTpdxs
wR4rYy8hSOfjAkaStD39gBh7wbzZ9KN5M3q9jDZ4KP77zWY3uG6Ezj0+XTUI3A1c
fGyxV+z3DKiQ6Jgg7WIuzb68UMPR7CAeMLBL6hpYk6ncyiaw3NEssTLt90bvBlRx
D8J2HFJ/3cXfGNvxHu2NUTckfrVP6IcwwF55L4qU+3kAxLLDQtF8PoPgAerMK1sx
QOHELtVm+zhmV7Y2X/xbATlmM35oTDMVwlcnLWb3y0oprBAfDd3Vrx8mCTxYnSov
Jm17J7p5a/cqMvKDMeJJqpHhDp36XGynNsbaDPcMBCXoUi/3ojl6GzWD84J4sqKq
V0AZ8gxYYDLdbif41cxtI4nmPCLvQjSZt6IL//S77BP5XcIV6AjuKxpmdWTW/bUq
EkV4ZS3vQiutwqzmI70kjEs9kO3dZv1Sb5uxo3LU1qYQcg5PcefCMuqECWlR4Blp
Cj0Kc8HvD7H3U1ubh9j3cGyiAJtvNLUjXaisLujcYWd2N73hcjTX3YQbPg0pc4lM
ih5K5jwhtr/VEH+lSssIotzKxQxf6QaaCySHvPNxJjG4G+0uEePfhevM/tL9gBFW
4TY4p+JxkbGVLloubGTkv6LyLbXYtMJVQsELuteZMda2MuadhcuUPhRkF8IFZrwy
/UxPAI8pVVVi6RZwFzkKRBWYuU724pHjdy8r6DwTyjEnU2fKaNLQFAgrBBZl2QEH
p1ptYcxUfQ7tvLThiPNLCD88oPcR+F+lHmzrUMTPsLU0nQXmdinAv8AE3Sqrk4UJ
bAM0k+ITIQf/7kGiU/sxS/L1PC3UYe7ohd2w3ErbWA6ipkdkTyC+spVL4P96ACRO
fRE85/ZuRWJtqJj/NhaTRw/lOUJVUrrBB/2N4Qxu+eEYzbzSySe1jtFF2ri7wy/c
i+XOy7t21m9k1O5h2pNvgaLgSPpYjn7CQ52yRkRfyvPBS6yeXbBaRD+O7eI7yDcG
rf1YbG91A/NMDLviVYo9c/Qz67z7hnPtaowxo4W0lLM+uuStY1MOU132CIiINz+R
s2FDOjfx0WzkSqiaiyGf/xj5LifN6vYJ8S8179yFlpz9ne4P9Yk8MhiMFguMrPXU
Y0u+Vej2zfQw5hIiDigKyl2z/KGUqbZ+a9xm48hU6E8mtmh5xqEVcHv1b003Yy9m
+NEMoSjq06WBSu0c6uf6ezkL0Gujga6YEDuuJTmZfL/DG98TMAlEQJnP9BrmbVzL
Qd2UZd0K1J24JSNmsm5hnPxo8TIo8xO4eqF1EILT+10BXTBcIr73nThNVk6vYbHa
YN/7/qwcccswKpNPn34Z+zyKmU64w7t8HkBARvTQUOxNssMXDCocinTQCXMqGH/a
fMWkrHfWbRZ5qNeFK9MPKn9JSVlxhRw2jhf/gvLZULjDocnDr7Xg/Hkb7HheZuia
MazmW69Bhr3wCF/pKaCZmOwrVhqBrSsSY6wuvYrWTYei1dyvzT3bnoaKAPLZWa9s
plrG5SgRcBTYnpj6kwXyzEI9kSxeQUaTov56nyRrUsuulJ8frInPS/cewuZIQNme
K/GalSB2PgsNzQi1a6CznQtXQv+RKeWjC1RWv+RRwcClJBSf1ZGMiDJjmNYPh23F
3a/2Hy5Dz8SvheUCvTrsYhahIExywACn238br4dNT94mBQ/Xj7w3+gZL+oWyoF1g
3lABg59GR83h33iwHomBRXo3IK9q9uOnv78zSRUkbyldIbSALSWHvo6w8WhI1mo7
eplxbmTfpUKh2UKqg3Y8dIo9widfyZ6QUVK4q0OgQkCF8sSMsdtyLgg8ZM0LvilO
0V+rnnBX5KPVQZDiqO1VK3zzeKJnsD6dgeSfEvWX/tVKcj8HwsqSnidNqtv9z9/j
7Jyw2AdlGpSvMltRu8d/SAEcsJqM+KO8iOSiT2VnK+rQlvQpar6rnztmPMoCsBoS
VlOUtcYGlCXI89TsM/GpTfov1Ah0UkAGeSaPU5B4ZPHDwIGDcnCg+K5KnTFlKv2D
b5Y4pwDxWGLvnH2m6xuCgYSTYO0FKM1fvx3HTqfxSLsnKrHSveHUze3worl0/8+v
ANVJygxlEdAt95Xvr+S2t+VEmFEFW1EG6cDKReR+dhyPR8K1gbMj+FIDP1+dINFy
arBdvp3mwxa3hOQEysH7wxBb7e8SAPIgNJeKvtgSJIgTo6U3igs3N5+kGPh5FkmK
JV26J0UX6rZsVs038Q0Gxx225xtX+AkC70unt4KyFcgaNBlglN94iBgW0ULBBsLJ
XGdgUMkI9lD108i7VR0nlIZ7nI3d05dFQT8qqLNvc7hMC9GowYk47sFYOdT4ejf4
72yAiUWr0mJB4q+Bsxg7eT0otIGqJ/YOQ24ayR4hoCeGMe1xVCmQdXI4QNYa22Gy
T5tnL1NLRGuz7JLRjgvaEcYHDjrKhvRIPmTq30usoxkaqfSUcOTjckjDah7+jC68
4o5F4hizak7AsbgllnzNg+Yd7Bw8t2ueXG+5U/A+v4UwipCGDGfXbWFlI5KRPU00
goa4LPq77SMjLP3+2N8emCwAsohP/g9js55YloHrYXDXrEdkj7YkoZ84xvXAvEiV
kvhZJPi4BlkEmZw9c33W26UF3s1dG7HN/khdu2UudVQLrGnlRZvHO9GjHMMBW5Ip
9qdfF/6ewADCEJNMH4CzVGKHBdEXEt2CFy15xgbl/6W5sioQvH/Iu7qutV7Ptq18
TxpzOvvwhrFksV5bfg/hL4f4CWOkmzvHzEUTbPC+alveKa4+HCKcA4F5UPmDeX14
oSisKA7VmKOfMp18WSbgu7uLHSPOHoGZ8GIVUsMg+aSfZ9ptCPF5q8Yka8sJh8cg
hTYRmXJv2USvHF/nPUJyP+LZO9tVNpeN6liBLe+iiXr11W9Ptshyv7nvhUhDtUH6
6zfD4P/KL19p1TgTcme4tRsh/WwYVflLPS0903HuGd4P1DGybT67EXue8TvGdcp4
8XzTeEDlB0gg64uOvzN/iwKsbJQz9bQJgxF9X4PNbZKxn4J/UBekGNNv0US1czZF
t0Qy51YusCKDvj0CFbnFOzrv22193oXgxge7PpKowgYJAhEHC86DWs6hFuTRpfuH
OoabbDJNUd/SE8LDwBKbULbxsKYIvvhXAIVvBcKwDkHhuAPMdAsJAaiu+e6XcXVf
P9Uyef/xuM4cJehkCiiAl70n/lPelXGqxSYb6Yov9uE1vAx+Hy2OhYaiG1qsZZFZ
FTeuMx0mnI9ZPBZcOQ4SBNYeunBRGDkatA2CM8OsStbmNy/aV+3lf63pZS0Dnfri
1bKmbAfkv6IHSmurgXPsFuQzzIkcPmnYWq7xee0jOoI6TnjxnWrpqUCOkOrjRkMS
2ttQnZf634x0giEm89chxPWIWjP94rooFmKiHpgE0CSxooUkrSNFaEypy/DZEqS9
Mlj8fTyFT2dfrePwf86gJEFjC5wOsh85cTEbwDUNPT4THEoMmabsChMn2FuFwQSi
gao0ene0sNYstGC0gGmMmMNYpUsElOsbo+Ub3xTuS0r5OjrVbaj6Kcuqv5G9p5y3
vem39pJTgjcdIJtSSodOpMkDp3N/k0jgC8JO+x2J3dE/kcI9F+MFDwfAs6ymA0DQ
yxLqr1AwwEUjWpXyFDQ/nkKZa1Y2QiHHilsRNMOY6sRiAUHDsZBMk3Gykkyew0FA
k8URops4e97t/yK+iaDnM3jhwG5zdzUc6OP7SF8hrAb+3IqSOB8gqlBXR2zB9SGI
eIdTr7BDv0A6U4ke4oHH2In012u6LLrAFMP7cN/C8RULg3Asc1ndGMaSCej54DH2
my2bRX5oUPuKk6m4jXwDZyxcyqRafV+1RFqQG4qk5YGkD8PNkDiX///2+3LY02WX
JPT7UWtvzo41iKx95EI44JSC66sg9n5nwmV66puk/kK5bwIdJ/QARcDnahY1ez8b
w0dk9XX7+8urtiioKHTsoarXtFOuvj5adT17kc06UsF/GaULEHocbwYcVIqfDdVr
apnGflRMP8PNPFly48kJnOZZRahEcdPeTHV7IfVQclRJmYFaxzF7yuSUsJa9bSy+
5WyNFPaCaB9wOhEJO50fq6DWhLy2+FF3DAB4ZbTmhVk6m23yO3857Lnhp0RRthN9
GsznXRgEYjUwsRYBZCRTsn9C+8BW+MtgZz4AbPUn1PXFM/NtrIpftf68IBUjR5T0
VjIdTtMJ3cocTqtgu7R0yPdxBkFrglP2mLNzi/D6F1zhnzXkCFk03az9OMb16ojP
4NyvtynUUhg47VFcegMKEtWQOcfP1k0WhN8hO+Wd+gOwhztpVeYd9bYBGD2R8Z68
oVS/floaFObC7z6CTsNxNlpS6r61M8ZoMC/5z60Hdch5eTd+UWIggFe1RilJBxog
ZMqf7YnC7lPZIG/YjJpeAnBdC4d27mQdBMrOWPnt6zFxNgtig7Cfv7w2muuw9QmO
Bf/chjS39r66Trnl8Hx4jEFcCClCmyBjRa+cYLWVgTQoRmqRjnL2U61kqqMADSPp
SwIARX1tgOy1tNTq3K09C/HUx1YHmBQWpWrGK90fEYAqqO8w3VmSU2D6vIlFDs9F
psO51kCaYBAlvfjEORsEXXZzmUGSgEFBCF5CyNaip+zWN0R4ZZJ+Cf3CXs/Gjobp
/cND11mDZvOcirjlK3WZ/eNFK5w3zFRYLxBFqGkBiQ5rCu8LKqg9mIYpYiOVK9pF
Nsn2fDFDRbLE4CZIIaYAk8LF9eeIgIxYZZiwoeHEgf9+O1DfT2vkVYZPI7M+TSbq
483G1cQ48MYbFEqUTlU/j7jG2jYn0spKR1NMeSHDv6ClILgIpMpkXZjATEX2itd5
QBhXEswmLPLE9wo44Rtg0SAUkjUpnk49nPuAxE6U8ICiC1LcPe3wVO2DSXFleqVh
smERU7oLhQ9hmqD1mfRhqbGixLujIsT86OkBx0fG+UmGdANwB6im2U1jKYb70lpZ
9vgzIaBlvp2j9GnWZh5aVeMbEs4ljUw4E+PCMVZ1BJH99ElYwap9/tRi16WsFXHU
uSRr3Hd5jxz6orgj/lTwoGc4CantoxR1m0arecrsEarUXSWl9Blxw9S3uHPNqfTg
jjuj2LzdzTY428xOWs9TIjeoEpJpSlhpnPo96xbo2O+adpvgkE+nPGFGsRuhfzGn
a1vgqlUrO+o6wASBL+rP2d6YbpR3zNDAhcLjfrEIwZ2yi2CORbpiaLicZnZDFiXc
Wvpx9QJCAdWxM57Ye7W9K7N03pf9uQ7zijCJHdrGSsFi86ss9thIO+f22/sNCgRI
4lqGuIDKdE8hCTE2zDj11X7UHRos1Pgp4ELDoTBfIWrbngIsC7lsWAvguItweE+Z
DgBBXgtpyEes/p7aS34fhR/5b5VvpyLSQt1sWpqo/J6UceNcD/wkKsMeU1EH9dY8
iE3QZlrJGYHGKIXOVU3k41wbn/whL62vZXuyVijQoPCJrAePE0KmwTARfqNm7tQi
1Ysn5P5mEFERuY+Oagr/afAc7lbF5+ODl26+6KmEgMmNkpLvtsw0nAZdSkPitshe
5hk7iaoISQsiedWoB9bCrZD7uT3RX7rsLnQgDKo98wQjlebnHADYSg53DY9ZgQt8
sAWfzxM3NidgGkdCsm869b1wdSv4NGHI3a85PlEKPm/3+DiJORe95ylYr6I+nInp
k36DIYKqjE33gsllSzgQ8CgVnhbj9C8iJjhIrAABepL/wCM79g7P3PXBewBBlVvM
ypEmFmYaHKV+yK7+XWWvKrxPkO+Z3JtZ+rrcQIiKPZSKecIyxlFg2oxwktRkLZhJ
CAWcusI+TepQKvKOnoXNyiLdJLPLp8VquLlnkdrosxtCA4jEwDxuH41SvEO2sc8h
DoeVVsFC7cX2ED0oEJ+cS31ZUsjBMWmKi/WtVByFm2C3SaJX4rAD/odpwOP/UmLl
P3nOCYQ+OFmvj0uRHedk3mYnpeYcJ2tAjsm18k0Fd3VgsB6KIXkCdZCE/9asoFjg
SzSrnBkDw4zhJ5eXqCKHARq2i3hi2YFxfY1tQ8h/IJrRBMTSw9Dw+Y5YCvVLsjLU
mWi2mRdlZ5ZMo/sC2r5rII4Ey74l4+uVrjU0NptHRFfMNTKVx+OmT2dNUkqmO/6s
B4MCkab7CPQjxUpdS8dbpV5XXmjN9dixQgwZTSDeT/LYhGe1JqJ9OFaMxuCH7aFb
PQRwMgvznLzsJvAVCMAnA1skiak2gtZOxa2haUryyTfA1XZ5Zvn3T2aQKKc6/7z9
PDqtGubo/JDWYc4iskXHK0WnJnEngYoJt14oEdjefc8taLAJz1F6VvKT6XVTayCW
1oFPdbYm/v12P5JAizXNrxN4xREccDomWg9jMAQqV320gqu0ZNXsA7C4HcEZDAXD
WeEdhM1/FEN5+InF8thSYd/ClHIFTfcWRqIXMd3LyqW7Txc+ueBAmDDvr18UTqzk
5z2rUUaSqRP0AiLhAgghTTjMi4jrZgsbIp7K0jfdFa/XVSVGSh1DBQzICwRHj3Ca
16941befQh9kgfOjcft30x+tZ+sjtssw9rO330TuBYGhk/K8WXrdVRTL4hkR7ttO
IoKNLBVzFXDVblk5kWqHbkcL2rOfbD5tRv3CbCpnYz7WJKhkj32kW2vImbp0I/qx
nmZ+dp/cecBWFTbUQ6Vn430IQz4fRffn/q5aOJnUxjLC5kivXAWjfFiBWGBuGI8T
VrhR/AjGvfAa2WYYF6hnhH1qNvufxMpWaigWKzvBdD1MtvNa2CaNgrOUaqe6Zuim
34Jtq+d5KSj5p0dFb4MebyMEh7f7lcKhukjTy99w98BvSYvlC0L1Mt8WtTA0Zt0x
tXGXcrAts+EB4S8o7qo6qO3QFQc66rESf1YxI/ki7sigYjfERDDwXoZvG8YMXn9w
71Mkb9O9aiw02Y4qn4ZCTO/iX0esncDq5TzsKIHeIV0aYzcQexZvfv+ZKRb8PkTX
AlDs6G1ULOC2wxarsIXD2dfKo5VYoVyzx9RQDN+PReccHYD2jUrTkxfzgloIvSy8
nD5mOZc9v0xVXk+qGd03r9vyi9sKJwa/pcCc25CAimGe08UgSiIFWO/SlRsHMdey
Ne6iaN1HgoflWrEvJPEBZBm10D+sL2yp3uhumglevhpxeqk2oSDRljEOSfjL0kCb
Vrq6Y3krcwtzEpQb62uZO0+tgPj2faXnmv7P63ihjtnaWZtnwlBX3DLTQ3iiyv/y
pBnfEutFkYbIDxD8CTwDid06ArG+WHhxa9xO56HV1d3VmjcHbBNLX8dfZq88urDu
qPbcVXHKl5lzCqS23v3Qfq6Rft6+CCFwHY9o4oQH0aw0JydsUEH832Vnc1Cz+yby
J05gPVUxJjjM7JZ/pLyW8gxgcIzPKjK/P08eH3BMWgAMcoYbm6M1336SmDlc2lkx
LlXb5et6Ft/QkbLI/r6TNDuT4nioAj4Sx9SuButuQ9weoVcOvz3ObYtvLxQCqW2r
QKYVpGIBtrd6eaOHq1rim+/AWeO9orxv+1jkHQQEs2Cfhw18OM6CziLtvOnf/I/Z
VifOxWOiY1H1Qk5xa5M/l9SrmANM6aQjPUIkA0mIhxgzTFEiNoz32UzsJPCp75rJ
TU5XTvM5RuihmbXsDUVgeucxOdSrGTpzjSFKsKRc/TlZt+AHcQ9ddBSOkjPeoNlJ
i7EzLHNI0JArTJJOo9ZTsDYVAFVKVooXxPBGeB/tABEBABFnBgAzAdGDcx143IJ6
JGCf+ZvFfNrK/4I4I6NyUzfNz+uyaWdRpfwIllGo3MRRjiosxyoGfbBjVazDiFNy
tDgLM0FghMR2BQF4bMhgXTrbYQPZ0FViOCDoN8eBEi2+0NCvonYHY5jXDMzaODin
uaQBy3ZEsHF1WByI6MvvmoRK/YdspXL7UIK4ejfNPuv8iCpKmKW2dfFIFjwXImMD
17MvOHPUe1F4aEqZBywq0JEzQiEsoLMHelG1oXOKK8IBF1FqOpDYAe8WYh+zP2WX
gr4ZaoHtOVz9r/UN1QKen9VsPKDOM1yBAnACWitxjVpajzuoXYJTqBlRGwpbM7l4
bakTMlQKva4er4nO5g7BY9OGlr39LSH6WzDxO5r1MasWwfiqiCuLyRJRYLjS7tpQ
JjUBUsuOsH0eV+KO5f9obZjZp8QtgnbYMbvbh6doe4oeYFdrsbYyhVtmQshDDDC6
0sSWXgAd5yUiKxNUFwd2ZUeD7yuv6Wk0vAqBSKia21ht2SXuM8WyZbb9tvrpsjKn
R8XMhrBSb/4DrhQ/ah1vsf4Zv3kf8UzxUoazSxVzOZxMzays+C47sSWAnW+Vo7Ce
UTlbRFl8SuCa9/6me16tiC9BMmaNGOtzDgyuxgd98FXmEvHy/TqIzZTJ06XDNW9F
bxSE0LmiX8bAd9Mciu5wNG9m8kS3DmSmWRLI3OBOxqKztqGMbn0sN5866uayR3Kv
1cewTf8ztSa4W8yfraffLiaoNtcC8AgmY46jW2xOYTgZHbAXk5oR4JnRAvUWMri6
iFwBAnvnNmTgifiQPQ9pYLyAAhvZnoFr9zvd13VwzPMS10uFDN3an/kkUVJuyxkM
jBrymMihmt4Y3eJ7ITHDoFQ1N8811bdm26HJCwVsoi6i5o3PF7uUYjg5x/VfKoYD
7rMg4pMYPres6CyOYsSMrRMlWxyRuvMibVehbGGa0CE8VK8ou5t6aJrsE3Fd/qCn
7Sq3mRgN6WNAEF/6z+S120c47aEPfQ6aukBSuS+FUijRDur2dnf1Sj+wSZi9kFIc
MzRrxQvbi8GfFL+dwapyjpE+vmvPHE0LcbY333LBwkgfc9JN5bbrNTCoPCvOA9Y6
I+BKxIs8nLLzg1PHKLJ6E0TAW4xHmxKBxeedgwoY1EMY0RjybQX5NCcDb3v4qkB4
U+Coz83v9+HOKtKrWfsXL6E+l1Mu5i9UO2BxhhJ5wnONpBQQeJJI4MKIDbvjy9ku
Y0oh8cKJyUZnUDDoWpJ2oYO18Cy++g4mFoi/0A0E66hh1Ru9m0TavVvsuAsRV5VR
qH/ByiFDMzkWt2Ta5DFSHdHkNHAe9MCIgUihbq9+B13ijU7ldJFotk7pO/xkHIml
Jd/jgn3I2uCNPt5fTYwE94/0gjJg+Xbd0Xfmy2g4FyyuFJ2qZDC6lpOzbDwXDmWJ
K8wri7S6oo9SPL5ZXkSGX1rJIe2MfCgj5WwVAsvMkB3U6BkUgT2kmaNgKxCjuz2t
QCYKJn0cw/3GhNariVDVPVhSxX/pLvxE9Wp2iR3ReEgnNSHNLEvLm61sohkvkUnf
Jgfd8qkWrpU38h6dO+F6sRTF1Gr5tnvsMuYwVaaaC2zPYBq3+eCmef/Uc9z7Cdb4
uFVfqdSH1w/7vSCAN5Vlsmh5hLmnguTaSdcwsIad1M02lRhuC/b4cP0kh2EoRJ8O
hRMfO5/0r53pINhcGHWB0rxn58KbJj1RWmxAdmZ2KZ5RvmEZi+sXoMnJ5QWPi6S0
8zpkhLRRMy3Dncrg2YJNnIYlhEzGoOCZm64U53i9a4FL+KK+aAB56XJ43kb7fztp
7KuL8ia2oKVhjMMlKf4CCyCuIf+m7agkLE/TctwvESnVqTS70bbdaXtkgxKTIo4L
+3psO8X7Rce3lt/I2m0OM4IcOnhISMDOplIfz33UowDamMYfYPaKtPOPKzGDJhI+
02/TvmXCnmTr3vwPmnO2T7w5uWVVBbDC7JDLhIzWgplxCVhzMY+J0tb1SYfUOZ/D
gxL1PKbW5W0kG5uXur72qmLb/M6+T4ZLzNQ7Cjz7HBxMdSWTuX41fvywX9wkdHKB
P7EqNOUt/JbqeEV+wL1UKqUj7Cz4IcGfBZ9L+mDoNpp70pOWb7010ylGknQy0Rne
QyNoUag2HpxphkUmyVxqr1y6INR9k0rGW5XJj5AwQOjSj4Dnzj5XMJTz2dOuFgzB
EG68FW2B9th3jIZJlaVSca+1PQWkhHRt6GeiC4KL3Qg2GSlVYXbSn8hDkfAJe950
wM4O1xS3FECqokkkKtF57aB9gwoUS8zJN1J/1AsCoH9+CK2j4UcnHFaSdMow64oj
WXHjMIeCJhNB9b3zG5daDbPF5l6OXnn1ml+DUsx7TQ0QbaGVqVdA9X9y8d0ltZ2P
/EOKHVDbaCYKGHiSYQV8vHEIR6Oes5VE9g5mbYGeAzv/anO6+HWrGpAmvY8GoEH0
uPFtKFGNfyHdsTs1yKoJ9+4aoas+qGq5QA7IL8GD4UCfmiPiYoy7g3kKtL9V+gSL
hAdTcVfSc6l0uCmr0SI5YsnJ6dbxGMsB7CXOknWjmB9a+NME9yrGVz7Tzb9BRkoU
NFvIDRSQ02vX71YfM5ZPUId1HSWbNGxMFbP1Eud3JH3UZG/GqsEqUZ4sjkdVxR9f
lCxDiGkqi/yuw7sNsW0hc0xzb8lSbe1aB0oD+vkdj3BTGhyVZMtGNQaSXiMmIWVl
HnnN5JfLOqlKAjOF5BMrpJMkvQr3eAOuTMGKNlEQVF4VjQjcOwiB4gQ5i1+Nuxq3
IgrFCMGf5k8nJaIxhAcWzi4wmypTTGo+FlpUYzPQLZNrZn+QCLQSErBvJckytwrY
EAyDNd9OXefbE34Wm/xoNr0Aky777aDvv605CquzcTcN7YANDcwpRM8a8kfsQNx9
9jdV5sRDWTkMVsFAhCsq7JZ1vVlwB/JYJs/L/sPOv1n8yhfAFR1YKqVKBl8szPgm
6smCzi4S9lHnMJkkbczSJCzab8uU956DUHlnJKyBycvuZGxJJD1y2P2ydWXR9EWF
Kf5E1w7DCeh2YI8+4RWEGqJmPEevoW5hc7eOK21GH9A3XOPm/uqjLodT9EBhnE2X
lsdAI4con8cEsgxCt+ZMUON/j/QqRsgA79cHHuurKW4HHJRrlHKtZmwMoVfSGy+N
X7A5sAbX6dQzdkeP1hb2MxMGBWZSLFkAHOJZ5YjdbINzXDbXhvoz0C/CSYMmefne
2hiYu3d2bSGo4W7zmDuAlG0JkwrVaoBVfczm3IIw0BT8OUGjqLMBnn8ZJ0XR7D4Y
CL3L6yiAgjGw6UN+SWn+sfp/IaE+abjtWxXU349p31qRlFaeuitFb5gquTpNXfr2
k54GSocRLIQnNISEFvlvk8p5z9CVCI+zKlBxePj8CeLCsk08m7Exp+bLk8n4pT7F
Tb4cLs9iagXFTjIZLBZVqUqaTbl74RgMow7kE9JbPWLYtJsRvNx3hEg3Z1zXeGw+
MDCwu6sCA6WlQdk7Xg8UAtBUJQEGEWywCzshdMI4TbsOHW8GPkxq3aA+x22eY9TG
tsbM+aSEN4HPSyVg9B+Z1qvNPNs9vNJ58cmYXIqoXcx+qvUl7dESlAyGY3FmiI7S
qaSmNmJooV4thHItkyLCR8AZMDnc/C4S4v6Y3kdDOezzao27/hctNx7gSv7C8801
JXotg1jisQDuijBr46orQv+KjroK32+XiQqPUvS2Wa53cjYLhgnHRuYtzvATj4vG
IgFjhOPnjQ/X2+R2JMqyM2efyKwkPfA6Uq4e3Q+Iondt24CwZ5Vgm9SDw2PwPRkO
1gvBsZ2EQWZ5daX6xjeGOe2fs3qCwCbGShoPVXQD6x6kRstU0X1JF61kuCXoIdhP
aHMYJeB8sZURVPOSqtPkfIGNFo2NCYM0QHs/W9vTVyT+bJm9mpFpnqj/HX5ZBJ2f
ZExsf1TAlYgOXrtqxP399KXZ6lD146myoz27xBWVppGCG4c/GCva5KEOhqC5gz+L
utTBq0RNcAHT0M6vOFMEklq//nxsFWhNMiivEfpbX37dDXkLXeildntH/Tt5pAXd
9NxAyokCFKqk3HmRqJYkT6K0d8RMK6A9CBh/CC2oWAxinY4S9+SCafxXEki4lgFd
JdReMGNH8Kvz1xKg0t5jaNsqG280XaS0VvxjThvtaQ6ZbpxxdXft+HczzOYi91f2
vxg3w6+oeZoXKlbC9Aj8Y1kk82xJRa3LeKkZlhevRYt3OnKdW0o0i6c9Cl2BD19X
8POFYNaO0NTPBW56CDcmb60rU795t28LhecpUHIJhyvk/yL5p1NmJw48/T6cugvB
S9FmqxLdN5GWzLWtONsxC3lBdu5CCbRFilX0Nqc4YFP1WHZSCN7P/BK9AnU7XZld
qGp/Yar5bxD3Iqm07LqhuO7W8OFrmOQAPyYo45gdlo+StgwLuxmyxCWAxj5QEJuv
YYAC/NvjmAHL0bQ/Apn+OqXNH4KWezDDZTDvl8EPeGbxns2S9V+nVWoMj+pp1KKI
5r21pPkXoiAOongPUEklIHbINMI4g9b4Uz2xNOtxYv6Y/V0+Itvr2hxGfrAi9Vgb
W7vj6bW720Q8bIZHfKqQix7UwbJIx7lIF7XgpuqEuC25lWz63pYFHfX7PoZBEKLY
4pIR7X30VOVAs5OvTf5qJu4NOZCvNqF0OWn8RvKzflpaRMaV7AQrj7GUkNjxjfml
A/+9N6QwlXYijosEpCMWNTw+QcjFkZTzHiprF/sz57SLg28v6isfgcPceDS8P6No
JeFTrsl79SLQLaFCIcoyIhxXIKLDSUnIYB+tIzteAJGUXIeWhRyZpGoAxBjFrdBF
A1DiGwwFsOfcWpoDOjPPKNzKhAHFr9S1FDrmX7EyWV6+WWR6wXuHltE5k7V3nraq
vJyKUB0YF0n0NfmGsAcfTZLdJGq7bdr/JMHE0/3GIxSBn//I0tApDrc1ui1R5YPI
ohGCfcdeN8yPU3VpI8APihegwudWaWg6VW5PLTt4sbS/GW6irzrZou6ahWMZShZr
cWZXIuZ9wNVJQsogxl3KsJw2bH6ryWifkA//2OnNO0v6b29k8ntyzC7QKsUyMAY3
giLnomidOADeWmT3lhJh51XTiW9NCrZ7oDFpiiiuO+8cQ1iWycpETMoTz9YauFon
cZn4oh7cY24+ZM4B3/Rgx6zr9WWPLkX9+lxWcSRohYgXECOevq4riqiXgG4sZoc3
uQwoqb1t7qfYdeIAqhPNzVnq31rdU4wWOvypkRki/TXLo4YxqSmghjAofAd6s771
urnH25iLv9ExJV6sk2vltwwBx15DuHxliIF1j4+OUbPwZX2ZeUy4ZMarZd+XbMvT
cbKKu4m8tPl/7lpwFP1MzTsu3IeSKLnaQwndnq6DAItMe21wfj/gVrEoX6IxRbPL
Fw2BJ7SOrFdSEGGIOF2lgFp/bK27ika48kzeov6rqFJ3JAgdGXSOcXg6OK/V0pwU
W+kGoEq8aZOJ4hxGfApCZ5ewb5Kr4eUUa/Db1gYlLqHZEvU0iEtpkgl3w+Dh6Lq+
gSOCLhafqUOUlNlN5RDY6U3mwCX5Pmi69Btzr3nnEfr8ivV4zp6ZuDeXXcAGgmwb
y/dyRlpreBR6QKkodEVerjaA3d4DJsyyx0mUJrqxezVqUSYVPAErum8zcFezg9AV
cTY5yJ6dXWTs4XUV9k3Ncq59/Iik+2TrzNFeRCkjPvYYCeO7EBww+3mnsIcXmR0T
ANMINsN83tVHvB+QfkwfK5Q6G7TSX6f9NQ+6EfKwVbWMsmxwDwpF1OG9L9BZ8lHk
66NlGL22iefo27Xm7myH4FA5bh08xt/yf3iaWC02erahVCyTqBpvsN09WTxDxRPh
Y6ujI3zsh6qTuOwV7y8wjA3h/NtmcnArrm9bl70FNJI8EsCdCkwU8Eeh5tcjmlW9
g2xfTN1qBmoJ5VmNDEwY9Y3GpMOBKruDrX4isvTR9+1a8eACMQDcJdnKeham+DMH
yDHOrAgJqooI6LJG9jOoKUBvnX9orX78tUPxfmyk6iXu62u0n3/m1QJceKxW3OQX
lNKg4ecxigNijMvL2clIu3aAk6nDJcuPel1YaFjRv+IukUYKGjnzngxfoogwH5pc
iVoLSAwwMQVxEsD1R2bjiuhOc93/8wPD/8eomgMDUEXNLFvWz7tKMQPS9Vi5a4z/
fToqdayLknr09V9nnAAy4DWlL5XBai1NiEe/w7k4LST/eOP20xc6yDnR3Vv8eMsj
YbMeIWFERZGQhwO/uqFuPy7Ln0mdM9eNImmb4fXHESPUhQAbjmJwlDNY7WwyBLDG
YS98QJCn34U7hTqhVIQVndwJGaWG8jvIS9N8z+mFyPdRRTohiwZcwfT5ihJeYj7a
brnd5yOfatTofzotDVYHIkdL44Bh7E6yarSOxy5e3nnoJjj7DB0L9rXa/y46wtpJ
h5bMivnluc84auB+zAA34vkN60NpPNS7YdP25cNgMxH+3YCWZPBHcEgRikBTIWSC
kRkbnKOCtvB2MFiJWyzqTBMXV4e7P307QJDqYwy5niN0QJcJ4QxpnI3QfdBuWA7R
ow6ZN0hW28th3gr1FXb/k6XX0bW4ZY0L4W2f7OGko7pNIIkeGC6OvmwuqeFcyrZr
8KqzrHKHXBsAbz8MthL0U/Y19Gcy4HqMQwvezGMHr5846xtj7KRZr/6P+Z+ltevx
hg6ZtYcAYh1QKNpPVfrS91zY3aE8gjIM9EvQUHLsISnQyWN8deGz2U8+y+pwRHd6
qGH3OEJY93iGO/libPFGXPJiJRe9RoW39aPiMR6qxIa4iKxauA2DqPl3wXW7c/Q/
pOmvIk4J1WhdRINiBXZ7pwq1QllTl7yyYFuF8OuX45hzz6nwzcHT6iTp6dFelYjJ
5trgjVsVpH+9EHo7S7wvVA3EzR8fFSO1/XDALg52H5ZczX4qERBPDr5ZR+EMxKfY
a28kyEVGby8ucOOK/AEBjViopZ1/Oa0Mv+xm3JuGHVFfUtsoWEnXMqrwzUpadBn4
kpCzW19+WF3gKGHbSyy7t7K3qwTEBOHuI1VNUr1/s+DbCfqROw0SQdgK2w9Y2X2X
85RQ6G/FXAK6dFQsCVmPXRiZc512PIK8Rk58M5ETfU2mYmiVuw20V8GbsuyJFuUk
EH/0BK4N23s0lGioZhP/1g1J9p7gHwnnOZwrKiugYqfSyBJ9dDA9ne/M6cW8QQxR
XTqHsb0Pxx43A4KN9IdnB1CUx0HLebWSQO8UmWm2sgNtbrJlZ1zx38tCm1nU7IGl
GANbKpQwSXxr7BZoNZnJT7BVMHbmmdA7OgJF88A5l0KVdY21MK/ifQPHAGkd/L10
soEDYW+qDp1RFWu+aVy1gejXXGhBp7ySgVUDGSjh88gpjNfQ40tD+hmjmW4jkA6D
wWKGekzmCJ1m9+Us9pJm3Hfvtvi389ju4PXX3dDX74PjQI13zkKTOfxSu+Xyst6n
uimgp8TxVBV4+Xep199UBkNaHlQw/su+xV/B1+t5YIiBAPzhFJnwTnxlK+ickzka
8O2SQne9SEcbLHIZr4lVTwvvQjnpLP3PbBfVkRdJnGJopTesVF+ynoiXzyoND9Jn
Yxsal6IePeaStVB0h7uw0sdY6EEs/bDKIuU3YIHbN9qovD64xf6wOexkqKSZaBhH
CE5SN10ae0D51z2GSiJ+Jmc0bozqG+IwYLlA+y6Beu+Ec5HHTOeD1VnHk737T69a
z+TflsWY3dKlZGUnxmeuyPK3dYieIwXlWqZPQMnpeEGeQ0+9oOzzzDedVESD91P2
vaWfjJiVirrq6W7bJ7184NUH2kQXYdp5JgllV+qvz4+JVctP1JGb/VNQF/PRaehl
2+rpfpeEwdKfJz9yz7YMKoUClzSZHQuZaCeTTxDhXoQOhnKhhcjAWvNRz9g+jt6h
OE22HdR9obc6DSp8XuTtkx7kORGe+MAqZe32Bg4rtkcouRTMDN5BFpyg1PThG0I2
0gMF1U3+P+gWdGQDy3T+nKGwgnRfAZ6xbtrD2OFWj7PUUwxQIDR20wZRNzEa2KlG
6sR8OekGGBgW6CpXOCD1ApteaQZxYE+P3aLSINNDT9ZD8DjmS4W9kVtptw3DzwCA
7vx5pH0HudcMkNwiPSULeHL7F0/Swmc9/9sIPTajMdm05BRpoaWTCcmFWJHORTjR
QlOxfCB2py5W8WfeptSzDi0jYq3nqXPUK0Y6CFz/dO8vO7kTt6nz+GiSOCp5h4/I
egxeFAnTG8vEF7oC5tjblYnZQlC+BDA05Nc/bjediVgVhlm2PmOGX4UwBjJgpZ8A
uSotx6Lb9pojC0nvbq99Lh9ofUYZfz0siuFiKaxbrg4LX1k8AcFDchbqzyaHjE9A
PEv/lxEIXRnCIzumPD9cS+v/RTNSOBumBIHrYdcS4HAnVvjW9BDx7HjGG5BpSyZj
8zegEbqzDk9Fjtx8t87jbClkF3/c/dwDqUlRzQA99tqv6oR2RGEAX+5WHe5tBzaH
dXHgXpQG9RSeRWh4WdBkx+a/MkbmIACsXURznfDeGNHlV9Y1jUBP7NscVAHzEH7d
PK4GBLwIJKpGEh/ktu44pvKe8r1QiR3d+WWcqANMzV+KUb4DQtr8Rif4h6A1v3pp
D9xVNaAP6yfI6uuezYKYIf9XThiOnkB+ZzRNl5up7jxfM/xft6D47qQhM2iBVgEj
CgwMe11FwpIZ+S1i/Va24zslF8idfb/4a1tWR4oKOJXQtN3LoeMSWYuAUQcCZM/e
QCjeR2RRsafReWW7kmrAh+ir7s8AGdwfWI//2c1pddbW/P7tqSqefoFx3HsE37Ta
hKfc3A/a2LwJLcO503NtQchcstC7enRZnIq/ggIX5hd17MBXuo/5BdSZZXHcjq00
MaoQHi7EzMjeUSzj8LdimjaBBtzlHRL+HEehZ/sumhRpX3B71yVHPpG0WR+E1P7U
J5khhmMdFH+RrvMh/b5ULbaPnHSQLTnzwYqXSXfgtcOeAOENTdTWYVlPKpHg8q7G
eVG35bTaMMQZQ7qt1GqNxMFecseNBRBvJwdc2rMp/TbekkD856O+T4KsodL0BxWS
Z0DRxy5aBy2MKNRXikB1mVPn0FLUXDLMcS01W2VA7xWcNYfjWso/9ct6ZITytAQx
xUMXYafyeOyTfejsYOLqa6kgchJ0n1Eld5Gamg4IopbxgZLFku7UUIV5VadB5PVJ
v4JNAozEFh5aCUfVAYg33sILKvvITVXv2ZfJ3Xu28Ufe9vbZSFEh53QfY0MppddI
77SPcVhdoOqLExwe+XIgWVO+nd3/W9Nd/IDKSPexArI/FX4/qygR/8tEtj77UWQ3
8KlVpwsvUusdkcLdipp+InxOqWLYazCGyuHtV2clBAkkW0W0ZbiyZuhvLVxK/F4r
TjmGUUW3x6auvqYg+g5qOG+QYzoKjDyHkxk7YHz0varZxQ4i4btCNYmoqRi2U+Sx
VjBOuvs5Jc9IgQFUPB8TRtAkmSmZqLKneASrdol2Iq8XyawNIihaslkgYKc5+5re
aXkzo+TruEznsLx7Whjsg1zBmxd+Et2H/H6KT6BEEX2yIYv/sWpPrsqJT5zX1B4C
VyKU+aW/YzZ8q9UU3cYA+XDV4yqmkhpEFZJcE5zHKlFz8qnLhdhTm0X+zQgU71X4
utmFcl0Jy86JxhpkCUT9WYjvNKQ6Qhg4h9QH8LHIcAhhIf0D1+OqjzrClnU+6wMb
OjXi5cpHJ9Q8CwZhu/9j0Yw75CfGGRnA8jW8XPjU1HBLnwbC+KaHvK1LoxWWPf2Z
ymRHfKhClpk1Eye4w6yr7AjFs2qtZYOq+Up6BjP+0oXUZKVLUBtRf4Hdrl08cbrh
Aw+cYBKA2EcVgMdqxrwn6j9onBIZ3LquD3MPtu2mZI9yulSXyl2YKHfy/C4vNasi
b9DT2/ZRZy4VgeJGpDz7wDPo0TeNxIT8SC1705xumcKHSicX3GoeX0jlQlAFL2dI
Abd8y3i1H2HCp2oPKB20QO+H5B7o6AYfGuqx6FEu4c5k8KlIV46MoN5dPgm4icch
VeUo4AS6qdAxZkFXAi42hDJ38AfQLf1RK1ehfA2yWjqObHl2XQDnVrXZ8oyc1qEU
ky303hTh+YnMgddtNCnlm7O//A6+rvmjL2XGDeaZAGx5Nfoh5OnRJ2ycAYuRtNdt
etWQngXz8rmU54kW2akN2ZsZFqbXgZMGghJtp+Sfh401EOyDNjObJJz06hDpA3E/
vGP+F6sD1qEpCyBDQ5YSodGRMY0GyK/H9U5GBYqH06CvRoqs05OTP0ykrr5KMkE3
kgrWK3VIf2sXgVEq0A+RMDed0I2cFhikn16PyCLQjgyKtK5IYK23py/EURL6aIFj
IDH2nCm0izTln2OtRXF0zCvvRK+LCWxKSFF/ShlBuZQpswE0pUKxkh/FkicQTGDP
Mp4vEHJUS4kPKWiLgveYGSH2o6gA8kXbYUYNwbEE3akpPvp37ihU/yyPzBX3I11x
JSSJox52YPM5r/7fSW361DtihNVP4+5xfZ8wHp9fi1ufZHJjlHj07gAGnOOTL506
EIIvNswczF2RtlsGzYfcHVtr+Jy6BLvqCOApuK91cHCExJNK3K/zVo5ETHElfQ2c
TcGHX6gDHeH42CT338iLMuWZoa6BLgVj4P+HB4b6dZpi/aMQm7W/PFaob+GTSOVH
PzCBB4ehC2OSnZmuPzsDnv9QWYZqNnkcGkSevTHeLYhLN8thKW/k2fdMjPgGq8aL
EzvnIcKz6FIugXWsFCK/xBltvokRFQGEPlKH72QubmG69iMxUgmzmgzYE/KshC3U
NlYyBjZfTw808chw3w1C8a0RPBBExrcWPyuzjvdBzNrlZ0wxEIV0wV4qOCgAlPoH
YSGFnfLnFVncafJtCVpSIBpZ00Nc47EzNMidm/Pfffdi2eJakkpnF1O1+huH7Sts
p520W8/AFJnRYxFQjWZrHQQY5QTzLPmbbhG+KSe4MYQMA1qPnX4OsYQbbQvAZG/R
rBcHCgKOjBzVOr7+ide7EatFXbrPX4nS03gbGdzZy8S9twHfUWe/72LFWTCU430l
aqN+29no9xXn/og3gt8VEh/TvtLBwWmKZeoM8ILXK6Nx/5OgY0B0ByfwGrWoGw1Y
1VtTzy7KdWVC/YKehHW339VR6cSxodKzyY5TfCaLybF68+BWOD/7aBEgM5u/7biW
YaYNhNkdfif+KZ8JXMuz8w+oeqI0UujmWhypWalVoSxKnmcUQJWCTaWzR7SGojCU
M5nrw/OJuj41Vcl8NMhjowdYPgvZ4uRpzn34uUhiY9SSu9yyM+ZN/VTJ+8MaSXkw
69/4dG033A2dtDmAuLLXLpKrIzIW5RZw6/8MIt/UpDaNWdr1gFQy40k/Qdif+Bvb
wkZ827Qx/T8ZSfyY+lhVHJo7I1OUJnbR8U45FLrLbOEGZEYUhPg6Fwvin5K+P4X+
pa1ulYmbuU/q4CppOwOLFPybbUfgaHWvI1vymtj0Dp9kA7iSZd2VdqjQISLclpO3
Pmr9j4i1im7xGWh58l2+nUKdbbD3Z2Dk5cAhVIztsKlHhInYyNkh0sSsMkxjA18N
GWob+C01FxsbqFyQ+uJ2XfWDcTTsU//rSdLqL9gH3AAeKFqxFy6JJ7rIBls9A57w
Cb0vEXJ3xRd93zra5CQ2NTQ0+gcyYONI27Q1AjvY7aCFBsPJdEvbn0YYg38yqJ9W
jytC5VS7CHP1jP1G6QPLv1JZZWFfHWkdc+VjKHmq93/Bjdbgj66MSksWvNNObSJo
w+0kguuCJjj57iLUhlCJJItQku0bHJ9h2aI4/qMbDySzGypeYUxRdinb5MoTXzaL
hhd1v85KZIEWS7pT6n24lE832UV3NLBHvqeJ7PWAnbxU4FT3oBKgafl+eNU69Lzn
SnIFL/sbwln3yrhryR+6dMUvCaT899En3pIGoak+2USUQu2hUNvADuMcTug3IPAU
QR8RdprO+euxsU5Ot9RmSrArT/slzp4KClSc3wz+hGxrB0z/hpGg7qoUEsG6CLdg
24iFZzUC+cf5lkWztIj/qY1Qe9NVWg6oyz5DQyr0MUoPfP7zHjVMEYpML7uJJw7T
peGhTrp/q82mpwlpyF9Mcx7JlvPk4UVR5ZuKZHyLFfUGytL52eGC5lkg6LF7npRi
W2Phay8NRHWSmmt6QS9pTVkLnzCSY+fjB/01MCN6ZR2FaP+M/eOjyNMF4ciZ27eu
QO8nkwgDXGGl6yPcr0qYdyMtaz0D88QlUjLhFfghIoqq8pXOVNBWWZJTOjLpwE3c
5sAePsE6XlGkmHnTaDFCjprir4jW9wqqkqaKIgIYTy+k0//fR1o3orogIx9v4pOj
FEOM6++BhyQ4dc4ERFXiMhbHMu7LnDmPeKTx1c6681suj5svpZbdWW1Vz9w7xWHZ
LQjStcJSoZNA4JpPkcZVWdgHr1/NIQJT0DMz3r1iJ9STZFXuQS0jKst1tDz5Ixfb
kXAh72Jx8XQxziy6MqJv1vvgesAnUinvD2GT6k+mDHlBbFIQahbyOcdfN26pgRDC
9l01/pPMzYosHbbxE5nwb9kGuEk7sZJFgMEqpb55qe+fzhXPbBPD+2q+7Uw2yck8
A8s9C27IBmBv3eYi4acO11iYWximCxki76YLgPTFmsajZIrsu0F8RTsKUjCRjgXp
yAvuDaHn43CZAib1HdfwbAvC9r6nGSc8JnmTZSgliA8dT0ejp+vZejw6+lPcNOam
lIVLTq4Nm9kfmAfyJJCUkdXRGUvLL2NLGrX5bmemzawL1V0CbEHb+OnYQP0SBINw
b5cVSY/IUXzwLXyhNh3USOlLY3tpspN5LqKWArr6X8GS4zg2vpQCTBkS8/LwAN7a
pxt7MPs3LhivY2wshxM1TzznCWgXOuDiZp60QDuA5kZoFXvdi9TLV17Y9WvpAJA4
N3N1BwGJhtT2g9lm0iC2jsY+wLgKUfEe9iqfwYpFz4OaZcMHVvvzzWVPTMvtSPiG
bhUCiHjrioaE1e2EE/PkNKqvYphjXXqm7SkqoKBMcfaezEsI//Kqy1yBsKh4m2jA
F6sG5Gg4uU876ACwyPOcvvtEewqwRM/as2emg01vjFVuCo9Qki8UPL+rwl+KGILk
4s6ealegZy1DanrR35plaYgUhbPAQ3Iv8LSjqxd1UGSgROdTJy96me/F28dNGGX/
KIDAasjXIkbRfZtxnrE9Tuf+tE5xLGWGibxYrYYSXiMSfUAPtYKts1KcPYeHijtQ
x+4W040pO5vtTdq2wT2tb1yQM5u9SEVo/tNw3ECqttvdg9jEnmi1tSDjCI7Km8K1
8bUwFT7KhAgmAkUE8cL30yr7un5/ZciY0UMCO6bU3yAPPGGkxu/GcF6f/vWztR9n
E7JHzxqd4GVCnqkznonlZBxwK+lOyff63Aw66PCTSC7/ZdaC7XTINw9bxgb4fdcf
YY3ea7sSXyRFHx/2WoqDDozqeS2jEQlILIKi/ZhfriSuZbuWbrz0N9N0XQo/TOkC
raCDw1T+nakBfsCehi4mV0A+aNxsnWs57nN073O7QXbwD8h/g5An6ReixVGs/Ozg
uDmTUlr05SX0ZU+YVP0npodYkwULmrkq6vYf/1TX0QUroIkGW6iIxM2NOUxlF7UY
VuCIk6LKeBwLUzoxpZ0zDeAfp/B5Zt91oBoOrepIi4LaJoiPukBYY/7jbuvjlX3C
FwFmx7X4gL/S/XSDG8Meu76vYP1wrKDRa6rcS8j7NwtpqUiup/s/HXFakoqVTej+
+7B3K2ZtNkfIxFhs2XRs2cy69V9b/02N/tfQx7Xk0wUTYdhZpsjZb1/vDqAlwdbZ
IQalYBQWIm8Dfts8z3d6g+EXGIAmoXgYuNkCnGQZ68/uV4ZbBiNBGNzw2z91LvgZ
mOmzVNrwGbvY707AvoQimdDeTvcQa4woAWpxFizIJSRtuIHWhkUF2ao3D37XsSDn
/rqN8rUuBDtMZc9Cz1jd6z4yBBxKP/A/WI9dbgRLJZAyqKEBbBVu7Aj0GpfLreyp
I/dsQIi8ZHfAC1IdlJjfLYwz9of+KAZFI93Y226y+Ko7IVYaynKgFCMbmTqAy+2W
w5Co1oN2tg7VvkBEFdOKphFXekbc2d3KIASKmGVQ/nndDelGj4uSdAzlHyEQWy03
kuRnnTv5sYQAmyHD77riX5VQD9kyM+eYVk4EAlWRocfumvDl+GuVPUeGQubE3VWt
3k5WvhPxb4B8dCmRcGi+Z9PcxXURrha+Oliol4Q6XWGHQ5nrsmb0chzUFUR0lHwi
MXNaaFa7kMky0VAjoWmWEOdlJqYAfUFt54nITLnnGaAlOID43AJw11u4cCFWUPK0
7mLAL7PkY3SWH0KnZncXOH7yxcijP5NmD7399Lp9snB+5tYUuPuBEPxsGJam9Vro
bSazo4KdWwxEWbjkgjCVP0Fjhpt3CVW9a0tWU1bXHvgR50cbtZsBArD9jvmzSK1f
E7vYOXl8FyIpGkVpwZg25ERTHsOre65GVxj3E0hHZdLOfWT6YTaNLz3bwVwK0fNf
LSdEseOb22cuHwzGPYmDg+GQ6TMJHw8XlW1hjEbEWxCo4biTJVuEWMCnJJrtl0EI
V2JEuz83KoLbsAFNpSI0Ch5k5NCXXPxvXxgaXxLXVsPyRrWuRzpIWdDPD7QhUZ9I
1APSbxDhiQdvNccPnxJkjUvhMAAkWQO62wvXsBsOnEjt5o/d4pmxU4ibEbOk1tCb
UTo81AfcJNuRuXL1jkvkD+KiAu9D+9RtgD9kEU/5/1UdUpYML75IhXetbbQLAew2
4xNLF6lwAahjLE58PNbk67a87THlxbEGLF6itxNR5qzDqjhKDcAYzOrHm8XY95HY
xJn5cim0tA/tN074IfDpddAxBLxHHgvk+d5h3O0vtKVgfOkGgrDxOJsDcFgLwUZK
ouI/sFEBs8dewjdNE412hALxZ3IFDSJ3eP6B4d9FncHkloKSsGHlTDqBjUU54D3/
wNvUrRFBCh+X8Ki9ntZG6zDWjAK+hLQAXsoo5WJkrptlGdZbR7mm1MkYe7Bo58h/
avbzbZDiWYh8Y50wfl+ZnNB27A6xfHNMPDVS0UUSxDhLRwrmvRPMHWU095QO0Ycy
qkF5BUN3ZqVTfmes7k0yK202vmNPqeKUUCl9erB26Mfuz9mDsA+W55EvUpbYKeQU
FF3WXgEj8Atz68B8eGLz9J9tU8/RSCDtrvH9VlZETnj4PIPTvNJsuSJnbO1TxqZ1
DwiZVC43yUJ+BMOIID8sac5o8tFzsSnHlPfuFPBJRkpxwYWLAyNhTFjkrDNfSRC/
VTr8BZXgLH0l7n6xH8LCEV9en5fYnKZVzBk6zf7NMLLazpdjlY/t+itwK+alvCTw
wRapjMfmML4ezMWgpnIX5y8BshTqPh544Sp8T/yEIECkq1RaTYvVXWL1aihwWjKt
BDiSwU/dKRYuBMdkHiiBwxH1NUDETyhCsDbc3OTIw00mZfQhqYix/IWtCG5DE67D
b4Csvka/tmT7BIDmIbJ88RmIeYnZpXOwBa117XoThOWIiQeyY/8FJsr5vvRUqiK1
+REyiGKVSAayhZHHEU8qH91AX09aEfvStuaM53Shj+HbaS5n5Jn0NGNQ1oUQlcMj
7aIdw53vRDllT7mi9KkFYHROX29O8eXeIkIBAoDeRTVF7inYpetCRluKFuC6kIQc
c0/pKvjzqi/Q40yFAHQpoK37kN8q8YCfuIhlV8jDcONnIGZLKvPUqhZ5yS4sW88F
XzDAjw6alhTa5GFIzdusLtRjoMLoDQw0CbGIW51SlG7NIVUE92etlYFqruOTG8Gt
2j2nVkw9GoUTl4rqY6oQgiwPMVYRXoh6N75bdWxiB3jdoCedgpLRwoESsRQ2PUcu
ykALmdpPJbvmYxgdTIMkotFLmGBqVb8klSArwPHClJ2t1w/1Udqsc07RxpAf3Z6y
SzxLTVlcKf5rHxqEO8uaTNvRASBGKyuEblT8zvuDlzsm1ji8J8wXbRBA4sH4GirU
6x/d9SrBsFsgJSYgEeRK1aRAvO83Om7912+8DCZS1Qz04am4pce9JUAmwivBJSLK
9mI+KIKTvzh4+6+nsBg5LBjbLrICI7KSzLBX2Xxx1keRThVm3gv0QBrNWfK7anoY
lsNjPs7PgMefQYcDf18EOSS/o3xBMhgYj+dG94IV/7+IMRTE/DqYBFUxCi8LSGuz
NTsU7nJyAlebRagFH2yPP5goCcMsekABjz0t1dwpDcWyVbzoQT7EQBiVupvim+6Q
fofpklZJ89hBL4g6dybJ8pyxBNbR4XhMJ4x+i9YGS5C+gpJaYb0DdWYB6/SM7xC0
g/A6Yj5ExBK7+8fi72VM5YO0ORuLbU0QbqsaQwNdPsPRs5wsj3rDIjJhz0kgJswS
LkhRSc5E0+MHlcvnGy9lLhxsCgS0hql79Ra4kT+VVY6JN/gufeNlEIqsFv4GjfX2
HhykOk4h1ZixJ2XnauweyxKfTucrNMoMOS/4uNURQ/ADVliPfBmA4uAkf1nsnOWZ
WExoaA1M7lfUryXvyaccDzs0BAd/RKPWvKVvSprN9eRiCH7J7CkRwfDLQSYOp3pb
G0cIZIr5K/ahebcsGU7GVSNOT41f28sfLEbGocyqq4Qh58S4AEfdGKBoDnEnfI2E
9Ww0TqzBZLInkATMfSTEpa5yxULfiYoYvXqtNtM+oKSczdhlv8jv1jsGCNVWc4Iy
vEzJ0HBWg2/K+ZA5PC3U1KzjrZcNpG4EzgO/ZWlV9nqMpkj5dHckoSqZET4GoxQA
AvXGNm+pg2gToZyvWJjKJaj8sspqhUgMI/Q/soSdNUOpxoQ2xfZlQHEygk19uMQG
Nn6bPhbGAqZzQpPqjrqu+/izgDCJ8NwTE4k7bDr4Zhog3yMfuu7wipqpvnLD4MjJ
7tYBa3LwvSP5Pm4Rfk1Cu8u5wOsdGJsqF8UUYQeo7LnuvpqNwH0AS00bO8yitVV5
8LmcweEqm/9FqCIjIco9XpIxnKpko2b+2NUwvkQ91/Znr1VL0O7iaU6cEbjeyY+c
iM3OXieUlpHqyEtbMqWL4eDzCpz/4gBwM+5c2ExFI3ip1bdh+4fQ1iDjoXEqH3oN
4xIHCsD7uDuVQFYub8fFtedHVW5BmkqZR6vllXuH0fPOkeLxUCXDx7gkxOFKRNRH
Q95fDpPXMuB8WIAd2sBIxZBMiX4Elc6smgqxIwhoIBmNaWZweCoZyuRwtial+76m
S7p3qOIsDLRdgVRNF3epASW0UX/Pw6SDTebAW6wy/FeiDNg68/hHCrNObbT15CTR
LXFCYmYh1krG2JJ5A8HVTYHkkN1pjMhzan+8CyuTfRqXOG7EVtJjRG1ZwhLWvSc3
Zy/3rqbBT3e4P6vTHwM1aRqoLC7K6KleIWQuTG5lbhqhY03LwDIeBRdTkUxRx1dy
nFvSA2fR89NrbSmJ6lMoeyWIoR0YON4YYteQC1EkaqM8RUyr6Ta/24pQXPnsfcmz
yF23+//nqaWXNZkgvWxx6gc20T3GIjAfczS8AAnVas44HguNG0p5oPBZcCe8XtEY
yNXVm1gRx+9CbUtDQSI8ncwePSTWqTZ/o1KxnntmKjEAOhhOpXOlaghVIyRkVVQh
E+7YqlOyz3HyVVqC2PPR8xSuK2HDEs8V4xgY6802ANktptY167BiVzrlKBJR560w
8L/IGmx4QLYYsjfTP+Oi5fWVNfHVXiJNnMKuSLYaHSXegaJnyto0yTR52Bg/s5YF
qoGTL0zfL4gdama8V6oy2wOoz4X1qvyz6yk5NxO2K0B1B2tVW0CIDIoVnb7KV5k0
EFBYb/63GR757tvBOsMVCocW5pCkhVARsN+QajTdL0ytcUzdmUresEDFLMgufatc
Sze2CWqx6wgbRF+qeiuSQB0iDKHaOZVzojgY09LavpApIcDdIPMca47iIOzgy74X
A/EQ64MsVLtunMxtVXiJ2GI1iaKNFPlKsDK6U/InVnsNKm8Co2SYzy47OaSgf23B
nEhzX92274LNAAUMCAOHVpe1rX4lDTfzXj8rg9opehO401xPDqpXgBgSz+SX7F9q
0XqrRvoyG9NkxqMGzgcpp7HbJq8nM3QepSKQ0bI/m3k3BHRyrHdFoups35u8859H
fppuMYSNnf66Id5ye2oTPTx8n1DxxThDS0tZ2iC/+FNznFsbubwqlpArPZlBZMoZ
WPlr+6uNue0x7K9ovoDeOuwwUlWg0RM76Hft41i87HhKL/dT6jQBKcC1TTf1htFg
5onV/2upWNlH2gkOcERaP1KX4xGbL+ynXSmW+cTfbsR/DDekT0GdADfufgPCnSsv
3nH2BfWBgJDK50ngpwSJnkVu+9qsRwGNzHu07WJddh/CH3KHjLWN5irdqSioBPVf
CMiS8qCqOGKaFg0vds6vM+t3rWRihICa3DyDTsjA2kcWguHTT/Nd+zskDxfU1rz8
ISX3/tPqYIf8z3CPRLzxxBmGTZ/PNxlvbv+dtIoimlMB8eHqJQ690oj+QUGRjd6I
ZzjkukvfbM1L6fTDqe64ZrrRN7iGu+h3Ip8PLS5z2Zp3YXO5k1MlCpjRrXIO4ZBh
nmSXi2S92y6HLkWoX44KrMh+urQOHqRPkDgF2PNwlShPcnunzwbL1unkRfzASeyE
yq0/aPCCvHIQLnDHmks2vCyGzF2xzvdgXx5CVN/UMfx+Ee483QFoUWsjQioBEAyS
eckYggsSUzIPnHZCJnb49KbFRPwYNQCFgyzz4punEiuA7oAhRv6E1zutxmXiqukC
72W7r0ZE9IZxrbeMg2hCqhetDiJxAzgy/aK5l78qpWEO3E2FQsZ0uMFR/T9bVGV6
hdG7vAGM8C3uvdjVZD547V6tPGzUJnBs2X+EdiikdMSJx4bVS/6jbOJxoOXXVdDN
2NwJjI3pWFBTcKfNhZP6V47kMomzRUKfYaXbyvgFSxs47k3zuvFJYRdZ2vUnW2P2
bKzjVLiK2Z1YL7RwGqY7TxDod3tTzV/ET8Z5Ah/uS9udBmnoMWDlqRDHPqCBH49T
lW6NVx6IGw+m6nKbGwRYxO44biPwIwNximN7bv7wczeLmYtbCqt1LF4wXumtycsn
N8W9DsyjrnO5e1UWKz6ybzrsB7tPdjmYw86uO1HERlXA+KiB1PZNCZu7+vg5xD1S
ufWz8h0+zdTvkhRK/3fB9GKgZyiOKm/57qha2Iw4BFc5CRbu9bIOMGkgTOQKcoB8
6/RQp/4LdjvtzDs5yYdOHXIBG2M0pcxAZPVvVkKSoCr0J9e5dXbiRl236z1o55+I
kEix1zuo+zHmnvTJCZ4dEc9pNljOgZ1K9RkcoIr6VoWqSxArWXcxL7GpEURsdQ0U
5dH8u+aEhxE1pewyhXd1csSm3Sox1TxqxDzdedO2f4TU//N4lM3vJoQcj+bPSyE4
pvluJOvfDNkCEPVMzTiWO5rL4Fnd+aXQHjeQ6aq3/woq2al3TTh2HypfqzFKIjxt
xWE30EJsP76XeTeue+u9rcGSczxFF5aLHQkPq+y7HsWoSBqjhupy+QS1Lxkdhcy+
7ILTyzT+oyPjaffKUyRf4zEyALf0u2+kIiAJuCJhBIArr7zVXOdWYaONlB2jDXMy
vxJcdwMzgk8EA5pZNjsC3sGTyNVlUNRGQICAcASV4LjtFeoZcJFQsRCP8xAvtkcM
HoTegKjRUsWtk2c4wbuA5yoMdGwAslDQSykRLPlTFq4jQzutnjmAb8yvjLSiu2k4
AVm1KZnZ6d7CudiH5PouebRh8kekNqQgklsly6I88nqAAKKVDLRvxQLSKekMKXDr
b6QfZJsgaGg/MDpPRKKTH5KOX6lsorOt2Dae0QO7nFM5xp/8ZlJdFmYtP+z1puIR
YWrcz2qrW1o6ZGwcYqL3CCTLd9EwK/o/E+M8UY8xBQmdqi96JaVGiXRHQhymo+8X
Br4ziXnZtZXCTY4kP7rncSixVJCNruIhospl4xJ/LM9fHrQ2V9oMS391Ly5+9pec
+mliYdp/f8ak+6Or2rgMrDTh34zZ5RFakweGapOUdCS4G3kcyimfhhygLQSQNZ40
26tixU8q8KTfva4R7ZqYVj+2xIUlZX8rORBgL9IYVmgA0IthvVLRPK9OdqbIvhrz
P5+1IL2tLL3Sx0JY+u39MAF9dD8bzk1F71tCjkXKGVaxiga4DTCrylspv+nEKQFq
SYE9sTgq8gR3w5KzNFvwkWeT8N3uTufn1iPzjwLG2dUgbhVOnVENYd74bKegS+6f
DWhNTyW07Yefa+kdbx4LtV6kwFnsXXgPDxk0wcUb8kyLMUdWmQ/zBq1xNrw9oQlu
seeLsYnPHvDqfLTJ90DjR5jKXBUTK8iRyuyE0PaY7UhHzsxVzffoMK57uyMyBBvD
Y3LQgORGGRo8J4zRVn6F/PxtKZZGp7//1ISBnHD0pbPQVjWJqImxR6t6dpqYmNgM
svmKA8c3vb5w6g7OAjsbM7ijVDDLOsORZO4fEcpjcsebSd0hREK6PICxL1BPYvua
9ZOzc/qx086zkg1EI5AV+8nNUZr2/SMjc6e3SLUPt1+kd/t9DusuYUx0jaOy6heA
gCSvT462TtkToAlArCiE/FDHXTya7k3wWFYH7D0slArXFM8L5LwNlDWfDhLB2DM2
mbB5FQm4BpFN99/+0nI2jwEA3wGPmJ1zaCyiRru11+TLzkK0bSIVQc4J5PCF4oN8
wt417+120Mo9GzSMDAFFp0j9FIct8eWgEYVrcpzdGjs5cxHNdam2POdlxgB1yeGr
Yt92bQndFF+YOXuSxVrAxsTL711rxzs3ssOJE+YhTccbw2ggCxqR5VPo9NFSxm2c
pBhnXxKzewO479WALJh++AIb9ZJgCEYJbSNw0g6j/marwkMTXb12/0Vrnwr2z3vW
8/7/3hKwOvefC9D6poBvc2SBtY7s90TAvVAPKogZD1wiW9pzCO8sdtyX7ENaIaoz
mc0jdWQ2CaYEydFxrvn67Oy9pkjUbeyhSAnU8lvWamk6z4DkFqb8LHV3cEnV3B+0
hfAFw8AQq9dxvgAVXUNoafPbUwS66gCjXvcVJM5lpkEUQnkjdm4q7yQama+mXZ25
fp+IzlxItAiXwleoZVhMY52JO6ySKuprBb75OQ8HTjjGVKRKyZydEculVZmhkitC
8/OU7LTNLehy6ys6/2BAdIzLd+oJ76qbWJGKggoj6xHCzpZzSE5AGHqUVDw5js9S
Htm4j7md1nxwFC8dNuuLfeftFGFfAehb2iCvoGgVsLqpdAWr0nSfEunEDVuim+wV
4IofEbhoKUEQjCy0TTgkofagNtlhNejEDxOT8VYKYtI3yI64Q26gZK/d0CPQa8wH
U85NUj5kSrdLnFc5bZkAMlgA0C233g36QpOLBJ6L6Ku1MzEnX30Qg4e5lBSg+ZT5
p1S/KUEAeez0jhftW5wTFIwvr8bgKrJFFcnqrqnp87L1/obSm7gkY5vPlnjXkdQ5
8GqOQIDfzQ0xKe4ZUq8L8rvc9nURfWxgY/vgUZxkisN4LYQvSQSkjQoMcCOZrk4f
bdwghkhJrqum/z7YQxN7AhrapbDy5HzAQCtovpMgv42FhIkDDaGZY6SWVdqnjOw9
aabQyXWxm12fB5tc6edRT9Y/HxxmC5iXFZMUzOMNJriCCyIIbBSVyOgEn4AwOFlU
9om8ze9jKWRtfqH7+OuUW6Z8hIvzhmvJEKBd7Danq0JEC8hCvPylJkcRhKPuwmGB
cfW/XOITt0mV7UVRwnfPkAmf5EZksBjsTfpWqlnfjkUtRKKwKKIX/ANZx4X1KWrD
V1WtTAN7c7mXYvCShrez/YOHntNK/0LBs+Uch2bpHeeI16DQY7wNVH5zbrrqOc9r
anW+blT9rKWuomnYgpDtLfRAmVNhVv22V9COegQzRzUZgluxlZwq73x2xqQ5tl0s
+hcZc4A9S/lPctBb3LKCiubBCjZTvzlDJLCp0ZimfWMpNLn1povPrSI+aZW1vT4B
2QtNp4fwrj2kfApdSKKyTuPmgL4ju5xqaiD6TbYXcBH12YAPXgwmzkhBLjnyIYR4
ArNzzxKzxfTNvSfcCdBaD81THfiCPk3JQCe+OwUgpjBBKuGBPNbaWSiEI+WEsxXp
ZDNHuohStjIG5VOjjVbizOEaWZttTO70ddP9ccYfh80NOuakJMal6pfmVnLieW2H
NO86VXnfr2jRyCfxpExAnNmqjJsP7bsNYWryxW8LrNLHJ3XQOcp5G/05UgbQkN6i
y4xhquHqm6lOzm+cad9FLhIcbEGmuyoANFeRR0LtjtjxLFUn96b5YE9YHViE1Xme
DFFI4hony8aPnsKVhZY1DyP7aePrtWwpStsCXM6sI+6xMYo8Z3gn+PyUgmN9nO58
Kx8rHew8MQnv6fU2k9D9PcjPNvHrCjEnR6uAmsPqcm+OToGkQlwuvACQVjbL6GVA
ALJiS0tALuHCysJ+mH8u+hPOOXlRuQuhgq9smUH5ukMsrxcBP/CduiwD6Bg45Grw
++jk+XsF/QDpitqDVuQB14pVZGRgk6nNJ7Dxfjs9CK5I2Fxcod0FWEaNzchN5BRy
SotW0AKT1OVTkwZoG+q1VeAaANb3z98WbUmg00u+rqdemAA3AQPsujBpAWgaxZhe
dj/EkS58RFTKbERY2nEj97EB6q2VlY0RrV0qc/OG+ox3Ss6z6cTqUl2ULZgwl1VR
V1dt3NFerATMdsXVy2nlxGmW2X5VPk9JQ8q33Y0v0M7RqTT9TmaW39a+5Ze9lUv9
ED//em7G5V5zdrutbnW9lP1m48GBva83OXPBa0XqK48Uz94HV1YUQqMy1jxknM5c
+dqvShcZ87w4D94JYvjCB58jFc1n71oayCUyjbhJSgXhyOflVISkL+dgc0kdDxqc
kJVC6aQeH0TIA4ZTHq+nCwC/SFLodLvTPCkssMd03vEaDrjMQYgCmAI+NeCkNJu+
7FSEjZ7ar4P62fzj9dmjldJJFM+XxJaBkbwr7IatJYg/Clq8uUFeXEs3gXFdAoM+
w6PJGACGVaw5GG2Fg9VTkuh63tPPZxSgzCY0qsUYj/BILLi/r/9JpS6tgXG0knEb
5hqUTUE/BUCmOeBhVmtuNDZRnVlLG9AU4K8isM81v/kSWpApiJJrYnsZ98wD+bhS
faBmm+M9JjlK4qfs90kYSZ+1Lj6v+T1xzJDUYyqeJ37TLtumwXjZbQCoz3vIfhnM
yQ8T5WKziq5Raf3m5dgR9NIhOBxGj0+YMXw0pWXiCmhw25fxpcMvlh+4K49VMeZ2
PXzhrUA/m/alm6QVx1bgXLZLZsp87wFA3KDeRxyFPfqGyxcB6zLYqA7lmzaHG1zM
bFOIbUXUmN7sO+6gCNP3CRutfVvb3gciGNbBJR5Goi8BF+eY4FRd8XdGp9g5aj4k
AxrKYGaFsLQqqDy7+xZZxQMULM+C110x10aW35YghgNX0iLh8FB0uP5+GYkeHxLq
jPf2UKc+wnju2EfbnHPAUOEJW7aL9KWu7zOEbszyq9li+FCdFf53pc4sSz6I8tNd
Y1rVnw5kUPgAHhxYbHaPMfJG0AU6WrAoMLBd+AJVWs0rTDu04CitInCfGCidG7FF
DHFcE3ImLqiVpbZ3eCRHRksRWH0g/Sp1XLVtuSCCxHdyHKZNK7Qvz4fo+Mss8Yb5
GGiPlacXW0S1TNBQd7pr74nVgRqWdKY/yGLDhh8MB30ya6YAkdTZLWUrpRce/Jlp
0coa1qQmsSNus45sc6hOivoS/aXkq3wqJE24wyAbjjtbXiaHXhmjqQ3RoGZGc7Zx
uLfKj0rRN73PsyJRZp3HUAk0gG2eVeg0xnO+Axt/uDTjtUMv5h68IJdsKsFQIMI6
OuuhfV+aZBqtZv0m6WHydEB3DnoZSTmZynLsuhtpAUTwA7Y8EG/xRWwyKnG2knAN
CzJcsF/0knwrYY8XeBx3yyxI0X8HBNmWTwHn63a933vbfzlKNQLZ2H1B8lP9yvzn
+lCZnCBY5b1wGu4+8lfNUSEPyHfxep6ohmbqDMh7G/Y6ZQf5fEDH3tmOKPahzIh6
O5AmwqVQ4bzESp5G+iUkspzp0cIMsfFLk3g42KDLRi7PB9OWwYlhn7WLDiQYXwLb
3lTdQ451/X3OfmLrld2vrACSltccvkNyeDRZFSbJXxwcVahks+hfQtGkO8FyarFV
loUTHw86H6YwwoMJZh504n9Ku/zWz1pqRgOIorVrE31HwPZItxpsWtmLc96OdOhS
YVQeHjp1VQL97P8wF7xAZ3X6NoWS3JDHvE3HyPvKZbhf0Fz6AoBfSJkclTqYoRZi
XDgw9DDmhp510zGi2bjlYmzpgzSkiOQFUQOaPYG4Sb/uYjMpUZC+Q11mcxR8TNP1
lsebgQVaJGDWCc4eKqtFKFneIU+mJnv3m8irc+XfxbXLsCBLfvtd3WTxjb9gcYRs
w3mBG26Kx9+619UORD0KmcBovbvDR2qdDRGMkeAU1ft4Yyr4lMWsiGKVwECrgrUy
pceSQ0pjJnKvywsNMTC9uZ7OrULt9DrqzF5fLI0PGLmNt6A+MMv8BUpKUTf3jAvr
KogIyv17gFlSFxVuBDo+PVRLis1Ng8Q5MUlxhmT+GIDigBsiXn/fxPp103pCcw0n
eDQ6apRb5nUhEjOUeYxb4j5RLUHhtl35FVhR4wjFhpiPsueIoUVxnVoDOr9icAKQ
bjw6oqb9mcMFdnZDYlWyIhUxUpxd3NAaDn3X0Faa3YCXZs4/X8ofi+RgkeYCVd2I
kmNwxQev1vlv2dGNoKOL+krPCSTZK8Q9qyNXsUvGQV8zOSYQETQAiq9vwgOd2ayI
egb7KdSWdgz047JEnaoZZA2iSdD5ZlH0QAZDM9dntlHf9RNelopL8RClNlpvuXWG
nRRoMsfwQBVrCZd0VLWD7ENBub2ApFz5E6g7sxwICyqMaUsVGacUpcxmgoEpXUOK
U6HlAkkTkE9kIOTcs6n1FuhMh+XiwGDEUrZCTrgfjOIDDfPcpQUsLMAAHQtfP4cF
futz2uS440Q1lsx78ZjYYO+TcXIdnMOKDfGNTFFt0x/zKhrMpsL7AE6dAH5wtthT
LypVWGzYhkpbil4kG28MAoTxxvndy/kE/afqEmEFNxiRWbuhZQzYLDorU9PxTim5
B6G2kjOFVGz/DnL+QJ6QMsSSH2dp/24QpoFU/yYUYMsougsQwPoJBQTetNirNqbC
TpPnVWZ6vqgWdqqibD78BuppfLxTKXHXNp1wsGcnnb+YPs2NmczIgQn7Y5NZ9Pgi
IHbcHGedzBNWe2LvxK4Xrde0A+7Qa5hTQmw0fPQ0++myXBeVi8v8RvRVgNWq8yDj
2385Wr8IEgzkke8T1kG4TEhDL4FwAZliov9K4yhbBqBE3teRbvU3uZ6S7+1YDXEB
m42k8PWrBiwKlcrt6tgUxcQKJ5UXMyK1lGFByOAdv3Sy764REnPeZ0JgiYONKmaH
u34BoUZmAfdO0NW7Xvtlj3sMaIveFQyUNE6txrLUsGZDbpAUVU7XH2ZxGIvHRtha
0NQnQXmont7EKSgAB4pDzU5oQAIdciuOzmdfKKS4qN5jcq0OgTYL1ImBjePG+rJc
Jv5L1MtqFvm/ZkjjnmGXmicRKbM4uPIT3Bc7w0JOhVmG4oRoIwsA1sg6P7eL2BJS
zktKd38+XoCjxnACkclx2eXZsaoS7T6Zb0lLjkjkBapNl8xLLW89SePUkfxxoD3g
tDM/p4XOatZmpiEAul5/D5q1cX6/s8i7pgZI3DKmbqE1ipC6FJQNqJMWCiTU6MA9
sRijH21ffRKiM/Xpvhnw+E/AiD9qSNqxTw/PmgsXVEM/FWLuSLY1xv+tEJMFyRPD
nUkb95IvSJzE8n0Bu2L9tUflQ38t1zvzibZ/MrHK0mzBTTz24lW+LbrDX3eAZEBf
9BrSMitrKcWy8EJ6JLaTOdymY+KjDcxyTN7yOB6BcJbh5v/NexKN7jAtMlb735SV
16H+KdeUetynxdadU/2JAGGF40KsTQKdar6HM9EySFOzps7jyasraSMckolBrQTQ
IDAkvdLocjbG6rYcOqUPGrGyE1DbaAzaKhUP4B+L24FU/B07sdHUMv1knjtRCoKh
YaTsE8EeEz4WLLloN90MUnib5VEnTTBKVEJ7vgNsFLXB+CGfHVS8nyddQkUygdak
ghy2k5dYJ3DXlZcCKN9VBAduZY5J3wheB+90Z4l6AdnMy5eD3RR0Hxyg/GMn9UU8
Kt3saMXyCPZO+dELk6uPa1dKzrW0BICUoOrGmXbVbWbdk5nVbl3Q3PZPhWT7nyqf
972PDvR4faeKXEcwoW3XIRhyvDpTucHIrM+dMHL1wc7D8Kn4Kyp4DSVbma7tUp5M
/SPvzDhxuCuhq68y+hp3M3C9Y9BO39rqGA7oaN1fZuV6OBWpFXuE2z2vHxDvrSM8
Gh2/isc93FfBsrFmSD1oDdSFSZSFv6LAvK1B7G/DjAMt+DF4EFlEo5mgsbP7i4hf
hfXl7+gcrlWUuCMpiH60NdWb3DlfVwLtpOUFlIuPRmQ9kfm16WPRbIn1bn3eDl3/
8YJE/YFTl/w8LOk8mOnLTyl2ln4sAkgqD34hk16r8n3kMrpXkEvZmMzN7v0knWtr
34NuWC/beAHxALoiPluRysEwC3XQTjvfDY5SMAhTTxHWjvooY2GDszxtbJxT3sfE
0m79JLi5ZYOBAkJYotVu2dbxeHX8bmmw+9cMug8SALIjWMR8Bwhe5pgJ3qRuCzg9
QiEvuaIrvlSId+2S96fm9kt2WarmCeyyXbZX66LUxzbMmE/HsSpxCmxHKYIIaA12
9c2F2kZITJGqZAj+IxVGvLqd9mtTHlexcn0P1tWiEPLDYfEC+SV2gJexV6Kbr+bU
+20URhIzIh8sacTMxBBlVSilr/JtyBb6AFVCRV8dfqwCCKzqMebynoFN8WEhZ9z9
nleIik9f4oa70pk0fvbpS+emzqx7BSE/HIWLkxKqrLbGZQdVK3izjGDaCoYGx3ij
2/Na2y5nXI8Pe4naBModr7BxNxBxnAFDC5MnqUVT31x0n9bfqaq9JBeoh25FVseS
zJSlqbirjI7GPxMOF+PmQnuTCVwWpsczqxUpBBODo+c3a6/bHaJXxoPrz11BFBgB
JozSfoHU6E6iCHA3iTz4ttvaj3/kwDWRriyluwUnJEsIh1LkyjgoC9uxCdFRGbe7
VgmzzJPTh1BD90JeFqiA8lHsYHLbp9IJPEdy+/j5s50gWbGdQnf0ZQUIZeiz2LNx
QOXo01C6nNDi04HKpZC8KGDtlohS1a8iG7LI0me5L3rZSp8wW7YvGZE0e0IpjTZJ
ct+19U4bFZO+xrg5dNYsg59PAk/eZWtH+xu4ZJDLNTVExUWBupkyCW4SXm0nROYe
Ygc++YzYdkmZkP8t1oBUyZ9gg1CFPwyp3J13Jml15Y4rboBFAW2uFAUOaiyk8yBB
3JrVX2mHG2tmy8SNyj7d3dDo2BFmo84pU+IoBBTMWKS42kDxv5XqxJLKcvwAQKz+
lTbhDPy8/X/GQGrE4OaQ/YVfGq/Q3y5+1T6wbGlbPhPPg985S0dnCk4RtSssWlkW
TocDuOwsEIiLiEwLQwgL9duynl+dbzchov27gCi3Z/ktOVu6ESlnaOrJJYFzNAk4
O1QzaVgOZmfwYsydjZTMODX1lE23OlzjISlSCftpWO6y5VJZTs+v+NF5/KRmwnEh
6y/M+O+Eg/Yf7yzzs1Tta4tUMQj1/cLDtEOEqoaRkc0TxkhNH5V9GIuUHjKT8BaQ
XOf9PMhZGF7sH1KrNw19S21gpPD27Tw28zUqYTjksJIxf4afmcwFHEBzK0QC2899
hsNZaeBXMRpZeDzBB+GfcftIpah5r0virvwEqMMncxllEM513BBV3SSFPUeP34jK
49xEBu6jdIc1mPQAaF33GGeldyXkYjXCaNb0ET/EI2gMp60+ixgGmSVq1s8CPKeV
s0jAZOEvNHn6IDFxKLbK9wFDAOUvorBgshAp+KllLCtiDlYcc3wnW+a0jROqKcA2
fgzpiVhBluhWMgAcqsXHMevG5xyiuwiFSzYIWigwuJkFWNGnIahoLu3dNB8EBNk6
92iBguUbGGuW1M76mZTvQow+B/Fhs4n3Dv10O84xCW2uGzg/DhR9N3Ey0NLbpJM1
/tMS2J5rfew5hIXUSsRs067e4jUU6CDR7Giij6/7YYZECCrQ3wJKb0OsTs4m/x7p
fZE7rF0hkVpnGRjw+qGS6Q2vN03VoBtKFPXQawGKBm+7lpxiYSX8je7b655wcQCW
7VFv4LIOp479mFo/CRqz1Fq68XuiqSoReTfJeEjND34EPpBjBTTWFgvE7ZeTOL0l
+O7UvUgue9ZG8JkU56ACQ6qZTfu9dfIt2t9/IZVzCOoRRXqGp8igr+uh+QI2RItN
vHW297GhLlgfGG+DtEOOrFyuaclWfixpeuYJkhcLn2iwjwXMZQOzTG1j+68vbNcq
Hi7H0C98BsQ79nGwVKtd8Xlia5t960QbtJig5OxJH6J65019aW0uJXV6kk6OqRdr
CHW81yCgFt5p5GiBPnDGPn6wzH3ZBAvO2f1EcmCZbM/cQBwz4OKkMY//9ya4HWUT
Iy71cCL9A0wv7S8YQ2JZdzrPqIcKNgeF9kn0aqQfnykIuhQ2OSWTugdHIvpYFzHM
NT1JZYglaOf9YFb/hzAzqmEhCljP38vnTJuCpQLcSCYr3YhDmEMMHNVbzDztkvpA
TnB6gPrarDxZVApJoLZVTLNZXKJj+Wub84WA1rfthaM6Q4Plv4zhnfPANO1GI2N8
aWa9z57dsqTbFAa62Q8/0P+crcqFZFDmtp9Ldx1YDXALjOCVRM0MIOGzmSa41hxm
kD2DmABebAS9gmrr4toXTMy81VCBUuh5bTgesVzHdUKLfaDVbwfEi+HvsklsukTR
7GjlGHjo/P3BZSFzK4S+qwPzV/YkhisfMnIlSzW8p+jjIG4q2PnU8QTe7iV+WwDX
xvsc+zDeCFPti9wqMtSqcKLzNvrDTs27XY0ASUGaqo5LWeNciMCJSlbquL05Da8f
2S74anGkea8sF9ydUNAFcZIFg3qPalYdVHS06mKueqK3iWRtfhZuqplhCaViTHlC
XXA5lM31S2g/ffnNaqspAj+IfarbocAOYaU9N86tmuhiVOhYLIRi0PY1h2wsBPwB
Ate5qdCRK/EpbYLPc2onnHURyPAIyKDAWadKvpO4kpzgPGf16sG0ogobby9PCgNO
SMDoUK79jKfMsU3iLSF9JIae4ZZ/5pa56R8bceNKL+D61p/Og0UNxZVDfnl8l7EL
Wu70ZZPQKbcwE+jqiuwESC2KiYHWdliu4ghBladMarIyuwaNVSWqw7634H07pKus
NKiNFhBe5CeOTZGSbrRII/j10hEDXeA3MpNEEkmkA1np5cSMrgQp8BN4scva9toI
3JTQpHh7Z0QoGzMDTBxX9BYj/1FFhojCInelxM7il0dYZ6OJvgGcU28ABORe/bG8
2V3bueRXR9Vlpn3yWzaZ9T3RyHg7G9IW7DnDRw6MWK0P0jrJB8ElLyR5f7ORhzFQ
SnS5yYd95l3yzcAx2K0vUK+YqAXHKKYzVL5sSoFn5er7HpZVSqfoUrw7mvg7gRkm
vaugkLf58dAc6IbVvjHdqWEv9yUM2E/UW8RA2TFCi5hYbEdu3tUos5tdwfzItadg
6MO1W7c5hwWtAchqP5nZCGibzcRe1oTiEwY18qpnR7gDlGl8nC81I9MrSAVckYsn
lByB3vnQUD4bRpY+sTshcb1s+ZwQFPv5YWSDUmWo2sq64thYCLxcmK615aDlFePB
EhAZa0cXJpHyJ6pXivfiRcfXLS7OpzdiuA4VFgcdNrdRmsgLw6rkjunTzoBIWIOM
AC0O1/l8IM6K1d5xKjkV26M9sdqbfA1qwaEJuEnoaDKWTeD5RKl6sQ29H2KrcBiH
N9v7uxmzhrP5AHY0ThZCfIPeSSEaCGZtg4bMtZmRcSvAGAUFg59TlDghNnBdx6CJ
0u2M3i92PyObeQJ9cozDWsVgNGkVyRqNuTN8s5QNSKkq2Ub2QsAihThYm2yfYiCp
92ty9B9ALD047MvsbryYui5yQXPanML5lGRTQWYEOuOUzPGqZfBMY5GjHLtOJuSo
i+ljdnwSbpjUp01bk8DSXUtk1rwoRmVC+GzR9IJiq+8IVg3FCdP4d+Gu5xedjCGQ
Z7z25FuQQDOtQzO2LWCsiUwpufNppc+jrLIIL/VC9ozTw8EudeDiUi6D3J/v5car
0Zwr/WCkpk2LAoeczGjD7ekP1AM4VoAIpq5D/J5PibT59yuEwfgg/Nsp07EoN67B
CEvqNPI9fJZqVX3o8DX+JzY478geaeHEPxHtJtMMqbC2NX/PyLJP1qYTtjsQoy3q
BoR/yAlBvOghV+U9d6RI8EBwifP+xtMtfcAqG6yamd1bHNom0BSqUYPZ/41DPtcs
XUVGGLZcIoarEbTBL/F8LU+3EQUT3iiLOGV5RJoudjG+bNxCwq3t5oArbQYC1+kz
tDt0mg2luGdlfOPmRq4QO2zXvkF3yc1OXtJFNf4N6QDnXSaIIMhBrtYrQGLm4XUo
5eGSyx8WqlJNRe5Syp3ECeDj+EX5dDMSWyTI8TghiuU2VYOf6Z97pCg8PV60nddq
BdB3NFdy+ESPMpC87c4R95RoJm9EHU6i07ZNCsGa+on0VqtLo/oBZJFICz2gPl6N
IfKFiNXUec3y072iGFy9jWkOXsEPrIaq1e65ywil6/eNIgAlEZBq2wgrWZlU37Tv
rMWHYE8BSluSnXkrUKJdzMPiEdRiKOFApb+GsgPo82kd77EDLMqx0wpPjx3FUxZf
/305Mjqp8YahLxbBiXbQs5Vz2RPD75h4GkE8ccly6qdhD+O/P3lOAz8zL9RKvYv/
dOKd/HFSoKz4T0K/SymadZAkzEAN1hRDZcKfBIJi100qO6MNby82Ccz4jNCiwXD7
Au78C48Q7rLavHLUn/OIknpljKW+ft2mI+t/X1fah+BTfdqjriuDHaZvljahOhOU
sqcLXTa7Z8isRrkr0scNJtiTAvcIxf+ryz5TFsZz6QEiMVW7HQoV/GL8dd5qVrh4
E79X86XAd38nbsR5ZE99Edcoa7+enEvB/wJpFxGV+1GuGYnQ8cV5rRU/SilYBbJV
V/BLN5gzS2ZLhzjy58ks/MBtwUhyfAZ4qRh62kD/dv7odzZUvv/k+jeQAqdbDCW4
P/UhEUuBOMhhN6+pTdOWNKcZ5Pwsm/Qyfbsd/biqvih+1OvVcjPxoGoktI3HqILl
ch9MvlTern81y21Yh/zEHmIEUm7gCRNKnH6O22NzLS7NK2YsKRjMwiyVTbdlB/w2
4FQMO908ts9FeVs6dG9++iiXlOcCfvAaCeckc4NZQMbGbozWYZqmg9iyMr/ocxxZ
RoyPIbTF6jAhvRMSNmPdm+HyyX5Y0NjpABWqTjZjv7THdOBtuG5v9M24sIZwZYvm
6XZhxQJRQiV3CmSmETd8NNRlGFsFXmzdyRNoUSmjZVfKWfzaTS2bBxWuWZr0Jy5m
Mqp/3pFRhbPNzB/YHbfI2aQQtwhotEv2mDPJTuWZKcki3J5fE8uMSJp3Wnp6T3ev
E2+DxI9rxIWLvnLl68En+NnUSw74AVb+AVEejHNdpTuhmbKNh8I7SefHRiDmxICh
CzGNoiPUAFXFvaPw8CcXo0Udv6ULnC42SH6cDbO7qTNUffE0RkdFfzCIio2XbVWm
Wd0WGGKx3c9aBKjbHwZw0a+GRVlt6HriPplqrC5Xul9hXIkC9KZYweFWluouncA7
zrBDdMA4VTh6La371kq3QC1WNIM//VUcHtZMNk43LjLpI3HzJH5u8nmH2o1caxVo
MszGfk6XnXMGRT1teCLF5UtiFZ8D90YXk4oVHD2W+FhORQDz2Bkin4cwd5kOSTTx
k3cIccOz1+W3viOltMRi821hRg29A3+PrwfvxnUj9mOdGUeR4xA0mSovx0Ky8IfF
MDyJFPFOKpD3wYPBX2v2bPRV9K5McE//eiujfu0FdWHSUIwyVUjocQGUUBc7xHsI
dR8aJiSb+2zgJv/HUUe9g3mMnIgxq8uBYiBuNT32ypyaJt24sgfuTYk4iLH5EtOw
87y/49ns2XIshOhetP757xIlK3kRFKZjdpXGi5Ie6j6yKbQPYjKTNW/kUg/8Huc+
WSQgr+yHJegjkXVqKeGOILo8QCqLuz3iI1mMSpI4zfDuWOwMVoHtg+QS7pJznGwu
l0u/Jf1YDPix/8NxIX/KPfPfQ+Cchqxe11zCTEmJ1D7DVAJGco8ECOvk38gm5rCm
0WZ689UF/TO+W0IIPQVobvuNGbZKDZh0k3iVPMyKqHUIzIb22XCane0MNfXOR/E3
CYbJaAjqDW76ZdpVQtLe/4mRjbXPbG1JGbQV3dgEgCHq61vwcSCkH/ej9fo1NGHt
ESHjXggpoa9cP6ILtpGu8cGtYDWpDtA75oheBFlVI5YbVMQFG+pGv9h+QWaWywvW
GqJFPRW5jWwu2wIS8NUPemRaxBW51Nql5QSEJL65lMebt2XcKmIdGqe5ajmOPsbp
9MtpFt3+DRL1/gJhllYik9XGXRYC8LDwgBMWU4dkkVej8fpTHu8Ibatfqb9cpxa3
fjvrm1xVnL/Z/5ZzuFCiQicm80iy/GMF1j++MxtAjtFnKpasLfNKZyP1XGUWcshz
0Dw0TpRkN7RhuS8/3Yvvg9mXJ0TAsd/D6SjiOUZNCCGNLPde+jVA2npcc0gptoPQ
BGXU7glwfuqc5eDiB9qvo7QgrIyDQY3LcfRIR0B8NBS3AVpVTB4ENLjMWMq2Orfc
DoNHT72gZhnRtttOmOMRoAbBPYhc+KLpJZL3s/0yP8xIsSDvm1+ihJ30pJRi7syb
LmF98PZ5L3p5x37y4PpLv8xCTAJUdWuy+qeOr8owi4CH30Qtjke1OSejUzXiVlUL
TSEv/3c8rOsA7sq4zWlRzgRogsNXV1Z/EDlRx+8SMvLG3ZR5OjwXrbUrwDdaWxom
s7IiJBSjnFCu1iYh09ls8sL8Llb4t9G1itj9/0Gfus/8iq1BIXZ9dsGJb2FsFSJk
6sF2xMK5xEXKUEyE7oeOVbbRsWS3hMY5LD8uDGUCTQpudjI054x68r4ky/3uXTLS
OMfiDs82aAhmUo7VGHxAugxcocOmJuRObWcSk4wiQ8zQiXnxOZjPPNazdOhGu5ZE
Np6CnMG8sAMZ8p6cNzBFdFnmp1+loqO5g2p4LmcWmFgz3Y2xYUI/YaDej4b7C4Fz
+9ZNmukjk9cOEEMLnEFXKXiK6Ca5aUaS7239AxFc0SkJ/Gyu3blN/J9YLy02Q3D4
qYejQs7ae3NTe8aQ75fsOt0Zhm7M+FQez9a9hUS1VtFMeqp/9c/qTbf3Tk92RFj3
iXyfaVmSwV7uzcIWvBFYaw6BmOKT0lNk7ifWnhzrAjxQmGBFzCbIcbR7Y1lgjK4d
DMy199b4AFKpJ+MWurbAJKPF3EB+T9TgYavXfzeKvOGcAjcvRFUdJSspJ+C6VGqD
wrr+ctWrlfS+pI7mtFhjR+lKH5JiXITjN5ZZCtIYQdT6MKwReIsaPoXfqK/t3bDc
RvDJByUPh+C1kVmcv792UA8G0cmt29MzWJOR0te1OsHGEypXz0hueMkFXBpzwvkX
9blDUsMGTBi5ON98QZtlNCgB//OMKESGIFm9OdCALY/hdKdtrfC/m7dnDl91HIM/
RLyma7ycvcavFq0eSY28qr4dmkOx2LJ/WPlvL1VJOe3D6x+CKXiM9NvY3Th0dtCZ
mDatcTjFJ8zDcMlG2ouVk83aDrhYotGWnUDd/a1FZrL9VhTgDChtnM64YciqPc26
rjx8AXSAQgnNOA46dAlJfn07UByCd/eejKcn2sr3tIMA62IrwNPy0kej9I5HR1rQ
XBny9K54C20vTnMaMCcMQKPk6A9951OuxMChZq9nLnHq3Dyir1qBEySZfePyyAB0
jirlwD8q5D1iOJm6zpSg6/jpHzfTR8s33CPuDER5bvutuG11GpIFEkRtYNktaHPe
Fuqzx9tg6ifXcXKwiszLZHgtIgwYKcKVQ3hggJShf6zY8zQ96OpjeAUBaICrPM0d
lX+Oi8yF8Ay68CrGPffXWkwcru6pJGJhMcrb6TKuuU+OyA6BjTapwaP5wIdDRFQ2
J/bCpEhK8n0y5kyw7GSsX71Xyazk0EP5wWo+2k9tqszp9zaaPpuHs9AVAHPzpsco
hD+EtxJKREQcFgy8tUPv6h6m6FL56ANV7tl7mjSQbC7H+ADyyEo/KIycR/h4xyMi
pWB9of31V73cQbMmktGH/+ioPdKk4QX8zZ90IHKRjgtJNXba3t+5+KtKNIG16ilE
u4Z9WPflbOWmZyiBvnT18aCkhSugdTSiZaq/DYvV5NdPPra1RRQOY38jhKl9bZvx
mS55Wj6R2nQVLi/92zgJrp13xtbrTttz3yQ9Rh/HcK5iLmu1mzigc1hOmLycuKMO
mEvgAE+mj0RSZJHdXRD4OEVW+WfIfkNbBxAOnHuouc8N8YDuREmDtPeXMNZiodlY
cXrCX46ApEX7Z/yjop+RxS5rG3azzNRPyq8KappIetw6Q9/EbG9gKJAnSlYQwQ4g
iFrB6Jc3bUL9cQb6EaCWrp/fX6aIfjSkKvDa/YqHabq+K/tEd50SLHKIDrWwckub
j5xN10FLpr5ghCoMjuNA2tUcAZlsDh/DiL25VnfUM7Ryb0R9i40htIfJQ7QUIom0
m4xMeRR3G2QpoHKRe0pNvlb8AEO4FIXLU/ny98HBE9QUCZqTSNo2sBZ6wVVG0N+o
W6ZcPzk4z/wi5K9v/7sIR+Hba51uPo0ObJtQhX2EOnm+YPZdl0hWjS/Jfu1PC4KW
g/di0FKV8Pg4RmZRFxaI7Z/DDE28bw+ix++bAf5CWsMP3PVJBm1AC2U32fao30mU
2Oi4CYAOuMkGLjNmlmT5dxqUGAUxSQO4QXKD5SoWeN6VgjUtsmjA31ljVg/Mk34N
e2hAEcd8etMX/RyYSIQasbMLg280FKon1wbPGfY6WEDl72bbAPlIGj86UUxKDgbB
4/2xI3x6yWEOCDwiQlUWqYL6IkOYFJxZnCP3obEFzIuAyElMxvFCxfNPO+ZRAuSI
KnR5nMABmsIKFOD5if7AwBpNKQYQnHZa/P06zh5dVpjpL3bjCFxa+kDw4Gp+RrSi
3V5u7wrldJkoAWhKXHYzWF5T37Shp5CMahyr7z+JO9UIujyz+XDAqUX1T2nchYP6
VOLgd//GKZsbB3yXml9LDDjNnICK5VfYe36TynhYD+9MRLQtSUmQK++ezgIjejEs
/U+kdMHLZ1uFmyfa/YejToZpoJa/BNIy1yUirWvJVjnwznn4+kzMgu2BzpqHrMi2
1YtyCSmlRsMF/21aoRAZczlkoy7uTaoZVOpK/+eyUSD26HtpEwLZYcPeHrH/uPb7
iScrmhwtnS4dJMTpkCNtHqulCEXKUTbqoCPR2Pjre06uDSrZ8CuUpcL/Q89Z65A4
iqnLw5YxCOmu9XrektV+l9qIzLrDQ8ntx7eiHJoxglZ3TWn34578llMTDpI7YRnW
+OAJcFqj4WlNs6RTIKxAPxdNVth1zhfw7ra/VQBEBccHWQtfOCYcPfeQ4iwHeF7E
K9CNHummSFxsPTr8c/O8ulC9z+wkp7BfEwYiw/DWSFnxPaeWG0Ob78eECNan14Xk
rQmPn9cG4c+TQ69oBRzhzVan7cKNyEpVLUCGJNEni404cU5UpyMlgDkQvXlFyQZQ
7EVS+NLGSgireFivzzjkcWQ/WgC2jgKAHQuk0IZbxxPm3MnTi/kqhGzwPqXlGGk1
LYjawBKMavm7JYllPA6CkPRhkp9e9V+UwhOWGghXBbFUEJvynEIFzjBI1HoQWpq+
qY85bPiYsrmPFl80j4Bku95wgpSAD7dRx1GZU0imoyqDitRKbHV5LskqcOKWFmvK
6H9tWZGgu26vldcZrokLOjsi8yZItBEL+Jar85x5kh0FvQmB30ZZ2PtfQ83+3qED
wmGO6vGXHZEZZhQiOkBfTVZvS5qWYF/1hi3yutma2iz8HxquRmmhYh76YcdPWsHR
9dEt/Lz9XmOamQmwx4Q3LvOXFssgeLaA8CXkMA6ro6AroMFYtOs41tmLlgLJDjex
N0l89yJZ5aaww+j+Ei8AMb6Cejpi3byicFdMF4Tm+KIUtcqfid+k25ocx5hlXw6q
xf9IdI28KfGs/9AAZImOlq+rYWZDlVRADSU58sGJf88jsPpQxllJkli+t9kqQTb7
yzpZaHh36K26hHBkTa2XFOoyQjuN6i4nZIhYFqWYWITtxEW7R7PvY0Rh1XqfR6es
9IygpSMx42fr/rloelb9C02lpcjvfQFsswqJUOEMTqZVCul13jx3BjEe8ux3KrMU
D25CJtWWRQIcLqFuFx8GvYKBCC4DbXLZo7aSRAevKbjm3eX290KL7WlIQS6T6puu
zBdLluat/yVwU6LxVSLwSGyiucV/+65TybRAOT+gfoHtnMmiZwrScIL0aPkW+fOt
ZC5zAS6EP1WZuddPdHrUMdNInTq9Kpl4+zYex6aDAFlTmYOU00gUY3eLM1JLpM04
5203z64uSQ6D5Zi3Tg07ZZdvsXQENZ79JZhgdyXM8mQlzKZKRXgXdUUqMVzyh9lu
QHOgvuZrnmAUkdypZbbIMwUb1DW64DjqI16Yog3lbC0zj5QEl9+CwnOo83SqO2Oq
JJHVOzLkdnXNQdR6T4FuHfOU9/TOCiNDAQ4wL43L4dKRJBnhEVmcgdyV2tPWYaov
R9gWqainIqOB4BqcfbispUGkQ4z7Yw4qiC2CP34WQQBngK717TWG5Yy+4ZhVV7X0
w3AWSs0CdRIy5f2l3KiMcdT6WzwWiUsXsnZce6hyNTpbPiZHsp+Vm4MxDplERFJh
0D1bjx3QygvEB0luFlyQMC2OzHAWcBNWwBsIVvTPDk+MEM6KA5Lkajcdr1j/mqNo
HiKHCFsvwW3GYB0iWXOQeSOR4C8XVrN3mrbLbOeySR+H4slyRbeCVbArJbyLRPsF
OW+GjFkawkCi8NjxWhz2XLMkIx+qEDiiDY+KEjf2NsVu6ajo8Vkg12VSOR6cc0IS
Is/osxIvd5GCNBUYTvTXhA9zSb3F4ibdZFoKZUQDRHXUzptffSK/3zAIayMwXBuz
Npmic5NeqsIUKztij4/YccVQP9WluUuBmHgBhC0ROA+L6SfEenKz5cbyLZHCIYsM
nzO/MlezlBI01AwjR5BlbprlD/smFgMwvs9ghdJdbPAlRwxGpGp7z5QdzazLT5l2
Xbl0lpHgCdK2uBwiOnZtqivVRsRrWaXjzWrPTY9CQN2bzlf/rTYDUDKOhdlivrwV
FBjGv6mIPp7w11vEo2EL2wDSSERKivk3hEyhiXC5qxQg7K07piJg4G+9+NB/eEMw
Py+2uA0vFO81zHqyYU3Zccw8FXVkn5EaaZPGNAldJUBy1u3J0LmBlJIiz6KyLCIc
vPU0/39gjMpvANw/QhObxIaNrup6YZDXbYdjavi0Ofdbcpvfay8W0BUGKjfuM5+4
l1YfUiZl1CR5yx9uvapNAjPJX5hFPESVgXQ4Wta6+yafsLzum+72P/wGDwmNS7ix
Qrveg9Xne0NpneRqjUiQgqtG6AgbgtRnEA6MTmKJXwNvrCMjN0LBfWkW9KDwmRrK
xq7vmmblLuB8ml/mclE0movoV2vkYWEkZDMM/UMsUD8EtJVO8sIGV3wYFwS8Dhcn
ct3HZUMONBCNv3LWcHd/mdPvHeclg2c+mtNlC+YwNP2j3hsxvNC1ONCuYfwuNiC6
f12XKQ51qS2EByH3VanTFfFE+UeH5xaz5wRUmeVkQf4CBnomLevYk0E6cO/j9x2x
eX/i8XC3rh7mwk6t4L9sBsXt3xyazTmj6KgQ6xPdl68RpXQm3SJwVD8EL4LB4J0N
WRDElCNwUIwkV8vU9NMlSq0cUsrHQ8aPPbveA4cZ6FT63tYTSYIt12RVQkMdYu8X
N/nx+CbUmHgqFaY/Yjd/jIVfufAyKlUW5ycsVtPYiIqtAFarYOH39t7TuUjNlnox
qbuc35pON/nX+UCYOG0DHEjIVSPNH6Jat+ymdl6TvXyB1/YUylvk0ABYeDoNMM0y
A2CaSbAtwjHvgUyaQemdr+3z4MW+mG1ajsQW/EZkT6aDiVmoTi7MSIpZpAMZ5oX/
pSsD5YEuBk9CXH6aUw4/TQ8cn8+QDgqcgZwk7GcjG5LjBe0hQNOZovcpL5ygh9LN
0ce9+dUD6V6YcmNr6I+EBGArd9f26MN62qoMrrvT5IFxHhNFb+D96qUrF/Ri1dxk
tuFsKZTrQLtwNLBTHl6mXUKS73eop8OaqpaMLh21gVK8wnUi7FDwXZBMBCP636d0
rytuCoCt420ZAwqgnCECT974EILdCWH/W61JMaM6jfI4o89ilLtEvAj+JWH8rHVL
HfurhuUDWuF5b9H2LkQ2Nr0a482/e2pzrJSM/nv8R7O0nlw2RIwwt/4SkqZPKbnQ
fVb3T5pvuBjVXkZmBy6+RWfoH91z6RnK1caaXa1o9OCeYi9+s/mH1xLXELx9n7QF
LEQHtex+pM26ZFDpnLBdo0mgmLVZ7r85b3u0corWoJwQF2sP/ebItf3W2LHFDI1I
qdEI8bnumFWI0WES0RrG18DjLIlHcfybpKkaiyRdlGYNAlAuOWb16PN4jQ5pXtUj
04VS2RC0W6WF7cDDHv3L3xoANYMHlVvMlhdU8z318Q8qoygTcANNG8NHAn0nvvBe
LBQMdpA61pAfqlcB9e2UuGnrjKX1d3lp7nWPZmHgPRArg/nzgRnDD4Byhro73RLQ
vYBdR4V0O39lWDxFy2C7q0XPrzd/r1jr62VM+FN3wZcKUjNJBLpUssnkTCb0/AU4
HX8+LHuy8UgPjwTI1KfBpRPlr9wlos27uQT2suHWSIG49iYgdbDf+SlI1V33R135
hoNqqZRbyEQ1p9Tt5BZUCTo1oicgpJ6fNa45J57r/sYej4JFeKapBLsJvviRplQu
wiwebPYjWQYfFP09EUfm6x9TcNMnB5XAnLyA99OQzCAjtBnnX4GSrxhi5B67LTxO
KUDyasv/0f4WxOG9rhD7EvvrYjHL9qq+3dJwEZlb3kq7kK/s1ICMZeeOZKdzneSR
eCCeh1AYpHXvVovsJSW+WXHmTOwHX+HlNDDAwVnI35Zt5JjAvvycyLC0AM9KgKjd
fiCdqBoUruFeB9jrwcdWYPKe6nCxR23P9WCHCttd7wJMHyq4EI/A7LSncuXIOYoN
4lx6JiPYNUgLCHZadsQ3iE6Xx2akhfwKa5UakSME5u+LkpIi7BHg9gSyxoLY/Lv/
EjN54eRblSFKKfyUwKYFMG4z57h+/SBK7kiWfdgaLpH+MZhvwW5wFZXW9aqApzex
tmKycmHFzEIVuBoUX+k5/4KL7KaEUUcj/gEvrMZvaXCrf4wnh70G6yEsDplWIpHX
IQTmckun9PCfrznzNpr9ji8cZqRAkw+MkKhbJyRaEH5lUI9kwT+vvGvdjPw3lIPW
UsnG80QAXYQxA6o7oZJefNllAPR+GFIKLPFdqyQ8sMYPj59yoDkYVegYGUag2gBd
VvwPjN4spHXlj3Gpj6o+Bb+5p0t27b9brXlmqKJ50W7vv4vooaBHt8Ez5RHC40dj
u5z0a6UUL4DKbUMhj4rB+8da0Y83LpDjebY6EwQgOCFkmdTXtV3pThRr2AAppwfV
YnK2tq2LudVOH/9pic5DLn1kbf95j5sXREn8eX9Rwon2+VqYAw00uJXi45QAiWhZ
d7FDo29Li6lyoy39wrz/XA8w0AGyYmX1ADbcq8pUzWpwKkNBF4qx3lmgrq+ow19r
A7XbDgbjNXKEdwlp7e/GlfoPdRshMsScVblzmZ35+NDOjqdpR/oB4kXr5jzo2m3G
7g+FDGiSVLfdy3OD4mu8RO9xnMxWBaIMJH8ZnD0jzKraPwjl93i61vD7QvAAXBHe
uGxT5fw8VHRzEZrK3fwhttc2cKwRjP2xVDgyY40/skdUHgOOZzCS/hiAEJ0yqebT
T7B4jPYRrO/TFs3pHEOzPLNJuZQnjR6NezILfBmCvQHfa2+8oixXupfARIlAzTBN
zQIvVm/ezVytsJ+KlxX39KffdGD5i8FZ9SRjwYIBnVsFYfcYSQJnsYb58Paf4QfK
kyPj1ZXio//7UYs4zuDYpBdBaSSfL8y9vybYjnAemHge6PJZ6AV6rfPShquX6oTq
+K9A7sRJ9zdvUjGCCj4qI3agvnpPIdL4/Hnk8RBWbhBm2nsVIv9JkxP6TNuv/L7R
bqTDoHKhRPnJVccKWywCqpthhhr9/26q5SpTIXLJfOVagiN5oi1TwsVbJ1cWLLa3
pv+nthrsjXAY+JsffKDucD0JOfn94eqXxuvPn3yCrcd8MZ1lzOVYbW7Yyqj3cHPk
cJKjXuaFdn2zK5EfpbhiDZfpnvoVsIpq3/1oMgEb+4ilzRf9CQNWB3bFv7bf44jD
NFYRqoM6Y+0o+PlF7hi6lY1Q0wc31WBaWOUaL7fHWTq7nZYFv2OL+4Yp0x8T/1Gt
0BAYZmYJrD+1LCsS/64I6y49/AYuI4t9bUeithtSFefnboxzpDHWr9/NGkDKWFQg
LYpTo77u46tZKT92fQmtsghSmSeqEvdQZjYqx2VupsklcEdoQ3wOem1pe6BNkHKb
BeNR08v1T3fLUXWHf53bWOkLA9UsEOHvKg+WwsUzYXY+BBzymKc+uLhww0msCB0w
hs6R9t9sXYl4bhyv1JW5Z58rrmrHQ4dKbCdTgRMyEUBIkpHB8JYnsrQzo3Vi1tda
QVqJsc5nm8wAZHyptvjGcHGOKdsoIo5fZJJHHfgpLHuAmEQ1xaq7FFq/GXKyoRLF
nsGsUqyuIMmOoB1mTch2wTtpnTRn0DyphyxkJeHOtRygdftXnWavEf3wzf5JP+CJ
/eYGVwwogf3+8sWnLFyuyMIZANkqoVRy4csWigQx3lwsL05f0gNPL8IAHvfjIvXq
/Qx/sJyQnvOzqvvTiov8AIU3XGdhuKM62sQU5nuhTzVlCh2OVPqbWxRP1/YuiJPW
c9u9NFhMrV6PrFIlq3LD05ZNyEuhIQRsZC9QMtLdV+PxVMQFfgMK3YVveSrQlK0K
rZlC5xmgrHbdUil2WssDECsmP8uo/yg3RGkRJOBp8qr9epkcpb2MZDGubumpOsD6
9yBrMVNF8p+cUtrYkR5YYjjtSmHWFKCc3PF7Y3kTGPbtDBlk/oKRPSHWaNUqrPNG
EDe281+O21WYpLTt9Ikmqz76AUg22WEw0xRawu/hgh/DWxwlZUysJmv5rrUFE7fR
5vo3/jhqKk0IxbvVZkBX9g1OVatEGWN65Z5GPEMQOYExiaGogyzNrJLb7brTd0XW
+/QUl75zhKi1tqZulnJzccsoeBQpP5njR2iR9JxXvhnkFZ4lUSovCBZ2SUvj2an0
jSicWlzFD5425Ngw/Xz3aiqKJ8z7sF6YaESeHwCa+2Ttv+0r1xmWKq1CZ4rvxZEo
ieKTxrFUo4/YGxT4J3jq70reoEUhsJQD01/QBmPi1bAYJE2GsyeYt9M0p/q0qKZ7
6mykTxVB5JO1RcfDzOt4eGE/H7bbrGX0K2zyajnUuDkHx9JG7hjYVfcfyw67u0pK
9TPoyCEDM2HUrqh2h2F1YcgNH+sCvtn+AE/JV6M49pSC9gDYjCPBip3IFRfgZiLB
DuNBvbDKjCpZ/1zMTUtd4MHxEi/ReqDQ8p43SNjo3UPiATC86iHkh+DSQusAVA9N
qgexOvWmTsSueU/q38e6Yz2NblZHSecT7k1mX5C99KoLaBS0RkL/pc44TUFhVtqV
ZouiERVOfsv+KdZuh2VToEY1EqLUjOSRlWgwhtysygN/5840CCnW7dRYOU1e/pMb
V3whIGZ+LY5Jd4OC/Q+kYsFc1FS50dTUnBOZYb7qtLuqfTiy8U3O22au0eneEBVS
a1YgJe0yQ5M4WoG2NgcvTBwGntxQnZ9CM9EVuBaAjH0SyOULbZjImA+Z/glamqAh
kJa9i/2ELYVxCnOmVtHYqz5yYOJCJGHY3Epw/zD1miN8xbKrvLF2AY4FC7ti1P7W
8++cUxKti4EvfMQ9P4KZww2phs/6AqvDJAHnIn7TcbS1f6VfrgUye9gnIhj9ZCEi
9Gqxi7EY5gtx4xBSIn+CJ26hMUyZ09XWza7CZ3eoLuhNecT1DeDsdWYj2XFv4BQv
d5h4kQTiHjgi1G4AfE5EztXzmK5NTdYB1UCP2hz4R59LyAKklP5tBLBsqk5LqYek
RS5ak54uU0y6/KIKBdWsRFfOtKZsyNjW4qC+LWCu1sU7BqoWoEVYucEWty13D7Vn
CqStROIX8SlOm3BUzX5yoDjAPumyT2kFcViagGnyXwCmKNJSAV2lZg6orCKZvePo
OjRx+xGithcNbUuqHuV32gcfRVHAlTzq83fCmBhtOjU6PXe47DPALm6GqDJbWnK/
Fb6AV+Mvkry0+TbDUXizRbys1c23Z1shoaTO482rDh+9s6a0xz/j7PvmOduwJhKU
eFobxl/VZRq7G8rXn0d5uWL66GZ+k/GQPXmxFso01gwH+aVdiqEvQi/PDuiqoibY
lyGmf3k0az8oLEPoRtcukPfHpZUCr2p/9WUlI0zyIpzPWXOCe4Oc8UHaGpJj0HeA
zbPBQdz3j+XaU8kjWZ8dGTwL54F5zMkm+SrwOe1nJZJGmR9HgZmuqg+gyHOwYWJh
Uybo9IhbcWtypHmSB92RcFACVeJRcaQaubDLbapfODfItfpERx7ZH879eH8oYjZp
8S1iD3U1akUues91SCoMDj4otPlgeEf/oYONE/M71E5eSDl8TgMqPHiTap0XSUBv
fHP6hdcuau8u5h2jnOFWYaVEKUXm2ANXVRK10J/k1+aTIh4yxOKRkv/sjdVTOXf+
mEc+FCXyild2LK4M2JTT7Pqa3EfFcnoTVoDOuNBC2uTcfCINh5FCQPTsQytnioiH
MKpo1MpXl1bRWisLyvEmGRsbHApLPDCPY2wZm5y6kLj9cSzG4+cqd4QbZ8tFDxF3
NytqrAek2d5CaSB5o7AJC2Ey7HDYNqSdHfGHkyiD1/KtUugFhZi9WGxBYRP5r0k5
JnYdOj5iC71YLS6fPL1ZFp4FMQtwmF/MEUjCuUjasu7FA4WX8h3QBbdCyun+1k9O
2T8XYxNnKhAk5pTCZndC19PxyjZ0/q+PAvRIRvRBEKuZbZ1znHbbeLCzIdgtisTq
ED2KkiEtBElywEtcRg56Wy4vP12vZFJanu/AlPaBGm7cqe3lJh1sVuAMpRzEP041
msc6lQNf/TL3ZwQ1UJ628DZZEzxR8XsvQ99KrTSs1ZZqrYc+zi/F2KMEigMM3K6v
F50OSN9Izf9xh/T1JpsRgtPsEu0if/7voEREM5HCzKS0iNXZHcflLSotRX0n9HBl
1oJ8ruOsmNoo58x2S8utMX3W8VjK3f/474mHlA8TZyL/IA384aTDwSdGeI6D/S5f
60HGnMiwLTQ+SPsActj8zWD0QQ9321mddxQV7/1Nnv7R8rHOME8yLZa2Y9Y71J01
L899illyoccBupNYVGLVJXYSjl68y9KbicZ1g0Fco1pcJEcyqXW0B+My0+6CTAq0
x857EXdFJlExIJLlYABEdpRcatb6+U5Z5IrR0Bw05O7Ip0ecH6NWVzurkkRWDhzH
ionxxr2kDiMw5kuPcPx6qIaYf1gf75MW9itHHDxkMEkBHg0WN9eZHVAIvt0YEjf2
FJDJhirS0iarB4Wl1KhDAhGq/II4vn3NwBA+46emfS9BhzxiAJbbm3m1jjK4UtbO
rHnfqZ7OWz8/Gh/N9t/+YnfVIYvpeEVj0UX0VONKpoljdxvzm/AwRAltBUU2CDmp
paovJ1/RIEkhKkJRBU/ZElG75v1YLSLW3fVCPhfX+aopRkr6frylpHcmPjia5Csf
24gwU4SrrvHpYNflH5Bz7I9E77GVEpUuFiZSLb6HqmtM1g6oqkmwX/DijW54fu6+
z/mBnhGetzr+akIpXsK5uELOY2Pi7wSckK280Htjp+0ToDxamiio97TI476zZWck
yceHefVbxk2bnKh2/oaQD2jswQgWHuZIFJMqtLAbiwPputafH8pHCu7UIpSedX5Y
uofQT7mnPp9LDxXSFXMX+djvN2kQDiypmju9RLTFdd83V+68UDEP/pVR4e3peRM0
uFGAHhCz04SA0pjHNU0MvT857trEJwMl1hrjHJ/9pcpGqKs19FLOibuLgxl+7L/6
7SPcnclqZDul3WUGTI7zbKDn4aNyRrj5PqMTKFRGfa1iynwew9G/xXHBhvPLSzde
FzXSV3YelQ6XohaDFG66ZsI+tZ8+lF9+Gwj1ylUQnyjFhxs3bAeBN9VmhwL4WRs7
QZ/dZo2nnK6HyCkl3sYeDDjFQEUmB5KQuslinG2CAjT+j6lu4HRpI0Jm6Qo43wjm
koVONf2jaz+S7XWGUDzHK204h1zQpxyFYpI6/uzTCpUUqv6gOUebKU1r8r66TgYu
PvGMM2Dg4Pnq5uEAY2as4SNraVCcj2XCjl2Mjzkw5ybClEs1XTU6TNktcb0gLghh
r+NxsakUkUdyZSJrU63C9mGvwhWAh5iG48cR0Lu9T3iCryW+dou2D3q9/BArl/N7
bcSyH5czR5H/4aXo83iqFkhK5Z2ehuD7UN5QC9zPQhdZrHcDcoDtOsxPVmxFvT7L
Bauu1ItaKjV4p3eIXTOPUYzA1HyEv6HdrlHu3t6gAy9y8AJzB5A/MeeobTM03DYQ
K8ecphk5ts9f4LvUD/D7KxnGHik141g32Z6aAIWh+oGVm+tTBDGCMH77mPq12Fy4
/azHn9pEHv9Ph/HLnDa6R/yAVEAukmiV61kggSp/1FVZHLJnpMHBZ6sK73Tkj6YE
gBal4DxCO3pw9WmvS0RyMTGCq2G8SnRvpzV08Dvm5ad/+Ff9ZPv8vjfEUyFrkr9Q
llY8PJb6yXwctDb36m6sZGZ7hq2ucp4W+dYuD8XgMBXmQbqQvbeY3avGUrkOykCz
5mh4Q2I3iddFWkSUAHPTp3jgsQ1jwq5qPzhEXoj2t7CzRjItV/qW5bhEcJxoeSkb
pMt/o0KYh6XH/efrHgCtOci7uFhyrPTa6ZJOWCCwNtMdiYxGJtFUA33nqO423gGS
Vz1U4FoIzh63SyC0l1y0Qm06dZxDaPgAK/ox80EU6ulO/47p+vlHErJrrJqKG2CA
n5YmfpJNxaHDZnrqc9FuVezFo/n6t96kwi6/3CTxGW+j1Q8qaghH00RNlKJOuged
yEdRWw3l8OUQjmDdW3YQfaosc5c3WfU3LEqJ/p9TELyV8tNhKVD1eOeXQ7cUqPYH
U70PDlQW5gzxfHTzkktgK36Aegx0ERtTHSs4TguQCIAT1EjT3etWZg29/DVB+nWX
BXtYIVDiZSUnFcAoZ/wAdvFlPy4YoQnP9//q2Oi5Js0pSZr7wj1JDr93neoNdBgz
WHBC+nDg/ARh+RxJIVIJUW4P3K0KwPgkVyipVT0uiJI6eM/jbk9i9/OFNqbF6V8B
EdZKscauUrH9Q9G8Tuohfpy2+c4nvd0WZUYuxfHnEc+zhSandRZviYgYnr9T31zN
KMuWl1lZNACJsPeicT+uDDcYY0K2h91DhwI8hpBe6zn6f1rIl9HIWmNZizzBO99C
7GHD5DHavy79viah2K3Fbpg62A3pwuvG70ZrtgAGngEWxDVE0ybhb1DtiSVriV7u
wuLqFaZiLKZ2p82XwomZ98aF0qcDUaHBmQsQNM/x9ndItLuIzQVjxD4fIdPmUSTx
4P+iK2UZpx+JZXQRMoAUSLlcY1idphGbl1CsdtmHnJSCixkvrfw+0jRpFVChPgM0
GZAY8QgFh/WUqkzFL9d2kbk/szGD7ofdXfutqKBlCSrzjczVGy+qhUNH0jwny2dY
ObKmrhavk73YRvvxYf16XFM6MAGUy948qpoVr6x2N6Sdr5VBIL50a1p6Sgg14uO7
SKXq2VgTHVCXkLMkNo9Yg16X7N80f5lXtGnwwEDHOWEQlCr0n668YxKrdNCpHiqI
z6SCaJbyc8nLWyn14VlLq7qeNP0521v1ARKvGXY2u3YDDPBgfbzeysNsCKMOTVTE
PJs/LccPVSesuCjDBGzCHjPppuJLuZ/QpG4WailsYx8pM6ZxHD5zDAUh2Qjpsq2x
TAAlTWp2TpCrMXGB2fOt8UHyS3TUsfmGdCT62mNGyD1ZWcvyzXfP+dAhSRCrL53i
Jzrm33o7hj3l5LLLok6wvlNpt913jlEnEMu9KRvaBFHdNheVlWeLkuG1/xLE5P2y
Q0yRjhoaRUoO2C/JdzezIWcy0m+XR7VntCXFfjugLGoLiCTvIZ+JT4Vtoim7jgy+
doG4dNuH/FG8XB51Hi2DiabbaPKSfXr6WdE37aNpNl1iHbDDZg22wOgN1z5FQT7/
MUmUQ/04/Cfqv1JbegyhjEpJS7O3nDt079htodAPaeItiSIA6wA/lokdLmJmZ4QV
m306AiAiZYSvqkBDC1cjey44djWK+AveutesjvgKHRHLUvEWYZ9V3TFU4cmxwsot
ADXbCTR4zROEzSDL12MRtRSHZtrF8wgAnfkujQS4khNEYJvCwFl73wDr3PI1QJ6y
Pq6hPnv97JiCFQgsyIXaDNhMLzk+hOcKtk5NsE+ViyjeZtK/yfHWtXdD10CbLOcn
xGKVjUaP4i0cPGsOA3nKRb8BjlHQjDHvKApm5Tv7V0phLOdchkgAQkjc/itqD1mA
ygTg9og9eDf4wU/AICbqS9gPj+m6gtq9d9PXNON+LQYi7upnYhlo1UGDXqv8yn1r
RP3K0ddXv67t0McugMi0VrGa6S3jXLKpVE5a89CjbNhAs0Z6lUGx+KYsh8P9ttwd
DgxzV3XIsJtexsDPqV7GPMEpmf5TFbkEKUbQ7qDxvE5CjDT8AKhkAtHT5mmL3c/Z
Y6Iu7rUyghq2QTMaiHi4khLqa8xaMVMnPX9Uw4AiSa2gZUW5JvMrSjQrDTQGA6Z2
Xdv17kuQRDiu7Kx8bH4uAacFyN5IZWio5XRbFKEbs07F3UXm8RHrPktpVfKqMS5Q
U5qlHaWTb8DwyXcJ1bO2MVZ0eRqYmnGXDEp2bCNn14wjRkydyqo5wXb9fdhkAUIw
AdnbFnmAY8PwQIFIbJdFpsl0L6UNWAfxhfsQgA+Rvfb0w3E12gmCmY0huq2TlXQ0
aibRP54kQxOJZNF9dSa8lfO0pHptyUijy4RZymHK8hYpssrO7OBg6g/joPEMMG/0
4G9U+f3FitFqwG39psJ5L4yfTnoeFIx7wQmhYnVYCR4sNe2O+UaQ9aAunoU8uuAE
+b5CtPN5bn0eFjW1584x/BZtK2oa/9KrMjzWm5aqCFNFZ2AagNeT8konzvpSsE91
TXobC+1t0jWTq8+Sa7GaSwLbvuxU4uQcwBUK6r1yJ95EGqUT6ODnhn3Tyd7+0GJo
rFQ6sPTUK3XO2PbJN27rEYMdoM48u57TvsezxSsmRUdF9+CcSKPcFgDzhr4K6+HA
1VvbNUsZtwgG5WWvaITkVjetw2YVHwGfaD2JN4pEUJeA4lq6TUhydDyaM0q9miUK
8ofTBAx2vfTJtKy+fj+pIDyXHSBVfJyldzP2nv1CuQH1QEYPG5WWhKbnANss7rFG
uNDcHarn10T75wgdpS/iSVYtYEI8uPGh/eBdsmDyzqnvQ+AcmIaPsBvGWwElGus8
4BFJY9z1+t32fPmovFqThH4Dgg5xr89S5NSPXCqyvdq2/f6+VhxSUD1UqkJ7R6SM
iB/CFyOMTbliI3Oso6GfVuClPu2MjSUTBz6apPnrrPH0TAm70Kqa0zcH4k0tE1AL
1542b876TD3Yr8NlYCikUFP3wBrk/tQfi/d8U585xzZ+SkdS1n1Ji+XQTiIXwDgy
+ouiOP1zRW5MMa6lox4Lwr2B1q4Y5dpJz/vb+AKq0ZWBcSctm8oRruRyoyGHiIIq
R9Zxv1p1cCZRm1+tgnvMCeM6sqwxWRqjidv3inguJkjXZ+nMnjo6EX/KQGscDpBU
Hc3cGRUfpNIdhsl4u76cWR1LjEDHQODKsZyhI4afae5m26gA0u30J3VsRYH0tuA7
IWU+7Nivi3/KP37wx0eoUNQSHSS9l5ZMJF8oBecH9IX3ELIgATDGzEflWWMtKEO0
+V0INq51/v+li0FFQcn+A0R25nY5lI2r6etQEbuYbJzX3Y9Bp74CibPZs3qB8FZw
VMi8CQrDiranmpGFpALgzKl0H9bcy1LS98rBOdB0AMU3U7kii3rEOv+G+4gDSPO1
OziDvp0j58aAALs6CDlbP4dHP4wff7Yq0yhivxtGWkL7D0I0Te42tuj1bWHn3FSW
PW94dG1qZgE7PZEQ3zFIZAFGtuV0WAmEBReDrvnja1PjUKM8a1Mhhi+3/mIl0xTh
rbHIdF1jFxrkdkBNgchPdrGyAOy1ZjP02OS1UmI5fSu1s/IUOlywK1v6J9DhvuN5
qD52XMVNbbeNheQZFNtwU568RO0ODjfCt8NGArWKXB3dnamAOs8f/xRs7PslVEak
t9WKQDWO68ml5bWGjVkSPe14Pg6wNcIZtlUnrOzOQdhtppzJ/vvq6C765We9Bbce
sVIXwKn7HpXIufvG8p/Xst9VLFhEY0EomA4SCtS2+9QQAtfEjFntrLkLRybuiO/E
+wmAw+7DHePP6DLqrjPYp5YyeJj9hg3w4mDfRb1YSilMWqUoBnQSIZVWgvRtsEYQ
fN2cHIjLbxE0pZIp4TDyVDU9G0bYfkDk+lBAkIPW1e8bLoUvbc8mJ5FKxPGrIppt
joJtIbgKnaBkMP8rf6eYfQwpQaBKV0tuzKyUNft6LkkWybL0H6NbqVAn3RLDhZNO
TcjUT2S6Ft1RFkb4Lom0yY8tQjND2E6P0d8oZosTKJuSu2VnB/4oBMW/d6IaIq89
v3+LvEsXWugFhyrL/6Xa9EGgUzrMDAddSaCiDeI2o6jlil7tPYnA+YegBrNOfv3N
1cGyq8yLd+3G1ngbdTj4dJI+W5fjZ/O6XNMotFfYmmYUGdkqkPZ1YPsh53g37++7
TuFKnMrAiW1bEWLkg1/07wEIJZSp1HmrqHHKDzU57MzFZ3R+Mca/ropMqCYsoBSu
//C7B63XkWwXwvzSlj8FdqMuRboD4NY12jocz+/H8oPyz3E5tJN7mLlZLFLzLkvY
AB3RW0h0Ai0LiVqHcm23Mv7itZ9aoeAuKfmgJPPa1fb1J8Attn87+Vp0+0wRFola
k5lej592Y/pJ59pyGuJLycjCH75R5FWYz0LhcafYnJRKz1ncLklcFlj954RR4Dql
PC+b9+O3lks4CX+wWnS2PraclNWxqQ9W80rJ9ppo7GaHUsyiMkmz5ozDiGLVi+oA
z9AVTexsMUmYLW0NeRV2lbQqUe+Xtfh5busa+MBAZ90EZ4L0cfwaEXE5CKNEqktV
C6Ni+kMnmCFvMk4j77K7BXrrbmXr4vdXePiRarvvp8t37lmyzqlaiLE9+TecvlcG
bw3vcd9sPftFQm6M88oysSNodVNi9SoEZhTe2f1zubfrGi2sa5CE90oNacr9p69o
kDQWWzpuci209rdbwJANJwaRUwU6g6wrh1tXYZ0l89qAuXr5S1GeUc3WjrgRxupw
N9q3KBELD4KbRq4s42XHY1DkNKFPQTIW+pOMvZBTfMzVGgbtnr98h12Ia/g6QyYS
bwYP+swEEqidGH9p8eQFrDtPaiINvQpGivDau5EU1wNIfxvJ5fVlvczqTVwX0egH
MF09/z+8VkkbZGuortcRyOWK1J0e2iKXiA6r5Lo9tAML+eGkeiG6dCaKmvppTVTV
tGkcnhbUrgkpBEk50ogVTTBVy70In+90OcVWk0wR4kaExW+qmtZ6tauX+kqI/oKE
duotb0dpO1s8YosBWIdg2fiz27hPiLvckDLPtAMlycOXVoOiChxNueMbVi+aXMgD
vGAVbB3wZ2IUP/TnHpe1b7U4F3NKNdVrfztYX8PDkrXNGaje+8rk/eUSF5YOpQu0
+pb0CqFm2SulDirxtOvdfOa+6YzQcTOJ6FnrupGd3W/q9X5gANZwt4cJ9SgU72sj
usAn4JwtoLl+yk6PxTWd/xkWc9wOucp2S7oBnxTka+rEhwG+2rXSQxBy4HFljXMo
o0Ta0esaYwRHTstrVfYYY9g21WYeWeMMwTwtjYmEunzbJ+z+UlMRv2HMSJHehUqp
qdGskpdLYUPi5mlCYGVNpdXcohW4vk4IFcjapXIVBDSIz7rpfmCBw2QnXI/97IhG
jC+CnBvcXxKqYMNWaqK3Xs65/lpIM0jsYSTmNCJOn9/nRdwejnhtEd6qX3zAc6YG
TEdc5NrAY0w4oMp1ZUuQW10T43Jg5geVBkQhsqb2UAmrtCH8ATtNbnA5FfL65/u5
8GumPtKR57TnA7bAoKw6j4lPQ5+h3eVlweJmeXLUTINjNrgAqxJMOJDHdqzKXfPi
3luWyJN+6g5Agomc3Cs2twH74aBPkcoxyjDO5CWZt5fEUWyRU45nvdthdHou7uQ7
+9jA4b0HEp2VQqFe8s3GsIevnqgKxEfTmVaDcH1KTSP4iQZpMNj9T1W458LVaRTn
gS2mnWkJirB1zPEAYKrF6zixyVlOu+hambhvtlAolPTIDnIbSXZUC5Lff419eUpg
AI5cx6UuH5o4UF+gsYPj4G7ISfmwcUxiImUnOtff3mc/lNj2wyVkabVmea5Xb1Ao
VIgk06VBvg+qNzrL4XokOPqDkXRbkIXk/+fS70llWymR53tX43smQ++b0zr81o+P
xnSz17WoNu5wCwd3SrlqPDaZzwSxy9EC6mQXnbkDdAb0vBuOhlLHUzwghDRVzDI5
rO0FAfpBTiD/p/ZpuvpKCYKcsmcEgd7Sl+D59j4fptVww7naEyaT6zbLzEQcsHKu
3USa9ew0NVJPkk0WstpD7n7mxQB/hJDNARxKzrTV6qCt0VDDRZFnKSWIFWovwEKi
tk020p/0J5luDB0QuQ8I0eLrw2aBvcQmWkYWX2rskMtgxMtwyesG2oJPy84Tn9S6
fFxnRPAE44Tqdb3IHuZrSkZui48USKqcywrUNiqnzqG5K7xqM62jURh4XYqOqETA
MCTuGi0mgJYPhg07ugwvkVXrx+X8is+X5Pb2vTTC9QUtx9vDBHJSYsZAWqqdn6bE
D3EEopEaOoji081h/3gdqr5xssGJgESTlmzlBqEeQ3eg5YKYWOnbLo93yIFfIV5a
nQtLrSrLOL0vdaF9OjMOSKad5iGH2d6WmSM3rnRkTt3JvD+gXroEPK2jc9ShWOoy
J7cnvn4fjzMbsjnwu/NxkAEv+/P9w3UjCDxY+MerG/8kkI3VjVwSClbNZ+mPUZ0T
x6zgw8yn4RYxd2U6UkkSZ7RDpUJzVy4bKFolxkCB+z03Nyre7IKWue6JssuRUpJ+
Nk2dqxnIEEhJSDd10GaLY/+htIXL2Ql1KmtmAyWQdu9AbxuhKuFuFcr9vLmXyZj6
4b+yPX3+lsE95xq7cDOA6DxVd7xL9+DYe+pe6yAgEcVAVL2fiqIBE4afcLyYH4Wh
7zRd7Dtr85kXCSJDqSA/VN3YIf/Qy0KdP6uClY1bvD4175K+h3lCNGAyfbtCvpju
OQ1q+T5xmzBL0qf7kUgyOxWBHimk7XVaiUNwY0iaJRYy/iM4rxd8SMAEz5k7FI9X
eIdFb5aPLS5lnMRoiMuikrCGtkMNwrIT+Jamd2opfV2VGu/EjAa0l0F7Hz3sVEJE
G8sHB0E7QS0kPAS9rB/NFWRaYrWwDhQjwjsGhTQPG5xkfwKMjZdB+vLVqblLyatB
9a4y3LzF8JdM+FJik1X+SESTtP9Ug1zxGyiEsNXmuX8Z4GPz/Z5576ru+1+mGF5t
7TsV2CIY175BNJ7B0OEgQ5t3T6EZkb/jsB5vpGvFPDR5Wsf5N9BY2Lhfsmn41LuK
X0p1MpS8o4sNp905+h7SNo0cZHxjC2VQFyP0qjUkeReBJrLQ47Z2U2DFH3SjMPs+
n5aOAYLuR46+llRp2SgLwF28yDTbWQwUifLcvLEttvUXLOI5RpTnw9AGmjfoJRLa
to4mx1nNupn2QOp+fFdJPPnWoVoYz/QhX5KritWtTx88mzN/I+6OF8IAamltjcHQ
B7hkcxgb5zQNiMnYwtkqVx2OagYvdjVcIfvX5iWiMDtT2AnS1yjMh0ZDdMQPQpQR
+jVWgopCFcnUQlXeTHZHyeyPipCO1NDRTz9k8o6j2fh9lUVbxRdkGFHsAvy63j/d
fbsk7f5jAvAu8e2keWsFfiRSMBcL5TF2LIvO6crN/CkK+8AcUzmdWRtUByXizm3d
sFzwHWUif3Vd7dOQ6q0W1No5FrHkTT/nyI+tP9RsIonurS6XojHfkl1KtSHXAGm+
CKD1AeOt2KoxI2tj41pRo35dgScDVT4iOhhi8lAggfQAIItZSNGmK59M1kUxYTTB
XshWYCwr++y2Qh1pJh55vu6MBICenhb9LESEFsO2HHbJSgtSsl7YXqFERkOT8+we
qptGrSp/ru8wf9yureTvpZTtx+k1v3IsTM88Ym7zw50UoMvMDftkniRNqIH03GSI
DJzcbdv/sQygjXugJZN7qWrive+1Nk37tgjS9irkiACFbWscpWev78kjqpcbfDu2
tuUQPbwMFu2FvoE9+N8cDNjBadWCi0kUnZAkZZwetl/YCgNAkN/jNZV3uyGM3LHW
CQP1aFcI4Skn+QzAWk5Euk+ar9EIAtpfRVmI7aJFuUY5U3PoKR8ESTfTrcJKm3pb
/Gt7OlEDm4GtfZNGfeR6FVnekAtMYo0/M/8oFyDHBXYt6uJymEpV9+aNcvXebdM8
6BMnEtlJcimB762aBZi0EwVx3DC8GzYJq3AR/9tZzl/k2g3tcFdDoqP9PI/k+C1U
MZzmWQQbgXBNOpsIn29bVizNVCFblGGIZoql/ARJN6IEKqDYNAS5LvPEFfwqyUpk
NFc3F6w22sgfvP2HHK/BzfLY0BYHjx5Q5ou/YfGMKE3Y/3j4WYoBAuvEThvvf1Xc
UTkS6VNy3X7n3jBm2Vi8R2xXfXv5ZNg07sLGxvEO5sZOLsl/7ACfXI2YfeCLR4f8
Qu+jSIhsjt6rVI2bS5Gwnaz6d1FzbYTYrCSpwPyMeSJlTo4fHaa9zrTzx6gxoFk6
NThaz/wDF2c6q+ogcFx5sNGDsAMIcxRhz1YUYL2klKoyFhb2gJx30hG8K+akHO9v
Vxl+sa4Mb3Xig4CJLAib9IAL/rlvKSxAA9ykIeOlsZSQ3lV4/C2aNBNb5V2S1TPy
M+p/LJDx5pz7dOxCNTn/AS2k6grlcKpGRFHgHz5ZRPpsBEO9rQ1kEwsu3Z5psGj4
jgxMEi6nZbd6WwSBO1o6ralSNvABjKZgpzqbWlKxKsMCHRT5zYjbqMDC2ID70o6G
ZMF42j6YW8q2VFzJoBPMhCEaOHvnsvkG3NdhXjtwFsBQXusZM1PVRWbLgceOZqR+
z2hSpfNvfBkCVzKs83ruECokUesM3doNPqniYpLV9jpmCtmooI2cYBqSaYcdO0fg
Y5MUKd6Pu7sgQcFIcMhggwctrAO8OcumIwvTikwuaAlj+bWpzrDGy0JDMcg0tUtk
0Xt5fl3jWJ2yjnBT/qV8ObcAngMTrkh4XEfjHU/QTCn6TheHuiHr4r9gUbH92cBd
CVq2H9ePQ3aNeHQJGy5BwhB3EnJUL4eNV4dbYqVCjL6Sv2KAfeV+V19TO9h4FMty
AgIjGC+Smz3h53c53frBQGEZQR9GeI2B2aL8m/8TOJwetJYGUL8p9AzLUp+j/34D
hoaqHkL6YkaoTlqDS9JchC17IpdAaJ7E8WuxwNJCb5RVlZy4BS/ixX83u1+rTsEj
538CNwKgrgt/qTg+Q5hlCyWtMzaax2xoWvBqGUMfOWo+BrbLYwRLqN1RK+jOS1+k
+/oTIpcJzMcOmQ80ZHwhR5n0tVsJO4R50XmKgdIbN+op+jIHUk10h/Uv3mgFaVlr
O6qqDZzEsALoMme6gIwqr9KXAonCCnXzP0TIrXHudwthSQ9UlBI4sD/SgfaI/0Rp
yn7RLGNssQbZePjHwO12h7NmT7tuLVKXpaaJH/8SzwId9U95zYR07bbJJ/iqShkU
mhk3NH4LdDmd3ljDPRrQ77NyTHNmK1fG1+JTCMNBB2h9or9ZsAVSAHbgYL2FJtXD
lGck4FsMRm2sVFPmO2DU0HLKCYsqY0ETgW4Ne0+7mCuzLPL3A2BVp3U8yzLTIllD
Z3VYLLmwraZVXfo7Olnp+a8q2FurnVAcLRiJ1kLVsdJLhi9IZs6R8X6RBgj5J6Hg
NtGna0uESm1uoZcOA9k2zcGwiDLzEKf0K4XBsA2jFy7N4JD3Oymr1IPDUqBQqFZY
/evmIpw+ilMZ2//tSPpz0QAbLXV+DL2OWtaZnfsBhl3NpWoPpwq3YY3j2oWJJr7B
Pymiaq0JoJAlVDbB6P3O+G06mFg30t6Njh8f9qORUY2kcjJ49eVzxFCPkDVYmVZv
a+g2SrC2WC9Qx5WBX7J7FiXlm1A1+5S0C7v/Ug+UTBHHoSZWzJ9w2fGub+9Jwhrn
ckb6fIPAAN2FuqnLcyDR7nQNKaWpm+ABW+0hRizpZYz8LaA+Jdm8ZwCmYkHj6u0D
d9WowJycH1paStyWrfAkq0NuecUyiRs0zG9yyJHBwuNzQzSMcNHaGXQQPitpbGhi
uT2ipvG9vdx4FjnEvHb2hFEvSZRCSzKshhpAhEJ7l6D/vd/D9W85IdxbZ0wPYVFJ
o/Sh0XfxknTBa9gHL6+wxzDOZ2O7wHksfM1DoKCkd2H4gpgA+FKB2sZldt71WgbD
k6aGII0IjBP3036q0AD6ZTrm5x9WH86MCe2fVzbKyvr8v/nKMDuh+hHOFscqsb0Q
YnFGuoD3E37MOXiVB88tS/WLU4xGDZ7d3F6UPe4saue6HnalJ0ePndpu/2hlb1Hi
emsOd8zGxzQk9QUoXKATQuhgfDRzHiZliPlxgjw7TPbMdo9yDm04Zueyr8qt8rKu
ybarJqdoatTwh8x+B22QIN/adTl2aGD7gEop1MWn4aRVz5KIAIhoar2dkRO56GMq
MDUeskFwvSgHeTn6HaT+YBencx/CstmTXBS/r2rqMmptgKtkCvMpEhhuiFGf70FL
d2X71ahDbTvCoIv6P8bKUeORxZfryB5pOzYOqLM0x8CAe9M5JKjyCDD451NEwvjD
Q4qIzRVNUVJlZyjbTP/DR4nSMPJzkfIItCkGSUf7m1sZ35UPi/qq0/NDcGmDKsJd
gfdfH3yPYGIjc0BGPJU9R0A5P8VFPONv1e47dsqCIO/UvDRZCvWtOBGvE0+yDnP1
/4igu9NyZQMxr1vgomMusKBQrpQQhCDhHqdgEFVhsRdHmHKAvwJpcXMrQoJtfuNl
VgXf5PCc70weRIt4Sb+AgtVEd9U+PrKaR05YMN+f0wIl5mCOR/qLEHINGF77iMf4
xrfCU4/2HY4qB+Lh0wyrGOf5x4oj4Ic0YO/kgyQY5aekwccyeBpLw5jaHuAHYxDz
ERCBNiGymjmVs0v2rZZIYq7XfxPHVzfGg4Rf+XkP+bYIuaI3fDHQ1l6kcCBkIUVI
p+UE8cm8dbs7vlvA5OXBo57rnCOm+Ca28qx2ttw2DiN5juZxqcqG7aOs8CyVifCr
oexScwzvgGDkKDLfM1Qxb/JW8+O4DR13JrufV9IW0hn5PpzizS7FnLwQvpQxGxrj
OLrGkgmh4fiUTI4eHKYuAnWnpqDi3/wtsRkd7Fca6U5oKEgxT+f35zkGWl2HsO1/
NeXvH4g49XRyFWBNMd4QqUlpsMHQJBLfk3qEh+fygMc4WW8uvpGXXqahlj7bFU2x
lYGlG9iyzpO+NLr3rsnBZehj2xfEcY9WaF6DrHLuk4QAVxqQbLqnOtQG8t8PYXKn
AORbOXPKyMwMcBfTtrMfIquPwVpnl+pk2MXHjw+g3uJHDltElMpHiwYge3g4V7WS
G8APHLEaD3RPJwNWPJSLr4Ev8dulwpA7lduIYEKNIs+1KhW9Z4cVbHe2GWn9vacZ
iBccGd9SevITq4ygY4JxOIiHToBO08rQwnDfVcve5gtMcO6E4Fmo+HkWwBN6+jjz
sHkQJXdyGL2WPIuRUNydAftnFs8YzcUBqMPVsbw6h/WyLYS9klz/j+AhAhuVuCAQ
FqA/eMxRgxh0oJYqAeDMEsOcPqH3JrVKYn+q40p78ygcASHB8n9ZxFw4gaiOxw9Z
trFmtB3yQHMCCmCQTKWyp7rjYewoYTb3sBDxuh8ITBFUsiIZS+FsVVIJyN/ex9QN
r5tM7GGjZw8I3bZ29CWyvxbfl1Ve83GN2vz12S6faV2U71/G5WU6E+Ay2MavrGdm
RjzTSu4ToWhi8sTaSnrkczfqLgKKpmP3jkhTJwt6FkGCqdKIculbPP4YFPHh5xOU
ipxdwJ0aSOpdAVlpNg9H4xgYkhL5tk6ACy7rAiucnTNBp+uM8xoBJoe6h/TvGWwf
hphnctzn6s4RlXr+jpjLz2a2iOufvzuHesIz/xlrNHFhv+vw2h5FpyrMMEsMyU5T
RM0weplI9XSl8gnBvL1wWoIrY61gsaCGQUaO2P0atb6fNmY9J3lu5Kn0oORn37x8
8JfOzEM72gJngiJjtCoItOQIVBOD8iroF+qO6qqH9ZEFhF4pEFKspBqjNZsc6OJH
5K/F5IgOy2LQ2p2CPx9pcXq7Buyai9N/1Ih+E7EZ5GOdwRexxqTdhB6pcWmWE/df
EFQWVWObIoQtLmta+fsFBVv3k/7OzYCfqAvJvNf/vNcnqxxhCfNuVjifnVQU3YjF
FOU6z0cyDZ71HVV2rcuH9ZzyqDUMS95G1J17b7mLauiKZIGrJH52owKSmegpJIvC
6WxpZdYEnbJPwrYw+6GABc7ubGK7V/1jzWSnpbGb0ufryOyy65nU92BwkYc9haR9
MCzWFx2wRyChXZUqSlhlKrPDE4YqxpOTzfhhlI88gW5VMW64915YxLUU0DY0BLek
9phl2z1dIJtOmmCVxdqekqhx3O3dECOH9B9qPWPmysVLWRvESRxaF7wivjMNTdhj
N9b2RqBuNkP2lkxumClw6KFmsQgjQHx+JFK+Oelb6Op84o+9RrL2ofYmn9UKIbRA
utIZPVu1cxNTboQUffpS5ZG95Wsedcp8WbMXMbCUkLLjgO8U/cvOE+1B70F41iB6
SaDzufiBr2lSH2sDzEz75uVbvfY759zLaHOnzC/UjoRIj+Rt+uJjTtlnzjJZYM/Q
ydn0zC84r8fJ5S2TYyM7gQjw+BPBLhKs8OZQPTfwiMu8SfU6JZwtAAebKTVMvv+R
eOD/AUMO+oXduD2mTnik24DfuD0wJ8VsW851Y8PGc9Ip918BOK+n75ce+j5+utcG
nMcpznbnMkJWs6WRLHEDgyuTROPEinWeL0sVg8aa4ow/wPfH76UtyLbJIfHgA5UN
NRUn4b9YLn03ooMbGGCURGNeJBVVGOMtJQdCxu+Z0gHRtSLfpTmajLsyh6FSr0gl
rWY5jYm59ALRE5T+aKgmJ+z2SbFwPdqiyj1FMYjb0TloaprUcqJacv5//QURlk9V
nXT+OHrP2RJatNdlUgFJRoilqnG0Mn9HYIzbFQHn/pgGqpyB9QtoxXgKtotgAE+T
PheNTmzlNIgq2Se6kB03vryoFBq6ofnTPT97HgosTy6xbSimpxeq6TJMmhh95j/o
UETOZ0f2GrjuvUTzED0dv+SPd998I0PvbzDthkerXu50u1RJYtaWI/6OE80hjUBs
PBHpfZODbz/0nhqxsBRkIkuZttWOwdBHllWIrIDrAkaxu/7mWBTYh4kmqE4SRPWe
fe/GF8uH3q/rjc/ckgYVwPeKD9WXWeOm+NeYprxAXahUg6VaI6L1geNyFAH0jR7v
which8Y40bXWrkQ7csIN37j/Ex123jTxkK95hkGLVJUExHwlCrS0jZJM58EMmULD
U/mk+9NHspUexP5pxQVP2dlu18Y/n28hQSZY7Nv7a93hfkGyJ1YvaKqwGinJcuAY
SzLAzwaqpfVhqYmzlz73CmmCRDdUlHQlm+/Wu4Wyttpkk9CxW+cEsc1LyymJgygy
PQlDsEkyH1L/yw68ATukyMQSWlBc+xwWIiyKlx/8XjHwIyxJdWug22bUWwMo3WYL
1uGQXeSI3WH0b+wKiUZiEq4GCyGaFXDUS4KydceL5QtZFAjdaCWYHF/E1UGim7n3
pOsqp9tD4XqCO1apeqbX3ye/i2rIGCY+UJ+4t7hv5qo78UCXSEw6goNj6b+yHh5E
DMdy/bhiDNca2jtWr5nAYDymWwqKzKgOpD+GbfnZ1pARqhwckW3N4m9Zt4znKy8Q
uGneWwKuz6VZlSVTf92lreMoPM8ipX3NzhIsVbMQ/NielAn4K7guojSnG49g23iq
GSoQenIbvH5XKm9nuCxDcPxauusuxTgNEIIbHDYW0AdLdUwsl3mww3k2+T/oIU9m
oWxqA9PN8f5kL8XJAQeqWpXjhjo8HUVlrOuLGupBj5Rm0Lw2igiWIyzvunpoBqU1
eWlLFA22irUvFWiOXpp2hntRVWFBGL83zEiWP4jWbwTtlEhL6l0Ww19uJfBDX3Pi
VEy35/wu3vMQukXjU3lPYhjrBJ6ocngXASacaPaktwWR06mDIYfKzc8iQlK1/3zc
hv/s1JFvhJp+Mgad3mMSmLSvHDXdmvoZrztF0hRzdlzE+epjNJWAVeoPUaioCH42
Pylb6OItlas4MuEcWB2SS+EzMUGPmRGXcIg5aaH6scoI82t/4Ei+ckrWD8t+d8zO
yV4DUKWT8gD5PGeyjKgpwxnstPypPNkgt5GkhyjaDLVYc2UyZqZg3pE/zjc8zqx1
3r9dr2L83idYBOHfN5EFCko2qsdzicqOxoRUU/CjCMnra3Bv3DgfxIRW7Iu6E3YC
Fo1nlCk0rJUB/BGfvu2jMNkjX2ByPlnMCSZCSv2d4b5jnygERmUl+KaD/kakQhIg
d2YiGhJ3CcTEl8AvQQ6FX6W+87Cdtiz3C+NAN/zRO/LjtCWNqv3HiBxUPIcuaAiK
TpQmAB6AxPkXDv/gTaV0HcqC/MRe3+OTKjgmtHA3v8/83Uafr03R9R8m2AYpjGyY
WVp0SkTnrt/NKpKU3U9WBOYO2O3DEBPsI5Tjuq2fqLchm7bMVGJhwuDu3kp96RtB
YiR5FV+S3wV0XnyUWSgbo7ZQOjwFCJ51FrtAJzqrp7w6stYKTXh7ev0q2W672XIg
fl9d72OJvvgzvOLqUka9wIwQxpBiEQEx8wwcB5phPuC7fI72CbkTKU4B9kqlYrcu
A2GjA2pnMiivwQ8POTgnTzrI56sH6UYS6y/22KsAjOBUtNGamTbJ+yNpfZM20LXB
3/4M0dxd9X+bxPUDuISBItUx12Lem9zf6JD4IDXqzPQkyD3dRe24X/8R2Myc8taf
LuPtI3H3ajPRiNbNZRO+OsAeBqYDDT2VhEDdYgjjjoXz3TebZKS8ycnIIzBWcbHt
DXJLYHhMfjavHP+BS0XutSlMk5GjsSxMVk6pSERVHR3UvLL2RZhCvNBHh8pfJEQ2
lLZT5fInhcTB2eerOS9FOpQiYSGUwIJTqkzmn5Z+M3bd8vscLUPFwJstNDwoxWnC
6mfpX8QSWyHzbTmLrNj/8InDJxCl5V/drpZMbIvnERypgOS1Zw2sfd6MSIwVYqRe
C9XEQagxUvhONrMpJ+vV0yayhCz0cxSqYnbCXxWB434JzCWvaoMYGqeQV2bsZy16
ntrXPhAAwAUXM0Eyscbs/r357aU+G5Lt1oYFYZdB3Qj5MSy9ZFVFvj4pQn4FrmWc
kI5WXGuRPzRuFXc2Ozr5Jm2KYFe9tl2vPiyulhURjaFEdYlmlHkXsCTnYLxT8t7l
oc+auyBpaZKdnMMVsIlIQcwQ78LdHDGYvvNzOX2cTdFavHsQj3egWsBt9NxLdMgv
ecJaKUDm67C/8W4l+6vvOtJM2Nq6bkvlpSLo00scgJFbMWrRZ4zWug01DKlLcv8d
G1gRI73uTdu7zJrlMJ8WRxux4IGaqG/V250aC/FREx3iLl6D2IjleVj7WP5fHIHf
VqB5LQuVEz0Tpt9l3bX1cBrdEGSWKHC+qHnBYAs3C0qaloBbAJ3qDguOBiP4NVBA
2ZM+c2E1xfw6YLSjYtH6j5OIHnv0+omIux81nw+IUnuLZy7s5lZQEJla60zEI239
DatLk7AvPPI54b1q8SdGVyQMbMbk4IZW4iN9pTwtSmXMA0i+cwFI/Z4/72lyNl0D
hyZrRvRUbHfyNRVkadhS9SBq/IFMTcn31+Szz+djEuVkEZwGh0d5VmSEwtnUQ35Q
kZ8K3i0ZVWYdB5yFkJGQcD92P3BKQz1FBiB7LToWTHs99KxF5RkYoU16LHLq86mB
ZUQgQEiD3bl1Xh+o8e550eoFx2xCPO6rgvKVK732ZaPZED2NjwBflfFXrDKjtiu6
wtCO5vL20YcUb60RUMFuR2OgvsagUdkhB4Zntez9BU21n4qGT8vffddix/W0XGCg
0N/spE1/ftj3fq/uXRh0Wa4X3DSYXPvjqnjB3polIZPO5k+ox9NCnjF7RsmcU6/m
hRfgBcvIB0MJvMzABWcVWy0q8zfPZi09w1VEiuRLJpgj5Welo0SCV5M4TTT/dXso
NSlEit2T9t916H5b3+m+C0FKFWzJYBCu8cWHQynSS7yzWnLZcfE4/1ZYmwEl3vhJ
sF0Z7dMnrN0/yzUYYTBRNCH5sz6V6BhDuEEjIb7k7Vcx8IGW9RyfS7SDHIrtCZuo
kI//UGaNuastV6mDMSyOZ4EKcHrDoDMmE4ka2ccU5gZzgcbiNJBmI6vWerav1d9f
Ye38dYNfOchRuT+yCkLolFH2Lkxv5mYyd+pS+SOBQZ9rLqkuqasIJxUqcSILbUBs
lKSM2y/zpcanm7lqxjqRipMBLOEZmE5s+SyKUiu2y/Ne5OLtkJ8KB2m82w9PY/1T
PBTNzS1iu5NFW2aOYBtibl1sexEgFRGV49e62DHYLrFsDrTV+riQ27xdmiS07D9p
3w1Zj8njcjbqtx2yA0VeuotC5K75kt1NcywdSnlJk73eeUlngyluFSa9aJ70q2+M
Ed8WkCNd5gsAz5CjGrDtwu970eiJjeTZxtgSry4mpTAeeIjutyInwG1O1F9LZUWB
ovv35L7ElGcX1Uv64tlrBQMlMMi+j2uMi6l2kA4LMGXxPf9kddEWqTnfDTzRrbTf
ipwAz6sJO9YeJPBOe36cuWUe/KKUNAzYNYGkwtC15ZPPMOD1JkgPFV/FfgmkJK0r
4U37KkcjTib1JQG3ghQgZtfNkxuVqfaxMmWTlTC8+FW/4QVo7hu6yxR68/z1eWi2
KYbX7xp56ngyJp6NZdwXJTP1tQV83nK+eFa6wej3s8Vg9V0oIYTMUpFnFj89Zvft
Q5aVdMCG5+M1/wrWfDNmsiiM2kZD6jnD+pGCyW9xjITAnjZfAEJma0mIVYGoKq2Z
2rKLAyqV2269tUDV9o4jybe3fHSFJjKCTeqOzsBcpgmFYt/ZTrFoRd2YPbBE8dpc
6JE6FmB6eDqmPonPRJwEXv9UMShkkK3vNMT+pDoIuTHA2Hh3OThMC+qKv1C5maMd
gLUnhE/xHDQ8BXqH9keBRi5aeVU5xnLu0TEOl3FskufXwoKPTgwnh4zA/sJ2+pcp
RqkomyY54N9XJDHwvVV0UqA+K+J1rfZdEAeL8sNrMgYYXlFDjM+Mx+EY3XNy+uZC
0E0SowPJ1+qS86Jq+LmQzsDrs4ulyR1rupKkJV33z0qLSPpmsO59RViDRdDdX6k/
ioqZ8jJW4gYIf/uVgAsb+pQh9YOipW35T9fXM7LgjM3OYMdoMZOwHS8zG1zTy29r
TrVlN94UqpfDf0DVmBdZl877UBa2o/k4mGQ7FOfqyfB3tNSDnBHgYIAixo2nJ/r8
/INlDC3wFyR55YRoUMuEE57yI6gcxTVhD/TfhaKcr3MFZneQRFLKcc+Jwwcq66WV
ewuskT1jlBrbDwr5uZrEEVc5sv237i5mC6h+tsZWmAuDhhC/HqZAt9MrJPW+7UKW
9VPtcDYa6KvNUfnbqjpuVDrL/3UVMUYb3m+CvzrP0MW/dhEphfFnnB1rijo/6xFM
nI56CumbP/LGN2VFX5p7PIcR7BU3RszvGhCnpPdU2wetRyvXC10LkKzlTuoQ3ty9
mdpvizp9uc2xUpPZnbvzfgyztYHi+JiaQ8fX3lPE7u8Zt9fz5v5tO/ZEZpuLVLxx
uwHOoKnqNWLlDU598IQYapmsKOGRbl+Qu8eVfPNHvp73wOZW6PKvOXDusTzEcnXy
KE/T47PV5F1l3LrCJOnudUcLHIBcgDWYD+SjpY+ITv+GLsKTGuHOjj0V3U5HhCbk
7h6lzRnF+sG9CTaJFq4bNjXDBVqMmyVisOsDoBPYfGnO2ZcU/MJQZcze2dOFK2vn
EIZOj8i3U/MEGrelRt92hQ==
`protect END_PROTECTED
