`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CPZy7JWKd7bJHKqKiIFqq94+Q0dOemx1025JDoRLzb+ijo+EfnHpBGgNnGxg7vQQ
GvWf+OzBHPXO/8QKF3loXlej0rgPI1Q5Y73fM+wuzaZY5yCwoJ3uA10uskV01N2R
Z988u0TMUqDlXdqQVmbWX2/LQA/hndk7WeUl7Cyl6G4KaMUmX0O3mP7ulfGdBUGB
r/KqXalekP/OfOEGEHSYAYVYjR12coXbISy0Y3Lm4YbH0ptq9PpdZNGquZqeMwCL
YRR6TwwgYdR7+ZBmd8jpiehQ32s3sc3yT+0p1bQlRAVh4y5gxB2sEmfKDfyWS83T
AjSCDO3WkaLpmkWTj5rY2pWIS27oxQGVBy9fJ9DQLCZfuf1papTxxJ1NKVfJwHC9
4bQR324CZGKTC+wgJm0irP06kmzFngcpLXvrIdE6ZlJTAZdVBUos3/uSRzAm6dix
`protect END_PROTECTED
