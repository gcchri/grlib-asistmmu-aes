`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dEJYjDp5oWZcZPQJpwrb7wcyH2JskPD9HcevP5dOzlrpnEP/CcbaM0sFo+P63WPZ
GQNKcZoFtWCNvzDC7e0KfYhifxzd2N6kKMoS6J1BQcKFf/7c9VH8EKddrz06kFOL
CklvIywB7D2nYLU7J7JFeXgP7WNA3rf59n3RAYMGN28w8NGi6CJTfwbt3z5T1144
hFmOdvqfbzDN8SDNNDyaj/0buAUBkcN3IBj3oEZroRTg7zfj6AwFbjubB4WVpSZQ
3Pkpnq0553gmuUrTcTJujRTv/SmBc+SSRhRNWRWBcotpYJKcL8Zflg00vVuCIdQ6
PP0zbeSEDESqieBkJf+NIA==
`protect END_PROTECTED
