`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8sa5Oyac9FwCWPTenioKkNdT5BbaIbzCHSbg1oROCu2utyxxd0KaNdXrslLdwcNW
4RiWH/P62oPiZLy4E3U4jgQv4AVvt9VSaxrQeYuoS4U7HFgimGW4N1bD0lZgPOZO
zYDhv75yw0PyovatDaynDI1Lx4d0kDSyUOLUi4YcZNWghwTUFGnu7gL1Cryv6QW8
Gsyqwbw266ZlLgdsCnEfUFAHBwEhO6PdjMbu8Z9CU+MRmBI8L56b7uKT1Wez+JEP
l2U0Y+X30/i2bZd3yf1n0mwjgO/FDcuomdi6bwTvI5ujDQd3lBxbJwRa6ZwmNaz8
/aPOPFhK5GPYS6MKv6Pck3odB6nriR1kF1bfztmJiRdKoVRE9TEVpA4iyrpPOAG4
ApKWi1Eht+q96K5vVooxmc//6qjcaVhOXJ7GrWW7e8qQLp6wgrQQzeHfB7NjeCXM
3HgQwWggBqIJ66tjHjVfF6hRWls55XhLK/n1SKbM21jgwwBhtC7xU8rXb8govBkN
CIIcCPo/3cQF3eje/uGSwV8HZN13XzbE08j42KLsdmXYs+dAVgLtazlD2gkhM3qx
5YsYzsWEBNNxchaF3nMvpJeuEXVntt3qjzhyDruu65tf+rhVuJpxCPDX7RTt2ndr
h/5Q6ElgqW61CoFEc+L5rstBjmj2VQxifLS2F2mZr+52d3btPbWh1kZdloMDV0VV
K9FwQSrMnZKK24CwDBLLwcDI3NuDRku2XmQFnIqtIBvfi1tE6RJ6t3Xk6RvR02m/
6zxPgFZEwBDCaaKSiBfgNA==
`protect END_PROTECTED
