`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b/DzuMt2jK8lQQ4FhoaE8JzvCTCXL/akOm08PPUd6w6n+WgrNksJuxbYJJAD5IHR
dfAcVNWnnK2iP41k3T1phG5w3KxGPO1kBbFXsKnkdy44D/pKcU0zD45EF+Q0Dl7F
kNf7Zt6igUbmuY7DU86k+NDNohfAFhubq4XdbowKI2ol+YarM1swBhKW65l3hkB/
BYHkwRoBbymU9c1bs/bjOepe640+h6LmdWAlLmKu7KfSoKhQfHuSauxJjfw/03Pn
Dn4r40mJACq3DuzcNmmaKyVQirE2dWT9sj5YXBVYlRQSaji2Tv07mqHbkakEwpb3
6cMAwL+q9cVbnRr4NZELIQZOOIajHC+56gxVYhylUQCHgtBZNSCymC0FnFP3U8cc
GReQuavmAAphZCeWlunCbP8HNCY3sILqqnjSabRB9fQYq7yMOTYrwtAnumAR6sP6
3nbDWXKuH88KjZX23fKf1obfwAAgKQuu7E5sLFJ9NRirZqABm6s8/sCImpqbV0US
BzphUYLw0AUjMPbOZqpH4vWf+cEE1ow2RMMjs2yXYAdZE1outsU8O17gGG8Ad/cD
PLmNZe4CsA5Lvk/K2UnD4jV3Qg4lrJMCU3vARUPOCbMtkJC2F25amhhrjdrGkJEc
tQSN0i0ccPxZEJl59dhqOfBhBNvyl4FJocKQYLicGTwB90w4chQRDkhcdmDHMVV9
USgBO21dyyyeOOM/8oZBBj1KTjF0f09GMzBk8aYX9rEJqUSArIxgrbRzGM9thblS
2TT68EB0H3YRi+CwcRDb2RWe5UA/WPKnAaQ3RNXQB6lytWtBwHMxKuFpbKNwvcbx
ai5OwQuWQtqk1dEOhZlwSObthxA3PJQ6VVJ4zv6IBmc=
`protect END_PROTECTED
