`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G/p3sDKwJhycpDBZLRT5G/O27Arm+f1Rjqttsl6Kh0bKY4GF6EGEVQUdv1k8XF0/
29aOK1ZAfASsJyvar+uLniD15/GkdLqoAtldVYnuvZUUCqc22hYWF2bbMxbAPflK
xqnuV3UXrT/+9RFKvQ5ZmPBt+eK2L570+/zhY91eqSe2DD6kYpWhPXuQsss4X4SE
VcjIfHeX1+oQoqncoFb9CLW/A2IgmCETMGUXwC92wUgX+2AeegDrMcR4ShR9kvMD
OZkWeFKO9rCWHU+eCB6ejWrshfklMSE7vRC0QUcliDhKLYJ4i1z06fFdESLPTpI5
skBUq34j8hOkyw4MWMn3sSmj33Suq9h0/wvhNqGzphLhNLr/AB3kj9VG6Xq718ov
ogdVSKa+pDmtbeO93F5fTnZ3wr1LJbzG3WKrPwYfGx2cPD6Yhtf6mXarVD9jdnMP
LUBRzBpqq+FaQPl83tmhuqt4k2CQg6iWU5x2o8SIUSk6/SDWtEwYruv7jCNv/j0+
cCC9m/gZ5JgMljYswMkji2vju3Ztohr9A7lDokFiAfdATc8qSzfY16fW5X/WHfkv
7nTeNSBp+zx0WgsdoVMdB96RhEgJ/2koPum2nCEFR9rE2KlEYHrbTl7vmXg/45X3
jRb2bjp/2iobCScjag0cknZ2dM2VBKNV0qIXJfPUYX2De5El4cSYdSO3JMCpKQZ4
6BI7fIbLfP9e0K4BSM++XlvNlweug/A3wP7qmVr3b2QWGNn3RqDC9OqdZ3fElku2
9LMyr7+ZcDV1hErfW9qbGTvLtPEF5qFQPeh2YeqInFY+gKXorNi5P+P02XBfLf6o
adZi7pm9KegkxAhUS2ROuj7tAPDDw9S2YCIn1Ey8KmLnIMffuvuPeCh7EXXLpFcn
ElOtoh4T37H5tfeEbHkhhenGxsL8l37wbtr/8yc5rDcImK+2vRfXIOIEteZqbfO2
`protect END_PROTECTED
