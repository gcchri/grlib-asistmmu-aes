`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V4mmgIhjsTGGSFdVPO2xf+zEzjIkkZ8fSIcwwl8NMzt68l5Ak+/or9W5wZzT7YNP
8q3smXPDa59UKqr+5zgIiE1/U91ADTr4IDYxd+ExCEjuH4iOJubBRMSswLkOTr8Q
am5A7ZTqfS5jA348Yg0WYX+XSMzkUoCQmgigDjmAwxwsNCIG6EzXkF08ifmRWqZZ
lTF2PIDCS1s5/Hqlx9nPK3Vw54wARpHM//ynlvgqz81sQmtjpz7KKLmEwZ9G0Lpu
8gI7Rll2wR1arEx2N9BCiQ==
`protect END_PROTECTED
