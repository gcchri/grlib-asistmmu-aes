`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rosZj5qnpcszOqsrZiuPM88prpVpGM5cEvdS66v8gWTH4y++vxGVpm7DaLKcJ8Vo
8S12E94stfGp+qZ5zetH1O+DUhYHyM4kSFehw4X7br7GVMoi2Y6aqVQ7n1VnJSdJ
/RtayhGiqJPHBeEzd5XAv2pJnira+js/NYcspcQDARGJHBI8K5RAox6DiJZSH64X
nfb7ljIoAZgjq/gAidEwMDu50Bffg/qgbrLiZwFHk8Xj2U9+Sd4Tyw1D9aFrDUqY
tVGrsDjIRvfOFYmzmSSpfwd5gtB9iDzJKAfHNfVg6Bz2dA0f4eCxKVVVhhrMEJNq
wYwwOeyHA8PNJO6yiLFSANJCYJ2KaFI8YrRicXqFaDXkM78vgyccJdrpMWaNA8FP
vRUoe+DzavATbRBGkz5XAS8Ep5/B/BE9mC45r5KT3nlMBZAaH4GP0xNoM08NQq9u
`protect END_PROTECTED
