`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Qpwzi7wAWecu2I2CFE1ygeuna6z6sqQk8OC1ZJ0fiTSo+kvMhjxknU3yrB4Ipl0
1n3Lf9pDk5cfPyWrOmpCEevGp8s4j1yskbQzfNepKI0Pdh2VRlKTSb6QBFR+vmE0
WQSxI0GLtG4Ml48c3Uee16bkAUKpc7044mHdpWze2Rzqb8dNR3yz4bd5KFsSSF2h
aDNmZEWjiWaDpGqIKcK4c5cjVKegmwhfsubAGtfDVHQ3rWVJp3vPU4ioV6ljbDS+
jZUCPdXUtg3axTGSEzlk5ZmfIdz36ju7aQKbMYzyzTE=
`protect END_PROTECTED
