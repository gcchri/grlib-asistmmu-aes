`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u57ZM6fiOH/leetvivnfiVpxw7z7JoLPtXTXc2rAUpuuA10d7MvczjjPllqIz0pi
iVK9pmp7rM0gPN2UKzAcwEue+eESC7PEpVFtFJIwh1vuaUkp878qIXmduidW4AKa
SiFgjTbGi7zhg5H87t3UvZSh9/vvalzBuqksXZQXsaOXA93bW79OBXYMFlZ2ZNf4
WkIrpvLw8+RKPWjZ2Wr4vHQ5frHPijoIhs+Icd8rdmFBAdhAjoeJDcgvWApQHR/l
dNux8RXLwONTcN0pBuiePAoikjor7z4kU83mnfV3YgcmjqH4UA3bDyKhHKhcqZA9
mv2slPK2pCDrhpAy96xeRbcTl63hfYv/7vBdtYY8Icc2ijrnZbXmO5Bbfj36OePf
YarturGJGRpT/Mt2inxfnIVlGx+9Ojf2yssgEGvTl6WMpCg4AHfXV2Dgcu3uEUj2
vflQmOvdPd6APoxuT2LVT4cm++vItBYZEL4PMnQGWI/dRFMizoeyJPbpGNMUQD4b
5Z/fOi9PA4huJnSKPTDSfJ06Fyz+IcTf7lkGWlMbNIwQGVPh2FhHUbSadNdmEmlx
WA9MkM+dHOj72fhb+IBYX8QGILIktsF+bcIGWp3ruxciVq5E/Aatlag6DvVtFro1
HWe1sR6HRhAW5wkzdPhiznTsy5O9ljkB2Nj+s5FQs+Bjp5lM2hFPr1BWByClgw1Z
xqxcuOi5Xc2ytm5DAmOlmrfFHAuOwwGXjtkLARJ6RV+WGsljRMgGFwVfvQgwcR+B
m9PAP9tnYY0pVq5wLzSscX8JdOdU0/kETXzqX8Tq1sd3t1JdBCdA/KO5XYucQXjL
MhZ8Z1B7AoTwWm2V8mmMHnXJZ8VrNu4iRMeqje6n3p1VUWbTeeCY4I9u7cEQ+Pc/
Fs5jqY/rtcn+2qTlWAhWpUUBbTX4qdL9DSaz+KI9nI1g95Qs0R0g51OzjeD/3MA4
7SxCTy2ToUqPQYRdWVdjczMr/hh/fWayzsefD0CHHr0MpzpoXZrVWaKRNujbhWqw
qHDngkdkMPAgHRChxTWn0HitCWsvl2+xD2j3frj2qK1uA/ngp+/QVnR9ZW7IYW7+
lFFZqHjsm5MSC82/49R3jMK1i/Z6+yFs1vKaqPjOC7dhcnnSFafNqhvB7NWSANd6
I9ZwiBi4qESgnPvtjQZ1QUXFLMuQYwaFxNBaHXL4MBdDVAEEVoTnN9CkQq3ggqYO
0wzrTXjTSpCwUYbDygrAMYMcRGYSgBB1Y1ybMSSmUHwXdy1uhvCiBPm0f8qM3uEB
`protect END_PROTECTED
