`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JKBWLqEUHibmu/utr35zJkCtqRWGyHsiUu2w3ag/meZ+TmPYGNzAYGFVrZa0uC2a
8YbDS0wfz2toQyjUCM7wBwMJlxA/LxO92stUyLzVJ1vjv8WGsPB5Q+wu0sYdvMxy
C8i8BePnQrSjWvHJmiUHAGR5qMizIsKaPK2Z80PB6YW0EC25QtGgoyP7vPzsrTij
RBCSE+e1UkLdqI+W36H8RUn9T6HjA0i9i0EzReV+1bgCuWMDoFvtYxGmNN1Pvc/3
aWQJDIHdqAuyuGAlXoxJgWQBxeIU7Z62vpRJE7/VsWfnBxYlm0vUWOo6dV6j4LXL
s+eJsSLqp3YMFIwGHrYIKhIflBjsdC7ip556G/Icmp+kvFWEKsA2zn/bJTWbyQ9S
SiwcD6t8xMQmxXKwKgSZpJkBCDeUqRiKrQ9ag6QiQPq8Ns5vGEi3lsqk3ahReqRM
kqGthKRpyHNwpWojP+oKSlkVNfLhrJXiEm2d1/ZDFolgDbsz2Xr3sgMg6OhMiYwc
joB/PJUQnHb05prkTPUvSS6VOXiHctyVqByAtAof53P+yOF4NPa/kBljh1Vz1irr
/xnCON2eFXr2nczwlvekfSYkWv42HyC3RsIuV/hsZ7Ot7pPtJqXzFdahlcBTBpm2
3HwvgsJPtrhDkERTYsh56bJ4fBKqkH90Henj2WsSaKw9iUGkNxVgdNdaczTpUPRN
`protect END_PROTECTED
