`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
99N/Vf/rjEAwWldidTt4cAqPUBJNPoKTYFCbV9KmaQ7jRKDAvXBBSfFI0B2pjz3w
obFI7uDOfW+a6xVxO3eDv1UasvJSbhyhJNNz6lUxAL6/E5IZqjfoLmvb58kBCHr9
Q1UvFiPnOC9PprpTiEOkgytVTgA4o+TkQ/PT6mQd8zkMmcfEdXEDt1niRXeSKn0B
F9iniLdQkMinEke7FJZmPc7qeDL9QtbDA8LD+KFcF2LLf1sas2A8sfwMLDlZRzz4
t348adgMN0fu4CY2i6CRAQ==
`protect END_PROTECTED
