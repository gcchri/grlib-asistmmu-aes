`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NrUcCNua1vyENQDJ7GgO/1STwKHp4eC/QZgDoFVAXBgQe40WcBgZyDk9Y3DXtco9
T7uuuyffnfYxYnOcJ2O3vPm00hXopnFnyuTLQO64d+nRMywq8ug2a6sDuOVueVv7
orj0DZYWQ9wureAhKq37slL9hlPRAwMHgd7hmJBW/Af4M95G80oGNdoH5vtxfxuH
wZYkDAoZOln1xwGY7klWRpvdvKQnJ3BIwsncqao6kaBNBhRcIOCSYGnJTxGu/74u
8/Bt666zKxbHMsO0n7rjZgJoL/50gAWsEh0cOH13Lk2paNaTf/b761O9rKnUS2Jf
okJalzaAsUPHvbcQmjU2ehaanOtDDqvWyW7yMF5Z8dvPwXbOwF7vSGQsvFWcBk1g
d1hVTDtJzW7Q1S4VKI10jzO6+zm24Ai4ltUY7TbI7nfPzToM/GKOvBqTRfSApDGQ
d5SvKx99/OQZNEhCBurg3ejINxSbJrmwc1X3uehkBZ7Br2NYGtnu0p4/WopsI40x
B7p1jltKvo6YdEGrsqXGMKpvx6djZkG4+XENrNux3pnrYiGPuRdKkyH7/vS2sDN1
a5h2CsZJa8YxvU6YlgiM26pLq1yDkHCD/7/VxQa1TpCbOHWR/ZMROJmthxxIqMYm
5EE5fLkgjy00s3VZU2ePbDjybw/BckiJ995Gzh/uj/9UQKx2/B63OmJAVp1EsYQr
Ts40jXJQyQirjvmH4J/BtDcQixn4sXVqGjdVJrp0Ct18kdf1491MJh/UMrEMUDDh
kRbzdPdsHbo//rAvdHWM8B4/6FC1LLVzzCUEQUVe3BwscNTsBBI/FYIeiALKkaT4
Dq5WUZD6hTENYq0M86fWxkttG1vRg4tgpYEscPPZ1uccf/atVW1R4LLxaJwTcFaY
98NJLd1NvegYQBY19m0tp7Ie4/fp3ci0pymbUHWRH1d5y4bzEiaeT5XDdjOnu7YY
XlZ2wiZOmhKyUZfHQbEW2Yv8CDLrvWqlA4r3tfV5k4VU9cHccfEeR2m2HgoL9Cho
k+Rz7dfHxOAZcdC51QckT2cRupguSdrQfImWr9ei56+aukiEhPPwfuIyYRUm+EhD
NQCiycHOWYkqK4Ha6woP1cuN3/A4dimNDJv7Of9qkyiH0rWsLz5VxqxjFUBCd/SO
ohbCBouT8AQ3H7K25EAdv1OBk/+4zqk+YRlQS3unTEQ+u1Nx6A16ajR3QZa0JJyq
Nt8Vz0zgVTEP++dphOWAWE2c559qDwLLWOIvfL0aIXoGWMuJlIbbTXN2aVq7osMa
1rKYJg1jikxnzZUdUX0dfRUYhHiH72lkcoJRMpi8KGrMdAcsME4ZuuFVkXjlgYo/
5VMsjY3su3DDO4UkyjfhpfYDqgBaST9jtFfKi/aq3f5wUYr6V5VcUWGJB4PdLi19
N/kdfovIw2/NYMQE1l3DAB/NkUDifNvivIpG+Mb5YqgqvFaAoDuCKlW8JN9DHomN
dBhOLXd+DcHDZPBqk1QgOVWtS9sw2STqXLUA9DxqluJkgTMHrGbXSZNN0Up6iW0Y
7qECNf35iMtadnlu8Ozf0J53UXGis7bRnE9WBpdcwg492xdvrS0qViqrc1zOoMUi
2tV8LU+X4pjHYJM4aS1mMTsRtL0jHwTXi8NSqWLRPPNFAW6ZC8614Pq7uFKxIVtE
tplBtHvczx+PWkvZ3M/aow4G5jmh3Fj//TfGVeQJW7rFP5CWTStIbnvxPjfU/h6g
X3rLRvvKBMRgA7NQrORyKTJytHfQc1ts8pEcsPG/gQKk/M+Yj8opnbwoHpYx3wbn
dSpQHxyi7w4uN35VGOMkaWo2CMlc/OXutvSx4rlzIL6zpDbB0SWJyrYU2c7kLbDG
Deho19Jj6kckBOz+0YJTHeIpg61wdxYNB6CsiypMeoHkJ7YraluLdl14xh1FMw7g
nfxDIxkAGfwcZ52ZgI6AiqnrcDZ9WxsBI1CDZRNC75+18+i7a0QU1E4k8oztzThp
UIlxmN3janxZBtgtSDpUeRdprYmW8iiJRRAy9SSlQ0k9EOpCDB+UKijVHJ+MTCWa
bgznAqIrpo4XW2uzjeNLBVk6m2/vb3vRUNR3Vv0AddKE7qhVGvsX62jfFcjnnOzV
fbctd+J5r0maEt2wZhtf/hnTXeoqdlbqjiUhMLFfcaO71Rtpr5QNRv9nAHJJfACX
BWejvosEIT1qem6v0MZs3WEfnX6wqTbItESt69xtgYYzm4YD769CmWLogWdDuuDa
ZZkXdsjl6Ag3C8Ycoqu1trK9ro5I8rCJPSOLWRB941G2FILU5rLPcxk2nUNGXokA
y2242Jk/ldcA1eQq+ecYAw==
`protect END_PROTECTED
