`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OfmYyFh8VT6YzD6jz3t6SaKnA0VDyhKFUm+R/dIU7dAkrHAN8KEw+bkPS9pTB+x0
ezb/gRIfCoMifYK/DFNb8vLAfI0Jv0xOirJ9MMnxyb7gA51Algzk+9JF3SUFaCBX
50+1y3L+2OLychCy6GguLQhli9JB06BAvpYHpw4X6Oy3RRz+9uSYBmPqYfci19Kp
fvtIHQlVTeY+GHAR4H05ZxtWqS5Z0tjYZc1yNUkFGacoInKgUsq3pD3F4rnWvoCp
qJaOn1yYDtmAXV9exJ4U7g308IfwksbOiIRvpVws43u44hHtviXTfd/brWGUbflT
PIbj/jof52uwBd+jeg1Pu6aQWLSHUYT/CCKR1ioRT2IULhJUUS9kZTAu1IGsVDhg
MUTFdfJzkInI4N/R07INsmuiPSHZCIZxAAF+bEiOrZiEfblIH1zcqTqLHdicUduM
Y9/gdJyGu9+/bmpWx5beAMmtIn+iw9Zidf7YL+ONU9ku4+jK7sVZrJ1mIqEPX+/9
cuxDpf9KXOBz/vMqXuQnI2alXyOB2+sUMic2+NYuIbiicdR0jeij2q2I6bBoKjsz
EGr14XR86HXysnEMqU8nutZCKvg7f7n4Q5144Bg0k6f023bYxMqaa8ZnBid0dcDq
6bIvFowI86wckOEmfhhsEGmDB75aewJrU9PnMlK8vm4aQbZOu5nbbHz6wdmzMQxy
PBsGvU+MJBcNSX/yYfFohztCxiLo5a0HCrxEu0bqAyY=
`protect END_PROTECTED
