`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M7PLs6m644byQ47TJe+Cth9QuZ/vDpWVEZh3bw8BVcXAaH34vgy7uJDa7fadcc36
xinDqe9aGt+i+DeM1GF63XXTMVM+MN97PCCpUrySTj+aAmtPlpi9o5MVCQ2VzBsQ
/zzb+WBHNzrvc3mQQxGjtiShLyyENh0J+3ZqlnkK9ag9zfMnvaLazzEbDs13MDZn
azdSm7gt+P2xVX6wHnmqO2YTEFkDBcOT+yIg9y9r3xchCz5q1A/1vscnycUTv4xX
`protect END_PROTECTED
