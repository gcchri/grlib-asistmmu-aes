`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EoIc+87Y/zNYRIFAnMmZhU8VoEC07UEhQVeeT/mo4ywujFKUrazHixFdMVFQbD1C
Nyd6Q922dTUE67mvlC1hgoiWpKy9YXE01o4a1PRSmhSOIpMvf3YFRkSLwEQbcSI7
2x+II+EXqw4M/C3c4kEOd7vN6C+DXCV0twLNhu7uoPNKEjop+VCbTUFqk5d1WQ/i
P9+//poyA6YSbifPMHotGPc4DOvR9wUVXb/drhGB1v0Il/LGnqYdtbkqPeJx1LyB
stqYOdNtGP5vaijxHklDzLQEJiTehX+GPeb6bT5MFAVAbajUyTQX6NRdoJKp5Aia
LiAsrNAm0D+rAgMrwDPKlHjfm1vh6CfBUWdywkOztxt1Wn3H8Xbaq2xwjnlPZ9DS
VOeH/GtOiYCOAr+pb9ipxXC3to0TnXZs6sTsWTRn45spzwjcIclC9S1GPlPTsDH8
gS75goHZBHZo0R0XQp05b9IrmExP/x+dlEb837Kf3e5oKiEtCU0hSu3rVqagv7Ja
5lUphjwWNbiBv1yPMF/QtTUqp1DZlFH9PFdmlvm+fsnYPJIHAG5QC7j7fVqOS+Y2
8f7XS8se0T8jD599PZNvcmQkRuuFkfLzd55AwAGbhpFN3hkdkxosdQOptYKi3fPC
4JcW4IxQn1zwVzjWX+5/qwuQyfY5cQN8q5vEXP96FJSxmNkhsiJcT3E9Pvkk95Jo
5GIkW+GpEjcR1LQVsrOKeDMkj4O8ydk12TXIWbZKuQ0bobxPlSujX163JcuDaBY8
pWkHdXKhhwCYeevdtv/V79ABi7qW8qFjkrVh/dIKF4nGTb1bGxvUwQg3Kut+pZLM
/cdCMjbIFY3tSQyM8BNBno+pNULcOP3WxvuaH1CdaWcpaNVYd/XlpMaoFwWnAmWu
dm0ajqlS5JLmujGBa4e0UjeyBlV44rtHNOMy2foKgLxVb91QLMrcveVqS5fOU6tk
Kam2+OLZ08/rzdt2KY+44QMOB6wEhM78cwPxlozb8NXBCtU6B2gwDFG3yV2D/Bxu
1qr7JmgwNhl3cnd2pDyTcISAylHoK1QiXwM2XdXRvt2DDGxuAG2prhsj8Jyforkt
urMkxATA8DTPkOtXne94kBJGKEw81tURT1Gv1P0RvvGmLIAJTNM4Xsapqevwc3fM
3rhZbafac+1LokqWUiJCoMuycQ6lFR6BU6a/G5P0qHftE05MuVjW26GC7I3N/9IU
V42FEu8mUR9J2t+J0RhqXnmBhBvwZWcTIcNXJ20NfSCqqW86zJTwbqV+v+twlqHu
OOuLUR3ldT2BJ/49+ApC4LMrnJ1eOzwQLVT3ZlFzboCmbD6JQcZa5VJUlrH4TBHx
HWsBBEbAnl1OJ/r6LJw4UtE4L81TB/Be2G3UhIVzPMNyJreGg0lf0bbqxg9lK1EJ
1m6dtzkBieO9jw3U/clafpE5rSELopF68NQRjOgU3pHI/6LMwTDXIvGUcw1ijdVF
dJ+hfeahdDdd9ke6cdmNe/tBMTLBdJ3SYL/EImyArUjhUO19UE/pNrMEYCa1Z8mD
wnMwyogW4CJdD0VXbr8AvQ1Y8VA0VWsQx/9JX8bLw64eybjHwoPmgYcZ9lwd/Juw
Ok/8mMc+uWB6Q7nmHfvocjUd8FQmiU38guBu47/a1RZNRU4wr6aJZzvwPVkK0VQP
QFoXGOk2ZapMSET0sIpDhYCxHMBp4EpDetX6TvyJWUMy7QF/ojvjKMD5neX/qh6+
lq+ntPGkbOSH+/9arWItIk+/UomC2a704Ss1E3QljswZmPfNl0blo9VRBfuTsMVR
EThkWDiZfdS8WOQLorNsBV3uWjNP3b2yvIoduo2Fbalnr5wxIptKZ0b89oJ+aVO4
l2Tn57Un5YESTvmv0Fptb47eQcKhbPQZyFfkv5I44f5F6dKSoGbstWHH1F7jiqrg
vqE9LhA5LkZm7SjWirPEKGaycjaOSyixW4L40bTRZEyWmIaNBofp2NgJtC9km2ti
6vxBHYDoZIoVvTlOSjvD4mfghNYIx/vScD++MhvxPhAOW707Tl26kR2V0NewUORT
uH7JuOUhqWrEwXZXoklE6Zik0mAZuSUwB37i9FComNwXWGvR90PPScqfnLxcmu6Z
Ij3EJ78Eqgq/d4RFc4r8Ib7JZdqZdlWh/04GkmFfYDqKxIWtjLUHtOBYZ65HAf1y
ZocobkvecjYERvClCqo/yVRrQNq6w9pvbb74ZCpxJ9UvSH1DHVuRQd640mSNgDpE
vot630LOm7k0Eg/NloBySnhOWypyPj/df+6Yh9eoXxvqYlj4qq4qSD9A/js+koRV
vE8VBzIZkwefaa322iW0tIcZkGQY0PEyCA9KhXx8W5wfoUUbICr7ra3lFJwD9Xcx
RYdqaoi3CRAJT5Rp+RUnc6+MTMvq0NAuQ6IhtFWKeEI84SN99XbT0bohoxuB7XMS
XHe+SU5CH21sZ3MNkIFTBOLu35JJKW5KajcSOregNjvAWA9wuwIMOfMxCmOlSpKT
bA3eVUJM38TzDbh/wIc9IC1Kx2NpR/ayq9NzjkapoxXokhtU+bMg/3+XCW25os3A
79FciS8+1pZRlqf9ndcgag7MDtjHVGs+M4Ooz3454lkTzHwbs/d7EoFHractx6aK
zXHXQVsHuzh1CrOKQL2ANEIkPypHHFt7ttMWmE2fDQpn1WEjerqvxGAGS2s6KGos
lIAFS133kNm1IXQRWAj+r11qLBTUgc+a0TYma6F3CUCxWroqsBjJcZbxIzNbShaZ
M/m/sqpbtk85pBQBSZL7TeH/ifOCHQcH4ZOctvlmNXY1oNTrs1yfhuEAOoGsC5Ed
pTh1N6gsSlYsTy8gAAu1qtKEBnW5R5TNEZGrkl02uqIr/hVk12SBn07yJPYJYBkW
MVDe9mdHQWsXrmNxfHXrrWtw94MP53lSgbTfw9E3Y0ES96JAE0WcvL0fmRTsIsRF
P9w7eLmNcflE6x4C8TKFLQJEuyyjEQmMryBGxDRlWkWWh/juq+ekA2SgNgT5l2O5
MG9kubwBDMvK1MN34BfRe2bSwGM2gRu+rpgCTe+Tz0Tj73Avuc8HiQ9e9nCdJENF
5otUUXU1/iB9lJxTlZd9zHEj/l+7kMFj+15aMC1/dE1cE4SR0aQuf7Pzp31p7HE5
/1r6QlSb7r9MYG9F3aO9av6G9JMqrco5/qlAXv0BSWZW4p5YqZc+CltStNY9eOcU
difR0U/LNkIfLZusFn8fTEAYi3Wt+AISkWZZpj9JHNfmNtVPdRv7N36P92q9QG21
xW3bv1ET1SwSS3fu0duXRlEjHL0mpH52NG18/SUdRDCHBb4SznTa1Hgc15jHcTfD
ZSPV7Vv8cZ9B1SQWch0X/xXZS9fs9NIjg8N2CFkpj4b27PnFYubwXHuBNfdeCWtW
R+oGhIxv0Wi6/ejWU/Dag7nr7FRCsII3nj37idrNWTNIxWQBAPOQj9vZBzCgSYhm
TooVJvsfWAfpfWlm3l1E6MxV6iF+0vaN7yfwAq29+UoLYKUs/+mpbBj4Wdhjmvlp
q/5qSBo+H17e00Cuvt58WvDFQO6O6qPy/92numLDM53vU1o6eWleyg0io5LRcztA
ulIPZJxsLu1oyfuieMg/RPyDf4NA/iVakAcTWzELt7mry3gfMK9l8OhtM4Q8Nb2a
pJacA9RAAYvqSGVhfTRUsvhPxr/pVgm/Ccf+Pd5SFKI2h+du3Rg/YkFmybu7xXCV
NeBMIZYmytUpLFvFgZ1uAQMtT+0EbyxNiorqqpw0FIGUHgxa3Y+bI+1YnOc9Vi5d
aokjpsXG0o/KLMUG7IhLhiOzcfvUPMVy5T4zjF5xFuFQZoxCySlXw5jH/qCsRWIQ
bWv168+4nBg0vqkbkVAtkpegxYP8tMrajkRrBPpBErVd0X1QKN8SqEajr0tyGjgX
RZn4/xHvvLXPlys5ZmkRt5GebRwi2Q2qb4P6UszQ+FZAzV5ZNlhrxWN35tB/4yDF
r5V2JAsvIowX9y9/PgtmY/7hX67eUkzN3mgscDSOEjITyaFzQ8fbvE9T/YbiVZVj
JP1O2IfWlV/JGJ9jQqQO2WO+A3VPEjngpS1d7U7rIcxoIWuzquFacF4Dcr+QqotB
9G/Pvl9aJqy6RiTP2EftP5eF3GtsD6Nfw2IOYNcCHe5xTP5P8zTkAf99gEewAUvP
9kD62nB+zdpw7qLBFvU5A/AJ+vWzNXPjUSJ+kxxjs8Agem64MbWNbRo/F+R4qQBh
S/YLR7sLiwML8ilywTmSlPsXbMhEeIjSM+/cU44cxWXVKO/XzQSvrpKljerUbf+L
UywQ/4BuTzEDcWy+aysk89P6FTXGxUrcx6ui3mLkYXPmwekIzBjGuLPiegrIbTS1
1D2Ujva2nCAkidlsv72LJ5xqDIPJCnH2Hu0OZYmWDFyc3jXL3AINvux9kaewt7u7
QQXbJTq6LA+mgGmIxvoeba99kCyt8qfpUyg9fb7FcKro6kW74/dFiKcSEFcIIQOy
urvo0Et/BVjjzU6GYgoVTQcUBBTh9rg04k9bp3e/j0X4J2Fd62ttf+qDTmn2+GCY
T1aGvMvKaEI7nv+DHf5Soky0JFMRqI9pm0PZwSqcR3MuX76EN1hvSYmVzr7d+LEp
qgAc8IQlgAQuJ2IAwtr6P0oT7RxArJuf34S2PPIsPHIFU59oE4wlCg82LFtqfvkv
PbLqmDxWES1VHz5ON8/08xh80wEpOrcLQ6F982tYoV84iS0pij0dLJXhzzP2cnTz
1tQRZMUBYt6GBxbfev14t8NmywBb4k0NxPYa3EzCgg+wxq2yugthAt/AVCNCEz41
x6JEF6j634HPPD3aebXwUrP0nNb3TAOIg9aUyu0gN9th4K5zojZI5LpLZIN+XrOT
MaUQ81NCLsdKNdKpGh+M38csb+LrrhFGks/rKmpm7KJCmFNCKH1noUC3NKOM1HCF
UlYPJAk3KhHOBLcc8OeAHachtEkBR6n5jiPWn5XUsF3Rb8TCgoXuV1ql0pkRno5R
fPINUQ51pCDvXqa3TnzqqGdRqTP1vwZQOFWEio7V7eYBEIKn0+34JDQKT2Z+EHhz
BeAy3Vjc05XG4Jzc8Vsde9AZOUIac11oH6t3uuvptaU5p6PtOOVTbEnwjTYWz9r2
iUgF7eOY7tnvo60nUYy8IO+yaP9HUXp7Ing7cPVc7Z7oLBXEkaoh/uZaSuKl1Sqf
fSExEFJ/gAInIX366hJcyHxIm/9LES33euByH086vlFUu47hWGSF3C/UzGI/X0XP
+6PE0XlvI64un9vbnYWnkjHU3BWphliCOmMhsgkZiEFGh7CrcgKrYvOheTLHHsmJ
Pu0vxi4xeNdjDDQYKnsoU2SlmNifP08njLnpNRznenl2Sa2zbsrjhf8zkTlCL48S
UHEcTL5lDVFriNLjwE+O1/6KuIz+xl5syJbtHHzrsgyH3XhLwMz7iWkpcePNwnG/
81EN3uEmkzEuhacxmUI8OtipRJ7/K48v2Ude/jltf0K3OE+Vj/40LHmcs8nuffSi
UZt6bN8GtPSYc94AyJLQBaowMBwo/TsG1VwyLzkcNhXvJHkL9WbEihdboyhQJZHr
wI6IK2a/9seFdfSeZeyPfazzfAhRpWgBBmBWnzssB7bhVr9hGohxSy2g4NL7EetM
Cat2B9OiP1RUH3OKEPSGNKotoIAHALw8TzYFp4MBJDBxB6H8WXI7Y/z+7uCTLRZc
P1G0It+1C5muNigom+v3XxSGf+BiAx1qcMdcugij9NIlNmfgkpO85Rwds8b2rtTg
wsxO9YQ7mClVycGcV5c/tzfgdF+l/tltji6UHws6NVhNzwLBWjFEW7h/9x9rV/bL
0cQdc42yE1kNcwzgRmhsgTCoTdDCaXoy366RmI3YnviE4FDtSTiyKcIWLY4Mp3I2
1SrDEbBoYnRZndGEX02CyXu4eDnlU8ghUuGtjdAZWRPTMXcIn8V+N/Nm+CZWoVSU
NvLiAac46kwYpUM9sYzD75MgAkz1Q3Jx4qBHqXjChpIRfLhVUv6pnUSt2PTggoyu
pWsyd+/jl8YsWTqWV2EaXPeAbG6T6lJS67ANYzBDFEvjcK80ayj4U4C2o1thuVKG
ZCUB/b9MEr26XIK0pJ4h6NdHACaxycaqpw+E8uT2K1JmrnK4wE+WGbuv6EZQ3Zyq
vxQaCggOYj9w6pHGTU8ESXouZ3/5juXMshP51KCDtOUQDHV17lb0Gu+WCg/5ociT
oSwhMcGEEMTDv+Ym9S3iZU1alG0UEwy1GqxXullvfsxN9RVvyouy2fTIexEujrm+
s82XNbWvPeDvu2A0gTLBtcEUzYFmIQLlRwtz/l9GDgI3CvOJDvy/TV9Tzzu4ac8l
k8lEUU6HH7eOA/WlhJDBFLIHY4HMYiQuldbBRy/GpDnUzeLQKMtUg97gaObjFJF5
a5ZgZX9tkoSGpTQnSpOR4HNcC1r6Uerp6B1PgLqbgiAQl/ZV3fJs0kJRrUdmPuNa
j5unr4uQT4UXwxF3e7u4ziwcH9VVzJQ7ISGjYBnEZlgawzYpC1oHNg9nzfYYLXll
TenAaYloxjrI6T9GRK8WYr8PnnjJVQn/1m+P8ekI95xwQ0MThx9XaI5QHgPS8NB9
5zWR6dIr56pSvqLNwvTKQ8ilpXzlXVlHsNBOuK/ZvzoRn7/wDN/YgyUZkQlkmTU3
f67OHIrbUcbT1pwm+0zVr+WMYFF4NTp3ofNWweaX5Tkf0of7tqzZN5P+KQjRzZpB
A/MslEVIVFGq6wbkHAqA8ZoR7saohEtzBf12I7G5AH4YPlGEZWcJmU7/W2rL1JqI
0gSZsPefjVPP44EBWLSNzckhtZudKBAGaAB5NjlyK3fQQJT3wR36b83xZSDxDTwj
9C7GXjnvNd3izvG+oymBek48tTUkxpdG4664q/MjeCbjWUDMOYyPmk1lHM9Db+uL
79H1fw/WWUlLuDe3FyyBlMGtv09tINQCubigTffTLH1zam4LifLMf2XM8G8lO9jv
+48bxDnFLSx0r0owOjkW9Aj0VcIDQUVlGRvBy4qJk5TH/oiL7bh+W5B5E4dGk+Dg
jKhJYNgbo3828PtUPI504XUMkfG1M514ImEVnFMO701+HKfySi3RDvevrZPPWkKe
D8HfkxboXF1kiTIGCVcKfPQxJmGFDhLEJ30SzDyf58fNvnAVsdw1q2eOeesygb16
O0idxtA1TrsFjatz0vadE0Y1pgckeRP5SlnM8RYUVs4docABNU+I8llCUH7IpBib
vsm19CckHP/dtyh50/4HSm6FzawIm1Nbe/bCG1cF4gJ609DAAGczFjwjnb8+ykLS
3Bx1eGqPzeWjpCZKLG0J+RJ8biW+UUysv4fKJY09i155jJKzDyWeBrPBdfc/cu3v
Epr2u7tKNQOUmSBfeAB1VsiYG3YgIsalmVAyEAyBL3KBz8aANp2i/TmjXHOrUR1Z
FsK6A/Ge/dyxHJDFgNGU61Hc6iQ0gFwIjM9+KZ6facTc6XS8VO4Ox1gQDyh9BM/e
WjH9E9oj01LfdFDavA635BKMY4lSfXFgh/7CnLGjhI8rNC/X67RttEdvuk3XFvxK
GSa5ebrp9DxHhRFC8d/Us705/VbBLbOOQ1s7kXbfs5puGfy+lvtINn+6KU7Yn1QP
e5RyY6NGMNG7JuopZE4meDuSBX4dr4xA/xJz6dQEJ0pAChN025gGme9g4IbEVrSQ
yg5BS9rHH/pfM1kcwIyHWlh1cmbf9nJAmdE4/A0/Zw3QRuhd72YHbv6VKfVzKaR3
2xenRe8bLfPN8fpXC19yAfnxTb3ZB7v4bIDfHCoQAKtUMqC619ivf8J5RHVWudDc
/ykTHebLotMfUFZqKESifcPmEm+0N70Rfigw3bCG9+MiC/LIgIR0GQjkaWeBLnJ+
46EOg219aDKZoIHvKS9hH238+YFeCc9ScOYDoGqz2+MNwFAe4jwUKFoYOfKK9W8y
Ip9+WW6ylT737JR/S1lx3wjOIGSeokPOmOzrN57zKripNbxpvIKjB8J2QLZ4q4NG
ki05X3ZfBY0myUVHmPTQzzSIhsjeveYNm09Ofp6ldQbJ2C0GORcTZeqVx7t4QNLK
EmC/0htyHM/+OlXWkHWQAl5278Jqkk/uvOe8BLJ0K3GbuiROnntpn98r3rNyiVpr
5b+uMKOK2iYXXQntMQXeD1JFXoQRorsWrhzbnWyU/uuwjIkQqzQDla7AeZwimxLX
LQSeWxFtQBoHOvZI94fxD37wAKgyiIjQV07ZJRaCsFjEVzvz0tj3waV/WftYu4LR
iloD7dmJ6ymXUMks0qNZJleuz98RFeMLOBQVPdTn2kHqVXw2tKj1CpjUclJMOUfd
Srs+pA6mhyk3zrlmba/oMkYMfJi8Dpek4BAn0B/LFbslHyj9QOIBW5LBmHrHENL6
dTsIsHTzdzO68TQZM2kx62ikghMgoUFNQiCxuvesTzh5LYYm3yAtmxKtsXH+ujUq
mC33CrdrqV0jnz3sN8DCDpAe4acuDfgM6+ENZ4rC+AurYvnknaE0VchQFThm6mq8
0IyWZzUQEOV2dcTiPmmGygnFQJgxSYCQXEHZOkQ9ARwzSKY2cLpgNvAH9LaAXO0a
Fp7RLddBbn2L/r0CGynxA/NKyvqHMXnjni9P4RnHsoyTS49uThx8StuhD6/xHool
/rg+w7t/floifCBsiYcfdHNvjFaZQI4CVmh8kYpLbiujkUndTtXesHdzMPBjr9y0
+adn7/MYygk0O3rGvZWdNA30+z3R8S/vpVX2hcYzTkPgGkxVQwuRD2NKuwaNU0gC
hPmGeIHmCYBhmasEi0r2TiXHq5QSv3gXwMHDfIPAukn4iIv5OyJ4xGmBkXNHIm7k
tjTwiFtdMSY4wTJ/pWACvXxee/rknWQAkezAnMuc3KzRCSh1BoI/1LEFWh6t8chK
bRH3WipDAnvW9WZqg0MWSNyR5BlZqkQWygcIaNEtB9lY5OlHUzXm4Xz2eIsJBjcU
CcSG4N5C6v4tu9stBp7MeNgwa+SSqPsX1RbaRgGeHE3MT+a9AVO69ehon5bjrCBC
5V5WVkVr1sKwBjWuiQMjiaP0vGZ8yqJ+X5L6EiPslUuhmOf5qUSevYExZvZEYpPC
t1gUM+Qv6bj5RM6D6DxKNNy6rlwi3UXQT/XlKQxg37bdhFGjI7qDgq1xz8sAb/Cu
4ZJZ2XAFU0P7kiNXAFSKLercs8SZonP2kWfmB83z9LgUIFf5q+5266osIZoUI3nh
sYeKvVVdsTdsZ1DieBEDHuA6PArLn+6ZjeaI04ME0skOIYdhl4LiNBoG5Ye3QDth
3sg2990hxzqXiSzDLdKOeJe4On9c+g0BpGVCx6MzHBBAVd8CY6nA0SHpE6gJE7iU
gkFCTKbaFw7trUkfB0z0J/pV3Dc3K8EcsHQaF/OB25YVEVDK1dJAXBYJ2wEB7hK9
J4XxwlFBhClvwBNCHBwUhNT8Gw1mUGWuOZsHvhKSc95AjUaGRz8dtA3jzF72gSuj
613miEbyVtufbJ18fK6PlSwLiccpa0k3phk7IzgkuJh66juoPRFPeMFRxA35vknA
FVTvXBg4DbXbYL6/HsIbrNmsLxl1no1MrSNOKLMvffkXNJ37Bm6BBFaFuFlrokda
8znfnyAa5x9ccxPcyrWyPypn7+yajVehAi4Bq8YC1SWDaOFfL8G+VFNvBEzofyH6
2oFazp/BFW6o8HUZ4L3VkWNokdaqYiTruxVcX1Xzv0IChVOEoBQqlzvTnVWRwLXb
sCTEuL9FyflGeMneWDY4zuZXASGvxW10nNVGGYg2nEFpGDzbQ4E2aajPdTOQQzMh
lL2RZTZ981/dTr2Wl7L924VkHKLLCyhD42PCQ9JuBBVdXZ2EquVFfDXbqDQ41lQG
mAJOs+qHWuzM00z98EFPUOuRaMV0jyqxfo2VWK7+qauNIMHFfMDBi8p7P2BglmhZ
0m0FmYwbdCBjYx/ZTnt75DEBSC4EX7xB6rrWQpjg1w6C8rYzIzyl7yR4imfmBs5r
/MxMmUY0sh/KEgdzgYPc5MKtxF8DdCKI9Ct9DixZ8SnmyfDOL3RNRrICFKeHQax5
WOhQOhIKzCk/0pCFxibHbI+JceDUNab6v+c0089Y6cpvrD7LpfD9Nxg49ZeLJF6G
8gBKmiObFz6G8QrARGh2/B4qhqi0TDpRmb2cMQG+AxL4/Q7vPtDmCLGlPBDPdlNq
r5zFRbC3wDDs6ZKH5cMUDVfvCaVcmxkkGdiJATsyVL8LdY5jru9UBBRSaoMGac7n
i2/sgP6I2tGz0uJwYfCl+023mhd+L+6geQAJ2C1MilDFV7al/d6ZRxjq7JcNDiti
8R9Sx7nqhBomnysqxVuYvpJe3F+lzIRz0XOm1PK7LEguwIBXD04iBSnEBSDr8o4t
dULrKWE+ctGfA90llN/xOgm0RkBBEjfWJkiJmEHtQ0PEiItNSjC02Y+r9JeGodJb
SqOwQ743s5wsmBXmfYVN3KKo73LvL/Zu8m5vQX9a+mFHL8MO27Vm7aBgOPDdBi6t
ow+4hw69ShdTUHMv5h3NnNkDRk9FpGOH4ict40cnB4Ot2l1BL1OgfFRJwXMumTLU
RWlxVX9s/mdHSproVz679fqBi1k1teiFQ1dAr04pEp0Qwv32AcHqsPhzclB52jny
Meyf4vu0HxhN9Mi9BZB3S86z+42pvWjCdCnwda1h5sqRZHoxu8bfh0j+fBvHGt6Y
55RwQLHcj+db/8Ox+U6FUthMFfJNqCONwlbBM2Spu1pzvSepemSsbdqSDy+JIvKW
WQk9FgbQsp58k6mxxjDDUNmrj/JOnS1hkmI+dOZU49v98H+JAQuMgM2LqR074F9Y
AdBM51HOa/+9COQlbTwyIvnecP7wOE1VmqgVIVUbUllVBkD4O/BiuoKJ/+j8WM+y
jLYIges1jIxcjMvYZ9VQ9RGD//jDGIAGusDT8vsQx2EmNRLG4H3OfznEbd2QXJe7
3xcUbxZEtTPQ2FPIEPiGojoERbQ54EHeAllctRIxBrtwTOXYrJmy2LlbNadA/8Os
gLskaxdSekjdRw2KFWCagCq5HwJw/2Qn5HiHr//VqIKrMqW7RW1BMUsFmpaHxdl3
xaxggc3LETWcbSaKHxsaFbSfV0IUo0cE5QLkplxNx9or7qVf1mvRQDijO0cUxXmr
ySJcQir9qitjIzulRmDb9noAYP11j9+hniHVaBj5YBh26DaN97NAvPoTx6xvKqGK
hRUbzukj+OsCWh+dVt/HrhPFliCJY9HLA1ZprEbclCpEqG2hPs3ThvxGDXLTLFQ/
4wOhEL2I76Ekuu3p0tY3IaRBKoXNs6Ov1KdTjxC4ASwUO2iCurZhaWRTJlke8pEi
bWLNr2nCmFR1jL4dzxY/ULn4omHIsfm97ImGM0SQQGfkMpnhsZl8fk1JCkCF/iG4
jLKHtZD7AMi9GWsChMX5WuaV0PdjfW28ORHbBKMJbhksRcerurnmOrDAy9Rv8bYs
NcfTjn2j7WVIbXZVPG4RZ/kxpK6HOTUUj/7rPuksxouLx11kwlG1nwQcK0XTMeAU
ZMCiZG+c0M8d1Gw7xTymy0AqMqzIEuQy2+ns+LWJiC0EKWDhMqBQfs5wBYLzlAak
FEfGOwSiETzyGjc+I4quCWskTsSTdFsPHURjvG0EQPM5nNYCKLWArByMgfGLmKIZ
K8aDPt4/WHOJOqUcum2uskca2es8wcrp8rWoRi5xUtBRTP2cEqyyz24YLQF/pGfB
jAVBYAEnboRorIa9x03Xza2FfLid63N33BGEBRfzKzeRRLirdna88FnUbgvfieXN
WaA4Q71jPOVfjNiEgG2KAekCoNQgTzXdIQh+PpfpsOMaAM9ZuJXhThaAwR5m17D2
PowX4d066evG8lsuqkkEMn6PhboPQTEKG4pvH77eObXwXN0smhwQgWpfTNpCet31
Xdn6BxEBIbgWbiwSpqcS4aPlpoaArjgRTBUiY2yfbGvjI32f3zpEZQ5rL5k+woB9
MA0mJ6gnvFc2kxMu44A2DioXmR4aEIid3Rnjn8a8VnCPD3702k9HtTBopf5lNANB
ssiWwuxZNl2l/QZKP98wt/Qo89LcnSUSEDVfBHuM6IdShM4TKyzyzEZBR69yr2M7
UKRvReYGzNG4QSAUFDA3w8q6HvxbFv/f9O8IWxBscYmk1BOW0ktAK8eOkEQjYyzr
LOj6UZd4UJPPG9dinKXoSA==
`protect END_PROTECTED
