`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0gf8kSOGB5hqs8W621DkMNu/AShh1gOcJdWMRYFqszb0I4quYADgGdtfOlev9dKl
ueaNKfDlBY9L6KTH3JHS89jTX6vt35wDmb75Pojy1kQY+zWMf+Cro6TwWCzw/63z
jqumM/2TKOrf2EnazyyXDGFaKTnFK6VokPrz+eyjRRIq+M7VWuIWmlZ9/T8UQmPB
uG8tXliPTA++ZgZNx97A3xKd7N+/rlVsJ4IVahOjBPc9VuHal3lDCuvoP2IP/GaY
XVP/A3hnWOBY4Ca3K6mPg0A56hqs/EhxGBjD9di92rD95RNyOaRyMG+ZYJy3xiIM
53Pm1reaU2bC/PiNr6GEnMHIZvUXTUAkOckEOFRLK2+iYscfNiWHpAtdVopAa95H
h5RkT59N5PtCnbdaSoNQmxon5fd2hl5oEfKA1uPl5IWSVfI++OhsDKrIX3Xo9Q2V
VcdK9u6/WfGOR1wwOHqDbcri7WBwqnBHOW+NB4Wtc3RYs5aKd1BGpr9vzYXs2yTa
TiZHyfz4R2/i1QfI+CKZmfUnz8n1WsOyOtcjBes6IRyox/XDMSLwJtlCqN1Ifve+
cbCg8scTPA7PKMyoibpf6BHNJSMt2LXbG1ibKgoiOnE=
`protect END_PROTECTED
