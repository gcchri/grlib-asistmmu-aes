`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aHy34D/23mL8zxrmsJnPXsu9yQelCKw22hj4w+j4PeHIsNIuHOo3gr0/qOopRU8o
RU7KpEaL6iIFfZJC6ypbDEt1kDVV4j0X7/5K26eIsqhhVcC3a9kfnyWA18/OvA3y
GJXdAxV9/Ih7f4svG1CtRvNb/0DnlcSMbLmQy5evJ2AMo4LMgtynVzAZC3YkFLSV
v/jHo+Mcrc44AdoR+ogM+J7dfYBdtrNYsaFTdG576xD02SU6YZ+yeM3mYHqBdkmP
flO3nt06f2BoS1vXvohpRKcgvRN+pRAHN2QbANRqo7ZIb0E/qqeTcp+SXJ/0FkUb
JPNZop2KST5BrUn9ukP4GBRoPp4MXItrFl+0aC+WoyUlShkP5LPvsZ0FrjLMNBLp
EkStG1Cy1z1ADl32gUw2QvHPSuSu2AfnjWXrW3Cartm4er8TjFOqr7kRTUFQlpRu
omGz4z0HEyEFgjuvpArue0nAYcOVWScNste2qaOZbu4YgLCfeqYyj1hKyOZrHJFo
HDK7FmhNDYI3+hVObR3BZpElxEYHXMBD4DRTrEA/dKfX1r7KIGtOVlFoscNrIRX8
hA8aZdWiykAv/0PnHZB1vLiXsOwzfhEyZfCvX0saBWu53dXhY2R6KOLpy3xkB0BT
0eLC+6r+cADej+X9hDIOI6Q4v3wytWwL7JaQXNIWiC8M+BhYWIDPz3Y/VNnTtqDh
LDAKXC/FOoGqb6F1E+tGwwW8zDDCRRoQtDThWsgyF/CqJD/Za6hO/CZdTwsmGlmj
ZLOntfif5KwBz/DeU7x6nuraUtuK6WlmkJgCkgOrqONLuM4mbXS1vPbrC0VZhUgp
RtwI/sA2pphWDubpvu3436JKVV8gwzvBzu/ivFrE9u+dEUJHggpXNEC+wtlrbs2w
ypZ/FPfYpPzV59UWn3tyoCMAN04XtwLh88YXBded8flMnp9jq3kKU2bWHiW+J2v8
BNcoqjYeF6Ozh94AYNFpeAhXFiqan/eGOOxYGpaQM+I=
`protect END_PROTECTED
