`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+K6tecC6hwx8b34jipvw266Oiu/n5Hg2x6nk7S7jZukjXVFO+uSrJhC3CqO7lzj4
3cPTIcIPc7/cwhzLvH66VIDNp6xKvZ19AtbqcsoDUicCXkV3GGc+84hwI2pR4vYr
lDGyVBQJBHqSCfiGW1fEtVPuh2RabU6HzF7sZwbbXMnMkO67HhCImVmg8kV/Yt9V
J8RW0DGB4hVqyzsCM4pyJaJl7gCVeKOYC45fdmD8ilPW0mDMQtaAb4N6672p6t6J
aQwg3z2nP3iNyMRrV5OR8LRSh/jlMnGGlj3OAxW5wKBu4FPPEMCV+t5lHmN+k2WX
2C2zxXh8uqIMnlrYnxjFQoRag0T3r1JXABwK7IEinFiDDNSgeWRBc9EYymYnTkLz
sKPiFKUqxaZVggsJkkeKy/8GLSD9KUEkjNp9eetAdAhm9DsIaLgghSJlNqU7W7Oy
tMNgZaIRxICwtRCpDj/BYlnbZQ4UjnaGB9qgsYiFfyW4dIlKyII5CtowFVh/80rx
m+0FLq74OuyVxurY/Yfjlk0CBE+1HWtW9dac5nMcS+BKnu97ONql/Mer26x4A7Hn
`protect END_PROTECTED
