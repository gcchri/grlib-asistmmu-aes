`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YTZ/PIK49AWeupJVdQUcuOu8I99VyUSjBR89t+CxPtyGDuU9iqe6f5FDF0AdSkq/
a0U9bn6RkoQCmifcclA97R7Ha4kCp5drrmvhH9NCWDHWWUVvXeVEr7iCspw6iySu
CcS+X5w3Df1bdfIYFvL8s5JL6HvaqY5rHDo5W1RSIwlY/FB9ipaWQzf4t9QX1Y3C
ewooTj+uZB9aPLMgqeAo2QRlSuVncemyRYIk3nfabVKC6UpBsfA5mdrtdFyiN/A7
FomfKw8yz/aZjMFJqu3gZvD8TwI5z5r/wgJ8+vThlG4DMDO+ulyBlQppajZyuwyM
BH2WcENHB9blRuXc7ULk9KdaxLSBujyBZ4SwmyoYptsls4vCDaCMbZUhFBskOYgu
FFC+x0nXuYDpW17c2+xQ7jCT0MzDRJOKlxt/uZFU/2wflTzkgLxfltFc5Upc3HO2
/TTGh5ry3bATBPOaRtv2Ii6GspJEz/+b4HV3FoC372fUbRXrVt/ig2Mc6WwMyjCt
jgOhMuOvXzE2Bl0hh7POa6Onl60A74mt2Ut4O5c+MZosf0sD0eNoekVKGJ+jMM+N
BcwF4KVnW/eipH45u81tTWe9b1CpMZDxoq8nrFLEbUzAyyl6rqN3ZhhhPgJ8D01q
BgoR30Ft1skM5S7sCFvMXDjUlNeyfZC1WvhDfqV5++5BQa9bPw84VhmIK16n4ngO
NJKBFcUItfeWfE1QLvSY3mov5pElsGY6jDboBrwMFEMluiTFk7vE5ta5BBcyL08e
H/aCmt2TREWY5x1hDybSpw==
`protect END_PROTECTED
