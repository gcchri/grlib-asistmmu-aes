`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Ok16xn3tZGv5UPKGguBESet7k+f3/QtIb3yc1JuPsKggt+5/L7qWNh4JoM4aYCO
HYP1JKHunhQ1cuIcZWZpNUhFBBZA1rm2SXLnvPBoYiHvpnwVsb3Uy23MpowvRquP
B+8r5YUT76M2scf6cXQ3QFqRDVnJ3m1T2VNB+icDKoN82W3fQds2pw3AsvJp2YnJ
cocw/XMvxxL/sBIW5WuPwWo0ZJ6KA23wN4HQ0O3R8RnpnXwU1bMqWMpBR7cqTFy8
mZ3NA0sB0KoMxp+sIA9GZ4chYsyFWXeAeMLYWF1JBDG7BGWFOXaSBDaqQpto7mNY
Xwhnh9+z54AkRNfYPw4ELdUShEfg1HQC8tLrWpsHGTyCtSFwmgdEc7/vMRjX63jP
x1mOWhK/wRJtTHAvwbXsrKdLd/6FPwbNs/M4aN2CYldGcD7MVIylYr49JmTATnkR
v7DRDuiWzMI6GDTpfXHAkrvbOHcnfSfYnhs7ncvlhKnzKaD7bsZP6PGfY+kuHw/o
c7I7sv45PAJxS8t9uY7uAAfmtF6tW4p7TpG5+NCsgTRHP9UcIAQrl0r3qDl/3dVC
EggE2fRpS/emGv0owTsus/e9QElHmVhpTTzg2v9FOvhJQRKAlNUdXAi3W7J9joxT
Yc32cuIerl0gvwEHY8xnm0PXxx7YpZrtDScJaP81Mvw0X6A6pquLLFSHh8lpRlqQ
Ba2sP7+Sc2Jqd/gq2RkkPTdIhUuWGEidf8oBHhyz/v34UMwgyC1vedVBGhy2Q9Ct
SzJ/LS4ZYiy2o6OGK/6zOq7hnj3F5DDrQBwCKYm7gZyAl5sQy8qkye4iwLAmk6Vr
qX2ObYKAL67WAgitkfSMA/y3N4JSyCdy6Mn2044Gnh0czqcFDbRbzoJ+W6hIaRqO
zjecbu5TDINmpqIWigkUgTTNbotPpk/4c4PAO7GT0C/ByLJ6epLbEq3fmhZS4gXs
SNVfQTUXpoXgRwNp13alp0jpdgl0G4WaJAM19AKCfuwpBRN7ukseCaSBM0wzjtcy
+ffe3FN4uf0np+0aymDRHEpFUOz2prCVmLvOwO8LlLO23rqwQE28a+yixlQpNlWR
UCwh8p+gW3OTG5cuAJ4Vt2mOBXrCaBVg8yPiPyPgXsw29k6B3m1jyhlFI0kinh9e
gQIzcUksd44rbtnNohRi/XW4S00+E9WWDG4i6xY3rl3vr/5FxIKTUPFIpFF6SKsu
5+ywcjjRE0ZUL65xaSMYjd8S7KCE5syUK8xiZi9aBirBtALdmrZdsqmJOfVS0G5N
V95lLtJu94PpctcdfWSsr9M09+iVRWkgf4ZmV5m63oOM+/H3xze2zRG17cy8oOoq
/2a+E9NOx3zCcPyMl+qmR4mhXPN23WoymGWZ+j0TJD1/vN/jQ/rCKondoyrhPvyV
10XpWlpYygcAbfl0w3WGrnOGaenciEXRgBVTrotCq2+flw59KTEZ8S7tcsjz6Wpx
jYzQE3gASoNsMD6+jyTnKGAR/lTJrWoLRd8Iy9pndC0J4YvpTPtvxUx9eBh0AULm
jhWiqEebm3/YEiMSmMeL0xUF2f0pt22OeDppfoncX76lAusO2YcXzC9lceHJXD1Q
09UfdztDii+Ok+SNZBAtbDHxPLL8huyW0ON8ian+m3CSE+i4HsSCEbFAybN4MK83
YtmkL+cZTlrD6vxlB4BxDkznE8jFmy+17orMsufR9R1njnhCGwwoqexJDs9ZyNoI
T1sP+DezpnyRkUou3NIk0j6H7DBp+seE6UnHXOz377+wWsJOpnU2WhlhbkqCyqyP
7pEuSLKhfG/LxNMrUjNY/887kMXxdSTXUR7x7kWrDMTHvdjrRO4PB2iMz+hCz942
DXmb6cGN+8iYjnH7njZQXA0qe6D+W4doiNLvx7LUF05uPCbyIsiUFddjnQUbt4lE
dOmtQKTNBUJKsDS3mZAOqa4l0UcycIVYGYUBBzqKSA9A+nPyri0VNFBQRE1GMZ4j
/dzVEUIWIRhp5+R/0s2qJ1+jiWU4lLebNoQRvBKT0mPpzApT4VhiWbd+JlKyBlIK
mIBdWiG1SFIA/WFDxwIQRyq+K+r675LEwdU0Zi8t9b74ccSfI7wCLll9j9a/3xo3
MSgLe+QgKqmqRGv6rQSBTd7v64Z9WT+/oBa2Q0FcQ2g1C5S8lNLGK93GN8RQFYZ7
UJXCPGPuCVEl8l40mRHPrUsRrY35y96Y47vzUzcI0xFTzAxnso0pGm9yK+e8j093
O0xnvEx4mdSJPGRD9mZ+lCvprdb+GHnxSvodzwWnJqhB0yGYC199tgbQM62H88Q7
mSaFHiU77/Rw9+SG102kvg7UXRTe8nsNYPAbUF2e3TSEzlXNfNBeKd48tKJBxmNK
5W2Tv8e0l7D/r6jxZx69PGrYjzTVeNJjvROao6N5ekkzJXiUIti0nxBdCLtoiTzm
GrANak21qq28ag4osAvQQzq10BcIhrro/7zOKpfGxYN/Ue0vclRpcrkaGixudyPI
fac6A95Fq+M17HczkZachWqHZLJvkKnZ6QTsoqZdYFKY7RluWhCSHiY345IpsKpQ
eE897yWXGJBWugqtLwAR9AQKlDbgCHDw8vbi6Qc0Tj4iAOwaTxJhgIuG/365a27M
6+1SWhE5JmHu3yBjVdsM24g1IGELI8R+CW++ubi7nDL5EUGwAWvS7HsO+lq6cZ0E
GN57JcvU5gBUUdVmJ2gOw8eDfjlN38/hTIgQ+jaqxfxPv94t/bBCcaxkNiKBtOh3
1Dox5DMcKQTYD55rY4oWibhvfG5wu8nONAzHstU/DLx7mIsrIO5MlDB8XMJ+PAKA
BGe4i7Qrttt9SzX2YwmJ9e2jLH1U1g/5pbcsH2QtbWKAETkDOkFGk6odOVy4aaWp
yaON7VUGhKCCX/XMADFXGzV8wNJ5hXOw11gVP1Fjs9wgRtrHGwZKLIVNe0/twtFt
slz1+7wk5YPFIeR1Hn+aKoOKqolBvIeBDKGgE0RBD1WgZQ0i78y9roWIcWOgePKJ
FQ6KbgUvXR4X0PLEP6oq0OxoI/2Cz5uq0LRdeJshbu/TAxWZo3tZNOSZVH3Lw/yI
a+cbk2guqSvtenGitEn9fq4kaTXK0sk/3smmQWFavu/BMDtaYTaUyB+t9uxZB+vN
4c8fqs55E/im91zhconIQaIIHpc0Crym7J4/ScKXVTr8YDUklixG2RXzEoOZRAJO
xzoFvEuItS7h2HPscxp77zCIlu8GE21E9mM1Q8PTMjeq1fmZPehU7RdiH1iKbV8f
QZvQbriKPCacNICzJvOOvp/dBYtKaqFiU6M79i2e+mNjrvdF+dPR3WFalMEUD70m
Dl3A6/M5uIHP3ItK1wgU61l6HEvnxCB9vUggg9RFv32T3SZ6/2sol5LfYsI6/EGo
wiXyOP3DHOXykkIeqDJqIoaRs2W1u3xZGZYQ7AuA4CxekrvawcaMzi+Bhb2O7P+m
SXx+vcpezYdo+gF+dg6Uv8+s4fck/b1/T+OBqst2pGk=
`protect END_PROTECTED
