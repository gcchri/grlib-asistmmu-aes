`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EvMa4gFRTwYPcWFLCVwIy3GpXzb0fVXo/6DbB6cTvPivw5bFEZb3HOCyvlYmdVf8
z5NQ23v1HQ8lil3ydAs9jIRsX/psNkWC69av+NdGL/byLx+7fhJ3oT3QUuUF17KI
6kMZ21z13btu+JLZmx930KcmYPxllNceN9BKGUWanqCPsbxKVS537vGy+E493ELk
W+GrJz6vqBfzJY8z/orWCulHDX7+p4FSGreJ+xMp1BkuhB7mLI1eosfAyXwkhH+u
v8ZEy7ynhBlP2iSciqwlPeHl8mgyxXvv4rdDWmBWT68e7wyvY7B0qMkIw7Zrt0Ca
KbzSn5ZJDWf09TnWSdx2SS2EU4vUUoVgpu9ygYhaKviQKeR01m8LSgP04ZeDSXJ6
BEVsC+K+hRd/iL7sErm8Bg==
`protect END_PROTECTED
