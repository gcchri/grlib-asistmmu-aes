`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ibZnwJd+AqbkBDXevgIozpx7N5KMuALN6dvBv6Czt1MfJ2GJ2TDW1gzlWymNzZWK
B627z6hYkHTmqSwm4n4MGLhpv3hCE0SIFp0Y7/yXTH3U4hwFPBCFKiIqfTG/V892
HWYoczhJQUeW+XWepi31ZEFvP2ZXFPM56CTAooMTFn8RVRsXj4LdY43nxE+FGhO5
KIGjAi3Uu/kC1w4SPcMNilGXwLzH92AgnLKSsgZCALhDGQ2eyO+nHoWLdueVXMr5
9N6pC3GvDBiaxXQOfbiLrKciXtN5jInkLEi2d2Kxyi0sb2LQvsO87JzXAI9DhPku
`protect END_PROTECTED
