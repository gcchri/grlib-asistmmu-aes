`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yJT29oYxHm8hDO/tkkcrmS32TRZplDMIVtbTcY0/br/U4moKAV/zjYS8huzJsoJa
2V4wO5JLR2taLncTOqPIqD7xj/lExlmMsd34lMlaJdxSHJfm05M1WhDcQt9vYB3h
hYSu2Hmen4DR21M5D0KMYm31iMzjrTK4pGBgcrzNcJuVbAEZ+DmF2ziDEYDB+g2C
9aMOxR04msjOLRZwPYLQdvNTQ+ovIgXYY/GhvhQKJwv/pwv+lH7fIgRZg/VlR6U6
agA+xLpVtkntu1PYIFrjOnBeHEpasg9FqWP0eRCL3Hz4lkbSn0CvOfYnPmAPwAkP
Sln3CIGkN78ZZEyv8S2TVPSsEFYAVLboSqf39NbN+fL8J8ivxuFNwBcsFrcwXmsD
opXCmItd91n7qlZut9oPRI8gm6YFXeAGWBioFBiveiC0AQbgANPls+QPP37qAHVK
0x71wnmW4TZZy35s7qeG5XX4pCDQFcppV1EgFbFU4j29TFoNLR9UjNGVwuD0sLeF
qzDzhZJ4ZEi4k20bs7oJ/a83FPMOGebyFWMBgitQjilM5mKIU3gUEwiXdg6C7XyM
aoyLPjy8TTl4u3GyWjOr7zgqK4xVQZqMB/GGkvU5tKvFrPogBdpaYNj0nMvvBzyJ
+SkdK2k2eaaZ52lkCeuuqDXQImNzLyfV3CU070dPNTM6sOsPgwYmca+mjsvonjRq
s/85sYdsDSuUloLpptV9tPqDbrq5K6z9xBupsqxhXqvbS0gn82WNO0fwC58rC1NY
GU1vGcJjxQ/FNLJLwGkCHDhdLucEqySANYal0+wwOBV0kmb4jldsgCf0HbILsgme
bJBKWwS7CfE9GqIfC/U2TA7dqzdFenuFxNy3BWRaf15ULhtwq80M3v9riX7xXcGq
nYAPHZ505LUGr1gMVrD7oiwp5n+yPDi+o6IkC18C2N0Y4daCohwzkb70N5Uoq8c+
/o8uEAcL3Z+RWKYkbFu3K90OsqjkReOJ1i/A9uBMxW/wWC06WkXymghhXj+pt4Qf
l1pmxX9V/IsOH2UOYc+WKXUpi6lNcUDObZgaV+l2PoyDBVXp2On60uvOP8ZFRCmE
ZMzaCRlG8EaBDQSWRbhDVyZspvGTKjWhiSEDqAHuaGaoA8CIiwZppvY4zM8bOU2f
oEWGvhDstWCSDuLmHAMd+F+P5+AkQmtCVW4j5qqg3okv3JecjNUSQNkazDqcXpNc
5QKtAvRGTeXq9KRsXZmvemIEUX+Lcj3C8eMCg4KncEPnhQzy/LmjWrStFAG+/NQW
z1i60FWqSJy9aMM0Rsq1KQqoR5Q7Wv0/9nMy5HmE8ys1glgdsSycWqhddM46h9hQ
h5BLRPQmAqCbaDDqOzsykELK3Hc4yvHz9+AM7ghdVoAVAF8m2bpSpS3LElpUX5O+
`protect END_PROTECTED
