`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AUz/MwNibh4e6Jmq5wzzG1PhgAwcoKSn3cpVf4nXGbZvShDaT7jirUloE94Yr+Dg
sNaqIZB++H9PNDOlTlwTxWmR52TTeNpbgpSTGEiQgmbD2gsF/OjJoyItxRBVA437
6nqN1I9cZqdgQ21O9DYQyuJK1WA66CI/6mOpHCrLcjWIPd/gCAjfL8jTvIaKza2+
AvqhhdNggHBkygs7UX4mWtxMd2rLIxcL4MSMniPO2/r4uLaOVGsJ55S0sIndu8pd
l1GJe4MoAOkBS0dQYfI1ov/LQzuRKRVZpIK05O2xKUL7tw4VI+2taSfYPRBB6uz4
Xe0OnpdKQNs3LbrrmKueJd9HhFQ5XpHjAIzLml/g/D14Cf+GbxjzAhv6VdTsKKG8
OxqaXUnNFvoYS3XwEomftFVy/BkMOmJnSQQ1fZYw6xc+NuzBKihfx/hOCx/kj5/Q
xgIDrw+AAen4dxqMoSMH6w==
`protect END_PROTECTED
