`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sJ7rCWcxIFGdBwLzN8VmFG6ILHUwkZ4rASn5aRD5YidEBnho9VTyuSIwOqA9TXD5
mSTB2Mo0VECbyAoBdaFc+3ZGEj+fbq6KG1oiVye8dXirl1bC+6K5BpPivSHDYJIc
ivBvxFaIL7ISgrdpmWK3NhinLTuxhIcSqLjUtQQFxWhQdwc/h6yqrieqA1kVMp46
2Huzn7Mf+su2JEF4hhP5zRCi6v9dLiYpwXC+YGdnSG0Ws4yLf0pP3cLwFl7Ke4pg
n5ujvr1jnJYPYcjRlVmullHXlSm5JViZ6xSL0sDOwHMQBfsYzZRBKAjTB2GezZp7
PT8EJYBBM2GB/N+MPC+ezTNaru3q1TIjd2qFXQVweROigVfPlsuwg1qDB3tqvIwQ
OJRKSi17wgFthfCFSMBoMmc8C6OOdO7RLgVnN91qYi6WAySRDcv9dgFCl2UYD+Xk
ZI8YYMWJGhV8C7qyAFuTOGPFunxXGBwkkW0bvPOwS9oa+BT9RyIU/EvsLdizne/k
bsHrRQazEdn9HfUdp+kFUHWxIl9RsorYxf3XwYdu9xXd4/QLrcJi8mQSBFPQVCN4
h0yr7efpyt6IarlAJXKiNdPeNSFgi0HeaJJYLdMZrCumq8DHkiXf0s8r5woHXvYb
anhq7dmIcds3DRlH62LugJhzwTEY3R4Ei5Kt/xqaYL1Mt1ZPWZ8qWWDddsJ/pAH8
cll4X+wOsJl13WdUgDXqbBgDdpUX15V0efAPJUpaOvhVSXKidH91EM2cdWj2qXXF
7VlOnIe5RK5EV+Aoc0+aLEz9G9Ijrhx8cdQYpacOLZiEjB/W7L+g8wIz2hSxeTOK
2boIu0DYCjZRX1DA49uBlHtypnHutqGX1XZu3l9Y2iU21+rchQDXXcm+g1J9YM6r
zNm/wAfyNTIF3V3UhuNbWG+g1OzmK8RmoFdBmLC71Kew3gy/EYgUKI7135Xvbq7B
MXQ2AdKqhwApX6IslL4msQ==
`protect END_PROTECTED
