`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9H0U6bKz57MbYhbXhVgA91HKZpMZx+hpTD2VIUWywaK9eVnKC1qsu97xlyKHeLcq
LVFzrQy3iOamo/KDv3PKpPWJnYjcCmLnMdmGD8eIelghnDs8NQ9tFI5aEzBiudHK
F3uEnGEcazlGQl1eSEDNVApqeD6UNJXtOr14IRfNWH1CiH6x5PdY/KsgOLBgAU1z
+t1mZIWViLwdvsuUt1TtqHvPrbdIAF0xtwgUn6gFQjG0x8+KxtG4VezWMMUTCjoW
qy7Fecy+yfU8ZY+HzmUSanvh8VFI9B+SEg8mYpUpoAqU0EdLK1wGdqjY2FVOLLrw
Tzg8WfB/BPpssaJGh1CKSU1KfvE9JmSgqK3L2CBBQ53yODhMBzhMvNh9dnmqWOZG
UCdg4CIswC1cGEexCGhZ8O5w+8XNRQP419ZIj8KONLv57ScbDHKkkWypi48pMeMr
eIgKOBinsycl86OJd+OMeSAdK3Jagirx7f4RVMnrA6z38XCLbz5oQKktxSrmUtud
M8pnsYi3u6fiYiEiHd4ATq/cv4adt3LlNvK7cTffLXHOf0fL9VvCu6UPSs5/G+eo
r9kij9hZGJr9eUwfDnzdwvKaz0DHCiKhccuv8mcmaihMV2HspIl67NI2RaNGzCZp
6RzSwKyPlb3lS+lZKIAlKAHzrDozQu4wXsKr10goPtrYLqdfwaIG8CnSccnz/QpY
zLX02Rd+7OQtPYSD7HHFaaohHo8PM3wm0E4+wUcGh9ioTRrkmMKY1+Kc/+58BbCv
QoGUSAswvoDHBXPvvDq+OK1/umm1FwGmektsZtEJMCpxDFmO2+Yr9wvD3oMYsP+g
Qbds551au4Wqs0vmZ/YtT3lSJ2TqOyLdj9mY/Neo2zSjtG61D+r28wdEi8ogqBMt
CVvBIAKl0rrZNR7XzHNaHRqBQcrTAeF8CF0KYdMggw9STUGiIcxh96mNwwAmcK+r
jXmj3dBqtBSLw1E1oCqbiO8qkNwEPmRX0mVW0HfJoIjP5tL3AWDtANPc1eu2ULCN
7+PtAW7eiXd6uIRtu3vqevtqdamhHGF9i7npCsfXm8FhXA5ssR0S8F6Jka2botEq
/PjYWaIf+CMKFpLluVHYea45SA75xpXIauofVfxOvRzoxE/mc/bP+8f+7xanvKkQ
ZOGXP3/d0EcFDFToJhTv8VefyLkBF1w0gGo9uytD1S6CEPz6MztEdl9ppPLNAnQy
IIVgoCkpvoTG/+Oagt0PFR2pa+gyhnB9ab/YFb3GKy34Gi3CsZBENcvl6IV0Lge2
1JC5z2LEd4GVemamMEcPa61Z8ErYT72aznLI40W9vTEud7U3qJakT/fd64YXdCQv
pic+TKilQlvpL618J9eTbK4NlteNgNUjMKAdra4IJx4WtUePhWSoDJxFZu/5Vx6B
Ad7ga5ifNzrk2lwpqh2Cjjl80yUOBEwjIs6PvrLW32hkWX+VRrVkag4Td6Cs4kzG
pA3/K7Y/2uAiNCQepyhvC74ephmptLsx5JYRm0wPA9k+nZaMb1IWLWZtYNB0rgp0
bLWp19oQmuJEAXKhUEj0o7FLJCBRh4HrJjFqiy1vRRfWLIxTV+RejmkBXGwZWpqs
`protect END_PROTECTED
