`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wDcB49I/37VkER5wRGvGhzMMoVmfhHeOE4lvB16lFyhWm5c+0P5oEEHeY947Eugn
hoIRRHPhDRlHfycUO9p6/RJCVfqtbkMGSr4L8eOW1FR8EIYhIXzgDKkG2w+xUQIP
GXBl6L5g4KMFq9VLH82DUWCUjs9PnLXFNt4Ovlcj/CUmwJZDotCvk8RNnznsbpWZ
5R03K7oyJ73vG/56zaQc5UfX5qYnPzg/i1ZYbm4aA0JSYBjibpNNdzxK4pa9YI2e
4u5cetGYON6J/nFNFUF61+RzBwGmpmbN7jmI17USM+a9NDJ/2EezabWdCoGCQ55I
v5c5Jatof6Bs4dFg0b/yhNSooxfnDVHuSFDB/22tvxfquytutwOBWn9vqVO2qWpr
r3qU0TFY7fCbYgPHkR7N0faqfijJgUXCyQrGeERw8+oDf49qDPznYUURLwi1rsNE
sFCHt0RdEeg6ut2vcExvjSahFfDKGQ5ln+u8pYWxEq6s13sL41luWbCpeWivWCNs
TjDCe9eaEXKyNXoPNaA/wnT0+qukL5i2vmo7VFICL3qcrNJ9oJHE+UrambdFOFuB
0tFToHxuF2xdemk+u6FhGQ==
`protect END_PROTECTED
