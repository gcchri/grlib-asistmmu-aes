`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ev7eObfW9JYKhn9pmLArQwKwO0rX+y4AC4/ycE1JAeliJRCd2lDdEIrewhn0Ppc9
vhmlgqNgFQUTBVVxqj6W89cz9xpv/eaQ4zPkcaE/Fj76vy0g4bL8bLxczHn2NyFn
KjIUrrF+p7zRXWv3Py34eTrxPStvmOQQBX1WE/itIgsX5GwVBocAP9jUXCiT9iDT
Elu4wR4dEBceiG3YFk1ZSAOFM4OzKzHsRUMd4InKh9oHkuC7LWAHNutGu2vxFog7
k5uey7iXVHt3r4LTeiPuZRj86pRuQZm6SZRqmZk+yxL14WraIXD1SOOfcyS3kBiv
iL74SiHEYvXmX3LJ0zs3RPTFnz4TV7giXHQJPVHS/kcBELhJiyo0/sFRvSyZdjNR
710ZFzHOUsqW0uPVR+LkxaGRwWeGsw4izZDriadBN7M2825HGmsjlqR3sk1Ews36
/SpFKt+BAqXtNP2szY+0NHPbcUOH81V2FKZwE1aTXZdwOmPUUdCrs8Pq7DZHs/C7
iSbID+bQFg/p5ubQzE9Mz0z7q8JPbS9PHrYZxf1be/727efqPDJ+qcnHOqIHNWxz
MpLUyDOI4dPFHt+1ZqjpNlGGTHP4STc44BgESr92WLU=
`protect END_PROTECTED
