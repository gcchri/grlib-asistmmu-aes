`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wAn8z6eKOWhJB/manyNPIClrgAkJZPgLZXmM7VTPjO6KZN+2uqq4qNr4D7qX/Be8
N65Zj+rnwz0YKVdO/HzuuOgYrG//xT8o8OfB3gssy+EkrhOIlRWBRItyBCt3Xt13
IJMMGOdmy4Uc9irtii+fhDOjoupTMs4EqNFNWh9ZYC9rlCyGUdORjuEL/oP8eVGO
7MflL22n08L1Ll2Qs0G7Kft3bspJQvh0sROHnafgRop+KzEhdkQqf9uYRP3KjHs0
wDFA7QRwRNCnMZfqJTOJJ/9GUY/xA2STI3G+VB3ck2ds4vJ5om0g5VYm38BKB85J
G9+uofkdpQTFPzIRcDPFCYUEr6zRpvb8mNZxWCLpSSAkWJ1LkLIguMumFl/tDVyu
`protect END_PROTECTED
