`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2w80l2kmMjrJVoX4N/DHgAO5M1vuiKVcrQv1zQpuMqOAgVXBmSB62D7OvnrF5eCC
6HvYuddc+bU86FiXI/QlMruppWmIhB5O3Lu/MptVtiNcK2TyAT5H34jmfqq5C0gi
uMXZ0I1+7c3HkZuwiqvdZ089mNacwrYGxgH6ioatdis5Y0pXdX8xrLgsCSnlOp7c
gXXbN6lpkcK3N6k4ekr5PizFhaHGvZyoRwSYHRmducD3gLlzYAMCcrol5Kb3T+Nb
BOa/HaJ5KLSeNU9TNzIX7iAHHOXOryDAB6UdGJJQs4sQZCAnrp3k+6aT+jHO9Ljf
fgnyeuUz8TPaTqSBwUwi1UFZwdwivnrdq4XW8rV/5P4tsbfNCW7L5ebo3EARPi1I
zbxu38UTh/bykNYC7M+lORTBK84g+s8PufLO0mkgetSJSkv05oHvOITh2Royd1oO
`protect END_PROTECTED
