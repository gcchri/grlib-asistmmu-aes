`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V3+uhIGi/+wBLA/afNLqafLv+TCmfveWynTEatlLx4/VSZUKIF511I9n7YClghR2
9dPby9WT7rKb7kNnOjD3Qt4BS2slF8DY1tcIs7wqrPT9Q3mNoBsbCH3aN8eOyaQC
roP+i2WwxjO+gj8V8bqixOGWHJm6oXJxtpo2PhokYdy0Fh3T2+7fNTtNhMQgtQjy
OZPnSCsxXeR/zva3cPZZhG02ssPEbFJEwtBI8IyEd0PeZm5mSvB0Cf8u4O7EuU3a
5qhbYVmocieW9MYDwQWJMqTXlkWgRi8+syP0UzYoMJO7DaXiOT3liEm4SZN9JP+F
KWwPq/jnJUo2wttzzD7ciBwrRTOZqggIAoUzpE8u+DOlf4g4vJG0LVfa7OYkHBZS
zNce9B2gCK0lJ6f2fwGUcV03feF5i13+k/LsbicoRgHT8os72K4jrgJ+XuAcyZQJ
VFfK3aZp1xhMvQoYnpjHVU1gZOVggJ2vW9N0iAEnEwDmTiXosF5hUGEbAE13Txxl
0XDorA39LDF+PIHL0B9m8SuzFvip2fImRco7qDLM3XhgRSSoIjcVHq/dPgJf1YcG
mv/YhgHPWGM2m9RzmENy9B2q5VDE7meNGL8YjyTS6pVabLnzI3DTL5Q9Kuh3jL5F
zxqHihSl25YqYa9YmoF8BRDuCC/KtJja8mbM8aJFGBUmvmFclYDJM5dPER4otM9O
pLnMIVtJXNdUJTgo527Ifg==
`protect END_PROTECTED
