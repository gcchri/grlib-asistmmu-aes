`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4GgRdtKHJTeVphtzAr8mHWtYKVSG9bJD7cvCvUCgIVmjH434SpcyXGskxHEG6i3t
eMqd48RRq/7ugM/jAvDhMaZjLff7Ir9KEWTXnEqBU+Aw9RLS+ClofA8ZepxAvDMB
b3PNt+8/xMr3gMhlakGnnwvN0dwsF86zkUQcYCwZS8UC8Pw9STLPH8nedl6ZKGbU
abF7R6RJEY532Ba4+jkCEv/w40wYcBmgTuDJfM8Hd15oX0ywimlPHTUJhQDp35Ys
Fcm68eh/9LME+QibS0qBdRkQCPALyG1FF5/4a/ShUZFCDogpbnt2L3gVIRK/tXKD
`protect END_PROTECTED
