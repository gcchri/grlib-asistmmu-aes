`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rBH4NPGqHoyrguIVBXrYrquASBbKwX6wNYzlJnpFdUISKosKKtnK0WsO6PrSq1r9
ljysJWy0ijOxTPvqu1rUeRuNuA1fqed0fnPTVRHaWLP/nvXkdF6iy7YS/jp7Ruy/
awu/YyBDWAFLM29r6yW0+5+UWQLWxn9DjYo+GeYqoclEbq4+fyHWklQlVLLKCX8s
Xxjar1WbjJkTUCbzUi/2MlkECJ6TIIl1R0zVcl21aokhMxzgM8YrsePrg8ZutJix
yDyWXYcwlf4L5XtQJxwyzz+W29REacxJRjifNvb6dkLYjmdIl40DJaOax1gBOk4r
0HZYBi2dLap9Rcu+jJRFus+iRPAeb+kBkZj+8NtLTsGud+sSfL7vvBa1qNLM9Wev
SZNLt+a5vbAFZ8fBchjDmDyR0pQlzE5JNL2OBKW3f3yjZj8MfJ+SqMFR46JjvWzE
yptRZFjDZxkLjou5ncsGLn9iaXcQfHFPvBWdpZi6RQs=
`protect END_PROTECTED
