`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CVE7tSgJwrYjyxmd1FzcZk+5jnnhK3u2oqMMapDvLCroIV6kzEuZuxb2XNh7uG7N
mwPJIQVuK36U6p+MjrT6krBD+prvXE6vLBub6cssHculb29I6AW9YYTIjkCA2K/6
L2yJ0Heio/RH3KCJBL4JMhjxeLG+pFatbcPA4nZwu6q5B8kSIAAWhUhIhSStem9c
B8t6Ex3+mf9rBQRowCfM6KXC8HcrdxWDotcc07BEH75QY8ESHcdxfztLJ6wtGcXC
D8ONtMDybzPXZs9eg2zF8p4sLz+u5QL7JOv5fa/ECofFAUdj506PpPcGubjf4+ZB
zyecTcX9aAv2mUY6+lPg3Z93ydDz3H0mqd0g88P8HlGSDVHbrl6i7VCbgVD4agps
Brg8nUZg9GVB21c0ApBybSsnjjQgIihsgoTdS79hsWLRRNMlcITpRrRQwvMEWzNA
O7502LhBxJnV6pmgpm08lnjZgMCBpXMDMLr+rMhe3iaLgixw1RgUGwb52Jr4UUJp
j1YH1M7A8FqkvAiFCD05xg//f2e0+oran5O4stN2hh6VS7VCQeVdHPNAj+oVpySw
NdukwmIFtwWumnpdxbpjpvsIuACfOTbQ9mG1MTScqVd9gbhnc+NkIuvc9HVRfLBX
t2TK3jEC2yPQXHXyeCxLpniyB7PMeXYDPXiV48lSC04Q+mRuVhlJj+rQVGsqlUBL
toU8I8q0Utu3IdHShVhPd7wRkJP+cCvVVauliKRW+Bt01Kx369lgFHHzyWanzL/F
`protect END_PROTECTED
