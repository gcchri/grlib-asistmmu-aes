`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VE3aePc+fGlUX+WnWopr5C5S1jHS03Q1FaTgl/gA5pjxj33tK50Zt2LfK5Pcd3tL
rV0yDCWprmY2RFOtEzNYKlTezlEh3oeRRym4CQAckthZ6YcNoX64rGYgDb6ECdiV
VGR7lDfcQLBxzhBzsMqOt7jbJ377eQevk1XYqxDggItSQjT6sGEbkeLfBH0z6430
rCIOMIveUGX4YEIem5I1UqmQfI/Azwrd97GpeF1Jzank7fMIQn9kvQxtzySD3qOV
TxlDY+LT5jtt399h+2Oqi7R3qmX8+Camzms48VMFF68=
`protect END_PROTECTED
