`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z35Jvzh/uVE4Wfakpclx0+zXa0nh7QrseXQk27KeCs6PgNii/O/JPuz2F26ALfAA
UvE8GyWf7g7LnJan63CQGlY8sX0RnRfjRAXbcnaq645V+RdP77zrfFYRxjbDeMJ7
iUnoRWZpo1AjnipXXPlhw7yxnUQBFyNx8TZcb8sdAWj/0ZDgKW6oFKpTwmU38FPh
gVZttlkivRzhSlkvMB+LPT5ObzTeD8pVLf8vR0Db9K6Upxc0eiLXfy6n//Vpzpsg
CKDqC40dKMsXsx85yhLbjnN7muRdud7BhQwjC1L6SEM=
`protect END_PROTECTED
