`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kKQaQVzkI3SSyDYkG/LAuu1qzqsx8emR0xkUqSfPI8sYog5+PT1FeUWJwKu+k2Mv
qqJK5j+4WlZnLoPb0tXwdKcyCEnED6jIgSxtEN1ZZy3jpa6Go12mnxidd8borQrC
db9mqtFRg66LQWHnpfdFcm5n/usRKJzlr+kVLibLb4DMLdlPSux0LLVnU6R7GJak
1zkMMdfXU/1wIvhHUaF+uRKmsFceIhESofLuu+Yu0XUkJUt7uYdz3B9DAnxKLQl9
+MeQkZW8ABmbp8kvU9TO7wZgjRGbPkILelq0qw5gpoenjL/NSbNFO1g4Z/17fuhD
Xr7FwmqBWOLt/PaFo3AdrSzXOMuXMuo2uqae+EzYCNvrfyRDniRth7panyR6Uz6U
MCrKh51Fgf/zA2pY/yNmpw==
`protect END_PROTECTED
