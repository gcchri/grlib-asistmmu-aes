`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nyUzrxtbupDL86ITch4UkkhOwwaUuSr4omus/fd+8VPLoT7a/FI0uyq8aMl4oLEz
q+C7dzS/7as5gG5oXQQBglOjb1DFrxFeaBeFhehZlHI3rC/dzKPoj60M+w0NJN4Q
It/WDYuKXdUVjtcILZgnOkL91v+xsrqQ/SJ5k91IxaM+xE3LLUXMxDQX9VYyiQqa
4tRJWBJv7KU9yqtwwj9MtLZ2b0OuEpSjO7E/nkL4DLq0WdALxrKstrFau0uHt1up
S0YVhKKlIDvz2esM518HiurN6St4pUR7Tf3XIevouFPd1wcu3hwGPViGqN84sygw
J1reck/51eBB+Z/4bkk3hLcxRsnCu9qrepsSBXQlapvUPTZkbeWvo3YY3KyKrCtr
rPj9Vn9nzgyZ+QAtEPoXPUeoHaoVXOqRBjAFrLv7xIURUfKXo3vRVlLPEKTl1ROb
`protect END_PROTECTED
