`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KtBHOQ3BrnV1nCDy8LbRgPwX7GtTqp6aqF50fOFuCPuY+S5sGIoDiNpzXLh1SG5U
2bg7grzWy34j3q99a3CRI2LxpYI47PREE00B/yk54Epb8Fkf00PXWQyI2blRGf9m
L+goRCVYNNCWi467+Wz3T5IHnLILzuEJsCnU4cKXMgP5RilkzoJ+x4qnQ3s6N//w
NXHZmUo57JkdcIbpGp0rFJnskOkec+uP4Ctt89kJ/D0Kneqh4rBGjhdjUUo3d/rR
`protect END_PROTECTED
