`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O8UtqO918L/bqRbmybtLMHtAV3yJebmfoAMkOjAdhM+E2Wc8JxRUpSE49N/zP0Ho
E0lwHi8hYVuYQ7fKu3V0tWyvrflZ4KVSvt3BTYoIewIMKINt36pa60TtRiSQWS8U
qiYc0wgXSnSGMtX6u4RH+6vvAXmh+P5QYuW/dSZc8JjIl+sirFgJQ4a+fxbrav7L
JqkCcXIJsajFOLw6QDyVn7w4jHSfnRTPp9e0L1bTwUbrDtCaLPcDxu13RsBt2Y8b
WT0RnnjwijVwBJnrDq7fgT3Itr2vxl1jWdjcyJbsEorWRClbwpWI7xv9Lk8dR6Di
AxVtAfj7P8P0D4rN8EDHrVar4j6Y+FuXBnq9RhcYJEF62CvTLMUjNJZhgj8RMMqg
VzTl8cm/wgQyd+W3+lxz4ir35kI6bTI/3GeA81xq4IRNPqu+4kUyIkk0J6WI2EVx
56B/38SIt2iayV+AY8SWEolH7D2pKEaZCVphZTb9lWK7ko6jnnxdN5QEgZuq59iu
jMpnpLhKl/d691Zhg5zBApgm9PjiqQIHExs8N5WstFnK8dwg7Kszz4mzN69oI+kb
9GkOFQGC8SMxUhIDlp0HPg==
`protect END_PROTECTED
