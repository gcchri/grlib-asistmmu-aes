`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
94DE0IV553mJ1ooXWlkAvB9S/9Uan+WtX+UPf3SOGsyhnPaXK4PDX7TQvnGe8Oze
+wYAWDriEnT8If/V/mG+sUFvGZJgawXycJfudOJuXN3f22VxtY21f+59B3/9dzBj
j9WGe/2cM0WjklSeiwPVvsqEOyxEOUMFQmJi4SGBBPQHZ7QJNOrnKZAZnvQkpulq
xAF22Ph2Pl/vLR3kl/gGMUVPKvIDpIonYLCVCnpziZCr1C4xLr5A1ZQwQ19O0YMV
l8Ps6FosWRlX0y1ho5Lz9Q==
`protect END_PROTECTED
