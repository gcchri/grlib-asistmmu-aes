`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jwNmnjHmiSc5xeW2GhT2L5gnGY3hx2Ieff1W3D5Q4jUcs3QQB1tVsn7FA72fcfUM
MEwhyPSkhv6/Nk9YkoTk6rSYER+j9jcv3tT4Bt7bIRT8lgvu6Q/fjHB57z2JTUvL
OsE2WpSjr3x6XYTeusvidAx71mpjmLmluISPG6owBr/T2awe7AkIvN3U+PlYkbd0
2wiw4cYY0q9OSfiDJbqpwrza8W0rDD/1xwxQxgWGvJm5YySHd6vMLAz2agLIQ1fs
27HALW9iRzaFnLLzWjm7gcXjHUd5loC8A4IxiAN0xSkUshVM+DAupm0Hk8gyrHFK
x5Wb2TtrsNSbxCP+VxaRnMeroC7CeJqQrQNCcb4y6RMjKYfkQVsfmi7kpcHn5OmV
LYKFBz5deImD/3qP4/1Z5jOHdVBJDkVnhhZ65FV7gNW/WIVsKsC2oowZqEVts60Z
2a7JWxRu3nqAKF5HpFSSZneZBLFFZqSlWovIcrpeoeRO+mCFok5HAEtB8sOz8+JO
X6ozkm96IDqeEfEk1TXOZ9rFEZHDEdq2dSIInV5j86T+svpWWwkt/CR3ceuNp8qY
FLc5qLxcCmDKfkLW4Sz0FVe9B8qJVQkCxTII3OfEgARaCtQ+91Hr5vkoFMDKe5/G
4BMnPkDxYFyj6p3Q/brm+g==
`protect END_PROTECTED
