`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BCGEqomaiw0QObujc0zm7uj32ywJHtcxx6X07udXWm+SvE7+MuMkNqAsqLxwtjem
EKwmYeZ+WmQ55ZwoTHMzsG6B4TJsOEqJQ9OzJDnt81GGIeh/UAtEE3OSp1kbMSPN
zDB/mmDnwHo0Pk7gPu2+PuKtfeUg2RhnYaIsyyV67yif3mEEwpIE95ZM6PTlhDja
3IXpNeNLoQE9waq9bBlodJW01etK5mTsH1iFkwt6TXqBhrQlbKF4GajHYxYEfqqZ
pso790Cogl1cl4XTY04Qqm+9kyPcjcpsv+tgDL3Zx+8=
`protect END_PROTECTED
