`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
exsiTBFEgwCumvwBKtPE0NoQ5eVoaEPrj/XFGIl6sdTSeZ1ZCnqoLqhA2inviJvB
9B0NPwoHhPH1cDfMTUGCIzzwBR+d+EWpODn5AwiuQOA2SuhtfmXfBDz8cM3q6u6u
wllRWah4Jkjb80wEb7moNvmfJ9Pgkntsv9kHxU/atHU/a7cS/iTRL0bKlmlOy1FK
9ePLoGeOgisVF+fI17TNemD6IgPmUcBC5MGTe68/+8Fp69zAg8PR3Zu57SAlpBZN
zy7OsJbtkmiqxBXMvGtGdP5IcCGKedGJb7gPIUjHD5od5cdz8lhYdFqnOg9Xl3uv
sPHhRKdDfSo3o8cqzhnKEhZXrx9LHBinZlRBdHICKaKNBzqCHNaQfgwvExrLV1dv
cklo8/o5O4XX4/ET39Fk9Ezw9o2syMH9SlulCtyDJ2BQM3bSzqp0F8qP1Nt/UCiG
1ZQEbkqKf9jIiHpN5Z73/Tl2sZVfZVomXfFfJiurzeDaKbZdC71x1MuczeMQfsYB
wJUwO1w7ebKYI16S/yIRg/k1TkccLtCrun1MjYhDZuiQ9y9TDE9HR0bVklfvqxlu
n0HETlpKkDVL84I7z6SloLmavbxw3bQJ/MPUlqlHCUrkT7k3e7aI+ivrmp76/kOI
BLEIPJ0++ikrEO/U8NerWCe+esjnh29GIuWDQ86K9p9GzA2DS4SfFTaJbYVFeH06
dmBUpe1RnT4YwBZI9tdOfDNR3D1v1YTWGlZm49G4kPaiC7Bj3MdzHjcNTdariS7E
vunvxUQIvatxrFSqxygBc7V5lMdHC6FKID5JnNzseERZvWe2E4ni7I9Jb74jm2jZ
F4Up/ECx30hujAgNNW/zGMivBp4aBnSAhPJngPz7xBbZwmCYc68P0+Qkly6lZV0+
F0+u5m0buawzl9iifebWDqsWP+hVaDAhV8TkgqEm7uJxPloT60buOwoGyGvvHMx9
UaHnP/nC1uMv436aeU3//T2aYS7VAlAvCYJ6fLq9a16XK6mCzQX8/eLhi+pUdlD5
Q/Vr/bMNUgrS6yPh5PtNlti7JMR8sZ77r9LGycegIy8MHsKqQb6roYhguz+LuaEG
ncpa6ykdiATfLhn1+6ns+DLOgF+Wn5TXd5BEOH9Q81zSmqnbSetE8vddiw/lV7GY
DIp2V7tYH12d2ghCjqsTDfqIS0ZlgtdnS1ngIzdKvtJT3iot4tOnlduLyPtuL2Tf
qtp+EnEFv1w5Dm9HYIFnNg==
`protect END_PROTECTED
