`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bj8F997CKgV0l824DJjReqWobl3dlbVBSn9jShEaoMR3HRXuAzQiOSoUcUs5HAkp
vIJlkLpsya/ayUfPsqJuHx85931wOYE+UuaaP2R7aNY4VV8aSrZuJ3oDWnjZASaY
TtyrxNv0qbydUmoQXbfHgzydIYhtNQ46zTkDuWEPi56yFzHhVdFxv4KjBV05oITN
SkO3NtdOAE19Iwv9CKDlnLrcCY/bcmaVnmN5Xm1fnbdWet5iHVV5cXlQ7rcxwiN9
zlRvXKh3OKL3Htb35VIfWVSLOQNfRQPhp5cI9IcQh8nHMaBIRcmlahRp8zPGg0mc
gl0HGZOastWfkE2i/BmEKvz71C1L8UYK1z51n4U4ETrmqvFgPJeYEzLndD9ZIKJU
rnsdl4qgilWhTx+W5BXiHkZT4Zptdn6064bGUmXuJwyXSlnT77mNoPA9aeheUedG
NY4kTx4V23b+z665llrYfeTLq5Rx/oJAFAD46ntnQIw=
`protect END_PROTECTED
