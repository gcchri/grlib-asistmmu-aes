`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
plWOAKvzS6F8Og2XoozlOsaB8dMEQ2yS32PE8JsCRMhR2lkPwlsn+mp4Nv+TWtsG
ts1Kr2sF0Kk5CWhIWuXIv0iyqIFzfqxZiS0knXaWNToCa+M7A/iGmreX1LI3Xg23
OVTf67PZSMHy/qPKQUentx9KudHIX/P3dXyJ1GOQsEzHIdr/eBS8G9KZJ1aUY1AB
Lb5itQPSTxVsFq3cS4Tj3Ntmhvnw7+Zr8qyIpJOkxPoVU856DiXURuBt5Yzjt4WR
NwmQRM+l0j+5yS8XmpYXXQZdyhNvbS9EyjGoPv6c8TJ/57YKmz4vPFgR5T+zUFcy
bAh0VMTAHxVf65aZMTH7wBYtBrALhVBiBQ8CYgjCZH8eCrWGeOIrSF4vWVF0w1RC
O1zE3Zj/Wq80Qi/y40vphdMuGJLMfllcYMQ0rRHBi2IO8EdLQHdzKRjo5476RkgZ
`protect END_PROTECTED
