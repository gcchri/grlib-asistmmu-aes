`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AuhjF8LOSOmauR1QV3nPjYTr+7EvCJDceoex5Y2E/q2rMsjV1dhSOqAccs2utMNG
i+zbz9GRM/S8aQmJJaPRt71TlgwtSPWYxnXULXfqn1ukViu+x/HJqntc2Ti8t0TJ
ZeHY0Zf9LSCjkZ7Bvs/qpMPdMMtR5+KTcsqgx2GAiWZBRYNjHlTf19AdClgMtM8d
pnz+AJCIJaABfs+/ifyD1xFIw1WspPBWx8iupiWbdQGtT7fOn/d7v3KcMoTMR3nz
gM1uSaQ9mK9ni3Duf8u/Rmc1LZcJgrul4zNQ8mpuFp941hFyLVyzaJmIly5ogyCi
2E6K8GqCZV4ZQAKTR5Tx8ghWqLIiUfwBrZsuDRUSAg/5iTJIfOLIAcmqGmTi1/a7
rrMc+5gezPv1wdkOsbNsWppZ9z1cmozUlWJrVqlQv05tNrbzTKk/8wxMMJrfRko5
Je1xn5ltspPWIIwbktmu8LGOOGKc5ULSy7pBQ8M53sfDVgfSbfsHDekPS2wuBVhP
W0k0YtfR4N86eB6mFShV3ACqAokWkxCsbIFSyDu6bH3aOkMTHDaArnUmtXZIICeV
CnXuQ8xWuFvmgYGsJ4U+GUFfrz5Qy779/j4uTkxcpvOj3e3VdF6ptpyevyCS567d
yaWK3KJZnE6LOjeveCiT95KFvtTGYvpUgl0jaN/u1aeu85tdV1svtwrso9+fc4un
EFDJ2IlI06ITTOoW8yCzxzPzojDrdtBJdnRaJyBiavQHuLDMJwfm9N4Ps07fU5UE
PAyRX6rsgSHdsyPZD3YQ8OFsFJsKsdlhiP/O1qagEQcRlYYbbZnttBZhurkwK2qe
5yO6GPPXz8/JY4iCrxfncBV18b+7VYuQzFjdf4sQQ93LH6e/olnNO/JL9WWMPES4
wY9XzB6kjpgPKJWbttzkdjqDD2ZvH2LwcusGkkKFriN95z3yvI9yqynFbuodt9MW
`protect END_PROTECTED
