`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5uKnn2br5Vuiawiywr5TgvFduHLKVUj8qR9eMxDDvHknrI1WlV6L+W8DuljZFQfd
AVMHAWvBnxYJGtIGlolDHYMIB8vJsW1T8UGccfLIVdIdqjY9g4CbphwDewryJ+a+
mtvm+Yk00UbdMrZqrivoMC2mzihT0KwiLvYKCBZaEPujGH7inzxQ3fjep1edn3n7
JUANwH2wJu1CKrGHHx+Q/xyTVJ2J/Kcxcj8Nr/SFkD4BKjPh/crN+opDJ890CQ3q
weNx47AW07jHYL3LmZcwMuAieJPoc5tTaj57N5GZtFa5GZ03lmrhLbToYbfZvV9J
Hd9FVZuLS+EaIASB0PDMuOMemeV12PbzObwS/rJ2PEjMXKFYP1v8K+/ppjbBxAps
/yZZ0qDuvk1aKHjXPNrb76AR+jQG3bozOscSsNdkXAeuxHYjINPejSHL9B/Ton1Y
e5gbGey8MwHO1hbf5ESrEz53+YJXaL5a9opmsFQpcP5WuZEglgtV9X6INUAN62Un
HDxQhLd2wbGg6+I1km5/dsqdvpsNxp5+ow2wSW6Yi/Z1n3SejQl2X1DkzRQbwnfL
0IpvS/3EGzEDl4BMM4oCEkHkZdZCM6g12Sn45dtWFWHURt+fkcdaXeVUGASuzT5C
p1a+7JSF2E+h60Dfdqho3tJODfDGXZBqzGaV8Pr0lJU6ZBhGFiw1VYzmfjCzV7xT
7NiI0U+VbDsNiMQ9XjFQFq0F3pWQm0XSci/iH+TrSOD4jJXzAJSTHU/cjJ6/8eBv
pY3W02DIwI+DUSnT3/dgUiOa9/UUQUNup/i6J6vFOIfw0Iv2sDVorr/htmmlsMtX
bYdhnMv2qGUEAE1FE2POx5sKcqYImNfOEz92I/YZJOBO1rDYCfMwRtfjzuLQX/7o
OosrF9nwwKxYUdPPdVOHDT2y4PcS0bpQUYnlbG6IGfo=
`protect END_PROTECTED
