`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TU1Zcgf7BwP5jKEACUtTs/Fp3UzK6KRxJ97KNZdaUMZ45HCqXVdzwdQpOWq5DLan
umY/ECWnFVDWCifM02jTa5aOkMfd/V2FpDcVlCPG2ccehW4IZ0QMM3bR3p4tFKIa
6lIG7cQV5dCIjF/2/26eqJhtrMf/3MiX6oJEx7pF/CK/62Q26C3PBWAxb578osCp
6CrnhapkqFljnutOZZAAKN7dKCszjTUI66JQ7+cDjfpUk+Q4VGbslb4K+b5cIKF1
l1OKi6wLWQxzre1/kR2AcGuUq8LK9AIrv6wrzf1SLjw=
`protect END_PROTECTED
