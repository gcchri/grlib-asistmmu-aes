`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qNkHtYuf7vQEPLKrR0d4f882VchWrf3Nl8I2DYgEafy4HSPLApqzqOJ9Y7K1bCBF
jvwMcGqcaC2U6g+pOU/LtdsBhGJYZOewx3z2aU4nF2Q3PAvwJ9jgN9rmkOHiNB4Y
+XjPvTwqRDqZYNaNBuGAw1/5kfph5zs8uyLDrJ2Lvn7dMO5xiemcya7fTu9s/xKu
44Zm8FQGeNUZUZLeGxGHlnRNL0TiUx3dQf3FfVMg8045uHqamnnl3jJQd6oQLu3q
4z0HTW6UA8tidAVMk6KI9+HQcFU/ypGQXSM5tt4OTauZKY40vUJXOLLP3PEXg6Mm
SG7SXsAiTE6/l+mJKxW9OuE8tHCg8sBAmM4vgS/FmDX3chkshMJDvzAdKgZrbh6c
UE3dsI5sCSUG1yo7VQfQeMMb5BdY+/w7qvGtkX4EELDUBvJSrnKkwbU48SQVVavN
B4tonhdJkIoP7Xlpz7h6++bqIL+I2XnK0Q87nBSdthrQzVOm5BKK2KvtasVrmoH+
tUE7BXrUax3XUZIEv8P++1523fhL/S+RkTcv+3Y3e+A=
`protect END_PROTECTED
