`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vMPdbKCe7LIbEf6a6qekl6EJ6pAfJsoFvzM7vBLDfbrGnykXVDXUwZ0UEZXSA3HU
VGpClvj5h8HYcLvJB9a0nfwDBvstLkADw/rSyI0XFw5WQVn1kpJbSZf00NcAK2hS
VrsUkfjpBhwgBfgczG1IdZbMAmr0Kfk38Xpeo0P3DpfXnmDeMzsGHJ/gGz0eznIW
HwT39e04kkWJ27ygghrB3yKGc1gsxqMpdzc7IV0TUyJt3ptE3bCCfM7HeettHWfj
unCBAGfM2osjCwz5pRHSceSlP2AkGJMmr26TKvRt+P/lxj5RPknYAulqEJ/j0Rsp
Vth3LaCUiZeY6r6FuSvvkiPhRq52S1cySj65uRWzJ3iXAxL3Ojw4oY8MEopMfHHQ
erzQIeZaDPwAYmVBijMS2uOLcmEiWzJ2WS7c7POECCgfWh9zY5YeqkEqLja/K4q5
sWCV+tjh/hq2KvTrtnYcqmLufOM9TPEoeRXdIHGIYYVHKTzhJY7nzFMJZabAUfu+
q8qT2KUsZv9T3cT4FwhPGeKpnqisFkmB89f5y2CM7LRzAwre5akWznXGERX0esiR
yC34k+5ACh80j3AZ9cci9VKGtWoJsCgykkktdvk2r2CfeTAh52Qi36Mks3t+iY2S
Z1HqDxRAajlcpg2+tG/rEA==
`protect END_PROTECTED
