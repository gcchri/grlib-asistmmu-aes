`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EkdkVSaqSz58bw1pcmOJ/5R3qmhcrNeZW+PXP4XVJbIzs/OT6Q7LFRK0YgKRFyKM
uV+R3X2qF+8LZ1n4htvJh+38t+4HSZmyqHNAyljj5Q3zIhsXGRfwXlAJInlhgExe
lH9+TIFM4R5IWbwkw1zfmkAsiR9jATcAoUIjcoYsSEqRsgfazrpUUQn1sVFztilw
jCjGat+SFyBFSuE2FpDx3pOXJ2Uo3rOqo+zw91efoxs5V0xYGrm2uEvn0uX8VE73
a5YvfhwM9oDqJALrqBq+qjsAV1h7oG7iDpAy8mClItE5lb7Irr1yfhtyP5Fp6DDk
RykrkiKUvOmCc/tv3wLo/V/GvauUZ4olIIwfu0PEdV5AXuqA1qRO5Zsbm0hMeD0m
GcwELSjvSqdLUKXtb+Y9gjucTQgnjG9xp4mNtFzTB+NHVh7Dqw6BZTHw8bAyVzfo
Q1UmErljdlikl0m+hwE7T7K2uUqJ8gesY7rksMKOYjXW7HKVvjTHyRA8ZX7B7Elf
Z7xu++1qu1jLZ+LrVXdotiJPyXC5Ugn+CyxPA19uu07j885zf4Q/+GmnY0s0FLiN
UL7m4KCacxsxduG5ahmejwq4jhWs/CV9h/uU7buUAOhmzAghrAaC8o7E4vfQ77Xv
hIYvk6xIlz0iLg1zI2z6TewPO/3C5DvADO+toiwCzX3qgW5lwwAP14SSaZQDZ5kB
Rykw4V64TCUO6R+bXuv8ou/dmlLQ+QnbzkqXAK2AZqI2y0TxR2Txsnw4Tdeo4Et9
08qKVstfNCnFlE2/jtcHYSKlnX4gaee7MNRLSk/wB4w2WE0FVTpvhCg+3iA0fRbf
kXMAiT0h83a9BLx3OnV0MA==
`protect END_PROTECTED
