`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/u+xf9spdw3EUNU572p+wCX+Q63uyLeLc1P7G80zQMz4W59udz/4LflZVQvhxmdA
qQGEbwRIqVqpcgqIO0bCOqN0FVNiJjnpikuaFPPlR38+6UBEx63RiMlKqe9NlrXA
MO0SyO96ZEthUDV/1GMztOEh8QLERD5Kcu44WJrkMSrpRAfxhVVSRDKtahk24+fn
RK5BmT7G1ifmox5KFUWYKz7RneVPaq8qcKOYGn9+QQe9W0yXlwMUZ+yrO9uaztx0
hF2x4yWavEFBLIlaADap8r33UgnHqpE3ob8jvFxoqAX+LOvd6C0Qw5ozDLyuHo3I
2fvZHYytWuVRQMFNj1xv1zs+esB88DOchgV3PZwdheWdpHxsfVfPGzsaV46SQzop
TB/FTFsCu7P+K8d3VtnM5Lj+jMw37Gp9l5dSW60il3XNdHqrw9u/Z8YULYD4ETS2
IDHLQw7OT03AXibXqyikH22EX6/70n2mkQP7yf0S3x23IkBa6B1dWTqvzMVkKcjy
pstg+4y+C7Z5pv77x2pkCOiztesak5kc0HS5Xx3XsJt7nwXi+jmjByonDw+oSmeh
KHUI5noHWeS2QyHKj0CFwuzauPWOAq3o4myjAc2IZw9PyMcZ7tNXrBMjbq+vqksX
2/e8pfLO8c4xI56jlCxXRhCXTZxg/UKSkhbN2febi2B1aLGMuAwj6G1Vd6WkoW+e
pGwHtLVkxPo/fvTtjltZy2oDMBpyUrKJuGFuTOp8IV0Bwv+nvlDcnEWTP2GBu5st
DSpVibjflh61+feGDSnmRxxNBSgQ5KdoikQPmdv0nSB1YdGbY3mPStm9RfBMFChQ
zpA1mZZmJHzMMM0HDmCmQ62h8rNFSV8DiF4Y4To/r9oiafTBs5KMXgHMwFoXUN1C
/a4q6Kd1H9LM7szNNCD3BxJLxEBpuNs3mx9eXUjyOmfuPy8hKj6/lfIheONsGD5F
ty9PfLFQTB4WBEZAjKV5u9cOdPFdpO0fo2SyTmaYlaByt6bDPkfCSE1eLo1FVFj1
kGyuaM9KOzY14m8EC6doHIt6symnzMiuV1acxhTjqsc=
`protect END_PROTECTED
