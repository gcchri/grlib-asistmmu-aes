`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mwnw1f8zjENkcWnaD3Mn5A3UNcooRqNjSSzVmDikDkH564TT8iN37JkLt9ewvlmv
Abq8I2Ksx2Ox2HWjCuyoU+GVXixkH97ths410reh5nd3yHP4CsmFQp3Fxjb4jVoC
NU0xeDj4+BXuyWtZjFdp6tHAll5YDdNuFMHEUN3/zZH6ZWhm5MC17RPYDl1SmM5c
itrCJSX0bdubrn2/2K4qmRdLiZ8LVamRg/qXZOK2zQ9HMCZTob9B+iAB33MZy1eD
JqR0VdHPY11k00hOU/e1IdM+Z5Hd57b3UXz/YH5n8CVTahQ+W0wyR8WmMtT89xpX
+Reyrj2WnI3JTgYuekZ6JDSbxIbEeLdOEc4b856wnInwa7bMcvqBXsiSMx8MUGVC
dXwNIFFw5lWzTXxIisTLrqW4Ix5wpbZg0OWZXTkVfAcEjw+RWhEB80dGjEz13hsx
luvdv/ArVjkTyg2SYK2DXV+MnhbIJTE7yChPhMPUtdFHFoXgqkLYqNBre8TNDWR2
87ssLjnOjukNdqQYJkTW7g==
`protect END_PROTECTED
