`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lyrYlvS+Xe5AJaDBtrPYMz6RCIm3JDde3GvMNvh5THx9BM7DKnqbbFKn2nFiiOE1
nld3/Fh2mnxEpO4BsMwYc9qS1ws58rGWnP0VepbAZJTt1H4ykW2rHoaKDZV4N42R
qrSAq9GT8Z5UPxmFJmAlc2hDd7i+ofu7O8cYOBcFFL5+QDCIDuo3GSLhVHnwIyRc
1m/DzOqTmdm8s63COJX7fKUbrJMvMWD2UViqJWBvr9qBY2ZiVeA5cZzb3jl8Yi6e
V4iN3Hsd7f6Z7W3YDEu0UQ==
`protect END_PROTECTED
