`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FoeWOuL70i0IoHbT+/UkEYoNy+8XQNKF6n5uv+8ZAWDHSNcwCvsQlIdFSR/klARY
5XnOnri78YUHLOABKQ1kpK85b6GLh5Eks+TNZj6tKZZNF496rmil/rLRO2+xbhYH
lpW/btEN0A0HL5Y79wvmyPjJ/LJgHCXXUG0vrH9z3QqKYiu4u3jPu/UkXAyzntIQ
91mvdJ1jRy+8r/44Cjt44qRe+UM5ZkBd12CejSncsr0gTfRg3QWVbUKuE2+EkiHu
BX+o+VlCPgPS3D2hMANpS/k7+kz/VyNPgoEU53R2MFe0m2bIH71puNFZRZjYSAOZ
4FRGiE5IVK3TP82hJ3bLHXM1lTxqgSyQXzRd986U8q0tABwQwEiWbjz+mUUL5LY6
pqcn97D+uR0T0GCUC6UFx/VlvWEna7akOx6qs1CDThFLt+67jQJAwy72DEsYjI2N
AJWSx+LKD7hU08rMw2TBorZlITufcS2Vmui7vj/RGB+nJ2on4E/x+a/oDV7Up/IU
Ad8j9fQUgKt7SoKMATPeB4XiCi38Nh10rFfp8J1ydEnN0bJe9+BdJJ26xFzXCAtF
6Y+EKGzwuekX+H7dAQfqChLogf6kmWrapNRuCGtwIFvOGgrjLBuuEp5Qk/ZMD+Xv
J7007ImqWtWFXu/qJzD2vtVVNN4YOD4yiFD9GtYJ+LvDAvH36l1P57A69HW/vM46
aPd54CBuzlipAXsl6VZl5WBPjyHHhU8hEo3d7i1J71rNvZ71YFtV5VvzVs/4RyQz
4/SD9+Cskk9KznTqM8DNB+KRg36LPa+BMc2DT9k+FlwB0seYRfR7wfZg2PIqJqRX
dVe5N+LRHNZ11lfZT6RVXzS1iKwwYLMo5iBFFVFq860tBTWifs5dipD/AI5G0Bef
SkPO9t8MPLs3UBsC5TsazFxzt+zMSGJksUk8UHFhh2Kxbr2BQr9QTcAE7xHz7inN
VVZ3FXoUs8UzITf1zLhNhXwcsPG7ZUHct8mdrhLdxtZm2kTiE8b56ku8IZmCCsNb
6HIGhJDJZqE++gkcYs4/7pTbMhcxbEXPZxL9Oz0wJ6saKRZpIRv3y4mqeZMH7jj/
jHgB8h3fQ5Jv2DWvYk8zr7+Y5sWnTPOcTyiFDPYVeM6w/08mAeMyEu9WCY96Rm1r
WqzWqC37t7mch80wt0ZyMs7TSp4kW8slpufIGUSaqNF7U3gdiPiKvrM5qCtaancQ
YhiksgkGAoEeg02cJuErTxDvOuqqxZM1djYFb3CVK6znaDzDtXAUynwI17hUm38d
Mfw3TNLlOhKhlQhNkprslBS0ZYCa00WOpb4IBHqn1HvQ9YZ7gomGFnCrWGSj4gvf
FL1lVQHTpXbKukFZK1asVRDJYVTLCSlOiZrA5FmPr6qzx3KWH3p1eVrB5LGmbhv/
MskHEnpO3nQCHGA6Z+ObYtjn+t8s/Xq3Om2dPTlDmH7Bw1Uc7w8+CKhN6rXir8eI
oAk4+i759bls/s2LPSJ7KOKv9OeQgjYIUv5fbHWwXVRchKTU4XCu9a2m3+KGVTPf
fL8GJOJ1xIE0xOY8BOOO/lih/zstjW8KH2uK50hicMvX7N++emUc7Q00Ic781poJ
wh+jjL8gfOBiA3xnGBJXyxFuPxvp4SNcTpLJJFMsCQLQRm/YwjrJ7q0Isk/+WRzd
dJpoBGCZTYO7HxrhK2eSU6U0My3zT9ud/drPbpxiZdQls4XrR9u4BcL0LbIrusyX
Oxaav9sFcCBDm6YkyfG6h2jiaamqjaDLd85/UVKH4flNrdSJ5H0cfzZZr22cgbjm
ZPpp/+ZHPXGS3cShvoVwgvm8MqAKy2oHUqeIkFPU61wSt8yrpv9nCuazzGr0JwFE
43JTLRNb7dCHzdN9dQgvZrUFKAQXyCr5pCvPN02BsB+WdVhy/aPR6vmGpACFMNSb
NHskcAhiyTpS2uBzVfx71u92E2c7OkT01vaxPl9csL6yFa9RdjcRNZOMorlJdR24
S8YhymmN/3JlxN06scPqAKJAXpwe2lUbGRCiYRpZxnbnvGeAcHbWlrQXuTRm2rzS
dAhFBxEvSVoVEAkznH3lIYLIxi+HYz+B5FuKGrZJbbQhFoTekBxGc3yKASDP/pI5
Xp0WDDs7KeQcb8MrCQqkw1DocIlhQFhY/mHXJM5+nCwCGLqUeROFI6eBEaR7TaYu
ACpe7kbKBpOKMHxGmv1RULvq5NX/9OfUo5lRisWpOZG/tFl3GpNXERtfoDl+Kp33
RV88ICkhxVmIUB5exaTDBgpJRjIIJuWWySaE4mT5XfJTyhkREXdQm5cXF1Qrf8Uh
YNBYaERGVTk+HNYFUE2vwyNFAy4mhF8U8TXDZ7mDmx0zKfWz5V7lhm8kGs82iAJb
YYtm5se6R17tNg0kxbwU7jCf5zGjXgiM3GXv2zLhvZu4zf2qY6be4jUolulkW2qQ
57Hi99gVNJzM3SDTQgL22zPzKHPS62Ds5+V9xCmIMFLoiyDq0Bf9aaL6bsSpfzZN
A8wyHoLa8MS8mFow65LMMLH/JvYFMzI91ZdbA6bERnFKwpYaM3At/K94CdBBux3J
7AzrbErcpRnn9JUNPNXEV1lrylqE0zDK5ELFHwTZTHvsY89V9n2p4fRYD3BKI6fO
vHTvPqR8HD/cDeiPqK1IbkOpY3D1w8EIVefXmmZpxw2/mqEImPP/Jo6f5x9X28ks
y6U6laLRdUTcyVfz0X0TNAMI3mEdIcT/xnV3BNpr1OkYMa3Dg21QxYLzsmq+U/qF
KjowxuQgg3/MwOxY2Bl4N7k8VqnwEWYZ4tembOCGW5CxKMMAlpu5qq3iwV3qI7QU
Xj2tOc05iRGhBHv04MEW5zmYDMgQdfFf5u8YZwKoeYRHCIM4QZZqFiTlxDLbEsMY
T9kOVIlEcmUxGmzXHU97ccF6GdcrUXTmBJ0fpuW1/kLYa2EVfNYaPsSq/SF7gPEa
H3I7QnypKEnr98YR/lo+VtMgVMcRxiJRCElBxjyGHwAVjdyf1T4wjqEcoKti0JPp
0ZyTaOOmeufAxbbNNFnE5wfIJK3+ncW4vhIggfZ+eqjFilac9A0KxySYO6t1mnXX
T1MhsvcC0hk8QlE/cNuuvMj8vWS+fGqI3VrHFPAvsWM5uqBGMkM2hpaJeWIavWlt
4iDR7xRrWOTR9THsVbn9KppXBU9iXWpMgD2+RRtd9KYzGfIxoBlQSf1QIGewgWgE
NO5E8PgjYFhk0K6l0Oqq2vZ4T006h39SE4LN0O2YmlTQyjsbqwLO9mMHzUx6w9f2
0lwK1xRKRN+s/heIVEgWcwuDksA5Ape+i8p6X7LNiXEN0xXywIO+Uixv8A07U+oG
9Bzv/S1JyWXUPKq6j6ldZPjW7FiZx/lPghgpQwnXZDJP4JxTMJhcGyA+r645dSn/
914Z46pJ5eYXBiAGg16iwaDj2mF+g/R1ceevGQWaEh1VaGuNHXcz2cgdc7lmpXY5
i5oREcek9aiHmd5Bp16uShSLNjoMueZR300SdQ3qZMcaFCG2VA6KQ7x9PA5UBds7
CwDcxz5d3k8LHrVs2g3QHMIdRqOuVEVGeUD+Jhl0mi/lHn513v9kecB/JgSSrxPZ
DcWwhdQeZ8CSaRsiytKd5xt1iHMpzEcs4qWnIRcaJnuTzfQyzNgJx+TpfErHjd4p
Whg8vBSAU5DkgMaXICoSclvMUkLRA+X7/mCNv+6Imvmh3VzZ0GC1EhE9qyOB4t3e
6sQUXXA3tW1kHYFUlOqa+iViovakgT6U6RPL2VXSv3y2Uz5/hPchkqrtkdxAPXcQ
dh84kJWI5s/duVCDSQByHZjq26n00cDO/0Xgt4PNEM+A8+lhq6gZ/VHZ4Ix4Q19e
tIfjKk4/b5dBfY02HLd1SC1PVjxY84q8EtG9vS8XVhMHrz3oQJjUUMUWbURAEWy8
jJ7ylIA6wqMqc7xcC4lh5rNgKWFQlRZxXYm18/tWycmFUdps5+Jpo680esF1OAeB
77qzMPM6HJuVzotc9yYtaz1h4mVcu5JruKaas6u5PTC0f4fvYlJpsarVM04yUssk
k4Ogk6Lsgn5HTa5zpqkrFQAbqK0kaxHxrzTPEI6Q6meyUzcC7A76ZBG+sWO/6eQJ
SQ9hlr0oNbJd3nQcWSNXwUd1koVbH+m+EIv1lEtby83Zr7ULatL8tOruVc7HYjQy
Zpn3X2F2HNR1pjM6ZPJUvxtHg2eRDgDSOFFhXdiWYmaXtu+sL0vMtR7sZgJ0thAc
1U33eWWNhuMnb22GRQ2dUWGyPlZ2FzDkdgFXXsSh5yO6jq4zk/6fYVpaeATLnc+A
ZbQa8dcEl5dKQA1XAJwwgaZgPz9XXpykoLkseEGADAo9w8Mrfs8IZJAd56KvE78T
jFMZ9LpBFoyMehN3Q8N1dl+iR9+jPN0lSbxlkj1425+sZbPxF+koHgPaN6gSGj/B
RnFx0O2cwZ2KQJD2bAgmkWO8jLfP63Pd2QouCvFGBo8bu3N+1frfpTi5dXIArUXm
/tSUzvuBNb6cNlhaLzQRXpnimWP4ex4vYSrpIMovbWF1xipt48jHS+jxnW5VQ8X5
EB3crmv5++qlEDZ+hCfRrptct6Kk2PIet5otHIl8icTZ+utSL/B17b3LuEqd/vdX
ZNsIrZoCzyJU1xdO12OAbazMLj7mZRsA6d+xoluvQbVTlM6Fl61Xx/WbEoxzQmUC
KP8Y0RO1EChbUUoQpiij7nV0Kza+vKFNwLNu/2WYeUWd3s4/LeiDy8ynwnV+SHSe
YdiduUXLA7D3D90+9z8uI0+TB6N4RMWBck0sVQvfujNGCHLpK5kRbWJ9n+BIy4IM
XQ9MfcTMm4iKuFl9ipH2rJenHsZiKJmZCDphm+p/sINyfI3LGAr1p3P6z2lkxpBU
sNzC35kSj5HpCebeD33BPUoFGOQvJZ0Xq5nqwwf0IyhW9/u1qDZ8XMfUa9WLUG9S
U42K9d5XBHZIb3RLkn2+02h+vBqQV3t4qPzjHfc6OKfbb0zVyVObIiUYXlGZkAjV
W2KGeCnhdTPQ89DpqiVf/OcH/lDuLqoQyjUQvURydzBVJZGnucBB74EnTJ7x15d3
8SpJA19bDJ6kq/J56kwDt0Hf9xB0rcUN1I9cVUaSqUb8Ll9AZciqXbFgFdFGqEZ5
L8RKFvUIk79ZsgJyVR85EAFXIaw9AkOvgjv8nHgXHT7X8e4L1MNHuNow7riz7+GB
3yzdiPzEpSsgH9dWR79D+BlJhYkbxZ9ZaXvJcQGFs/rM/ERMBiUQAzPPPGhzOglF
GA34jE2fCUgWho6jnVVfmc+pL3+vOGKvRS2b0sir0iOSbQ1jiGBMjh8SCiNNFanm
iVEiJacjoRamyQAfs1pbU4h8fA2Q24dWPCXbSf6nMNKyTd0Jg3oplQLLN2KSqg2i
6EPwkv2orU4ylWFyHimq5fAPv2+LIqB2rpYISu0RhVV5cqC/P6Jju+ictcuGa+8c
0mLGuStR+0qOBYec6lsRls5aZMFbZJfBxwNko4zn+kwJ03oFdP8+tudGnRXsHUQ8
ATEXg3pOb62MF8hqmfgHt/Cr5vJoM0l9rf8vrxiriIsgoUtCDPh2Gn0idMA8VJyp
s2YdZaDr050hCh441eDDvnINUuq00qEq5ixc9XXgl4crYL/V7tZ7SPqqI/Jc2YTV
z32q1pIUZCZLSMnkjtz5ivsswdT7RFnqTQfnPdlafTL5idTkqlaIE7cAkrWyaI/l
zRV9CJlep6x3DMNdHLouzREhcmENzYV8SbclY9hPer1CSLxa921+ELZm4pnGN821
V8w+wZOmtNB+3vbCyb+0JaKJ+vkS68GNYVu+FKI2UZ72VHO4Wap6Mdoo90oKFTCe
QhfUj/B8jDaF2XRFEb2OT3nL1MFpTvb2kHz2pCiYIsx/X3GmaeF9oprO5GGEZ6Js
m4Pqs5JP/kzKCfytTUN8hGmqn0tseO5HxxFSdqsHhu0D0Abz2iGTFP4InPj5HLYI
OnlmO1iey81VEk/hlnN7vF1sLdRbfQ1GhsPiISwvQEjJ0ZClI+uNjWtZVmvB0VSV
2xLJTUnknutTLYYsJG+nWyjNzcFTrW2p6NVdluvbntVGckVT4RgXjgyymUimPBDH
EnJCWFEbU7mVLtYA8eBw3PamXxtYErx5RAjy/HquMOkr73SMS/TblF5PnsJWcdj8
zSilJ7b8RROtuvKe0+B8I1WDnvrsFBQESFT710+KfXCnniFZ9Zons3WPCmzmkLjO
wQz72RV/Vqg+dmS8g3NuJSZqf4ATHErcMsSLKNnb2UWIpRGfk5MXc1QxAMx1h7HJ
1Pv4kZf6BrDZXojt/afqg0YQQ6+v1yQ0a+Iif7GHXzUcaTu11njKR4pEDZk1jPBE
Hrpe67IuzspO1O9YJBVEr+1D7up9ZPqXxEUX2TDWUWfFda8h4Ugoz9owxPR2n1mc
jAe1gB7t7pNQGJpNjNlb4QbIP2jN953G573oVwifjaYS/hLLwkeg3bNZ9FeBCc8v
NHIcZYINl9MEbmNwyBMsG0i6M6CUUnYjzNn1+h+OWcRbGpSqrZMHt9NVKfiTpJjW
eiV1QsB3BYv4aAhezF8kwb9wAzsdh8D/+MqLWrR1iA6MN9FQVWahH4xbJ/uaVJT7
lL/wxaOyw+ogfaymt7ZcxniLH/oDeJRBp622pvz2TaOriGM7PtwMhuCcsVgiIGVe
rMToFQOCdPs5WayLbXAn0e0Sy7p1n9P+/LmH0+Tm+mEoy4TOCze0txAuXYQz86+i
DIVLRskUMhmOPSr21uKpPDGZxt7Bg4GPIqOKOgKxcSh6ESk8NJgOnXDtBVVnTr+u
o6b7AXsltNxdBqY9o43EIbpVk9CO2Ryt68SaXQ4X+q64QnNDOODTQG8tGIiG0fHW
pJG27TaHa/OtTAyYs2KwoBp/W2fuRdAa6b/8L7zNkwtWdCdiuhiYxo6X2UMwP0da
2PNPL4yO+HdtYljWpBWLJFg6JYVbAftZ/lhFhB84caL60uKjPfexpkc2LMr2bOeX
c8LiGWW6W3k47UDCXGqR6hqXVKCq+DbZB97tf+XovHeCUJo1Ds4mx+CbAklZ0omQ
9IH5qI7eAcbsZpDuVbBmNmodi28J6MjjhGH1veKy0r0vEeL5R3OLAwX/gCNXPKQm
atKnkjL5rmMLErcCb4x4+xsIjIEHj9wjjryu9Zivx2jszVi52wKDRxfCG6Uf/qVY
Jz6cBAPW2IEpN7l8/hJk3Qxl/0BzoEephbbjNerjexTcPEqOIju2nnwL+jp2yP5x
663IMRsKhbQzbVcvvwZ+RKQJ1F9MML4F1OBgl7Wf9A0TGjmPv/BlHP1ITXhH65WR
tvP3nW3ldL09RZHu5j6GFtibTbT01FSR+9YXKojz2zBtPmFkp6CtiwZ2vshPF+g1
qN66kzfzDxTOFxX1yPyNabNiAm8/ooIEtl7tLeK1pr8U8MXtnZL3uc2NgeqExXih
qOc5mkM5uAJYwysa7SBvCrVh+yDzp4rKQAhkZNuLOtilmQ5NmK91B5UdwzuNxxDR
fHq4fme2gO18QYOAs5jMMwD2scXl2JzJpobFuKQSISLjpZ5KA9Kml5P2UD4GYLN+
G4X53WvyctOhC37eipL5mqTmGluI5gQkOUZPqPuUbP/CN8iiDSxyOh0dc4/8JW1A
F5fFRRHuoRV965icfHEbxV+kwwZE7cwGwQIf4+Z0/FA10M7pUqvI5rUK3u+1gLka
uFnvvoWmG4Eh8qxeHnwmUVfZeSqUAao/E/f/nY9VSoX0tghuyyWXS9zxBBRv1WNQ
3thp/2/1qaIAST5jNKlJl0HyN9CgOqzu8jhgvV+O+dIr4ez/ZIeYdJgnOcTU/HJg
HS0IQTKlBuxZIuvy7o0fZ3CEZFoKhmkYyjJVpNJ6mSEyHafPCJ26EoXowxqogMZc
QkMu0Fc8HvysBFRi578TQU/h95cb4RfiRSBqJsYpL/o8XFArf/JLVY93adwuR2H9
A5EqDtJKTKzP8ClWnuk+1bghKK123qNXLM/8k9wiSID/jaCFyLjO72fzA6WrhNAr
IluiQSA7vi1EviTLGyNx3dqhuxM/0tJdxbl8AF2oGRlrIC5h7BefpJ3HoYP+Ejjz
4qOEdm8XuKsGZVpT0DcrA0nxQDjYUUWQ/OdaHjq69US8hB0db0fV1wiT8/ZVh5I6
dWKE+lRweB2YLpbEc0OcsYFEva4zy1WfnvQJ4rqYEfn1n0f3DqiBwD1QKbCUC6RM
YSk0yygCKgPAbMMQrYNJGtTrs65LfcBAs3rl4drYMrK0W0KU+Zd8WxjxiTR5R1N3
oU7eW+HRme6z+B4/w38dGevPoMBGybS41lDYJpw4981ovXOvoWg6VVYSXWOOeu/Z
QQVTHRuuqU8cuqlPFPzBAR75x9sip+LGTuCsHdrRubMNjDGAM8B0g3li/7O2ydIn
jI5xUc6IZXe/lcBKFaPq+kF8P8aZCrnrm/d7HQFxnEICB07e0GzqOi5xULiHXv5R
SsXBxjHsUkw4LLGtxo2wo8oINwnnVNFT8Zn3Ny3mfZOPWm2TdUIENwO4wYeJip8v
M+T2wAUFgERvzwJIH0qozMAYQyxHx3cgfaiD5MHtj8v1ELSN0LjwFWe2hqj3n0OW
6rvnvEtPnw5wgaxKpt572OLoi6JBOWwmZQhaewjqzB8y33pAuBlCHd8tf8KmpdGd
hO5DDrYqgrNAsd729EyT42m1BLu5rQpaEexFAXbm/jxnWtp6CE3D3zX38U62l+mM
pk2FnN8IOdYranLePPqVXIkBlvdFu7SYSxsW8Wrh3+KKuGGhoYM/q73e22EKCCdX
WuIJ3G5Ylh2LNoS20fOnBJtbE5LVypiGq6pLf1MkugsuFMc7q7+KysaneW67OcRE
DgxDljDv3ajLF1SOd/FzOHT7dAfxOeWQcI+QI8D3/cN0jwuGWzMoYFUmPl2D5Ezr
LTSvH4dLzjpBPCaB0lFqb4RsUhj+mV0noYJyYoys5xDcq3d9hyWTjJGNa34butP6
amope4R50OtaqJGLW7yMOXY5N+YRXW0LOC24lRuiyIQMMtlzhevdEv1cBFbx5xHr
CbFw/UhTwnsyS5BQZlymOrzn4d2gCKnW7B0fKKksfiZLEj97QmpakfhGgajTZf8A
C4OYYtRO+xr22YXvxCmaYNhojayS4Ouw8UP+b58CKoCIg/rZ4as6UvknJ+rbdI9l
flDe9S4Apgi4G1hGqabw+Ev5I9QNG0jBOnRZgIcfXKWrhD6uNAaLzyppx9Wv0PB9
X/8aLsAeXg1wJqfu2fDbhMKRanIZwuaN6NP4GANPAHzV9BnE7nXbTiwDHnEJiDWd
WqKRgki0j01TpSdjen1T9168iLX0ggEvN1qA5btL62xORkjSYKvKDl94BMfoYCjq
jgb0HiHbp1evShQoiELE2MBkDmTb0aMM7cSv2eI3aKyljz7wsqbjo2ujTrdwC+r8
P1D52RD7nF4vv0Qy//UybsG0wQVKBO+BuCQ4wsKY+mlaiQwp79BzFDF94xy4G+wt
JzCy2Zu7nfI6eZyUeBXUgFQf6U32CtTdUzlR6Yruh0sk4cmZKYKYyYNBIttb908J
qpW5ajZI1N1+7LaF2Lp/hVuiTzicQwrEYs73WeKtDINZj/xLXo0IidKB9vo+dZwh
CAkWK/1cbedXrV8DGfOsS4qSqRx3pZ1xmsswdQqCQBT9tbxBLURpyWjSbslmrGbI
iL4RgQjprJL9L6qDRqykvs97HdM/etQUivnNOGNVUl4vWjXMRXdNG5pD64DuvBsa
7BqIrltILpuYxKDWdla8GrVTASshLX3t90FuU1Uf2Ot0bSRZsogQoIHWfnMrytyq
G2q8pntCXtI+iEiRpMSnHJes92e/6H21fLzYeo45TZA5cKuqlxDbR5dSXQu/M6mS
ZnhLaZqDAP95HZDBMoWrHdbDLo3MtZwMn4X9M5C7HhV1y2NHuO2cfNVjmMFu7Kwr
INro5D6U7xRcN0Rohjow7FD5TR3uC9UuIH9hIqs1+dD5jRpPy5875iXH0B++lLpk
F/1Xo/D6Vx4Wyhrc/G0qBh7hFMh2bKQZiFzwGhT//iYd5H1YGNXs5NbnNbjqvzIU
R6q5j1pWpTMZvqtsztilqaw/35JJSBusumd3HeAww/wb8YgB8/fSi7H9GQgwKvja
oy0EodStrmzShlpx4O/w9sugSx4aFycE6sKA9UX8FF9E41kFKjo60PABLWiGLJPU
kCP+fLRtWoqnMrhPlueCGaDVenXs2aHKBuUpoLTMw1OYNn5sKlcfS1zThzKNnLiq
+PWSAuGbML/nSBiql7J525knC5qWfPjcL0K9oiZ2T9VYA3ct2oUNOuaDcKcmcYge
YQcMkac4HHghlaFe/lix3g9m6S+633HC428iCrculekUEmEP6nlKKPJLcl71bKvk
LNd5BLcIV6VU8qJTWTp96jJxli7zgUzNOJE6wki0us17EmiQUfY5uwoF0A7ovsbP
OjIoGq+K1AZWOdInJ5P9Uxjvl1vM8gkhncPyJFDN3iv3pesj/1tpYQzkFEsx/xj/
trm3d2q/sYPLpbD2GKTpBJV8BSjE0mPaytkE4Ob5OnTKgdYzTqjxSpkWdbLHGdTr
JiwK9LKp/tN8u2uc8JWP1g==
`protect END_PROTECTED
