`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4MtRyVbd4rIcHg9U359zy7TrS+GzbBn2g3G1EZQJZKZOR2BovLbuf53P8fHFQ3me
QwUtbXApYqveh0jdjBXQQcrkuWmY4O34p7XYql/yEu0wKIgOv1NhtExUzFhPRn29
J0jIwTAcR6qF9KnO1RkeubzqSjLXibDRhu3vKdoYGrt3DVDnSZYkedEvGG6+bJiU
Q2pYp48e4psgLGLVzWO0k0WphAvm8DI3QYTFaG6Hfh0yzHNt9FqOv149Xhi9I+C7
ieUJzk0ir2ZVefc5K22VgEONt1aWUbbTNRXzVicjvgPWTRTwgYogYMFpL4RXOGFY
bSEaFzSpn5KZhY5jCsV3FFXAHiaRqB+aJRQoUK+TEr51PyF8Gq6LToftEQrXBGWU
/DYSYnoqOI96estuSijorcQTtW1ZNXxhBmMUpl8Wkv54dDhqBcJakVwH230pP5PG
ITx2RzVtDMf2AaVHDYYKYF4M3sQ93j5z675iYIu0tdgkd1voqNAtlDFWcWfbBIDh
WIaLpZRLtX0SLlBzTRvwoLOfDbFHHv0nfeB8ebZjQG1O0wjIx6egdTd8WK+EXx4N
jNG07CAKKYWwCF0olhVluFH8bNT6gp0veakmJaHjx45LP+Csvp6O0Zzs69QPZZ/t
BLwyu4QEJUOwFoDJ+jpQPXHziV3sSOyp4AHw9J7JtZic13ki8A3yNiK0Cp15dxEi
al346fjRx0mMMf3H6QIa9W8sSunAuwGQK6SPXiFRIMK6XyskNJ3b5qUKNQ1pYuMH
c8s7MDweVoqo0rgd1e1aVgg2QodevwfL1STZwHF4d/1vByCO5YXvKF6td0qKTvV1
`protect END_PROTECTED
