`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FyjEVfKfHnUovCkRY54dPeSfpcg/6cI3/m5d+B9MceI9UcGOicDOpsKVCqG+lM0F
4cATFfhCSDv8QBxx5SUHg0MfwSe41SDT5kJCcCeFHOZa2aU4+Ztxr7M/FQCfc9bD
eLAAbGs69vlb/Mp8pK5vwj6uoDxY55ltGGuog6MVeG34MW0nsiVdDCgH53tP/qnl
UGTAOdAZpMNBx7tuBSkspV8VXuMD/Fnu6q/GfrfjB5ICJgo0dLxxK2meMWlSYyy/
RJfQFvPNGUMrVHKmzE1ASA==
`protect END_PROTECTED
