`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UXJ1Htnr8uTnvSelAGPgWDQPMbW7g+6wIKTRY3R5+AFguKlmKIa/L5LXuP/75U9L
BJj6jl3J982wz2VmmRtpOMDMYSaXXA1WvJVobqKoTSNCrRBklDFREss4XhX0DXqf
nlnSg/ZjIH0NgpQ9/O3ZxA==
`protect END_PROTECTED
