`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HOISN2RU/XFLrbJHBX2O3FUdGlwuXpNYyiuCawZ+T7U7mHNoZrWrohrCB25chLsV
i0U5DqxdPzc6EpzNlj97Ac2ZVm8Yc8ZBdklwQ57e2UPsfSkHyFjncAdkRJ1z7TqZ
IAHY3ZTnFJckVHBLd6wzxWBAWVZ9PXoanCA0uUpIWGPxw60NiayJZNFV0jAzFs3N
pjP7pMj2yreoEBPmKAtrSMaRoEI/FWA/XVxfZezBgIsN2znXDGS/bBeSioJgBHyH
j+Ss+L6rTplZhKCx4yz3Qs9PgtONyRSXbkDE8J3bejnW0U/0tSd3Xi/aRLXdZqjz
xh2tAaKQYeK5uq7QzddTfT8tu82SJpdvDgtn1u3fN/s8g8F/flcdtTkHnaM9AiY4
TkJh7FHRuhSmJYhD/MNdPBD2Pat8Rb1hvby07EGSrEgYTDOq7/DmkThJ6tgrQOil
`protect END_PROTECTED
