`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WdAk6iAIYtb2x0MPE15yCn7uuzZVyS+8Qd1msuWr8DHOWLs3PJbfnGPdUFNvmVV4
RNMpihQRe8w535HE5nDYOorg5Sg7bNmvcS84fZqv0F5DK3ET9jpWL8RMEv6f8/0V
mdpmV0b2f9ng6jUPqhYW3aL6IoljdpQtfuLRCX6M4At39PyN0FSsu/arJaABRJZl
X+BhPStXwRFJn8Ish8AusILHaNgvQ6yLE9WlFwDzPRXaO9tnAS1PF5kRFGJ52Ixr
C8VdLzCyTm1fkJCMPanZND8THlEdvhw5XIVSQ+uCL6wqM75H/LOM+Xnhq7Ys+6H4
XEVLkuVUWrL4u8cQPNvvvw==
`protect END_PROTECTED
