`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GNRSPZSA5uM3x6eVx9pX1zducxXIDZzKS6TBMo5McnSJwQ53V5+S7DNc0QC1yvkh
Zbz6Okc5EaNa6EaIREJ2J/Y8ehBX2PfKkiZewFefxoI1r9br9KhTHZtZtgRiOPoE
0dKNAYgDQt5nKi69AE+1M59YE2b+qqoVhBFJolLWTF4BSGYWK9oZIZZhujO0WxY3
hD1kIJPWgNtmlI2f90qJW8vk9Ihk/UHIkA9HlZQsRjdSHGyryzP3gtmmiWIp/Qih
AEDtCk4uR1i/lq+Qb42C2FecSg2vXOsdhu/qzBJYftkwKC+kSEFk6VUtZr5+mxk7
Qg00XyrytkUgpo9pHrf65uGZ9KlPHl0CIdE2jalthg9ihyxQ2HT8aa3ASJuvzS8z
+F8nyK2P35cQh3Al2Xt6y74xv80CkDGqSE3A2ADFFDKt76AxZtFOtuQnoF0j9XR5
XpaRXqIcPXTkrQC2Gaa2nyVwmEg6MygTRg+pYLCTLQ5joIiyNw+EPAaddPfNlEwr
sZBa0952+DeoO3V1MNrJk60OqaHbrgPqGDovLGPWHdWkcKAulA0TBASRWrkmEVX9
5hoI3DSJ/MKGo1bFK5+ZqJ750XACgmDPvD/vM3W6LDjfSMMImGgkRdYDRDh5fZ0a
rYcF5Sxq2YT9OXWhAKnm76fPzf2HOt84gYlh/isAXyunkE4LjQxoTfgKD+N3ZP/b
R5VmrToDYxw/YXfA4klk16xAQA4KVYvZfFP8NxylhnU=
`protect END_PROTECTED
