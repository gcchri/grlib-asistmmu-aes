`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C+O9WxKVAAdlHfeVv5WUAsgNF/nvtu76YY1umQggUKDvxUXTBe6pMRfs0EMjuTlb
5IUHV+OSC+uyc2c3CVm2NImW4x++R34A9PUn6muVRl2FeWvW+sIf8jwpd8euE1mk
qLnW8FqKvxiIfvPCi/R/ygZd5Hg0quDWvFwRCufqijSqn3aRz/YOS/O9MUrANizf
yWDyU2PF1diE/PS1aaNhqOuutT3DI1KBrsxhx+MPQ/TbRI+9UXcLCnPEIQ6pYWvc
ksuH4BXc75IlhQul4hiK7QvJ0j3aBRXXXjBQdqPT2gDmUMdHtWacGhIBNP1uvDD0
PTO1ySDFSkU/Vw8PItA7xZyqhp90FzyiaUCJJCkGgd+gGlZvWfNfxbglh0T+l3TF
SKZ7HmXAsmZKalwdJh5ldtUWt8u+Gn0VaO0KAsQSkTJmY5iP7NQVLvfCOBUPVQho
iFXAeGzrK2BLwBmkB2cWrZlYATy2FOtNbqsblrlj5gM=
`protect END_PROTECTED
