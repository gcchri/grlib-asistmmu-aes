`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jATEJ6CT+Z4JB250Y0A4F+IIyxrSTWutD+40EuZn2lFcJxucHvcgZv3I7ZKRjxlG
C35HXXLbyrO85vOk+G1eAI74aXsPPu5l1plW19jD4VDbaTU4PI9XtbazXr3aQIA+
44VHgrXUgDI0pZ6MXMOQ8d0EKeihe4cEw9hEnEV02ziPCQPeKvg7k3zw4YfW8GGH
sFINSit9fAKLIC7Ez6lkiV3lxZHyU1rtmY5m+YHZk/A9eB1/5egheCfXhv0ppZ1y
Z836RxBB+OCEN8myyHLA4j6N2nU5hLf7tK2qXnz/Rtd1jSPE4bCxxkySS5dBy1MP
12TLkKlWtctq304G0jEqk5OY/e/guJaBvjTFM5XJGUCv/Qnf282pUwmCvnXheFk1
4IglqrS+s+no84bGS7F+klwR9oi4WL023qynm2Tst9Jdh7jzs0qMY8BU4+myoBNi
IJZUiR54Q2KOwKSfPugDCR3593vLDRj0W6j6WBm4uZeTPbmMICdu9sgoQDz4s7ER
KkTRoKaHy+iUlG05Y6rIhlNLO+69csNahTyVMWvbuBZKmFmnyvuudTp1nwya9jvc
`protect END_PROTECTED
