`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ic8VaKjyLcvh50j7wFkdDkT1B9A+OF9KRfApximIdEokWYDlFkXrhgbUWWZZn+FB
BV84VgqGYkY7tmQDva6mj5niefgNL6MiXB4sYHelwACdQtKFgzjc+kEdexvZPpqu
bC2f6+dslklgicRJ8T+j0yq6AEbyePDciv1FvETtET+UqF2vPEzN+Aw8liUkJjhs
NT9QMgPOjuk7ohL0izUFyklBIFMrd058BJs4O7FdG3mPzLh84fvQn6F0X9EMA8PC
yIstnChYMqygu7DGwGIuKO2Vte19XpEb9oMUG5sD1EgddO3/KJXMJlVE5EXiT5m2
Zgzuj/9iq1G3gPbjYePilH2vcbQbiY7TjQ5o6rGf3yG6Dy9Dl/Ie/OZi8LfVUxJp
j4q/m7BTm2UR9u21qyvAy4Zzulzivg31ydLcqDDY4iFMSYoQVrrz5CPIqU8df/ze
tL5x0wOAZeQiwcGzoYwMBfDICzkD8K0PL05872MBPmO2XjrVCCGUxj8peIca79cw
LsLkdBA0OXIhokBzgzFOuMm1i6Y1Hb9Iq2mO/7kHznUR4ir4fzSVmR6LNd1CTp3y
dDzLxC1y1+/ga/5VkedoGbIuo9xgt2kAIrI9RLa1KSiscbIbBK7Lk5r1rNR8dUGg
7nuX0h9zYV5NWg1MEzWlrhT9/8OSMWc7EXP1tr960L3kJQyP1h9O7CeShQeim++U
6oeFqfI5uBSAeuO+ijLGEGAet89e/bvaHvsQFCv4zhUFt99C20H11A0awxEtS8ph
M6+3eDw9HURaax3/aaXQIBMyGjC7vRtmFrCCdwxNk8DT8r6sckhRuXoeN2SY8Kbp
s2OyjjhjLRuBoQs+sWflcLkkKTggQXYKtgNdwnXQHuJ42gXypblptUCKcvO+k+we
RGADYp0XfUOvXONdHTjKQTPIkjWOhgE5WF9Y7LcrQX7IjJgAJYeC7qDDx4Eh6VEg
K6L3X1OfwIdvWo6YhVMQHlPC14KploS1raQ7oVo2ttMrGVT0QW4Ny78wgSHSc/zY
tBJRxj3R7D3FDZueY3nFjvrRJEDtNmYIblMcXtuPQfMUbuADH1eILKsRpx8V2trE
oxCipkXuWD/CdLOoN1NR3JOauXzu1Rm7ocRkuicoGb5ybgnjIwe5OQzdNHVuwqHe
`protect END_PROTECTED
