`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NlgYwp+GzvcdsMlRxs5eHvfyNt4/vtBlkfbPiFqxfjOLu0IQoPAO8si/Mwls1dk/
S6QXWgvMPQov+Z5Dpa4XQF67rDtB0T6bmmFqK9qAXvAnx/I1ku+7ktUfUku/3vrh
4N6SBI7lIrH2sMgMyl3Bx6P2nMM1fsf823AIFcZFKbM2maO147SYH5pM9Eb4GR8U
/mh+ImqigEmEWa5Cy9FI88yB1ZCeqgQvoxLO4WY2iKLPK+xb6EC6EI5TKs4qBw5c
zFHhVFojXaWW30KaVrc16Sxg0gQ2hpSOEXsdrD2+0PtBfYR7nS3hnpTRe9Y8O8lz
8JYxkkeilRyprfNEw2oCp2MFTxKEutnIYng2Al/j6RRcUOvrzIR+IfWWRMTAosNp
NQIcH3QBVXg9Py1LxXTSacRKQrwwzyUzodXMaD1q1IzDcjwzZ/5lczMpa9ceBJLs
GlvxvyDipIlEeRsFz/Dxnv0OmcEFsEtYW3Vx39MzBJaF+mHyWy36tqW5Gv/QhH++
rY0AHmiwpuQ3WUytx5S9CxF6uPbml8DjSs/+UM2Yv0WAGcAeMQ8f1yAfvmF6GgL3
SX5k/5RfYBHgEomeJIbq1u7C7XBRXFRpPiQmDHD2dMBiGeLdjqq070aHi8SqkMvS
lOv4lL7cdWPr+bmzkSQaoNTREeJLVfGLfKghuNWPDgd3XlV64M9hsvIWVvAZ55Wz
tk6XNE7jqmb+3ppJVDaSD2YFL6LSXDQ1iaCvulvdv611N7EOEy/87cWvffLV9BTX
g2w9GZxWPEyno6C3ozour0CHnw21cb92D/WVeUrNzGLM/pnYum1G9GoCpZE1yOta
6i3HvRBhlOTPqV7XRWIwVA==
`protect END_PROTECTED
