`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qU0LqeHtQISNMkEa3hz8jm2ZuzrDxnQLDXdksHErst0K3ELWJx07IWmECM5LD907
hmnxpwy4KAkndJDLivpnXOExpeboGi/WONb5ZGZUM28TyuBdZbueZAeJLReHCsk8
20zYUMeGCi+v2jNxs9iWiIF3VHKZDD+SBybqbceQzeqB5mRd9a62jXHvgQA/aZwE
za91SP2Kdo2fH1/Q5iOPjORSXT27629915yni9eD5y3iJCsnnhq7ehvz734pT9N+
4ZViUDy4G3feSPf8f6x8hKl5t8BuD3CA0YtaEDOYuzNUZgnciS9O/sC7MQMwIDqo
bxM+KuB87546yZY+mmJX2HSSRi+lBcqN2NuuONFS//ONHSfZisVve0RVJg3NVE0V
sJX6y7r0yB2+I51AhkvqZD/PgXpw/Ly+HWXEk4XNhpsc28iyhXO0r3dtvDs5nEWK
`protect END_PROTECTED
