`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Z6UM39v3CNuSTY9Q4Taqz6d95XrWvaNxT5yCOJBaieZEWMI90UrLDeq9cC6ABTu
jDrX0wLtGzLJUVmszU/w8QI36HEHESYaJq/8a5/3wP9FoT04qfO/b0o/ynJ2fEJr
hbKqcqKxycZ1tekjqeGTt3OWDjWjISqnjJFnDV4uf0ec/wz5LKjDdMvi3LY5BeCz
+Gt+YlG3wMvLy7RwTgce0gYL3erbYq9BprrLdOCEGut3RAIzZjK89XL/hpmDJH5/
pDdGbL/TXqxhLHzPaOeQlePZmWKo4DF0CjBSsGo3DyKKkzx3iDnZsifo76vQKdgS
iuXpB4T/zAaqebey1m3Z8Dhhb3f5trjov+zrzPKddcqsX+L1kN+7yZt92PpUsa21
pbkVjDckI+wf03l3UtVOmDKTCfJ2IIH0FC1s6OjkN1hbpXplGXcniG9pUqBQ790m
amXsU+tRxK2VsILkL22otAKdTSTx5Rn2GcE1xiHB8bAc4mg2d5oDZnBghDOLU43M
qNR8NsCn+/eEOcDujzIi9cY5cdIeSjrGU2mfxDzyduoeDt4t7Ztlsf5Ff5XZPGtw
gXJYypM8rslThaTJK3osLiJGPLAhFSxezAvETnFu/LzzPo4rdlP86nLucBHSg5o5
dnHddVzGhip5nlm8czzxsv3WNi5KjAk7l+UycQXG2L2VJjdoqlxMTMBY864qFJzW
a9pRlmoXFIeWixThYdg/6QTPp92fIlIVhsDlQT/4OjBnTf/ozQJPQNKLynK8bzLn
VwV1vH3DGSM2DdpLTfvKUsQTTtnsFd5p34AyTUhNouNAjjttRHw3vFavvjI7Fj26
I3to3VM9boQpA5xFY/Np6w63oKs7kj2ZYF+JAjTMvzJtrULwtBxn79/xC2AOZ/dN
adXDKJDbWpgOqHyd+Ud+sh5QeLE8Pt0azvR3s0j2YJy+AdNeFlt3IPhtz4ohB4KN
GNJq0TkPKA7geCWQ4a0Id6LM8I6zKpzkg1eFHE+kM0ea+dSH2U2SJVoXtKY+/g5a
nhvINNTlzwOGTEfaK4wmrg0ta/vt2/4xf6ERABtec37/RXXDYm3eYG/9ICIKwJKI
TeQdsjAsUVHGL44zo+YvDA==
`protect END_PROTECTED
