`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V57wDkgIcOMiBPV10vyel+Fvngag5xa27rM23nrFWWhfO+8pAF/m0MVkmeAPN5Zq
EQUjCJPlAxKT5DRwLxOckthoXBh48v+XbZxeMxnEvYcZlQgOJS1AzJmTSdITtmA3
dUA4hjL842VykTjYC1OFBWLMNFC0b5ONUhUAvdFtVejh9uPgi9cTF79BMnqM3S84
bBjeWggp/EOz169Qx+Ho3AgFrz671H/GKMhK7HqKGLjbp57Vptbwk7h6JlqTKf6u
y524k0YEVs9O22aOk6y/ZRD+zkA8uCvtWDftBlzDZE6LfkSXbu/95MiL9PCEfiB7
tTjcRVODRlhppAnfauaZMx9Vh4TcU+eQuHUSKOajiLEEaS09fOllOaptKfQwz9tI
s5rUfDOGkVct6k71+BfaQYfSh0IebExFDF2jknAgrh22HWhTLBhHZJAg/z0YkxsS
yuOXNDvrYx/S/nSISM0kOSBdiTFFdnnRlGhQ6IGoX4BbJmaPpH+Np+39MpjTKSB5
8ERO8H8lK84uYZgGyY7NbCPk8sa044blEI/Nm0MFmfbR7UUyRuhaUuUpa28CyH3g
GTBGjOppnQ4PDkjYTatFpXF+6iqpUFggQi97Qk+MykkLiwZmSKWMbxQHRODlzX6n
MJroFFxtQ/s9dHe2ZJENC1vEXzgV+Ty4IrViL4LmktCcYkPEx7+cxU+r9Byp+TfV
7cCFysJmPOVEJ+piad21UBX+aDKa3lwFtETKzUrzsZH3LJQ9f4t/J79YzQddpkrK
PJLSv4p51/5xVVF5+w+Mj7u2N7U6YWe7eIZtEgmThyTfLk7VaoUYUY9ugv1Mllqk
0ocdo3dMf6Hj0gGXzTOHMo9rZx0jkF6i5RqvDf+L+Oo8OoBiDo3bIcPzi+Z1bYM4
`protect END_PROTECTED
