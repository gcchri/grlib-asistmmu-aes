`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6VYT6dEEInCHISVbBN1Ccuem7ihNmxRNOLx/xX/17wrXjxz/49CscGYlPUy8URSo
SEYoHvlM8h+MHcZiQCyNBv8CUbSxAFtzHKKo4T5Ep6N3hiS3wYLT8TG4icUZEbEK
Qtuxu7nXbIjRtiySu6XkcoJGUlH0q53qD0Z+naet4ZYl4rU7WoJmy4Hs/YiArxu7
aYsEMqqe+lol2eVfjO8i0GIvjsIXRWiBqyR3zDanYuv2C484SzUJS+HmAvnY3GT9
n/0BICJYAVaWPWRTMfEG6tlWVopgvXKhFFscSbORf6ZPj3oILl/UJc7B/0efL0Am
V1t0Ivs3ZchoqSpA+oLCRw==
`protect END_PROTECTED
