`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nlgMcIpSidZC0J9OLSxif/sEC+m9UZS+uj5Rt7+h36T+PpK84AU5oj8lPQR12W38
L5VNizmcgAlCu0IFoU/kd2sSBPgLbThnb7AX/QHO4Z3ZaUvgw9ngHvM2GcF3u6e8
NeNL2fLrHNrxIvVXlyXD4hHjGhpX1PmoEpI3qIh/oKtYxSkYsK7JylJm9zPNrR/u
jU0+HKqTAr3vzlx44yO4N8ZHcZ2kbzJxvJpfTDn0/1T7MlAsClWtXxbF1B6VvhA3
Wr5Vnrgtb7EvzTTqkidToxpIM3KWTWHOCj8elayQnV+SvxDBxW/kD7FnahDg8HRz
MuSUNpAo+rl7xt9myCJKhWmIRFgQYEMj2swxio42VIUhQZT2E4LJ3Da/mFPJQw63
LxQ3VNqygTBny0++w+7s7nRf9dhd73mgpNXcYHVj4ZX8YSdYf3gNH5TBlJ/HwT7O
9gzFM1BbTTuMux5vAiqtoIAgRxz40li1Z1Fes2DhnaSWDVlMQ7bWiu2oW+ij3DRr
krwFmsEN006GQHKKdoJOB09tIKankpWztv+PIg26bJNY2QAr6/48pbiSkGLttEYH
jF12Ol36iwTBRvf/I2aadHRqUsA8uRzw/jlQhoZyrWGDCGNjKTW4t/pIyKVg2KGc
jM3mZ2tVsMrkuKuqUHp9MrX8DxCkIZXDjO0IJtmfbpA0W4FHxeoPl1oxcyaNygFs
zRVgg/W/8Yjy3Dd2+AqNUhP/xPo15hweLZzkkbUx1lZ3nf3yhv8faLvT3pMN3bam
F00DeSChcZXkUV570sMwXKmOqQo5tqedcUtJhGDbFF8/jU4qQ0+kAfhMaRlwBOc9
/D5pBfJ9m42o/PJ2t1snZT4vxIb2rab6I42SsYAf2QOh3XeAIioDo66HUzaRtqrO
4XK/BRyF+x5AYaImVuGFpO1c7oZ2p6Z0NTxx4/s0BWljBCqkGb77OlXM7nOUBcem
vyjeFF45iqVRlm91b0Th3Q==
`protect END_PROTECTED
