`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dVUE72Su8tRegzT3YOp+WCMxz9YBHhGwiqbefJULuzzKjFFPRSUwUT1123O4Pqto
4tfHr4hfE/qzAI9YKP8pLnEGItymObURil1/kRV06tRJ073AsYLao+E9KXCBuiJT
O4k1IYTX7OyHmX8QBnVPAncIssio3K4qbKI3G/I1Q8ZFwgI4qMVY2s3Ib5F3YK33
6XlMZOC3OLg6+x57UXN4cHdn8wLIJf71cFM5CyS+vLMJ559s3Nj5xqhuuyyQmBte
KlznRrk8RK4LEbli/Z75BfgI4N164sWPyV7JQwrTYE+PCOItgfchwUC1tPio5ShW
YNBQIcGFxPh/QU891KPwPWo7kTiK6R1WGTPnh8U3bOWyLOWJJ8r7sEjzDFwYBqj3
Ed7wJQwUXCYE/jiN88f5BAA2Ye5FCG/CaWc0dOV/02ubcihHWUlobnhkeXpETZNZ
GnQiBAP+bJ+HDKKG0luQdYCzSx4gR9qaiM9b55/mKhf+E9lE29GgYVCWhkq8brya
R7OOK5pgLuOWKZsQQWFxHOlIN+DlqV3/Ca/mprAOIfwbso4OStDjSnCeH8ZcbO6t
+nomy6VYLziaShh5ahHV8rgRvZMe9Hjfp/0kxklbBLueOf0me94VzXiy8V6TrWtT
Vv5XAVOT3oPMHCpVBF03IggQC4OkZ77fFqG2eCe3UvcgzDKAyU8mpKBbO0yWCiWZ
QD9GDym0xCYG5Xv04NCqb5PfTKdfoAjHlaUYsTtIlvTwhxwigny7wmI18DAYHxND
8i4yLWuuvK/D5K/woQXb+WfH/wnuKI8T+TD5A4StoHyMg40ru5fYiHbBZR9Tddik
uyxNXJLEF/Y+Um8Er5kAInKPDkADiZ2esGXK6w3TBbXZrlWHNi7YfwfsEMix+Ap6
gKiX/iulzR5OWLoxc3XHZXacfxHtxis8bkTXoSXdj06l+TR/9n87HYzZEfqAOt6u
rcEz9vviEld6joJaaC09yGuBXxGAw58FnT92ZMfuR82NsmwG5dtoUFhkWbZmjIKH
veZ+DRqbpPQwIYnbohsqOtXAUJ0h/JRkS6sz4ly4u3AFH2FiOqPUj4xWaIUpf1Uj
N3PmTP2krBxBq7ouF6hPFWV3mTbSd+KfpzBExGGHf6T+7HV75/aW+kdSOYAMdtbM
5W0/IcPFyAH7813dHJ31ByhEARPJ2vDdfh8ytQTp8WDPIuqUSFNnePSPjKFatLEv
1MfZhLlZ1/usDX9TH2iYxr5IumEWQUklT3WjPbAvEdobb9uUReXIAvewT0V8p+wG
Q84gl19EUxZ+naRglW93AZG8dHwE/nH4Sz7FDOynLZqdDTDW+sGGhjjhEGxOt0GD
K9xl9RcQOICbtIjVt77vV0xZbJl3AS/0i4A9GGkKPhwQtJTtRCewjXwrOlUmwcq3
8BPQymEnud+PZTCDgjRazchlC+U9XgvnN9MV/ULPGqQvGs2pgppnMt6RJdGNs9WC
egYD9+Q2g8kQS/mNFaqYj+ENMTwK9gXZot38frVf9QJM6fIbQmLy5ck44CL/4A4l
Qix49ihWoD4qZFb9Ebv+/xswY43UBfqldpB9bmIFC1KfBJMoED9iUoXqcELG6Ivp
`protect END_PROTECTED
