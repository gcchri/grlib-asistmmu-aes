`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6r4IPyhkjh1RRVjMlBjUVl/xcw7cPVH6YmbjNwZVEgviCtrV1+t3R9gA41Um0xza
ACncWBaqMstXs5e0M3dgUvw1KhdZq6QH7deolp+ZYU0COiAvoqZdiCjNexl76eXG
kqPJ/sKKbLciKlMwCiXHezHDn2qxK3n5yz2kiNYckdkqWfzfp2Il/xxrHvvowTG5
7S5V/d9fJ1pCMyiouf9y3hQom3zf9FereO/W2lpoL/yaVDjeUTNTKpiT/TQm2q7U
vSTo1obgWeuSFc//zg7+YaX+AR9WjLuJvwhM5sEI7RULeU0xSu2OEz/LuAJfQk0p
L+u+NOSjLJEldKaNGsfvK75iYuT4UH/Wqbk+2XLzagfcIHX1lK8B+PGGEkzWcKeY
oLzq9/IUlo3p5EuFNL/DA21R8RIW+h7qrx/itwtqfR7mgGu3VEVel23ic2p45esa
yzCX/l5BMcFClfcKdXN/tEq8qLP3Sv58QvNvUwwFrSkX4PacubP1ajNL5gg16dwG
xtqs069ENSkS9brz4u1qFkS0Ygxcw7MKqY2ZN5mBcD3RYLRjH+G/svwXCLZqj+OV
yZn9Kw/J3jRVdibsA14gZ9dPwRaL7DX4Ay/52AvpZ5i/rdwa7kfjIr4t74XrV+UW
ylSKQhRqjm7JAB0xbeEvxfnOPcRhYw1az/NgGOa6kb/0uec57V32hJqdjz85qXEm
Z6wh7mK16d1P7WUGFZocKMiKkuSQLLfQyBcu8nVaKrzl+EbMVPzl97Nl09+Zz477
EVK3fR1c3q5dYOpmgguQAhweJsHrIH4zd1Jv+7DEzd9BUxoUZlL0oY42KST+MMbq
AYyeRCFpnArYrhUC7eqKxrBPAZTtHwZTfJfmffOFE1rS6BelAcsae7Latk1aYnEl
Rf/p2v6y4hG6HO+MrFrilSJeXZ5qLw4LfrT36Si3n/2c7wz6bIvGagk/YeZ5vbKI
5Vuj5hGIvDEnWYAd4Gtla/TKYpolSqhA3H9X1Dh+Rr2krJwvvA6+pSyaSWRqmeX+
GvXBYORJLtYQZmavVPpvVq4Nb+FXsQ11IZPJrwdKJp9V7RNo2qioHx/fmSi3TARg
QzZB57jqsr5ZVeJVDEP7vOIQ+PsyyFmgR8528/naHDHIRG4pllBsl6pCOW7tO1oM
oPQ8JbEs5ek7yDdOZ43xLY2rz35GyH9hPBDAh1PjO1DrpZ+5CvJOjMdmtzV8NXx2
jaJAnw8PrbSGgMogrbeFPPByuVe4ml/iv1Rf/vd8wZ4Xr2xzjS4rdaCfHPuLdX72
Z0/13lETgERwtzc6DFFPb23WcrMRhKTnjKvuaO5aa4yhyVQLBE/jL6rD7mI+nk7z
5JYf4l+wI9nKmCWesGMQbtT6kB+P6oSv3M8R3NrEnDYLPw6iCNCPjbvL55uNY9wI
b36bCsK/AybnDibew4/dT51CRiF2ds51ALfKeY/T2A4S0LgmZmj++LbSd2CRQ9kU
OJp0p+1Geq8WixqRqM6PjOgizGbbSopCJsEvzQ63aBJBXx57sJ3P1Kw9i3Q53Zij
ThXVwf9pDzzJgpM0ucveVKQQIqUB2TVdUU14hDNHy46erm0WEpi849l5xK+G9uON
iFa5IrxNjzsjxnWAcxJExfuke3owk1RbwnmicDraUJW3FoMKpMKF4XMcAwHqTDge
UvKV+dq3JozRIz8hmshbfjdTF9izLHVh/vQoKb/l3Z3iSHCjv0JlmmQ6ukfTiRFU
eQwbsUPNM1J8wYzgQPSRvh5stu3xORHfgu8q7Zy9tbJnlFJ6mY91JisN2bo6hREG
olb6t4l9i3qBEDBJcmreZZf28GUp0CNWJsqgypHR+GaFd3nkri+9G5fn0KYl1xvX
gD8twfsD87zgCZ0ixllulJa0NTdZDMER/r5y3TGF52Bulr14wVmub4/qseVmb2Jf
XJeigChk55Y+pCmZiZxclZfTkGWmsfqLDktKigraTUtArm4kEBAFabYatFlKQT2A
g1lzltxdziI2PdA8xzHIsZhkTfjfiPp6xs5hQFzAdIkBz+y8jEsfgknJtPxBRlhG
J8i+bChpP18ppcbyqiibiyWV1qkkh87lowDj5I7YIO8bSJnlPOCY1NzVBBGkBtsq
VjzR1P+R4ax/ynwzoZvwtVtvrEWOj92Xu0qb2xcVL5lJPxxKJs5AvML3OYzHgJWs
WOe90+z7qviKRplvAkMseC2PJtqjCIbd+6WY9t8/XTN7ddr3BHQAGdOEmjDjK8CW
C+4rwP4O0TuixvnXAnnIvg755m+ZFHOicjUCqki2YEkZNUnnKzridCBjI/0CzV4f
c5IkoZu9q4x1tTPdYVqvu3Qe3/33VNlBaoys65fXDHJGKBsAOxgZ0L60cM9w2oGZ
6VabSQNLn/WYPYHnZpb4SWYDtr/Qfrg2BsZ7cTE2Gb845I1QFbZe3TGecmPiOr7c
kpjt4UXpldoOt/sTHXkuzHn3Zc+pbbACsKFMqdT1IizJi/mye+5NOEyFUGUP1054
v2y8OgtcnF8imBGATvHvSaqgVFjj7imdPxL1tih+0o/oqxW+pNP2pNbO2T73fLUz
C7tCQI3ygswwKQbZFkGdacFCYl0LLQwzDvTLY9TezVe064WZbkXo+ymVQCilcZav
6FYw863CQgUQac11DFbQm9LsLjIR9xiRy8+AaLNxfvSFDQk2xOsx7OgBH7Q8eT/Z
ZpdOs6zd7ojEaTuOA2uMw1Yn3LIr4bcuDl1SKkAGaqWBBwB9cMnTYRHDkX7l2GKm
AyHnOMIPpeCEUECto/r1xGonk8851bVteMWRkMgFu1kB8SVe97tzsVnxD0DPtp5h
T5DHFCyrd454OvL1zEnx3qbaAnQdzN7AOGWKQXWron52l1+jLAKSMWFEtg3EWfeC
nE9F3lc+6Vn3c2YR951cCjYiKc6Qk5QwWS6YhSWxq/xoG/6zjx1ibABnMBekt+YT
Ps+ZpRZEGf4ZygftK6uGXUYEK86BtwScNWq3HLjnpRKJxq2oApIELzXdB4g6G38y
3wWnbEm4jRXzWuwivO7GTgkYl1QIeI+T7CE+Pl22UNQdpi/Ua8mdY5tD8tjnO/3l
9RJ/tdajijx4ngia0pkL1zPBUcOt9udX4o0Pjbmg5XXiJN0DWSxrwX02cIenuE16
G2oBf9KTu7xvKrz6MeKdAnLwYHjrxPmNbHKzd62emApzLEOxqv/fEywCiJa8afQS
Tee52Nf+f6+JZCuBrF3m29Ab+vwUxRVSpaD+kurWU9e7juiKALa7Uhc2yQ+yzwr3
phYAUnHF3ENsmdX47RKIdiomQt0aXv2EPmfn7hEQFRFYthlk7DrXhh4cXDXW5/pU
HDfB8vREKa195g2tli7BmqmGkUg9aGyM3/3W6+Mo9PB8CLoYZbF1/saDq3U1m7i8
ZejBiF3WATZIPPuiiEg40KcX6ysjigw+I4jomg27AMjmgRWkAYOVGGcGMsrIBunX
wLKW45xE6rxns45YqoQw0/1X6AVZyuMuHCcrnhip7t1g48Vd6MVGF/lE7d2JFLjj
5ilqCYbBin5AaatOMgPRx8xwBA2NO4o9qEvWIvyI94wov4N5pjmSktL9L4JA4/wM
OeHNk0fayDUdutGbXESmTsTGkludVNtAiQZj0bVmWagXf3UnjiBkHOTYiH2zAUJi
zRD0Fp5zfMuUBtXtVFH/8L/cEjcvdn9omk87n3qCwkPXjo/4udcIbKfVdaJG8k74
O2Qtm2XquedNcjP3HV9MczKkryeiO24qtuddLN9eIBbKl3FrTUJM2HGmE8u4iW0u
/eB09ODOkT8i4pQT0FysfInFdVVWMVrLPJ+ots+wSfl5J1qtQQT4cduHaHEPWrGk
t79wtzBBLx7zanhUBdnHeA6SALchdPFYky9l+1mIk+HxdIBQ5JPRSRVEJyRUlppe
ugwns7hZkYffoHV/7KHGwtCniK8dAfFuJw5k71ncsrnFW9i09FTMeGivFB6akDU9
xK8Z3ZKB9vH1rvtdB47geTE6WDW93ryGvY8piSlE4JkKVrLCSuFIKE4iogGvqnGw
uKN+tcrZZf3qp3qwt4D0wUHdPuHW1m9Llgwr5EIiZJm/EdTCbpZ3nZpCwHrmDUcF
HzjnK4ME8+dQhroev0jp4XXKt/3829Fg0IVcXtTrtdWlZRGxreK7ABJHije87z9Y
`protect END_PROTECTED
