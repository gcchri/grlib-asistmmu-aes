`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GOIvECKIJ2fM1q52uYna33ewXLbxP5vAFUrmOut9V3OYzgHinMn0XAV7QZwG/PRj
yKM/2Zw6Eu1xt+5WCzyy8HG0Ob/hRZNOT4/5CAGHc0eUZmd87B84Smn/a5ONR5ZK
5g2Tl65QvOioujUAcM1NzMt/rNeUk/49QROq72VbGbafVbieyQ6JcU2RDZjfYW7G
o0qmdTOC8uOmnUmKrYp8BkuWpsiCFdLDendIZ8r0qNLR+UvatqEK6HUstUekh0ai
hn5ItMVgqLdFvRjwiYnaK75Zrt+MbG4xcQOF6cjCYGEmuPJ5T5H4tqGHDasliUi0
bG5J2yQFzq0K7UCVw1cHHSgwVHBaXzUrnX97c5AajD6+M63Agtc9n88Fy8eP8UJT
eSXi+ZZIWmEtrSDcA3RMfVq2nlO5k0jc+CmRLNRREgMA107/NVF/FfjQ6j8idx4Z
ON7xMg9guBLnkSaoyjnEi/N9ofS0Vw4ynZQCVbEWORL+jAd6fzgWbJbi4CktwJ4D
wWW4F1D/aLIEujtvNNwNvSn+1Nhslf0Sov3RxlKsgvp7IxxFhqG2OHIetLb/atLB
QeWbxs8QB7+i52jrYJ1GHFerpyO3WWE6Lc+nlUqr7yzJSJ/coYu61ALm1huj/X8+
YsBJlvAp6atb16JT8R/NwuuGE56315yQs4V3N7PszyKhwrnMLpcZubWvRlHtabCd
`protect END_PROTECTED
