`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WT7JNPUtGBQxg/v4yyJsoGk4hITdZc9lil84eBVBNpkNebGC8dRVGdTiv+0xdEJQ
y0WlguNZw/N0FuRjFqAUTw9/pAnPCnK9Kp8YLKjapIuVp7FUMSe19bHbSRYAnZPm
NNomLJqVXjqSvf0P+PARzKRCEFckB2BMiz1fNtjkhutHyHsdpWX9bq4AZeQ4QSk8
+mJ+whlY07N2YX5flD1R5iFDy6nploMEaAiIh/9EgAeVBfqtZJBkoiDS82YT7Iba
b5aOtT3EGq436svdVaV96uEUwjBtDP/0+eixQXQ0y77nA5YXEkEE3A2HKsUuXtdD
hopaVhbd94xUiiaw7KBnTmnnzCLia1vi4YB5qKYz4tmlS/pC9yuGq/SG7zm4ZUUu
tGKnwpq0x1btE+tnRt+QOLQagbWf9wNrgpKgiKq8Jsgv3CBxx3ZILDK31aXKxx3U
ASUdEwuggP4s8gCdcBfMxr68R1qqDqx7zEBKS3JgvLusa8cjaSKaYqmcALFjPpm8
PNqdCAYU9f37dYEAIKH+Iw3p/TmKGpvMCLJYykZKlM6byojxD13L2SGH12nxTe29
NS4yypfUNRntBnT67BNtK/58m7MBmFYQzagX9pj+ynr82YVTHh8B10/k5e52qq+d
3g63GKQ7Od5kPWtu+o3anQ==
`protect END_PROTECTED
