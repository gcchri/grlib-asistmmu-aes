`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bgqmepLzT6nfeazilH/898Pz7dqOQQEMg8EqdPyQ9cwXOfH6tMW4V8gxJ8G1ySFn
s+y0cPvX/W0UZc4fav47cXaog0uTr28R/jzPrcI0f6+JNyQ9olfCKrmn4itd6I4d
LFfwN6LbHGsB22HZdP3nyVunOVIwKQTTrZW4p0WPk1NrxhjobFRlvucbUeaeud50
RiM2CWyUsMkVfQLH74gSr3YkqXcgrEU5HFlS8oCMaMWybqHZC4wrW1tg7yh6zuNS
fesEgY//uKwf/Nq0dt9aJ2q648sgnMz+uZUEYMRL7hKqGumCVWvY+oQkp8dVwMO1
fYtl0dfG0jn8D4hf3L7/MCnAI4B84cYVVwHloZo6jWU7CRXTwORIe2djVIL73/VU
8mZJBUPj41UioJcHgNThIsLxPXgLa9j2vhbLIO/QZZkQefxue5TyiWOHf75tfvvh
NEi4KwWubjbpenirIbwrfL+PdBlcjy7W0WbX+bveGpbs6epmrUj3nrwsC1AzyY+r
vbs1t/TlkdX/sVLYrCh3seI5Kr2sQYN/rk7GYoq017+ooyku5fE3VyO9l21Zz+zY
yFvuSFkEeWyaMTZ7Q43MgawWD12FNWbyZhVWRp7FX/wDDsHGuCr2KJJuTtRgPkPo
gp9Vt6C/YH52yg+1EUw9V/zxYdLzC5vH2dS7fs7jWM6MtrOAt9TH2VXuH69/Mnh2
qZ4faYfZGh8yhee3xFydpwCKTr2zFeuBAgLRa8tYabaxWEuXj1DPHaBWIUdfQFcG
7O4xd0/Qs3e6KlbTkDPKnWLYShpKUi29c1k+3ODd+imKAE/YJ9pmJmsAEs9+1gWo
IPcz+1TmnUo0oorAVpACenoVpZirKc0Nmc3xtFMSgGMZCU5eBFPyMLZag/aPxbOW
4qsjegewljQjFo+Ln5UwJTjlY5scT9h6wazeXzKKVLbwPKSrQlf0EtXPj0oHqtiw
3dsoEqXBaUIIjnDwqiVC/Xb9zesxVqsrmY9uVtO3avyZyOnddoeydjy1/5kwFyvA
CDkFf6eNNViIbnJPQZedMD5zUoglLYC4SefUrFhia8gynxpayAR01wVHJj5wsnR0
wSVb9zUeQNEnBGzW0hLI/36ynA02eNmgL+xCP+l8c8g3EhayfCYkjP1CPO3QGuBB
5R5p5dSqBTgXos6FGwOCLgjFZvzNqp1jtXSpNihK/ieNt6/tK7OcYCA9SuEN8h8Y
6SukfViz5npU47B1gxuHkW933S4fUwg6+/gscpxPnXjd603b0gghAM63hkraDW+4
OqUQZoZf0HZZlBLFSYFNeQk5GdUhxrIF9F92YdBi1GyLAxlFik6tVbrMbv6jO9XY
UgNE4yUVnpJbihZIjMC3UGOEdVuA55sS+NJps1iv1toPV86I2v7EHBln2ZfeGPlZ
gUd5/+9miPKu0+DjqEkxEynhcFddXxM8QNu2aFo1JIhsi5yso1bf1Higa7Bh9uON
hptNO6+ieGi9pWfDx75SIeltEd6W5DDwXha3HPt+TAwPPER+XizkrzQrpjiL6VVW
7NlGoGVwKHDcJM403v8Poyy7u+WVjan0Gdfp9BTDgF7Ltghbw/7u1SF/lL2ne0mc
NrmcvLp4E7/uJsgCj7iHA3eJ5fZzUF+WFSZ0KERDSI1saZu4rCFpvT19j7hOZfWt
6xxZ+tb5UVXuzbl/WfdJlRRuiHjj92JmGV2uDgBn4WwxnOiFED4MNO9BR3rMzBxb
xMcM2Q2uigD8UqOCANcguqM6qnNECm7113Aww2RB/IHUCGuU23391RpH4E7ISDzn
E1xrfLQKvZNVS0aR6sGsg52CTQUXZXhAzRxGh9mQnV90D+7cNyNgCpiHPfshQW7Y
6sZvQ65DfdcFbkaeQZ4llMicmRMttaN6CR+D0KeVp/uH0/DwVrve8vgrfTZNxgYd
LY9jfbSYMb2W8yADo2+Fxteo9LZ6EWKGgtu8Bo/UthIhBGZCd9Q+epRrH8TkSNxD
2EV64d0v/IgSlml6UlxllnUUjSFcOeGeSyawcvLpPpNUL0xXJmhIgTBiB4/bB2nc
CSc7ulIU6ebauCC91xHkLVQd09WE4xb6nhROev1ywz2zhJ5qvMolgwxdqZeQSdaA
PHTNF1kdoCE/p49nyuqtm/hlLNFjsjb6D96jVjfXhgmFavhu5wtpmCFc1kD1uO9T
StxkTsZuWMhhPeZAoQdvfeGB3mWDEA3J0hWAgJMFeETlZs1icokuVOxboN4A0QkC
U3MGUSrt3FOqczNShh01kKiZFw6dgFcwIP9PdYlyBHmOSPBE7dgOTVqIRLhvQ1/w
WtEGozEDlmzvWdczUaCizB/tt84gcIPVZQtGnGHusIoATOpTXP34qrbJCjl7pOSV
awN6U0gXNyXPHTrMo4wmUGq423d3VxFOzHz5ZjwSIYO3Kp81jgbgA21ITJtG0caa
R39psx0Ii0Aa84hLPTkEldn/aM5GVHyZH7oBH5OChPhcvBXt87ZB6RFfdq/I96WR
22B6d93Q9RTIp2Ns/I15YNRFfxgTyWpo6gXMXZf9eXY4DB4Dii+EJSanr2JJQ966
+5O88dFDVlGoTqbOesYLjvFGDTq6oojYu4+nDdfrEzgERcEQ1b8BRodHXScuE689
7Jsr0o8XAi6dA+4cVkn/njfY54mgQpu24/0XeRRT5tUtaSRbdwvL6BzsLprolZVC
3cwmU7orSax1FY0a1RnBWVRYLCAnkfaFbPVnrvv4qF3BXVR04LbkZIhy7uf3dHc4
bOFDzIUHl+N1/hW8ROimCBar/s8zz7X6nJQsQwupRjCVMUz8HS3yI0Ux0Kmn1e8R
INyrfLm29ygfjkqgoTSLulp56pP3HY0qkHjJVQdKv7gDwnAebOa4Xm0goH+8oQbK
mD+us/n7wPNx66N4Byjpur3wLD6D1deVmxHJQVDHzkKtdWIlApRT4DipH90HX4D3
Pruh8ZQVbWYEo+TDFnby13yRHcqyGaJmL76w8UAamJo2cyW81FJspsBRIhHODc8B
XX6nmB95mgQjHbCbRl+oOMKHnVTTGXmd3Rpju74vm9mU6t9dW6ddO5uYH01uu1pA
MCuuKvZJljj8ZTdw2ReOOfr6Y7eg9Q4nq/0EDeJdrNiE0mwNvNteu1rRG7rOuAx8
y0ilaIPViRjFfDs5+3X90B/LGwyP82VPbr1fNJojVohRLEprmNocz8KsNthVv0WT
1vTpjZYnbtLhY6P54Da8WtsNPX76+NW9DcHZ9AX1jfqRYwa/MrL7oVmAgbUHDOXH
xbtX8OTgGaqhW8iR0xWoB8FEu+EcC2C1XCZjfs6y3g8nytHRVZxThMtPWjmCf3Vx
Z84s5uqyY2kzrRFyZqq8xKZU7tRTf9nsgepM8mEFV0faJ+mtxbsKpqppTlrMXKwF
bKn4PGUDYScZE0iwcIs+Nzv0crxIbSfDxAowJKpheBUkCRJ9Q1CHSS+4jmrbsCut
TUUjMqgcuRuumshvSBTDEFzXv9L7Y8aDx/FyTgsRqSc2pg5udUO6/rGSHbJOagjo
5ioHwSYifcBpP4Pwjc166xSRWxl0aJ39cCRYRy1cXngjg/Mkuf/5+Kku2LWzh5xf
NS0XvVIz39/ru0BaSItpfdizB6exx6C3kc9gK+cf8ez4lGqfEVhaIzBHfqGTyGZm
GAjkxpBxhglAay6Bo8t1BaX8PZhgB4hlWLXB1xu/wf31BWqwRHgs7T+hUOLKbTaZ
LhozT7EHBR5ZgctGqcag4hQQokfg4b5q6VT2XqqDre9BXTgh0D5zNru8xDLW6+lP
vnHU14G4DUnNtXTifJCvXoY5DC7bcohpCe7/FL0uUJZrrH850sMbO8AQj2xLkJIF
VNSTsOH8IkKzc6RVNdZZkM1T8d788tJXg+1m3d7TWPIWWR8bWd/HTPEgAkKv/YK+
kNZmUc0q5MzfWeoXfOc1lAYUW33BSStS6o68omsVrURVJhMNatI0ksaSrL1YgBd1
hvgIGxb2orhJ4jqTdSll0+24Pzz9lk2dcMbIYwSirGMGozMQJ0/fusAzLq2sieQ0
UOZOENmgiJ/gRXGVHOoRl9t1z4R8NAFQwG+ATvhT63wnVyIStgCnUzhrmLW8XAS8
GiiN0lOK12khEAaMCFqy73FXnY8yRBnOaAxuVkvOFNmbNSGy5EBkxJzBatdm7aeg
uEpSm9qCNlUQBsXo1NYrkXE5evzVq34QHLPQT35v86woM0GU9j63Qk665ol1hyFw
laf3EhNuYWAykJ2KbU75RGC4Q9pa2n3FKrQhkXu8XddiZuRPEs8SgVUDyjWjQci6
rW/2yoWi48syPr9Ny5zxkgh1h8sG9LFVpIWiUI2y1tLFp1GDvEqaNVMuinJfuwBz
fE/jtKpvWZ3cwj70228IqEFMfeKJup0xeOcfH+2Sxt31iXVuvOjKppsi9JJh4nY5
VqwvBLw7oILcfUqqFaMzS0Fow+HY6j8e1k8c75CYw47Y8NohRiLCigUIHfZRILc1
3SmXkDfDVhktBzlb7pteIg+bBkA2A+fCX9H+SvIXqn5uH5y+inyu0iYRlDZMkaMt
DxmdeS6eA9vSN0Y7iS49LNtiNTN2jEjoPqq3/9P6AJs4BG58FKVqU2TQxHXZQFpv
EWKBevw+L/gFKY29JZ1v8ul8ZryToY3EVzqNQdvZx88Ot3hZfp/rp97Lx/lNeXjg
NXg6lbe1s2pu58UZtnufUlFfEvZC2EM0Ul9Df8end+M9b3VrL6RaEDB3MKov5SbK
JM/imRzhXZKkklUxbqK4GF2EdMKegIb6lLHQJbxlrs+SvJVe1BfDGeL4KQ8CeMxt
H3X85Ah+cabG+nj89ZEJhcV0RZaBYjXoJPeuRKiT7ZPHHvvPHyj4b7U9ZiOYdSy0
v8lduy7MyFAS2jM8mvX5qBS9hxIc64MOKS0vU5f17CpR/gmk4YIxlZg72HPpE0bl
SwrbEGf4xqPGSMcQtPc9rBwfw9kT+FoUr654P/P/bxZ8vr7PdxFNwktBzvTXjWkC
UkCne0eEDPPmbv5kZs5Drfcd0nxmrv7uZcYG0C32EZrEZQjh4IRyBFKbdbvAvfOT
/z4AhRsJpeCyo2V2pGLZdzK3yR4cyIuiRl20uGZcHhjtf8rHWin0G82gIzBa7tZe
QREoBBeNo3q41mmb/eFh6vp3x/hn0wolalmf6Lfz31zOAYryhxnCsjGSftia4v+X
lmmC/0ufiN+9MIEyaIoyGm9yRViaZs+R5+hUralJGCHd0+vHeMIlZFf0yrIy3eTv
8AeFqIZl5+X198GXLpO/yDOJHzujp3knopvXTB+gqUWK7/6K+oP54/UaGhYqwU/2
0oI1pnSr/g10FwOWHHkVq10yQXCQ8pAKYuY5odJkJArFJVGFAVT6mHGFqn3k9ktN
GPGBEhblZSKaFYjAoVqRtnNViy2ZCaaUgUlak2it4LhVkeHTxZYV5EgOzoooPV73
lBak5tExaFF6RvSCtPx8DplN4Cp2B5yJ5MmY7Nrl9VkK6Ijjv9EFNim0bM5fWr4f
VIqZBrBeJjblNoQHTPt/ODsSEuBBTHAlY9ZU/f53IQkJrpSENeO5/qj/BQtRiVuz
HHbs48qIciCmlWhlLJitQn1ZushG6+0Q1HhfDHtT4AxzVO8ijuA+6exNRrx1EzfK
6xHVKv8ua/PvIOWNBVywV3Qkvy2TaGxWWMvS9XLMkCV13Vji94qVeKukliP9n+6P
hYnEwD0AbwyGTgOYYzThWBvGQJMbvxzR34T9dVrieJteWOcIdZhEYtHuv8NufSa5
9c0Fa7RLemd0yidAgrYw6K+KTaPLZxzMVUC4NLokS2L7Tcuv6ktpEYL99bdYI+IQ
fnsKjvRL9Y+JAyEvjYP4PaMtPpjtuTMIqfMFnA+trpyb+7othsd72sJzqhy5eifJ
Z+of43QUU4ZIj5SwAxjVYDjfjmHy22kAvDwszkowFCyTGrH4Jd0wmvDW28wfzWNG
94i0gMLMNsaD5oPU57hF+8AJeK4cS6xEd+TbQOva5fMyBxwL+tYttpIuFip/FjCG
K0HmQobNhtcPlprHuuRkqVhIrnhCYUT4OFSwc0slrkXw2k9o1pNtagMPBhEUvmTP
wZ6oiXAmRSmxf+iogelt3vQH28wKEgWG8uJNosxLHToU9UiztHwA5DfeLwcrI5d7
9ZU3OQ5ZXF1yLo6SKIC6X66lDrVg/4rxurZPKgjI6co8VwEQlQF/4xXgop0K4bLp
9QArPDEw4YWFfADl7XgnlZWr3HOszgbsnoIW4N7OuzwY7uzV3zY0dXN6z/uxifeX
6M2wTRe390mZ3NXkUq9ARlWakd7xro4ZYu1K0MUbaNzhPBHyyxPpv5JDEB9d1tAq
Aw7fHT+maGHOzXUbfOsKVciAQfCF/XTVf/XOwtVQ+uoy7/+aKIzZMxSlKxFL4PAk
XNAviFBhtTFKjJnV3Lqk7ENY59xjgpwm7BOg/n2wLdL9+mIJGM3FoWRJQ9ovARe+
Z2jCD69+CB8TAKQvGSzaJ3uEDzHAEvMtinFKwJ33lUcjFO4SzS+o5eEW0/FNKQ26
FI7iovFIlVTMylNP5QHzHcVzf9L8u8ce/2QZmmBPwZOzuvhn/FjxDlrb+nrsijTg
8Uuc3EkRqip7ew+BYUqVGqPwWNey+DSvPSPuVcYvQBHnCkYnIUraIqUXdV1W8FN+
wamVry5CVWci3T40K3LxGFfWbUMGR3Bv/+oFI8YWlcL++rmOHcLZqjvsbBt1w0Ki
DtGLg1pdu+mj0WWJF5dn+GSpUcWEUWEl/vNsB/Sqfc3HXLJB4LrdU9sLompGhrd/
iYMhwlJ5wKTSh3uG6mkBMwrBh4Q7dvG6MVcN8a3L6m+G3BYC2hyJ0Og5MmQYC0xp
sReR+MGiMgi87jivow0RWf+ndB86jphshkxFNd7WRNyQkhQ/6IVpS5pw8aTwSf3I
qIBOX9cmYmjnshBLSfXBdWfV45oUyF86D59zFcNK3/WmetAK7TbIV079skMc/Mc2
Yc4lb8iChGZumTfjy60Hm+hzAjr7bLEZXKBHKb2PfDhQVXWfez0Xwn3TsnHQQVYM
3qRpeyuYR3gPn79n++m8amuoSCSbMQ9nnM6Lo8BBIQnY5tuQ05xlVMe5WKVmvPgc
M1bJeJDSLm0lfa7g9/npf/BE9kmAO4+OKeL85w6BcWu/WZjTVpb6yeLSwI1uuPir
MGzA/jp0UsO+mtPdT838jqxEBFLuVHUDb05IDb2exyrzhtHYQIJ9hwDCW+HgnAwM
4i3C9mE1IoZh72QaF8dpBk2uSEW4+Yi9ptWCoewwP6xt+zX8TLjoTwA/tebwW0EN
zZU5lWjWAUBBGzDjzCpu2qdF1WNtZUaGuPYSSar1bbuvqlsKVVNTp/95xRpawm62
5ceGXfqHR1hyQuwpkcsFx1iupjul5f1IcCnxldeQGhLkRbrI0a6/pD4PbIZKlJII
fekoiKlJTWZlG3cB720iI+dR/f6IQcQyT82HQnWH8M5Javr4nUEekSvCgFQMZalp
vJq/s7oQo3PPlgj36Y3B7jHN0etQARSh4Haz5iqmGNwj3mw+VxVU0crS1NmzK2pw
pysZRgaLI5poymeHphhX/peL7Sjwry4QqTBO0O+fPSkL3IRgfA9AgXoiZwCUkNou
qpeSwl/946XJKlOpkW+HYTeoxiVNiPFrpcYodkJB1zkZ1aiDjlXoe4hQBkEpRFv7
c/MZiAHbm92FQdweJjOvhH24DAKGikRkVZH/MGcgHGGBv0ybOKGWkfmN0DEf8KAt
jj5hcf08SeGXZPFjO6cEm3nsVsZNsQC1xD8C7o9oXF5u2zi+NQgifCW50jp7Nsmy
ByUnX7aLl0oEkZgZqmmi/mGEDjNm4MDwPW7ou+A5147LU95P6bgr0smQr1hRmpMN
B13OA7eCoZhV1YpUIukK1OXYut5l50+1tAeVxIvmIPElcDmKJbt67+Dv/FJ6Gf97
xtO/zsxBCXT9/R8yynONSRDJEFkkc4SVZHI7e/jrtF0J+jaW0nwqz9NsMFIHWyLM
u8VFwRWzJcQaelHZMC5lNGM94Kd4Mx5EltlxX6sn26Zln5PlldI0d4SVBUDXjgLB
c9NV0pu2VbjW3g0fh2yU1pRRmIC7N7wpFsXjWBX8m1XCZi8Fn3/NmiVoR1u4CrGU
twZznQgdMztypX0GFmOOjODo7lrXHiRxjroUpxvbBPvAcMbCkX62lEsWCHc0iTHQ
TppZUhKnSyH6C+AuVl2rQvJKH/LtHs7CUL1c3MqqyATVoQyI2wqH7qa7l1c/QGNa
rbi3ulYt6LSLADS+9mGNWOQGMt8g18yK3tmupxihp62WSyBV/paVL4s4Z5fNUlky
lgBM7mIoP0pR10RNV5JcAe6zkpx8Gd+QoMf9bMXt4K4iiWmieOweM/y+pwHxioUh
e94qhxmxWmSjZoqSePyPuneneHZEpIp+S2N6sDPnt5Fj6EHzE+UWXAnFMsb4lCpg
qdLE43H4QFhirIrh+X8BshRm7XP6WxTtKWiLu79cWewLV86yc63QwAt3WSAzwQQc
9uixD50A9LmkLdndsribN8AmDaVKrt5w1V7ZpTMTxPrToBAp02RVp+OgRyswbCEC
fKYY2jqTfYJJNDLazfzAqNmZ+nMP002Ydb6WDM0NL72GSTI7qj3PFNJo/H3RTL4N
tLk0Dznks2x/9CSgGlccMIugc05JDCMsNJuBVhXcAN2x7nZv4OrX2WxTlv3LGxqn
jyreF2M4hNIGa8EYdc93PoSwY/xQVvprY0cFYqJVRn7q9jOhx9lH1yaAY4bVS742
xVI+hNeAWC/SIFeu6JFX1ZcHeJGYCkh7O4CjN3n+CyzeitXIvj5kLpq2DVYJol0S
I2IxB5d9c6MU+hMhpzQZBiZE1quPytwtXeOIT/veHSgJUXmt/QQoWN8QdMVl8O5Y
zb07zUaaTFNu828astObjFsHoqC/U8HC3wouOGHb0Mhe46wNnKBOIzXmvfPjlRyG
FySW4mEo8jmFv93/v+/Yxjv/O764/p2CbwyC8sH1PmqzJZV4n21ZmR+mIW94GKOr
HqlArXLLGYeHjPSAOB03BarwogZb6slBDIIttSHILuP8QIpn+/jeXDZRdbzQ9GVg
RTW7/LZ1YXh050poTeC9WSE/L2xGXUtrmjowK20XAUjyCpUX7zSEv48c8EZct4+W
9WGESVb2DMzPXb/5jBv2VxAx/DFRvK8W31aDcwirD+G0IixSLz30GVcbAjFdUWS9
9bHGukjL6xvvqlWijAmEqJzEq2I44DDik9k60iumxuZCNsnzjmvYqL4XW4AIaMVZ
VJqsRdqwfAEneBpvnuaaoBLavBz57kzukkxyRnytIQqzUWXRqBDD0Xqw4AdYyb0r
oknph7Txx12wVfVXfYCaXcRzJT/E6H/IFiZI5tkMOacb6V3+aUaEHQu6pZIMRR86
Ukn/ntaD9vwZtrnw2LPVlBLTyNi+7CIWEHSkBPajXsj+tI3CIWlHccVexYW6XC9W
yQJuk+ARw1ADAb3yexG+YrqU+oUtNLO05jWetsRQhpHnQBLGzlt7e1rAgoYwMJuo
4gx9RI7WBSzkilZWvU5JUWi1aXSlBe0adD8OJgMtNRzWm3g/4zWvUbiBwCPDAQW2
8wSV2QkTAOqP3H5FmxfcIElUB8a/V2NuHSZLrxxRMP0mF9uMvH8jTzHl3/swBrIO
nQyvoyMZ+gq0JLKIKpCSiLGUYHKvjSLY2gdBnDwaPgPuoqPv7crT0KQqWdJLYdXV
zvoyovLyXJs0hkuONZNdF0e5LUtEXwU0lUX+2I4IuFdprmaA+Wd7bDsWA0RSfMD6
FrntKoFO5YBvAaU92gcx3XN89tF5q2FunG/wu66/8m2S9s4gv0ChXMBfPkJyXSHq
YT8j10IIuGJ5BVx2lZfDlFE+41DLy/EmGPgbG3EbJkEEQOq1hTJTeIXl1il6tunC
NAGXCFsNJzhaJSb3QKyOjI/B1DNAv9sOJNVgsu7moqspYGsrMeAXtVU0r4FSjnNT
KZZ/E3Rt1S7mLjaCgyJf3zV7JQb0A25VTKqxIKtzeFNoWKcJ+g3ZbCuUf6JRPL5D
dVx4Crxuab8MV0UyRLWjHvQp+Rsj9vGScv+/u5TqMMbcZ23Wyc8dVpogPQiTVGHq
oS7wgPf9JOopfRzxXeWyLowx/e+Nf9I3A/G9FaWVA24SCYUXmj3i0+yTH3gbYkjm
9mJve5s0NklU29Ghl5lD1s3uxxXPscWXbUPwlYRl2bZMA06SiME60yOfj1xioS0Z
8hJZ6yiwRsk/FTWrRCPu7twYyZzv4gAU7ywIIC45n6uVBJTepj5ENbhamyf4HAQu
nQ7wgToxVCjBavFXYaIX7v7zoDquKpF/Kk7qFJEuM5oCz5LPHhFl+pdy+QU2Aa7H
NueTob4MafDuqN9wV96gnEj27yLOWKV2fmu3DcjgpHdEkPXWGlvzmhn6BzNCZE09
Pqh0loMWxFPZ2xV3n3qZ2vVtT6qmHgpQjXMSvY0l+NrVRLfgw8pZLSC4q+iUTR0d
02ZnRVDRPGCTpSLvj8lX2Fd8ajPdzZlvgG/8mB0hEG6RNFS4iM4TJiieOZsBVOFA
MuUFkGmCihla0huB8le2gXt56YkfqqtjFiI7MIhgkCBW5BYhA2e7ZaxShQgRmX08
QBDMscIm5hdivZQRqm8x8cB0E2tYUDNkDtdu4ukAqGEoevnijlkZPHKNW+MXeIwC
y328n3yG8D24e2vd14H6j0KM+O1NqBOkx+JsJ3kBtw4ygpCdoB5YASLkEFEeziZA
5Ct+IWyrIAtxeey9qncjNAC50l8ohidsAN619C10rtl3eeE7mgI0eIqIgRsOofla
irM+9/N2ub0LamE69bEjDk7EjIzhRtAz9hGrvxhzaeNeeTG5/HHUOoHjDZ+u13/g
3aJLyD+e5QL+UBCOydsD4ZGnkoRKYgFz58o3fbNV/2KLx3nrYeFhKhO4VyLoRjos
8eS/7Lz8oiSlo0QyTRPk/oAPUCm+rLcr6RMWak2aj+1//7JIW6Y65ir/60h5jH2s
hBpksLGmz7U+/974WGQEu5kNEuAfvmINnA6PAAwIh8+oO9drYkP0WlR+AmascTB0
/PDBMKzDY/ulfPjV2m9ckAhJ4C3/l1/F/9y+AhZ6QPWSvWQ/nSHJOx68VZOJOwCM
hOTVWLoid0WblkR338CNENzIXcA3oz1xaMT1tmObE7DSQthUvp9E0SgF16DE04fB
KUZJSjBwRDhJ/ZRs9WJRXwi21YyS728OboucT3vZx+E9VgaPoY+0Dg0yiWSfEx9/
AaIS33elTLGcpsMCQWskp7Ns8uqdBC9lxUsvt8Mj9wyNk+bGdYJIjXCke9kQJJrS
a1AZTMkVAZvZ9Vh0HBeRzx0O/qGY54tjcBXhXfR7g+zSaT6jWHkm1JqUweBf36Yo
NSt3A/NfYmH+GdBFvhx+N10Sl4kZc9J+X4jxxW3ftH8/jZlaBNUG7EoBED2zhOJ4
Hhp7QrB77whIOfO9feFjeDPRT+w1YvQxxcMQVB3gb17ZluZ9TWBDIDYKUKDvnt5D
jhndK3qV2mmPzwwzr14YPOUGv1xRc+D3+fCLBflbac9BFmsxS3ooYbOdJQt5rirS
5026Jr+S3QomI+IjWLVn57/qDwk0It4lBcKGL+fPQKFqwpXalDZKUdDye1iJeh//
nvHcJjIVgorbKKKmcgMYzcusEXnPKp3BBg5SFh6REZxQaqgKltLIEohbu+PM9odB
rhvuFYhfQzLTdF7FzUC4sUUqVtgWiDbARu3MMmK2aAqJvtSbCWd0NssFouM0hYdV
DPkD1IuL2uO7irFwmPggKWhE7TiYqhQKIxWoZJG0KXsMcwAG6lWwgqPAMbnZkAos
xpfb7+pEHuuNTwf0YEbazpTr81yadkMziuAzt/KK8l9NoNy5vqJHAqN9tnVhYuD6
kn9LcNxq2nSd0DcdB0s90//RoHoW2sQbgnDu2N6/ETHqprO6SBk08jwJmT4bnnRo
jSS1M8MjPB3amsdSr8+2ADqD763QNa6SqNlBLpXggwP9osmbp7CSpgJNdD6nsIiz
mBWTbPkLkEcqAlyhaTf9fQmcP2tf04sEcXuxmvKM6JUOYQZOqkxn2ZQB8wqjccs1
xMWHwaYhk4kYh1mgcYs+1wz+02BgWccmQqXrqcM5+1QHS5g9YoujV/CjdaetkBZI
rPchK5peIKPYlZxCePhFDQp2EvzVXrkpyP6yOztRcECnuttu7914NhGatBlM+z+0
5XuNizfSyK2Jqe4xjJTsqwXs8QGioqEau3DqtL+whmo12vMnbAFw3JcYgRzwfJpC
AFW3lJM2lRYpaw47Fi9x5XMSadTeu6AIfuXowzCELtAEeg6FjjlyGMAX/+cFBl4Z
7IoVpUny9S161Suw4o3hh5+T7n8tnuH+xkIHkl9VCP4P7PmE+aQVMYW6nVFh+kfH
VgoggfO23N6VviU/cSsld9lRqcXRAs6o2lY0K0C75QB7H5/APfLin04PeqAl1KE5
gIu0oTGaBbO8ViTk61YheXEMVHRCVuRoG5JtWj9zubhEJB9SKqHzh0B+ulMwz2b6
whkF5ooBCul0e/w2oXYXPE+aqj1UgHcScuaeWCKiE8nzd51/4dNT3hS53g8s9W9T
5N2JaZ3rQJSmTFKHE0EHPulRY7+DpTTvv+HX6tijlB9HfDf9Mj3+MKgcdWcj8Vu0
qiufX/Zh4ZkGCSJs39TRS+lSnPg/ddIgi1uocNYhyoGMSxS5Jubu4mps0ngcsKfV
CnDz9KuWdSUF5AA90pPydQXUxvCC5WsnUKEqxgcfbNyG5wlMw5LNBaCa5V4q4tx2
+U01vcej7h2oNl1ViTk7GjJW4nvf5gRe1V58qKR3oIkr0IhHuy0Ost/O2zikWlqs
NF2sL7StMYZHMzuPG1Hi/XHIGLoAo58cmBsLwmNHFgHuNqPbUvMQdUuKrwsU1AIz
Kk6/la0H295uhgI7EVzCsodrzK60lnx1d4lSGmjOi6U703tEBZhZpdzqWA8Ryu5s
AH2ojeo1MXGNThhJmZJ9kXK+WVgLkcDZqg63eH9dHSHKv8pf2G0/+SoHoGidq7TF
hT+UKvSsYCQ3kcsRZCwd1y2iwDzvwut91dsNRl+/7s4wKIzZoyvL322BfTnaY+Ug
/4XiFXM/NqVAw1QmN+7gwhaz8WtY9GuybX/PGDjU9jsm3xkIa1VhdL3HVW0KzSLt
Xg7ftn14u81ZyjlhQJbM2yKvu8ygn8zWbhTCfqMVjZ87YtwpHPup104yg378pOst
5ZGbFsJdEp+wYqy3bohxBxEKK77BQ1Od9lNcq4er8CdmuohiS3fNCWG7lP9kubKd
5Vs3HTozlQ/CVNBI5vGUa8hoTf11Iwz8N7vgZzjCOH9b4sG8U5+w+byIG7stkngt
d12B0g/uY1xApYJcjBDWZuD85woHF1OWR4vZGxqtkMUgGM7f0qvEyxmMrdDbOz6y
20BmgA9fQMH9tnWst2k2p32qzNTHKeY+he5G9Oyi1ql5A2zY/R7yW+3e/lXeUKX+
qeDUjsWwrJ+tpwWo2e2cIoFUEmyRV5zTj9McnJk71nzsJJ+JpdcaN2ai00T0B4yu
xdDvk4CRYEb4dQpKedFgMUVQ0eYHDBi1frggp437bsWut8zOj8iGKXL4C2mTXi0j
SG9OzwJynhGg1v6qUSMshXye7son8LElbC3flbWZDHs4F8suB6+YZy+hgJ5accf8
NsBtWsCYygG9BXxYs6QUdwuFmyD3YzCmuYvA+6cBpaP6LAcmgBctYYe5WJh6s7H6
hzABC4Dqrf0ODN//pM0MvcA6SQUT70iVsxfIKhJhkuj3S9s1OPSkfq/tzzwOzmYL
/+WCPu+X5l9I3ywYn1/vswsjVbwDfduYHwf5dpmMiuySFcqLurTAdoC7ytcj+jVg
TNci+Ls5cCRDybSnWGBPx23EkFuNdM96pC1BGgLlxN4yWkLR/cItLLQSBCv3mnWU
R8ZOxzgQ3Q/pb/Qb521EX3NcZ4ueSXK2TmeANTgLs//RqJ9bmP9a9v+Mhkf55jcl
Q0HVdDtsGR5+WLC4Dj8PvR0HLdISJ3ZguGENGhQZtEQI+iS6BtkQq8fNajaZWhOo
eCH6LJto6IoJ6F/cKTZVwYjuEEspqlPJrLfKRxOKkaGx3ftUdHOSpptcQgJhifaZ
grhGAUMAqLdLxNFx/4FawQzWbkB97TSBa1hyjCAwgU1wEy1BvGJOduOvWMV0ummD
rZMW4awyvYp4bdmh4TK5TWFwe9mFk9XaPvgJiONf97pO068EytMJP8LmI3dtVZ0b
VFjj14HgoK0nQ2bvQ9TlHAdh8LvX6SUSnb9FBy+aUJ+Pum1q4Blcagqmn9P6P6Is
5+DIXi1BqUYgg/yzcM1rSdxSbwmdICutQzcjnuz83dMVlrNDxu5cCINz8zR9OKvU
fiFdyb5jRuPeLFkGo/uXZr7igkjO74NFvCYofgPIvCayDJZLmbggE0FWUzUFApHk
MQtOYE7wHLRIKpjt5dGZCsIP3kvtl8ngLiV/Yp4xYCwnp1QVV5Iho7A9wElpptfe
Vjdyai24OgoqNTjASni//rDTnz0Pe03tbdDn/6+YZdZHHndNmxHRVyJwcSXnweSj
JOgUiFr9e0NpN/zyhTp/8GpjFMzCowgB/wQdPh0E9J9YfrvZwDk0ee8r3RYilj1K
wP7jotEv/ewmhv4e/Ywsny5j5+a0jXiwc19Jp26D5u7NTwiduvOQJayV2nvM3v3q
EYUeLZA+DaM9f+cB656QCzcmxOkRPpP5FvVuGTk++wLlmpkuQlpxapD63dK8eE8a
38l8bjK7qIwv0lg+zocPv7mNZ7TxlDnvfZ4C5yU5H7b/L/Isk2GY5LP0Y134nDIl
XEHKa9RWt87q96GkzoTFhiOkO9Ky91O4mn263T5M7Rz1sVJyZ22lFe/0vkLHeBQf
yxj6jdLu0ZK3jHmjx3qah1+d/hh27vTJnuoOPp9LUDBP56YZmE/kZM7OsOsP0OW7
Ghu2l1Q0YZ/2upVqgKlbqctQ0M4ano121nl7jCIy45VSm+wkPRiSYtFavrYtqedV
SwGBtKfYQDiH92QZD72lVVXOPFTNm5nSe1IX0mK8sItJJUJ0vIedm1SmbvXTKnsp
xM4ElSmT4IL3Q906PQU1SZkn2OnoyHXK3/q1bQERgBkaUcZHv+FSXft768s+jCiv
vLm47SGf9FhJOxvXlgSJvLRXT+COs3j9/OQSJz5v4uioJMEYgowxBPrsZMlZy1/A
YEw4Sl/p/BWLkvmvBdqYhlj84/jsx8Fq7eAVo+49glrapUxFvsuYPrZkyyoaemVs
+Yqb0yHyHnCkbpj0sFQAOP1xtSFc6EvwBSd0Nnq1wCVY2MxCX1aRgc4DKFx/9No0
M6bCNXv/q/axWVx+sVh+klgA9gD1S8T4zs3wGy5F/T5rUSW2sNB0F4/+PBYgc9Wc
/SU2SwfJAFuJg2whuCy6gMs7cWmvH1gTD9O2ENZ5hcv2Huj7JUIxsIuiX16Z+4Rd
X+1llNz16wYaQY6eywUQ8OZXlSFJfA48SY7m+SP7iG4eqTChJCrCXaGAyHyW5bmx
SaJ3IXAP3PGJ1bMgA1HjYawJ6ZV3Gn/t3mbhzunYCNVAV9XgCsYfnO7w5myKd0/U
DObKucCdQi5ZM6hpugYlfBRelwOx87iLyioDZYyyV5rSnijv1Nb2EBx2809nVL+2
TYgLbiM2Symoz2CpTuD+RshuDF0PawvDSnFJpiIi8E6vIOjgR0I8q7WM5bIiDAPk
OVf7QojHWhqNL5PRQ/CRvR0db8VohkpYg8+IEYia0zP7k4LOifK/vYtNV2ACyspJ
Gi2KLVRE8T6zJkZYOMKiNYQSb3XapTwnhcoykKI+85RMkvi98kapfMwh6xX/9gsP
TDv4RQqzzsU5BLXN4kbdvr8mdTQJLGI8DAeF7VU+8rta9cYAZpoy0dPTE9bFxyVO
1vJygetDarqoxbgsqbj6LexZ4eZ+/BSzTORjXFyaJTA7gRu744gtv9AjZUwalIEz
U3tB1djIHFP/EuydEK/nBzDRJ3hfNBicJtSMNzx09UJra03ASgVcu0ETNIjsU8kM
a7+UEbA2yTOovwFRCfeAcC/0OkaBz4thp6hOyTw5zBr2RZ5fMGT5nN4PaRB0emMF
UQsKVSZgfReo6gxosKpp8+TWbB9n7nDFM40IdOUTo4u6mLqYyiSfDIur7A2q3zgJ
p2WQaLaA0UZaBvsIxMUf9lsCcMulfYx91D6K1/PYIZoKbDlCnKYu/NV+vQdC32Rp
2stIQ5Wa525xD7tB7RB/F7T0UXIXquuq+IpmwMs3AaLVMioyRIOnzDVysmaSxq0z
3QcgEhk5URvKYakQi2DItuFvTmwajCBsRROOxgNJXUxHDqYGwIUV2Q116JT2YZyl
A2sBXbF2QgrAoTdgTRZhojJAToUCht3Sv5w1qWjq2/r97UVdAPjcCEDVGQpWAlmP
Hs6GLW6lowUZwzIhLrw0TpthBPnhtR8TjN4f1bEP+iTegYmvDqHwVcPy6qXG6VLV
fWEg8uxiaodjOkYCBH6TLN/CU8OxO2o3eIUKTOazuhinT65jMXzp0lXGYf0tBr1E
+61j2tcdPWCPhsLlUq3SRjJyLE3RcupMdEHVURyNW1lTnVlUjHuxoG9hvp1mbmIa
dGRO6VAvK6LFbzL8tQJ/9CXL89XRkV9ig9dAXeX4E+JTDbBhaVNkOMGPF1MSpAC0
zo6hySM5LVTOXIKNPXEaz8EGptXuFKlSYH0mkuNO3g4sXPhOdlX82vH4C4znpc2F
R4Qx0+HyzRPN39JmNaMgNv02X4daSnY/D6wP30b5C4I2vf9P1yGjf61CumDwbuOa
0XjiBEkX+U86UUhmm2CiV70EVBCL2leohV6d7GwRTYeU5eN/TVQQ9eeFEmllfbey
hLE3DCSM7+bY/d0dgc7R8SgH1Si4Aa3/q5O90R7Idv8uy8dXUNIHMFq3y60q0MKd
QpLvfkoQcK5finuK67IJmCEoq1B2dJCw4nU0Rfix29u2GLJ1FFcir6WkMt9Y+h5R
rRtPGHseJpB3Qibsp1xHeHISrwONk7KP6apFRZUflgeqS6+AXqNz+VFrJz/nOvUZ
ApvQia/UawYZSPOZHvS6PYn1jIVKVjtVXu0BTTYBXVMN13ziwwbZjC5jxYSkBoWe
BD5lCeREotko9idLyTIVqwW5ehPSyBCYGE5ADqTSCape8cvK4oJJEfsXLKVPVfUr
F0B78Hye1QpdGRca6h+pwR/X0msZbTHNHAmEQ9JAny99uGXs0Gtkjzs2Ia1pL37q
jg539vPl+WeEf4a15lUM3pu/xSDXbHxVLG3I5ZttLjs0T3/H1LnjhmEFgu2Iyr6L
J7X2lhEBQGplAcBH8VqeuULivlx2/P7K+YRnlYJ5Rvx6n0GFGsHOBb39mIPBZ+c+
AiKj7k+3OL/tlxpnFOiYzygH7FAP6IHMOTsnZRz1130=
`protect END_PROTECTED
