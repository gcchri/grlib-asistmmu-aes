`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
762L0iHftWPErmeDzikjshOdYHvcDuhdSyEBpMzbP/pOEKiKhNqUGqDPQ8hztA4f
Sew2OpRDcUUEnQFd+vmIVPpvLJ4uc06PzwEe4fO8VdWG8fa1AOjoYyAHMBflMEPH
0KKqYOJP/LyjJzHGKARYrpUn+3wxgPdNBBytmdWBJa1DVGE0bXP5OGlwD3L2FtzK
7IQZyIUdRpynVlwEWSdhImR6DvJJ5m02/lNm73b75c/SZ5I/bQQxax/MyuqOItGB
RcH5xJcuGSdy3IMytaEQkSFDpsqeI8R0zf8UwGZNENGVdiqHSYqk3cSTxHLPq2Hv
0ChVTOdDBDzn60kb63lM6I5GO8rPtajkmkq6Bemt/D8xsgJISgmw+oERc7yUmAOD
rmP7iS7VSyuoyqYZ34FGg6EhuL6SudLkhGcT465wMt95kSk8woYRFomq+YN2mmxa
78JcKp3NW/xsNj/Ve5LYve9Pj6WwQU0RL7Lxd4p1pLUgl2gUbuFriOeyd/ldqWNm
pz5RpF8553HPTCzx7cGdwWgtOX0ZBc7OiZc1e0FQWl31k6fnxa1ZS6yRXq0TlGPG
CM7mHbWDavr05UmRFpIJSitXfksz+H9bvmmXYz51so9d/L4iSO+nCM9TwuddCpPG
2MSQ8A8KT3TV+0ancM68g4biwBTtnQ1+z3BGzRgvUSzP3V+nJiMiD1wDqCEkgzTq
nnDXz7D92LOx229OcTqzQZPHcVWV1nEZqqNOhr+cdS5oMFFjDsQYrPOBFiMNsDA1
b1g3LYIIyxaO/DW1VhIToUra3lqeV0d4mlSlUfITX2ZL2UzNvv+V1GC1sZFP1W3H
K1TYV+K+wTrS0IkfplRuuQCnU2Rekk7V7nzvvyzk50wTh8Uyu5vmQvVO6wJKXs8c
9EsJg9IvNfgNyzRoPs/HtIzbEXzbm1RSQN6jyC6o58siRX+y0X07aKgt7jbvJf/P
xknwePYTosVyS8rousxTLRn+u57vAbNneR2cCLPELZRDWW7ZImVfzxxQZWeMyb/N
91z3FHfTrR/Hafmokx55+1+LyQliXs+3Q7S29rqOHFEvp5tCHzx8cEYs8KulzVET
lrDwrb3NGJNh2ZyvAaOF7UiTFrdNWhDSKncVtF1RbcQkubfcPeV/ydZLSnxAgxbA
Dk5EaH6s+jyXaHjvC7/T+hwW1FEbNmLqo19UPGyU1F5DT+HaF3XVlbx+ZYMXhJpR
3/QeATcqtraG+Msk3m4dtO+fvOU02Ws3A3w62eulE0mtyJPJNQW+R8OE3+Bs4ce+
zLZ3cPc00y21ZOsuaYoL8+ntoBm+rtklB3OhVfH/VpVyXY6iJH7R4K+FL0oxUphn
yxzQ2tlRX/cSWVjLWL2mE+Wf2JrtK5M/tFNytyLPM5B3nWE94Vnj6R6CRLNiqNHY
mWaqgaq1ZgpDO/wo0kQwMrBO3L6k+qKUNbPiGGVA9GEnJMkh+iDRKeH6JGPyeR/0
IU1OfUl09DWKsGyU29F3BVC0u7Z0MP1ZzaCbzE6SffoV6hOUOP6wgKpW0JoFUN3+
FwFL7MxIqZux9Y+EaJimXT3Wl2NlPHY8Xo1JzrGeYneWomL3o9r0V5LZkYTNZHAY
b4Hz3+dVrx+J7uj1ZAGVGPzgQXasXsWtenyl/ukN329c+fwI2Ae5xq1e/0AZIL1T
TVuQmLmCTWGqQ0q0vpSQaGDvjx5rB8tfYOSwAGoYWgnD8fzdRZo5cH1jEUwtFcZF
3JJ1iLSHn6/laR7tQuOdMghppLLV0EFeUGcLr7GU2Qq0IJX7X6BZhE2LWRcIo6dF
t+0hZGm7uTaiyAc+jahO2Ewvryf/vr3ELG9S2Av1IeBwaHGUdlx91OqEVF1bQb3u
Ybc+yTrChlHy07NI/wdzXw6ZeDBzp1eP4SQUJ9JFBiMgmevr8rUmQNO/ywjbXEvP
UBNKDVCyhkf4pbKWLaPHr+mLl9H2WuYef9pPmKQ3B8A7UeIJlHUTHYdu0qOjj2x7
jfGL+Z8uOh1iznd2PvYo1zdJTL8DeKJmnaMMjZ5b91EpFl/BdbODJGCxSKQAv1tZ
0jAKXqwlNZJ017sVih4+ym5BPcDC5nAjBTgFOKmX+YJz2D1Qk7sil0CNKYOD8v3e
Jm7QmjvJ5ect6tQEUySpCphxvKoPxB88CgH8n+wUlrWXkLEDcGaHe+v87WIGCel3
j2lByifg8QtRaPXtmFYXu/vE5lRAiqjF5Q2hQSxmogRfOFnqIFfYUok5RKNlN0+m
vZyoPhqqPHvyDMj9Jn3qyuQO3cskXgWOVT22Uo8YjMlI7HAbUPpmTYOWgNa7R9Ui
p7n4QxhxpepxQurCNBNL2FJ9TX95OoSvILn4Yy3fDGhXoDyYAT/TZgJuwqQ1xLx3
0/zRTlIfkyoYEhIhUQIIrExwUXFsAKI3JCk+Hw7Lydyu68q7XnWKEI1z1G3+PV5o
wPmEesOhX1S4knq284FNjVHhxrfin1GcB74K/p7kyZmeAeFzMEGZGAVQmxx+Q0of
Fi3l++RIiL2VV/CrIxznnxYvTXOAyQNxDd2t6ztwHCxnlQJGXTX+Awmw4Y0QF1NL
APSC/RKCkEJeq6/kibUrDq1r1uge1SlXP2R61qrXlDJWDAWoTTpLmd+w7FbZaqiD
9EUCJAFFO9RaTtwheoQGIaUV20cgrpnC/Z7lnWWgLWzWqpcWHoS9rv3CH6kklc97
ACHSFX1XxxX9zNBT1mTIVKMFHncc1z7SaQIl5XAt1JdoU8JOnUa7FEm6ORfd0fOB
7mtSSxwOQJ7dCLyng3pDCJjuOpRgLgwETgYqqZyt2u6jxq/kq75SDua7t3DkJy5O
yMliVKhuSUkLCRsGZHbcvMFIzRQTABxu6zSa//XacO8mg4eNxb5AMYq2fILYoNnn
oMNnuW7AxtlW4J+ungpk9PT0LO0ngNMXMWP78hoGukMP/XspSafDhhEoiEYHnTTh
/Z7uStCEP76U5rxbE6WZ0F+y1FZuBllVpDH1kWoQqYDpatP1HSOQPc1UYXsph3kz
yiqc6Rw1CzpxrtQL8X/BDW3QWN7K4xisQXRLej0UwNvbN+rIz/JrLQ7171YWY2r8
MKnHmFvJoaM0klNs/4v8aOD4HjB4eKJE/pXheUI1dTIYj9lPqruM+fHdCHm8Vh+u
1qYtC9Cku7a8Lfa57G5A+mv7YXbnekHv+r6eFuNKxYDkhXsBEtAClSeGwzfCygkM
ZQuiUoZha8lNWS+tPQY1EAqzGpQVnfBJPkPq6+oBm6CSG758RUlnSJkq0zTpkGpu
jHs+osQUDel7/wYoQ39PUTght0fF3SgsMto08wpo28lCY3LCP9DEpJflnFZMxuHE
zvpn2k/ffSt3yCPAbqgyrNbX7MjUJSlFoYgzg/vIBW3WlL4Xfca29SqtPNBm7sXH
aY3x/v1vYf869rG+2fmKl//rNXeE9WrTJz41g+hhE/0B3WsQpgkhlF8fyMHHa4W9
RyzfcchzZO96qRzXNW33hZDpuOCXFcYcY4S5BUy9JLKu36yQ4ujGZf3Rwl0hbiiG
GncTBW72KyFM/BVXV70d3m+hMg5scc3oNzyFSZ+M+wr7V7/PDGlfcHcoSsTL7SWT
BBrAWIZcmh9S3oKqX/XGZsaMj7pNs7ovI29D8bUVWIjQSEpAzqP2Ugi9syvdXScR
tQjqmB7MER9rnorn2wOUWelqQu7rOhVFPwSRdoRK0Iw9wad0ItwT0HVhKjstA2jD
e8qzxVHhJKiCEJIzHeny+1WcJZI1glCNO6ffoysLngORfzl0UtQlB2L0afFN7Ya+
eWd69jUKlpOLq3vVPzP8dutv5FkgY52DvnufzVVmc8EoLDRVdo0XELan1a8cl6L4
C35w1BH8qAKZ6kUZhJjAMm09htUU24Cm155V4tOJt3L0rV2IKyZxv72aKSOvREEK
1N8zV4y7TDsHmWIMYJ/AJTk0/qrGTDEh6QDfVQ+KQ4JxVj5/Kc1z/qzhWlSV+rmO
U4oOdhPzXk8R21yVU5d3MuPQ1r2+ZKuuzIpC5+m/NPx8FA0zjFLwJcUovn7ffTod
9WldnuB1HgzZqCEGZDMN7w8YX0dB+xiZPesBvyJ9Ok0GxkRQIFtzeTiiMxiJERDj
CQauHFpy0aukrdIBpGFL38lsdMztOsATb7xF7tFFXWXkjrr0kxGht1FXQ71enMgq
5zKgDdDM614D+ltQXFF7g7lPXXCQdYyFIfMkl0ds6NSfAea/fPqkhdNhHA+/dnbS
FTpj1afKRL/wYZvQEBYp1j+zE5DzEGnHdamvfl8zvTXvN3i7kuGTuVpZto8YfYrx
xCw3x6Pfu4DSKGbZ5nQHBawYsrT2BT7+IRPmDqvGQMjUnvsWc/KAXkVd3nEPURL9
rwfEztPD0WsH3Kzh5iEs9QxmXo00JG7zxv+u2jHFJjwxenqCZTuIYiW2AaHnJCee
jvBVpVLH7ft0rKFcb1wI1z3aN3JLrAYCyZMEU9x1FnW55dz6mI1lJaXjIhgC95Cn
0l/9CAjhF6WnSiauhNtgK7ixV/tswtGsAXYkWLdgXWaHIiBguJoBU8L3D7XgQNrC
kj3jxQTDHQjjgZpIjums/g==
`protect END_PROTECTED
