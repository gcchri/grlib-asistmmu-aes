`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NQdorfZMVF+AUshspyc+BxDj81ici7AF8vVaKjRk6igaULzWraPTjHsRcGT5TQSM
NCz07hUYpLtznUNJ8wNk22Uk8BIMiAlYxwYqRY1jVL4ctbCsyQsl4SrWZcWtKvtK
99gynfWcAhCsh/lnq++TZIHmh1CcX1cCdAsg85uObEzlVW0RWMIl6JVJCg1n2MwV
oA3Ip6/JI2of3/es6hTd2PdzIRNiQW32M7MeaWreYgH7XQFAQ55TgM6moNoYBRhc
UiECxcoWyF0sMBFPCzQT29x0DP51EKGRk1I/BsTVjNvWm8Lq8O+BFl3kCxU5BJiz
VX3jWz9D8FhzV6sL5iPUHZG3OnQ5Tp5TRKFEBYe/C64o/nm9SHgU0YwgUlon4vpj
ltCnsf11xpEvaYZ3H0J2G19c3yknw7tAuG54ho7eRbyyso81ilzEQZbSBA7Zi+GZ
AZ2yt5KiIj8tNLph28j/9bwVAAt53oIgQA7Rt16ysKd7p5sXkpICpJAHqEBQeRZA
bEUZTFVI46w5IAWDlPiKi3kw6PorOQzfKGRUNlYQfKidssEJs9gRFss5PVRUrn92
bmYtR+RLy5IyUUR3YPipZaIwOanINV5zc3fu4pcoQFttk6SPCKDlu+hwjkBrPBYj
QQJQPku50qMOGwQqeV+RPxJBJmgfOEAJiuHoZ8e1osnksCKo57TwT4iP8vlg65Jj
K+tG9HmMeQQIFxhxdmfQ/jzJy2LQ6AwNZpm/yG49mNOcoxaWUHg9o39Nd5MYn4rn
sxRtNwPth0GcMgzMahjIAE1HGg2R9mJuqhh1IX3DrAffMAZLiMZQoM4CGqA4Kp9T
pDio6bWS/bHQcgZOplnJCg==
`protect END_PROTECTED
