`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wVvvdi/vvUZ0q69ZwTbamYvrxlsc5L+2/5pjT3K6XtGU0Ybe0vgIDKyEk67Oj3u8
IEhtqkTdvyN80nXJUgdXijrpFmyPj2oODgOGf4tu7XwwDJjkR19hRWnomA2aDCp/
bimFc7D6yrZnpPXj7BHwQdW7+abpXw1Tr0raQyaw9+G51I7ki6Q4DUw8B5tM0mF9
ti7cGrEkFsXQC2tUIa1zc6u+dIHyZ3SI3OdCn2hx2nKPxi4pD8aZbOZ/ikvIq90e
1o7/Mz17OPQ7zTawtGRMekYhF7D8vCiCUe3Czf5Qs0ZK+uNYkK1ynuBPUSVCfGZI
pcL+6T7RGlLfEdRqVTF43qnxixvX/hg1X2ddPxt8hD6ULkaY3HRobTNGvidiqIrk
ZtuqXCeEXZ6Rli10Um2vC6bwFjUlUD0Uomdgk5YxJc/25dNuXzaY+jhUeMIX6SMD
xO0//zx2BZitcHzU3qRwp4vrwoJz223HhXYlip2UGZKeSv2tac/wave7fTZP2FcM
O+XAc7jlUFfkf4K2nmpxPE7BX16DhTNWlENgdtk/4MUPQy/92Y5ZQtScWu6j3FxN
MBE8MNWaqo9WWPYatLNmg+fAGsxj90zQj2gCPQsU41AJf2SFG9DNKRPFce5qB1El
JQ8KB5rlU27OYfLWMOdeLpCbb23rkhYzPhFmlTrEH70m3gl5Noq78JhieYJZdgBm
DSdiqt3yNmubmaKZ+3GTRaML3VsOqPa0bORJyjE7yNa88/rMGz+bk4mxYlOGtVev
jN/E/HcezDdFftH6S9u3CXp/Ti9vETUZqCdbhj6ESMJzNIR5ilxYlWZXbjD/jM2C
qKSJhWJqG1fzbsW+WW2QvKMQIPJLnxPLKkKGEmX9XhPbD4Kb0lychTCSiaL47qKp
VxZmmkzjjvjSOwcUfcsXcJeRlWMXXMr3eNjD7uxk0Y2rDCbsCg+kb/CJGXnqCx2w
iJ02AfvVKv+hPHXeltq5/9ErbtLKe9CNBUGxeNAHd5FItWzeAuhrFS/MWFycIk0i
8WVlfYlwGKHlHRCqlH5yqGpg62AqlwiL2WW73OK+2tBN7PZ50ikQzi2nsZwIxmqF
bnPoewxjqW+rJlF7DIkcMNMFmlKK0l26p/8SUfedBhrAqJY9difcrmHLj/NYKxOv
dw/bSzdbhX18ciBLDjwSgDL5+4a0VYyZBraRnc9+XDmLeeG1sdC/nN2GjH6oH1Ab
3hm+Z9R0f74P5FteDOhYrwkgbci+4jseMAUBEI5Mcq1HQ5Z6RmdwV96iASo56S+C
E3ME10r8DfupaNCGk2MnfWKQKrxr3333ALPDof0GsZqVitUh1ksei/rOhXapD9lM
UBiv3Fn4OSvvH+QQszRbHdletXoSdVXj3y3o8EySS03iqvKtDVt3wWR1uYUgg95k
Ii23JW2rW3wqG8WhddmXlYYYJcpARZCNP4i5w5beEqgp/+luxVQuhuc8B2vWSfZT
4QdCYUtv9Vlt1wvnHH+8HQ20vY0mhitRJyH7UTlkR/qbKzaapF6XNpdryzAcGJNo
nVbaiJrPINkmcZaPdxNqgEdEjIWGWFXZTic1ynjyHdaDcV68agXQFDWCUMEJpXAx
HEWUTBMlvQ78F2LmlvrWfM4fjz2hw+xfbKmGwdgL543Ox5600T2cQXlZiHz19I7J
SR8HgudP+a80ozW4U6/xOliX9hJgQhrbZpM5/hSHGofUgHKO176dg8aZhNUggYxm
8HPv456nM/O97XAXKpMvEQBFMAikslisxFfOONhhGsJ5gP2J7cT1Oak//z6LW/VF
J9uI2fpWwwTe0Vwt6KkugNjxcd9NbmWpuRsBZ2VwbZO1eV/VU88/YOepNRcpNori
AlvSdNNpYQYUSGgvzJWMTD56GqGnhrTjJZO1OL+5B8LC9PhDqpK1WVfDZvsDefEA
zkOFbs6wT22QXjybcSjCWA==
`protect END_PROTECTED
