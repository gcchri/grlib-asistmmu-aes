`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4IdYjV6J+oDnpCSPuje4PP69QpYUDmTiD0ganPl4yAzwnSBnUZOLpyq/tjiajF8m
te/6E9GDRQCr9KK3egS+ZHxWBjnon6xclJed/zOBHdRW8CKrL6YMQ34KD48MM/LI
1NYw5dizYjHfFLiQuIdhURR79GnTiiOM9AwAvp5Usm0P5ZSiMiU+A4YgGAEVa0Px
T4JXdgYsUasI2guWL8HUfD8NmZCXZQmbFEThqVnHKf4b7Zd9icuUYIJ5yZFBSvRk
97SVFkEDfbsyJpZKPqIvap2fy506KJQVrG3aUNOImgazN0l+vRritzz6enUNr0eB
R4oU8gah4nju8/huBt3SZQWyS+U0B2aNqFBlDNlH4Q/SQLfhR9tC4dWGHFeVdv8c
vtVg6blNwWRtf7Iw6TDLRI9ZPcd3QwZsCjR1yHiLQq5tStUYoUmtkDT1OWoa5wjq
O9ifV4CUnB29NPF4G4F8gA==
`protect END_PROTECTED
