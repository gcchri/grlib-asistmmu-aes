`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d2ECPHzAYHAu0Y7yA0nvDYgc510oOn3fUiOnK/3fLMN5zQrF0hL2/nXdcuA9I/1o
B/i4gaIiLkXq6L9NuCVF2urOwKdgmKYX+8ji5dqvOo+69yK/8725C/s3B0w/+GIR
behUfAXR07XpSSCS2OYJfQOpYrx0Aj+CwvuoKmFtNFpCfUSpvbEoxXHxutxBFpIX
aRqQyIW+6RUKL31zl06CcK7iuDp20guMmiA21JjXSzP0t32dY+G4wUuylSPQFbZb
oztcn52EQfMguLe8ZUP/kwTFbXdR6918OpCjipEbJVTQcmuys47/0oPFUaJxVFiK
X9xi11xRJOcBzDJOneVBJb6XRjarKYm1rqFh0KBBu2Ac5xRN1NeY4OM7LzwCqN4A
hBMCeqbESL0inajppSzpSrOvJug5YpIyLzg6APebowzQSUe5UN/q6Jc75haClMbD
RS+eYxtM26X41q6wZoB8ud/0ktQZT2yEhzu52FJHpdmx/RdXm7v9CLb8ZrsaRuUN
X0pJkXDOIq6IFrW9dbTCaRO1AtMzUgdANbIjthKQnt3tXuf/Rfti2dXYzLuc/kBf
g884Gau1IOiPhEEuHWlGsdoJ6rP2vSC0m3ZLYRcXGyowwCcKC9m68RWN8Pk4dgLR
BHoL+mKTIiHubmAYYpAX+w/ye2xCbJ3ZCsAT5it9vOG9ovYPmmCmpvs/STCLv/Mu
topMr5BD49dPX8DcqoANSOLNB9xgD3dLY+H2RaPK/rYKw7/MuJkcKYTOj6yfuthb
oDfqOOw+pEg7huI5W52JicR6BiFCzy/9wZ1PNEPj9l4P5tmITlWerd/dOmhLGV51
V9PbPYjvkTZbfkL2CpK2ub+op5vKD5WF37G+WizDOfqkNXHDwkqPMx9kvk1fGsji
UnbFz3ynTmprQ4h0nUQRcxAROdBoOhEOx1T5bmw+ZM36y1t8aiLB0T6zkTG7KnWy
Ho7ceDB0yShZfI29whg33ibZUP29NlFe0OhkFfE1eChqEJrM74Iw5IwRkFJh2EtV
XsNEsk3tk8T2CZ4PF0A0+g==
`protect END_PROTECTED
