`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BOAyP/OVGrB4UfSajhq+vM95XTzQSyNef/Nb5Cp/W41cfyxmeXfYJB+jp7vDMhh4
yN6++O6U5jQ9HSroHd6/8+kA8GqgybbCp6OoZ6yrFcYWz8usfo8RGzEW41fqEl6y
k6VuAgqBI2EGG6IZerfRpQOaIn/ccC3O6lEpjoL3YMHHoWhbJYlj0v/nIEPmxwHL
2PkBbMq+0YmuVmGkKeysPGZqYClMwL41fAX97w9koBvHY9Ge645tGOrZA+brXahp
tJD1sBZ+iieif6ha7XDQ3pCI4N2gsbBbB/Rik5nqkfpQRSev58Aad2BjW2RVouA+
R21PBxU8yVk0S/mNmO4tTmfz/SZo/6Z3bJCEcLHvF6gTYK3wN7BaD+jOc9TvlJGC
u2DoI7wSTdetJ5LLbvHRY9loXfh1FNwWD43zCcOobdwTovNwHmPmv1CGAiEeTuKF
Vh0QO+FMeYXec/H5QDyfNQ5BcS1WmQKXe6gWE9KS/AAUNhkQY7i1OiboBMcxpSFy
NkNgRHDjIKlKMArtxQzxHocK+yM3oVG85ptsNZEFnsU=
`protect END_PROTECTED
