`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IicOyX+t3FLnt0IObpC4pDdiu6hcSGhZZmRSvJy4c0GtegeFyrskQro4JyujG0i/
Q9EyOeMUokkGRgKtTUyT6tr6k/FmZ1Pj0T7//2uwL9pkWy1UZojcJHqSI37WsY07
jUA7PavVoXLLuraokVCwgv28EivaubzDI64/6gbozl4hYEFpguboxwuEu1H8CcpA
IrskDnxr3HL5t2twjVDsJ+2LhyYpM2RXCbc/sXnWeCcRxDONDm0ujwvMvGCjpOWd
W3LE15NGM+Iwv9PKRn6rPra4pfsjQ9SBBtvKPhChEEl4ZPlOtLs6QTvdMu1Qo2Qj
yjotqwP9RW93Ubv+waw7B4e0rrPUWGSLHCnBhESO6v9LfqhS3U8xIEFQKYQgullo
XYg9AuUNp+gbpvagiE5Vaw==
`protect END_PROTECTED
