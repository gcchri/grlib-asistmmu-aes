`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/gAUd+GA3LrBou85jQpOdNiShwK58uwD4gtAkHRgt/VsHqClvXBKVBsPwTEza4rF
rMrOhAZGdDWBmRUoxlGve8NfEXMf46JIHgP+G951Q1bsX6bZ4NXtNjqb8SdCBsHR
A7HKYsYDWAa4mq8g4xqXsPjRKopeTIX85krLnx0tA6QbJjh6Y9LGBhswEpLHRq7s
FEH4oSBIaFSegkYK1LyF1u6UYqXo8l3Sj3B2XluvnAACzOVEcy7ZI8RKMr3IoW/j
sBht5xqKMjOpFfkMOEImJ8N4x/a1i5PyTYCKxx30u5RBiltP0iV64OZ+J6FupK12
nca7yQFR7IBt9kvatQWCmMc9fUPEen+RNxRscKNkqlZJOgPrfyTDiG0zKKdwTof8
k9MbXnwWy+UmS3FkUKcQUOKDYe2JbmC+mmZd8NkxML9IYEYDQITRIpOSIGAJlasA
`protect END_PROTECTED
