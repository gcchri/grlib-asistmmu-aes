`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YueqXnOKw8SNom2MGh1t6OfhAjLgiYRoPMc9QPiMUzGhyfXkpex8V/xBjQO/hrKW
6m6cddMK8Cpbj8nfjcWr7ogoM7xChlJDynWKncXSU6obGp/XqAXMKX/G1r813taq
Knx0ZK3zjpq66JMRfzj5oJ6I/vMapOzfIEVjx/7MpKxb6pCLBnlyxq1vGp/8HkVG
3sVg2cRmzZ8GxOS1tkfOvDbQZWMnKWlLhFOm3k7rVNDJ2Pxc8YmNqIcz/gwqT99E
gNCIv4aQ+m5kA0Q3qtCnV/gykswsmJTKpg8NrNpVPbrqfffWqBdAf/MQS1j3LbA5
4wukM3MVH6ZH4LO+BITObl9aVzRD8auW3xXNqO6AopCbGxBdHfw2Jeok6Zuo8ocS
HnN5nSXUknDtxMHD841jcLoGXMeIiuSdfDKEoOByLPQ=
`protect END_PROTECTED
