`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
13iIzQ20znWZxxDOFq1Dvuf2mf/6fU+fU7qlOXq2K45s70GaioVSUs6e1dZys8M1
LRwmSw9MPB2NzBVI8Hrh9aKnuCc21oP0dK8XuzP9xWsksumNrHS2/XXjhxHgCFHR
liA4qEbJ6eeqUGgoMWMsVJ2+1Rqbu9nUzAjbxBQ6ct/bD0Yp9prRUwkXwQbA30E0
qy51p+bGnDXE7z5bOwy95dmDXAsmJYYMJiWjjuZkWygvxr9ULgZSCrCD1I334XHt
lQe88IdOuwm18Q7ysTDwz9iTh2MjW4VFnAMA18jjHGe6a4GD5TxiiO2xN/9strk4
Gjya3j1M7cgyg6aiPSzPKRBzo38444T4rS75SqW0Ww7n4//paVuSgjixvXOJYkmO
c0t2UH8R9Rp27qI+5yl/6UGaXEfp7BOrHbPbdXVw3jO9/h8WzGMescX/vHU2NkJ9
BDHFNlibGOXBPEKK7scOsCnf1gaM1L2vSEUTlMre28g=
`protect END_PROTECTED
