`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HCzO+L80BRehrMRzNlbvHoRx8bMGabn4J+FuE2dykE38teITjSxtSBeFY+hdYfAc
E5qk56HwOgVTuuoA2ScBiyY8eKPEeHO4wo4l1WKYOnMbonlYrBevTw5iwkOyp/YY
HHGVdKuulvjLWYyoCLIgHeV1uKNR/tzK02MMQGJQPCRr8iZSLGCR7GimIXspeu73
JcXYjjpo3rjbc1NnM0M4PdfaFP0CZaM7rPMJXAqcCVaxbRIwWUtI2JKAtuQbuKHa
PPevI+UJ73QomkCrNBayxr1Y6AWg40x98CD3wGWfr9s8yVzViijOFIzXgGpjzKzM
Ix0OwtA3W8vufK++afYz2VxjN9MSIQ+IeiZ871qusYXpi7Nyk8q2mprZD3cVEahV
ZSzo48AHSQQwhJVTkLPkM2mbuAqyYtpnT+VghZ5xlNrBKeJy/yJL/n2IcS4tn5cm
QCCd0pXzw9q6RKStU3+0cTA0sIhVQv3jL+juxmmNjJjMDhr8iQ61AkwsVcTKeazQ
2Flsk2tzvZqgO2m8E4YzbomnMgiguRDcwVb8z2RlK+7shr9qknMM5/Z2grOClkCo
bqXeFq/ZkrokHGX/Sc74mg==
`protect END_PROTECTED
