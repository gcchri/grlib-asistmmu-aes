`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dNOvleNbquE6gG53QzfRzcoqoTONVeXlLgkXz81iQ9cJsxVbgasxndua8v4jJ9V0
NQFCZmmJIeqXNbnwOifXnbSrsXg40xS2ExcZFB2tWQYJUkJzNmYEG2Xt6NWgr3p+
lieCnVbK9D3ND7hIoJZpk/f9UGaa3S+sCXkWoX1FT2valKvKcC899uex6YHG1g9W
4Z/uaX1esujMf4qmlhJ0yEYCgoVWofRqWiTyy3KK6XuXMFgnKHIBq1488zgOXq3s
6LMtlZQA+1GbsbtOLTvG+rcdgfDXHNu4g7JWwp/oYfvbos2Z0PeQJpBYwPkmr/WO
9snf8MCNvhCTfRqR7CeuR8I78sdX+DPvtxMgtQ0MUs0PwPgVNn5y7eP62RktYY68
vP6ayitroxsP+LNUtaGlkw8HZpR0Q2TiOkwtdqQcJdc+AvMg3cpEPx5Y8CYw5hHt
KnB3YltxTV4eeDfNOsExFOjWz8FkIgXnHpKhD9Rij1r45dhwCTT3pc7vDhBA17Me
kiSUwpY2ZCx7NVu/BUxf7s4GR21U2ATPUIGVNPY65AuPSliuK9OkJQnNSZh7BID6
GODqOjmxOhkwzg+UsBNlfd/K/T9Njls0dK51DHBtqSzWyD4r/RxQBMXARRcRhH5n
`protect END_PROTECTED
