`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aoRKvayywAuTzrSnLfm83SZXypQSHS6drqauSu0orqwMFkbRWbz2moHbwUu+lZPX
Edtb3fF8pNsWVF6YK4WPA8ZqH39e/mQBgd/h4vD3nutxMJoEH7zX7c1pv27T8xSJ
gPHUjOMe137vurQdNCY6pE3LWjBmiiJLU7MuYK2kkp3MmuKBoXLV1c3g3abyXocW
rKqK5qVkAPKQh21ZLkL8Wgwd88R2WdBGqy2JofIZ1XUX+3FvqxBGGKuTBjE0p2lW
bZlBew8RLIxYrMu1YvTsYNrEv5snECowWQiDoxUTd3B7NvGws7LfROQfuDKQCNa4
MSiSrC9lmGECPRRDjAZcW6MppOBmgi3rY0iYwAEn5Pwg97rmDqO98soIs1uvMChd
tVAeHbY0V9rYhsNGORVsDvm8hFS7PTBazgfL5kiEfW4JScfJkbPtIMymWJMC8465
73e+uPQiFjT+z2lI2zHTZetBKaGgOONmkZsbDqT+GqxFJZ73KEYKOvgxBKh1n+Ss
gwRNjAsnxkECOvzqvwrSkNuDTBrWdd8sXM87HtVmVYmCUfHa8NkUZ0IILv1nxDm2
tObCrbTdSTQ+DHzKfEFtG1FKs4fWD/g4F6xN9pCaTBTOq4Y62166/cSp5kZhWgvQ
Xe8Uup6wTsy4hY+qB9/emwfDhes5T0LecRKO8LGQFW5P6ZkCPcqgEiYJPiFkHI8V
GPh8ZHVjWzcBPiw/4IA4ZJm/Rtq8qrCykPUZUC4hodV5D2H4rb8CMNac/zDsxD2C
MR7eSGXUgeY6JbR2Fws3Dj5LDLZhgGAVmZrQQd8RrkbnRErSQOFe4m6IGWKifVIJ
6V4lb8cgFEvBlspAlIYg31Y72mgzfttwSw6fJ8onDptp5ue1YsG4MuQ1Raltgjup
1PIhLMhfg3H1OuoavoUACSDGxK638J+bUcj3yJo3If8WXSStEgi4UXxieW5UYC85
UwY6o1C/XkYI9FEs+T5IXPB9VbyeftPtwqeNkMwSqyqbG8MuO5xVEDtSVdInqtZ+
o5jg/ndZcpxHTSYV4NQlrlzWzgKRV7mLb7YyTQrepkAUMs1ZQOjN3Efg5bfhBrJn
bSzHr7MKUpKDKwkRxd5R7BOPXoZbu0qBvF7vgDHA+I+KEq7n9By+39sbtlAzWdBq
/UPW/bXQoJXvNmPUJ6Vm6ibcS2T3rjfLIURntdpJ7FqWHP1OG9TJa4CQci2bSDor
WAStc/VtVzcK3SxlaJuyTxYHXogaE/C9s3TP3rrkt+9gQN04J50i1NZNU4JjXYbi
Sbmf0bdOKeG8VHsjFp1zSg9ZJ7KsIduxKcmv+gl9ZYVDh0xVeNpq8/twbABNnc1h
Xo1KhTe3JHw95H1noEQo87ABW8RiVz6WHgsKko8tZ6QuTMqagrdR3P+tCx+SLabb
WY3twXgTWEb+wjX/noqv+c2qBylyNGoVqL3nyvtPoTmadGbjOLSI/4V4NzfH5rfy
sNmm1lnCiceM2pwuve+ARTKzhm/TVagnX/ngI7TNCgpIthJ9q8tXeHufTTdLVtF6
AMEa1UXjrKgARai4hqrOUGeEmfuCAJU84HVSSPb4rmDUk4qg1owGDGHm+d7OMrFZ
ZXIEJwnW05PQwtjc8BYJsrYsE/p4/wER9ZAyCaifeuXo+cDd5Q42rJTPa9WQJ9/k
1Zisdf4/pmNPe0LCTFgKgwqN6YUNqBUIGIhUSOHQnn9hQG9wbGnOXxVRaxODKrix
7w5xot35B7TIUptNiZ3PuwHQxXI/QaOvpkWpLTAmhbVnfZON8w8qHIxXyIRwACde
oF4vJPc0YYKwshCuQhNushv7q19w5PXMD2oO7E0g+8A2r9QtzrrWHIjFynzTLm2a
4z8KsAgaOtULMPlv1kJu3eIvCyyXJMz8nXdq+jWPPKFPIpQOdrcILnYRHmxEOiFH
v6AYYrgoaHyOUPiqdSF/U1vrC3UUwrETPTsBFZClouVU4Pd3bSkonYZamnVyxSBd
wINdGdMIoV44J4rHWBasabnx+VfwdQIjML4VGsMbaf2ghxZQnDL2+ofU1r/Ajly5
oFiamxnTOdicNzPXpru96mEXBDHwEycUZEDYliq2wd1eFVAMsW+DU3jwFOMr9D1e
q+6+KQ/Z45td93x0tcmDEHN8d+o2NZeRllVdF++RnCca/9ETKiY4qLLwtSBSR9KN
ff48hwASODuPNg9GxwcV81T9gm4ubKGj41BPasHscTjaDSWmCPQ19wxlboUHEeGD
R+pmyxlda7DyWYM2LkkgfI3IXCoZbGU69qts57XJ903rIo48fijfb42mdYxgzuqA
yTzjo82EcQmkH6mnDxbCNA==
`protect END_PROTECTED
