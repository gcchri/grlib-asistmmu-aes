`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9niQ5qf8feHHYWX2KsUBeGM0vzQYpmlwMrUuDyVSWWDzrlvAsE65XbeRwcvOm6Qg
q2TrJtfNLXcvbI3QFdu9zn5Npz/BmtqpsAEy0oe+35+DBnrifaqwwuafX23IRQUR
vGxpp2qF7dDB4l5GgF84hSIt4svm+1vb/hmvWD8AyeKMpEOrB1obuAN5U700eTLQ
f/DnfPPxPOYhVYZrTkXTErePGnjwrpl3lhdXvacEFoYwGM+7OxMJaAPRum1MWnGb
6nacxpLuVEdAvYD8dJHZzgSYuo0u4xndgTeHG36EEVgIcN2GGJY0uz+GDfeGe78t
gxrIMyn3X8DL7J8ZJVPqkcW0deRHEi8Bbf4TKwVXwYnq0kF8ETc/qs+BFEUPZo/y
V5BZkUipXB2Ye6EeiG0c5obTH2xewyHU/RHE6HXyYpiG7pDb5xjdWw5AJkKSzg9P
gXB9LcBkJ72TCmOWeva/uMthaza0ChDZD2ctkOhsBj27Gly92H8hqpG4zd54cSO1
bfjxe1HHZnTrAEE9elQS2b/CgSlEJEDgLfPJ2yN6BsJ0LkrJ7AXj6yP/CKPCBRyh
Cq0+AI7tdjelRekOfh4NPu+Uwsv+IMJWoKnL6KcG2vogVyF5rrTG9uJpiOs/WZp1
cejhZQ2mMqBczvBhvHfF/szrDaH0OdwBaxDcPzMjOaTacFtbAisi7F7E4Q/jWBv6
39x9X9HcRAYo0vyh2JOH2pm+Q6XhmeGymrR4ra8OT1XKaJhxD4TLKsg3H7s3x9Rn
LASbhXsGlGpHBKBN8lfkOqxJxLt8MUiMH2Zwpx2T9F8IQmlaVQ52bUVorV/nNvB6
O3YefrYk9oxotyieNcMymAHRM4SJPcyIbycVvY5xkytKoYtecRtrWuELlOVt2d0n
L+X5yHWtx8T2Zq6Ah5O6dcRDmnpv5tK2BZd1WpjLASGCSKJh+XHMbIzxYZ2XOkQ0
2svZ3xYWViWD2KiN+AZ4OVyiy3hv05lmeEvsmUkbAXcegayWy86IA66DpDTWI+/2
zkMYtGMi5uFCRPsFVSw2ISZwe1vpX9DvyiaBgHKJxGvegF7zEBGIMc7HxTi0vZ2H
dKc/bRo+Rig5ENWgvfJUrsGAPAPhdx1JlLZG68RYexwtDERFVfnt/j0Ax2KLt/bp
1qGeNjSRR6Vuph1kYB2ynuCsBpE3bkqEeYsCq2fqOe66DWwpOstpZXWmR0goSwuC
1i+wbmke12XafyD8qDUAZUmpvTBCBnRO+2ZZ50zRIzWU5vb20AI8Ui+Hn6OsEOJG
uXk2IJDMfN6T7c4rYSRtg6XyxIfZYinyXOWBe1OPFpZRYYfW7G9d6GG259O2YsVm
mY6G7NrT55W18mjeaHQ+sQrGCg805lOjAhjH3O4cnwQWdMfrIv/in+kMPh92on17
xMD005C4rLXFb+M0zNdW14UIuI5OaZc1IN9R/4aripDjgtOqZFlXdCU3Ad8ZHhvb
s5RIlQPIDTK4Sd1qSPL29P8oNOIKblMnWu0fVWfNyz1rnBoYYTkKEmYiwW7Li5zG
9/XbPYezZvOHmY+1jjLgUuaxrzz0QFn1PJVaVaHSyV0CVnL4ET/tVPhek7p1f199
/xfcxkNid9nk7tFdSnUuKLGjAOdyhJqJ8G19sg+t+vryZSwY7sf7yiyyusMGJPBS
yC9/r4QlVdY6m/w9CoOMvyXg5kAAfUHYk/W38JlXsBHb5MmylPbsVwtyWopL2nsU
FT35Bx3kAfcs/NnobNnZPFPRRLb+wI6qMWgaSlZBgh9jwxj6eVtBMS8FhZBk69gG
mWXUvGoda2EbxnQ1XP7wlhtOqaX+2Lh+kDXrrZo/LZgiaiXgkyd25wFJzFTRcI6A
G7tg/wTADGo7mdgs49Y7XgOVTejKJEEmZUusjTXOkzpFRW4Sz2LNPGhMTMuqGl+5
JcInRdi9AzkvT3Phzmlqe3P1vhskexp720Vx86br553Cley8Sjhw9C4A3//zASjh
dstiFSKtro38iaCZpcQ15pXB/DG5T68ztMLIi2Iy+87QtKgk4REqOpFN2WE9aUGe
S5fuVqCAH6/VZfmEAqm4GNJW37clIF90RFJFZWdPxeYrD0xw6VjZN4hB//mXRIV4
99FMQLTsxpMgt7suHHDBJwpaL4BSS3RwcxihwHEVG34b+XnNNsKcwU/wwAjYXNMh
bfzXkAqz++pjVdbllvWiA8KS/+iJTM/cBPiGs8XhCFoL3wtrF3qv2civ4eO3Rjul
6A8hRhDcHX88ZfJ7TqOb370QQaoS43CW3qF80jgkWq/S+pQsoN6ou/bSFnFv77ij
0dQjsMEJoIbPedIM5/w/w5jmlNsZMFOcigbk32mgpgTvlFBj7f+XQOvNbzb13JsM
2c4ym2K+jVmtGS/zbNlGm8nbvEmepFOkcImEtioyKs/lIOUnGQDwjFKAFBFNIA5+
f6OZnKCg2HuIiWKQ6fSZhlZEJ/3IxRnAU+mI42xmi3kc5FVWR56OzavQqLw8Xrgo
XM32gr1ERN0DxO5vSWHNYkUAEaWduzhe4oodIZ34QF0lqTxOy9KKABp45AC7Glr6
gCKOH5oNqtl044aFKioam7qX1QGuSPIOVYCF+VIu5eJfufgFejMvvwRDQh2yDFJA
+STspUEbnoFllYd8TrQFSsHo2msTQDPvPqJAAGkXp7XAR/iXW0TsFqUOqW97gUFK
zuTqPV57Bxf82epqU+GBcylcx0DMePhsozWm+mHJvel1qB9ZVy+rJwhAN2JCTRyv
JzhzIOTehDGj3RfoOFB6jWjJy1JRHqHNL3gCNygMcb+DLztlJjohn5mYYYLdncg2
ebT/2DhQt7Zvttwk7gjssb0U3VVrRr+MuoSFR4jglnngAeblz1DFF0+GXL4aTXaJ
/U0XNsakC1B4wADaOr/kiFTLX9j6xR8KLwuNKV2spakslbHhPifU7a858NMuajqv
rBFrXZIJy6ppcHPLCZUgmarIY7rJJ5Jy5t+8YI35+3FvHfx7VVVx0ZXg1ctHw+0P
uRqFA48/F/SSBkDIfnHM5cqMnulqNFLQsuaeWZeh50X/EocluZsKPb1lldSPo7DM
hGwOlP5YdzXCOa0YEyaJG2Y5mn8JIQ2mLRyelOw4yjRfcNizRjPFxc+35AAF0uJ0
qBT+iOHMMNzZKbUcLZJB9OcF1T25AEHqCRULbYEZtPw36yK6hGq/F70tJUVu7fIa
vAN+w5G31kwMBrh3qmjeIka1AtuWRdZkoMtgqQvcIOofhhVijDb7BmStwqBkM+j3
ZYa4h/rYEZmE107BtYAuHN2zt+03k8T0vcW9GFDDIQPrGO00n4Q3F3MZVZpmjIi6
iSRxWALiMZ1DocTBvaEPmnlZ6NDmcitF9PmL5BC17QKowYYO9heZUWtTqx0C7Yy6
Jb9zXHCh9NJka2I6y7tlSCF0D5Z5GQu1Y9KqWE4pIlXAt3eAH2REQaG2242EYxRo
Z6YVdFNkYgHIzpePhQJSw8RrTz3Wc87ofSm4hmQ4pr70Q7Q6VFS5K7CEwu64kqjW
xpY6ifhBcenW46SbaH0F65MbbfObdh9BkMjP4oIO5oN8z0ub8YlPlVv4E9TAfBMK
Isdx5lIoppPsfwFdYCohQaCzaZga8XehXLt9li+QVl8PfFA2KS9BlLLdHdpH3VJv
4suR465VUYDUsGPrwszyQr1+yDbEE2xrtQfpH7oYgK5pj73CtEw2OX4ISyjtVlDr
EU43Idq9MfXVYn9kj4MWt3lABKB1m7kDqT/5C4zdZdxqTgyP2gy/wd28cGH8BBUO
O8WMpd4+D66TncCKqprnnOnW+Qsv55wfYjI3484WGjZRwu6O+4gKJq67NNY4FfzW
6SETlSh4YQyGg3zBhAH51AOl/N/80rg7+hzqANdIdaJhIK6+8omYBSFZMl9Nzsn+
`protect END_PROTECTED
