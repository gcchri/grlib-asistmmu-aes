`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cXgipv2CQ2XwRD2hR14w1NtuOFpVgYGKqCRFApX8hCH+D/7yYTUkNmGOGVqAEfOr
5X9/cgbZhpXrJBpbj3DQ8NTXF4/LqloZoxAvnZ9KiOO0DNfJGJk2UeTZ7fGgYzj6
scCQ+DnizpzxL9dhjiRJ6ogmCYObYj53WyKY7Er79UVQ4Z9qGctjamgoiFhDyF1C
pFWcEz3BvG8YX/2mM6sVA01kI7WiykFCMDYzbHzE+FnlI7X7Jl7+y5xKeg6ywBLB
W22gA2hoaWT/BX4hNX+BgmqXvPgBeONh9/EMVwwCX7vLfZXQhSbxtcptpQKI6oMz
vLyfpD2lx4LcMCenKUbkAO//9TCq7oIsT56VOJMDWVnZEkfaYNB2FzZ+s8lYyl2p
aP6bTz5LbXJWkwgk1EHskbVYExlgxg6ibZWMB1PkfUUoLtpLgfB1aXR0juk2XbhB
Wo4qNxfyxsiqPNNuwKSaozDHSjwHZnst2HF6gOjCo0GQYRMlxwXewVwy5TzratGC
F4BZTfxOMZ7pUbsf9t7Q5m/LzeXn9PSjIr96gyyB8OIWU9vn5BXz+//3tSIl26Xn
OWqV489Y8aJ6sdrn/1lCkqKtz50PGAK2HlQuMpSqOjbkuI9VZIhxa0EBxtXNgo/H
LSts4BJIfGfwNZYJz27rqFqpkS+SYTGLqI03EOxw5QPSRDqNAUeuLBg6nbQfc+aw
p530sWvXLHxfCARssGw4comEJkSwDntmf9Txjf05BndWUaBsW6cJshGn0C/eXZwz
vn0Nk5/LgSfNauMf6sVnCO3CwzJWlmF1jjTyH4vSwv0F7jTRRUrXGBwQ002ixNEr
RnR7AXYtGj2Hp0GJVEwxlG83Q2GuPT6SCg4Og2E2aqC0tuYmBdIt0SaAxBZ9BDAh
efgqAB8zOTo3J3/NhR9Hs6nSAc62MfdWAV5xRcgG2fuuF+wkiJagQcYM4hc87pqQ
h7T/uqYFStiE6sF7ab2Q3eXVfy5QEbnWhn2ayv09roDxtCx3E5akIJxVkvTB3ygy
ItzAN2M177LAaZfYebhjc485d2rUE+RwIeG5L2yOuU62IzDnpp/bZxhkgXEv5dGm
EQVmOcwG8Iw5rhV1I4h8VIrvxpqkZvmjRTF4nSQib+KEp8EPxGhRaQgdQR06VJCJ
6IJG4h9BVQANGFlONCLp282iDKS9vGneEECzbsyt160yAXhrNGuRv+ECuyTMvIu/
MyzzVmyUygIlDzA1kyhqvKT4pf0T0xU7s6rJARYBeSSZva0MurGu4F8q9N5BFJq7
a+resxw+PDV5XCUIsBL+phUo0/3cqe38piO3eVV4bJOT3iCVdGA14Z+ITqboXOvM
TF21Bpf0TcDmSYxTtLybbA8AAH1wrzKF4potOanRZdJljVvCASTZA3eWm9H9vsWq
cM4l9PngczpemWFjpBDVfjOeCt9DTkslRedxQaj5GgfriRAuyXUWnTDofr+cmNM4
eLkBiBxh2BdIFKFiUA3VfWio4O+aQQrSLMImQEfwSY61A1ef1een3UPjri6LLvnJ
hTmstdCWUpicBlqTPfK0o66iMkV08xmNAIPds2JXjpdrYDuNpHJeXCdEjcprxsfi
HCNt0mqKSdHNv0Khg/pj0dG4FiTg7t0CiQGsq0qsWIfTBZfOddV+gVc3C6pKn8ZY
vv+dbjBFdLlVs5JPb8cY/GL09kk0GOjq8VO10JJkZSj1NqaPurNAV9r2S3AB0uQI
Jp6Ui/Q4bhO/ycq1+VQtuJs0Hqw2acKUoWyeEz68Klm6QVowdG73rklbmeabvArB
mpjmTHo7cxJiRGTFGDxpY1YyIM4dXCfRjHRQJkXGQV8ZaodIj3dC7JFl4BRIb723
UP0iCJsWNMmlyaoY9FalRyFjIPB7gpRtlXLN7nfbRpWyZoQ7tiIAFiwXYNbCdCCl
+VaNkP4cj1qC+RJ9oUfSun6xmzyppKbKK9GU3Hz27kfsEQnsTOKIGsxO3joH2nK3
7FePXl/IN4JXJ47QaaBD/wUoQxjKBHPitbHdu/zib/XvYSK6K10aGy5vQU3qdMx8
cUIMJngzfNRYl9Y2hrXWE6QsUdZl6a2+71L2XB12snFSwzDCivOQ9PfXNOe8gYdU
BygcupWhl6P1MCS9T68RZdF9Xrb3PMe4dyzNok7qXxquPY+kj1VFq28OXLVoOotR
KoTwihYtK8jLuhqF8MjeA+xylG6ss23MDF96pULXLWHMUuwnp6cJeEdttComj2kI
1kSKlJFYiRLxKRV3847KRKSxV+Zc7i7oSRG+k+S+yPSlxnDxvXvVkkqPMbJjLfja
r8Enac/PjrAwSHP+0uUUzfkvuHEVsaMDrN6REJveUHHaKaTGMBoJVMbQiKP8SCk2
VP42ih8C28Hl6nFF0GUO3SWChK4kbGOmT3cdQkoFsgOCX2ERkbngL5crMkM7armW
6sO+5H1WepYk2LfZ+b0qQ9roqNHClYJoVXnvpCBtNf21Ih3jSm7x1AwP2GGmbHR2
CrMs25YbbrYnxPwWWCgUqw==
`protect END_PROTECTED
