`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fZhhl8dkOlvYofv6k66dv+efCtoRkabjHgn1SEDK7N66ZXIvPgAdfdmTbmLfFT4M
dpI1IJuSHzBUX07T69xqkUEkMO2cZ+jGSn6kqxKBIxQpbYaQSJkyEZ5CqOwVqdNS
JlqaWoYO587/kwcwK3bbAu+UbZZEa/Dpvz+mC5JTzWiCdpkMyKhS7HaoF1D20WVS
Sq1PTnWMzFBvVD1Lpy/yxZySgx7mhdPhIKQt+YWYgXU9KyyFedLS0Ob0lT1QF/j5
RtS4s98FAO4dD1DCkqIw6s0ob6ur1X5jNpsmrTudtLcnA+YAJojjHPN8iMjyuKu+
MsVcDLpAS38cX3+9R/xzCP1od+7++/FPivIUR5A559+pPN0ZVCPciEuWz8X9+EnC
iRBKgpK7HxYtY3SGjcmgM0chPICCqkooJnou+PSKUIof4+YuEZ87gWJWjA/lEM1s
9FsN25EkPoGvpad55wIuJN+Gs7erVt4+6s9oOudf8b0OPdhjFPeXLpzcsHnrtIoR
4FolJ/x9veQqbkBel4eLAuif0wN9gtgmU0D/ESY+7RjwBjveGmBjy74QcsvQwuZL
ZkabPSwbCZlR+mhAjRN1cLxwW1nd6YlHVhSK3KaxzSaYYyM9iA8DwaiQ8+s9s3so
6kTCfoMDsrJVBCow8IYQaHNjAw3E/efOQh1h3Z8xt5POQeovMaLDz+hGZWgbMJ8T
`protect END_PROTECTED
