`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vIbZhoSW7ygDuS86tMRGBzu+qQXcviOltcS/BkZ58uyi6kb5e2AChMsL2OL5q3Td
o+kowkXlGyqjO0OfNTv3TrlBc2XIKTn6aF7AaATNkzj1o/PrpRamvY6tVnabYM8x
e5LebuUeJ1YkoHpLzsnZUjzPlMYD27mkav81rg4EQrrOhx9mcC/U7kFwL062C207
pHz/DMXdGG5sFbUnDgX9PkWp4OnChxBnMFm81XSwg4/6oRA/wFPssScRj+C2wZHp
36fdixNkbGbIMe48xpGnwUfnsocButtRN9NZfW8TXUzz0HI5BptyTlrsNtBWWiXi
kBiiZsnczpPcf2+QPlXAwDYsL57rhOD+PHIWw6i3rk4ZdHrZ71CF/3FxGdph8xfY
nyO/9+ZrIo6uwkVuC0CKNNsrK98Vu6ZWo0RnaqPOdon3LdYqXhnrC24G9MLuW3XA
nbOP3H7+ANAAi5J5syPWk4wVpGzZsgE1xuKnWo5/Eu0=
`protect END_PROTECTED
