`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YGcgL7zlc9dRbmMZAt+we6DCVMRtDwJ/qjulbT4VkRlhBk9RBALQVgGZ3bBFQLIP
UO5kxDyoW3ANh4FADH0s5s8uNruaPrg09/dWkwY94Dgt9MT0nRyNhJCZQn1t2daC
BH89Z4mzJFpXgoLbvBzjhCWgvF3cCNDHDeVpmRyLG1vZI+ZAh3ozn4x1TXrG+mds
UAcCeiuUYDQtVt5FDjjdHRhm8k+KZh39Y3va0kC5yCPhjoNd2RH4DPGD3pxFo9Kz
MpggjiN2RwCc45Kcr4DpJ1hpOkab4jIW9z4BurdtMvTm8GwJQuEV1/ixxmeXgJ7Z
BpvwqsaCCdvqCgTcBqvTC8/ikWNN4RNSBmcGWs+xwgQeO1UchHjYyEmI5e9ffH8m
PLlSbAvR3ZJtGm5caktSJu+yeldgWNY1yDBMi2Qjnm4/PqJz8jIcsqBd68mvZ8N5
TRxkw3+wyD/CbFwPMBxxQhteQxhopkoNMtpa0nZmUgW+7EfqtR50UJhjjaI8+DIA
tzI4wi/oVeyua9Z8EDOOibo8WS0D5BJ2owXKJoR16zljcgoSD2K07KnEJVBv9nie
IvzyefCzWeBRJ1yS0qn37bsythsQKt2cqwhEEY4FfWWfES3i6NVUvnjmWHvC0kCM
Ajnj1Ub094LdXgbcAJP4AA==
`protect END_PROTECTED
