`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gf5pQA5nzdLnfsa6LkjYg69FplAyuwf6G14y0CrkFhSDUDFGBXfybAxAml+l2JYj
wQnd+hnZygjdRqF5KP8UERif4s7gOG9KrRkTrYlnXT5N/egGgfBNafOv+YZ9NPRf
522c21lFmGD1XS8vLblW+nrO0yfSlKYRQ8l/HnOp/VW7QBiZFt1PnDXDR4TWCQqL
f1fVi2GzSXrqQ8FEYskNj4fcKFR750ofgNkUBCW2MfIjZIre5FP14ODnPJRnr9qG
2OnQ33BApFNwnbziTN0lg2CJ79Ei5mxKEdL3Y92fP+k5stZfy67jz8VL2+iIDada
Iyc1dpMsDYb5He/weycT2f+e3bPFs3bt9YIB8YZN11etRgiiqoTiimi+vqPI/ydN
S9/gaVpPmxhnEmJsPcp1IouleLBBpKxuZXgeHIKnI6GDJljULJKLJSpYfiw2eb2f
ScuBgXLcOVg5ICt2YkI9etsgaxrYoe7Td3DmZPin+q+/ETPIicPDrVQVFV/YhryZ
K3pMfNj7OetvIiX92z9+nKRqS6rYTiXgCNdwI6jbvNNDhgRYb3FP+LDGDRyfiaac
/gDtsAHwnQQiLrhUFl77FVsg8bGvB5FcTlZ2mWbcI0M=
`protect END_PROTECTED
