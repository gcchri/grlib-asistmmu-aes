`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b87wYZV5Dq6ctCMoFtoq0nnOI7M9ECG4jYe3xm2qP4lBfIiqyUIODnmxctO+YR40
plzTZy9QzUqJXFDobI7rVg+Qi1GgvYJi0cioA2B7Y9WTIhrLhulnVpopAMUmTRE/
wZjd79FvzmaKdALIm5cn4rpU4MEC/LRzZUZIoWQg5TeG9wVqZt1fqP2N7HI4M+o4
S1lfYkpNKk3/fcmdCO0n/fRWfN1GQz5/yWeuuBeLiGIAyzW0XZ7LTBFTLQAFE6sS
6RQvUAlakX5ZPQX2Kbf0hM1lZNNwlV4z8aXSq9TioWsaNpOdcPyJ5eH5XIEACRn+
wNwAkkad+lsHXvpYDLO4oKN3IlKSNHXhChC04cmBxulQ018O4mmmyj6Vq2hxwzdd
AkiGzWMqvDmsceREKdfgZqotISlQ8Dt+xWoyqKQ1N5obnBQayEhix3mDQ8EHLksX
0Nto+Tw4GE4XYglPJWRpSyWZQeprzd+zBQXf36n9EdWYMXftHju0yftAnW6MSqfi
`protect END_PROTECTED
