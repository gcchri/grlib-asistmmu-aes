`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5u0d+oD8Uo/INP7ZUTDtLSswh63EZdbBZrfXOCZQ00qcwpHV8m4sVp9AkqYsOW4C
qRr8Akqaq+tx/l/9ZRozPX/lWfviUv/eBt95SOvKMQrtc+YndipEBKo/WNx3SpSG
Z3nvoHEkRZvyqWqNF5SgiH9jXmAzSXh9xr4sOVRK8YD6Zo+xxWtA0Jgo6yFA+xF9
Yw7R4DmSFTwCASffwgDodgyQ0ujQMEJsgq+8rmR5L277aoB5HqR3intD08Hb3iyF
BmQrWSNJABCXl68CfZzd9aBQoKemcqKNYpPIiuStxkdoH2erXct+4CxRW7A3u+mp
rQZgJeichG0DCBP7g6BeyqeudF3neFh3hLmkjGxpQNQAYtgORX6euFSamQqrCcRv
vl5yQnZx0jzF7K0LGQ9G11YXogv5n39OdUREOHLkE7oNQ0eTxCOuzDd/B5HX5aau
4o6EVPkLTzx0o4Lo3iPAml8r7gHpr4W7PWvX1H2lngf2SL4QiZSJN69rojL6eCBy
UOqViWpTnQ1iLC3Vzv8dMpGh2O1xrxJ9q94rQPCLVvDyeSP3Din4x53NBHroFkzw
hbNlmNM6bzwwO22S7fPEIeF9L0pDdNystsDYHfbr2ot1MAlwg/OT8kL47MqkIQ/E
BWr3NPlUSRdEbL7xA2/luaPpm16Xa/z9OTS5XdtqcDUVSxnxqro25zVqq5whnVQU
eF1yFCkYjeVD6JLHt/2ohEdmgbUcW7BMyqWwYyE8UM2Ky7ko4Hb0HyzgeqoFlqE1
g7eeUMEi25gv3p1GeEeSVdKcV09dYndQd5QegvUZ5oQCdNabQHREPEPAev21Lcqa
jhCDIUo6kCW+2hlUDFFraKXUBc9a3dSGWZ/yFHc3mrdNP5yL0skPKBrs5wrI0nYC
6xEFWl3h+BzagJGb0opnxSUaKE9FxVwJoD3FykR0UOZsPl0fHIMKSetBBazCbV4F
iYONhNvUHFdcCp+wlHKryom+4xI9rAu1Is8dDg6g2FFvOOUvrLvRSJ2KzQvTYZvs
8XXXQu2y0zpf2HMtEp0c2q2cOZPbzNC2G0jzSr9NmoYfW2ACor5IcBGB8qJcz4r+
c45tkxIScSsnAcgIPrJSgg++BGNF5ltESgVdlyj+c3zqIRRnsYj7Xo3eNQfR8lL0
YKjmkub5txtsoayYAUrEMajN33Gmn2M0DlGv0Dn+n5vUSh812wWNE+m4R6lfZD6o
A73cW3pV7nJAGMMtbGGWwVQsnlFEm4H15OfN3u60thiWA4DgTWIVF8tAshqY/s2s
`protect END_PROTECTED
