`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5VbY3VyRk9ZybEwSRZlnbqfgBSJK+t5z9xxiTsJ0unsc190f72T7K7LLa3QEzoLX
w8lX4Y1vbI5r/SKgMkXqHeTXpfyTUWRTt4RLj8TWficQZVuLobSrLN4Z8b3Z+yU4
4a+htXdQXGe38FyfbWs34JyFQrWgRYmWmklCoZLAJXD+tVYkh1gP4KPkntPTv/hC
vOlK1qdRpFNFry4d++z34Afn0T5+qFTBpAoeRpxlxrIIG3F2lnwpU8Q44mSbxFQk
WBke/J0yP0qT9SIDWZd9Nmlsw0gGoxypoxE6uDM8dV5k9C3vwZUavvWme1Pk8cRe
PPClnFVKWhiogETX8KwtVP96dDS3NR0jguUnls5iP0HTHuWtL0jhbKb4XDBq5/pa
B6s0I+wEZL1vBZ6KAaFTH3SQBDkvoMW8XvJyUZcriLhk+t4NJJ3OlAagk2dElk5c
BgrLauRmbX/hRd7QpuASHusNShvo69IEslxSH6uc/1ItLEbzCpI4dNOJInFW7ZYb
Hpm+v0ER/x5Wr1KXiCl5rBRdHG1iqqpv1nWWUn3/EyrXdFYl/kzhVFDc9/i7xfVH
uL0rZuvOlAIlfjC71cFa1pSsORg58qq/97d81M7HrMtY4evOc8xbg2xd73qxmlJ8
/wioVboGGihKQKNC8nb9yhYyb/JVErjyHymcG75E01Hvenp7U3wSnMrlQgbnpgCu
FchitOzNys7pUPNXmeWjZSaxpJ4OIakFnwmNWW3McGly4PIkt5tt0oFXxE0fKroe
KpZjR29dBBw3B10JmjFEmaghdmXyD2V2X9yz0ihFCptO6UWeEqzRnJOX+gBLoTBa
NAtzdplUTNg4W0YAo0bvUE/7oWMO2jsFfMFzlQA32Re5YeiQSL3eSx6fr/rSp8Vf
EwQEISKp5QSiuJj1fy3+R7FxTl5knRHh+GYffos+VM+6MCxh2VZJHvP+7LC9U2dK
z0AEfX6ju2WjzF2vP0B+gjTXTo+7zTCxNlJI4OwXGxb5Kylghfa1IqCA3AG7guwb
tNATDma2UutAvUotTDeIT4yo3hDnGHXNymakTzyDzZR2icjI7n3uWilyvdQMGZqg
3QGeDj19W8Otalz6FJagBuC9HsFNPDfPYvmPQHa5QDnw/1GgLwiysB3MRbUJ2umN
xV6SMYmq7JIFBkVcmCuMsmEB8RuLsrlX/xkoIBpL1vRQzx1ebPAR8uyihz+ffJBv
g6zQKhZE3sR4FX5TQFFiw/PEyfQrF9SfCfn0HzziXujXoGf+uv0kElPQtmf392nL
Qkar8s+svXJUt/bttAgh1++aCRHD32ZwC/5YjoP68lyMIXwd4Vdw3AhIrODQzPYr
M3F9ZUcRSU8JIbMFriTrywZbZVKmbdaWkdKTDYLauN5p3q85Tebr7rfnIg1uYZwZ
jV+5Sp4v0XbignwSpWiBM1B3fPCZLgnaDb3+/q3qsJp9q2KISN4aVUmeRLT5TgyL
VMcwJfFGV+Y9OJ/WtsGii8SzdbOKk8UGqei8hvEEKwM5buiyKU8AVJtI1VCJF11l
p/vD1IQlCPR4OYyss4XIOQbranOCbl2gGPcpTICNXZhCYzM0mk0A1AzfeVEJXLpq
URWff8IreVGt0E6ed5iSikJBf/ZC458Ipi/Gg8WmW0epUoGG6ZH1MLzr77pIfufE
e1QJ5pct59k65iJrLNQOUvk6UZ4PsMOHssDqrtn+EAWZhgiiP3MMnLBY+roRTbPu
yu+Tqow3Cjqg5+73Mce3QoiKJAm9udnRPqcJb3j+0PlOVMeyZzbWoQAbXRbVHlNr
vApBjdajohoLCwfGfyKK9PMRoIzGLwi+9J5gnxw64rfEa+Q4Rf8uZLO++ycM6n3b
fIIoRMJ2s+LzJI2fY0SsM+OosC5Iz650cONQZlpSUhHmTcIpmktqQR76uq32Irm9
BuI9V+nzQjal1GAKqWmn0GUgoyr3aEhYVBEqfSBCTz/fiolUcOQZ00UrMM2ALshM
GBYX2IizR43KK/A0xCXk7x/EHpclONkoFPL6yBSLhcfE1W4+7rnEIiQMoxfmd15A
lfxZ5AVgy7jNaaiDVT7cRCyXaAyfgTsMbSQJb8+mzfLCoREwMT/nfdh5nnxAdowS
bc+IIeJ4/Y4YQYpM4EiOqB7nE9/GdFqMnvDgwtKoaJZoBAyCNYrwWvb123+ewrWq
T4jHZw/kj1E8ykC9Pu50k2TOOjhXEXuvnvpfDXWHGxizM3ElK1eOLTi8BgLEhUs9
TsxmLbWWL5Yupy0wk73oUsrrSwBceo7s/hfrW5cr6J8giuRLzkmDUHba55OubX/k
T6gHWYNy8dsvtv10jMu7+spTL2zlvdFSc176MxvHtot9o+OUoXWSI/dThuPx3dhn
ksgJCxvVbBnbZmdi+BseNKAOjCv+BWaDvT3R2EPD3ltxpv5Fax1qFyzkLermBisx
NG11QgSl7CAhaeaqhdwLtUBsIuwnMXNxXcgfR3L+EIe+kxMX2HM6CPeS3g4M+IXQ
lXxF1NweIUw7fryoMQp5IV1AHh2ic0+rn2GMDPSGr+ddK2A5/bG4tWoyqINvTwKB
p2rbqhZp5W8gOmLKaZvJPj4Y6WcN0kKju6gj0eN1/uy5ineKZiMrTFMcfMTMt5bp
8uctNZOJDCHF9uIuLETokd6apLvIf9MFwsV39NLaLmxtgeu84JVU02r0gWKV2EgI
LqWWlb2wfdXopWqq8HsBTqo2nqVvw6gxlTvuQK4bfnlSNocFoQJRmhkR/54p2HRE
cTFHS1+GD7IVs/vfzwt5Shwk40TJEuEYfujJLPJmiXWbGsnehSn+bJRCk4CbVY6r
/s1XnZf1MXyHoLgilN6YFMtOEkLw9PyBDOv0ebTW23JlM6/1BmphLRSSJscKYX86
0E/UQdz93CVA0MPsJlb9Qk/VzI8dtaXUGN+oHlSUJCwt9iPzG1uOrZmxfSh7kVtt
sLPcf7R7150LvQUn3w/83rn3tioy7WwhZK2zaJcWpJq+3WievR7O43+OALVrp9pV
x2ugIhORBroyDe9vUns5xrPutyyadAP055xU01StELr27pNnwtj/kE7O0OVQ3VoD
OXSpRoH+ty3zc5wcfSlcFYR3yTbQYkIzA2MUptE6BBY5YN/LlAjVyUTa5lBbgayu
xqBCVNg1/wPSpxHRsu6eXy4j5WGEF4JmakLZNs+LKT4JzrcRGrMHPGU4nOmsjyin
65GLGaYCQtsBzAXsoWxOtyOjwv0mMgZqsYn1u9HoXPYWfkH7+SzPgllS8HTH8hGx
HxEIOW6BWFAAQUa27d1/W9MnqVwXPoL+Wb3EKTeUB7/g52XzhO5y64VBRpUPUwlc
6BfL56Y1dj2JVE3oK75cHwNU7xFGQB+d+qNBvC7mFjmFuWGhBdPTHn6asUHFFfGo
3IEO0p/zKuGMLbCSH9eeZujlPRU4/UmGGeLpp1TFzttHtaohm2mzlThPnzP27UTi
fIaonKhI9zUaUdFWVJRyHlu0/DIjSYzIIbau0XvjZ7ihdYikZ/Obh+X7qDs6L2TJ
pFDRunwznKaXam0bB2jtV+KCu7Ff9cQsHSmmvj7iaZn43pqeG18L/fyHBjY9EcXh
wpeQobEggvTorb7rxOCy5emQTDCbvO1tgrUIhBlJ+hvu5a0LXZpjEJweBqFdWDhM
ENQ3OHm6lu6/C+FrxwGxT7rOL8QdT06PTU3a6bEZ80d+7hPoB6xnNAKAVSK1acvA
S8Q8jNh4HKpBTnxjA32WE4Ro9BTQ/DMOzpxY8jQKWsQ0WjYNqfbKBZkEZ35paTmx
bxAYK4/rc+0VhbfWG46JEfy0em2HhwcHh9Ge1W40D+Z0orTJCOfWiOhbtKfPAKmt
LnpJMpJ6D1vIdrq2M0UU8oabj8GD8TIFPt9iPAr3I+rajo82JzGbb1PiIa1KC/th
kj9NAyGI0gzbcI3owuANZXoK6d3TLbUFQEsyC5cFyFpQ25Va5eg19RbtIUkkXFoV
bpviFV001lYk2tusmMr2EnIZJWWAzDCm7aEoqzNpISO0PsprhyfZeG4iNDdQ5vY/
Z5XpYa1FGXQ5xlweoWKcgw69TmqjhYC0fGrgkij3rKz6zm7olwzJcMKc9Bwhnwi2
R9id8G3+xaaearHqUpFG2FNCHEsJv/VlZ60igYbvXS//VizbdGdTDoGf/0aFw2Yg
2FKPxzxSGopeE5jCDdlpFzF6v+tOJfFKRFesNsvUk05zdiVsMqNBAwUhUBuZN2kU
ujZCYmvir4COl1J/AN5BbaXCWjM85wYBpnVwHSW2WMXXsTGCuVBbvvKeuzR5GGfM
y9oa2lGEmbnWBt2dQqMvanZfuZxKYjjfMMtRYRbjY+FLfHOWKgJZIdscsbrpgpQ3
aJyU7LCXBxGDkdEYxL0a2h//xPin8cNOPgLo5x4cT+dD2O50hHu30A/gxNiWGBJ9
SzJfoHNs1pWJJemkzvPI3DFyYN3YtF8fZytaCq+RUKZ++bULQOj9VUPALO1QKSld
KHT3RUS/7YClx64h3HmwZFGbPGH7jVokqHb8jck62Ra7XLsc3TPI1f2Cw3oPhgnj
q6JTx77ezZS3SQXi+MVmUnl2qWXj1vLUaSJJU+nvQhCRhmbyOm+YsGvvOnkc2Kfm
CK3vGWRDKivDuNaSdJHnuXGVJxomCsps4Rp80cTzCVH9CTfrKQb7wZcBJvVmaBMt
x9KqXMcqSzH3xURTIlDRhyb0HAVPbul6LXidyjen+MNyFcREXTjB5Wx+dJUrPix+
Z3W0hQ6VqGNOMX+uf5KH750BK3Bcj/1EI0imWi1isHJVratgi/xD0ynrslL6vXbw
W0wuOYg7nS26QBl+CGX5M8TD/+ljtYJNImDJUveZF/bfKFNXba1tjnTKSArRhwNq
z8eZCvSpTWiEo1c5EYtt/lKcmocIHDKF7ANKutfpYBXDZiBV6NQZi6ckZ8K44JEj
gFR83x/VDysxESrBySlKtsmAP3MV5LOqkOOfo5pXUBENh1PNnf6hNRRzZByXIuUO
wUl9vGFeNMWz/O6ZPHtQG07x7lncIN14wcF80KWqlpiJsbzkMbC7Sy8qLYLDrtCB
j3fToDYtcua48RvD2EsKMrxDeFMQ7FLNKm1kZGUnZddIzfjO61khJvKJJRiSTse4
9OJf+m5UkwCxhCI7DmFE9KrEMHwUGb8tUKGHhpGbMeJvjRlOs8HpV5LOwLUwj9TV
ZZpqP+iuFlso52YuQ3XGoj8FUxx5NQn+C9r9z5K6PixAAQcmIi3xESoW/qfrRzrD
002P91Gnj13Y2fYxXwHVH7XtHgCUnxMcKmzinvS8NNQhSaJya6A1fEhl09sejCAq
HfV+msIpG6lMLSAtsEU5DmEgXoBdcuobyXaJlUYgKYWpYH1kkjOI8LwmnW6MBhWD
5dDdeNcjZIElosIZIVgAAfZaNkadA0Qq/enCHJ82Qje/KUxDfTEdgNJE5Ic49kec
rDJbiZQ7GADaE+1ZXTbX6iphyv+Kvq/Fs0HRXw/NBjjJlZC79Vao8qZon/zgKKPv
Bk4fhXO4n6hYx2puhT5V3JwhbF4SW3rVsCzLiI65YXAl9v29bYL/EcrSSvma7eKV
mv2HUFMUspE2TI6K38gVJi7Wf4zryy4u7mWm6OIo6Av0dYbGpPmMamO5Gdk9xxY2
969BGvfzctKdx+hhVhxO4FyUcZXLGMsKsBLi8/bKkFd/o85izev6vg4Rb2WlEb3K
XmGmtJGOc5HiRLG8xWlDGSD0Q5TDR1XKunm/tLzGOeLK3KsMJEv/Tka64IexvWQ5
nRW7l58z+ykoyq+gXXC2YOvKV4oT9bg/lvikBw9QGJojfG/Lto+Id7n3GCoZZe18
muH7AY2h9iHvmivVkNJuZKOruYfLle5Jeh5rOCxW6wUjRJt2okgLrgBL5JhdPPlo
B7lIq5htchJf7RjjFD0u/HIhn/uOv8X4MGXPqNqix6L+Nm0kepeO3RZ407mC3WDr
LC6f/jAy8PF09sFGKyBUo5ikO+wOCsvdiUvliGw5/7aQR4n8pmnQmEq9iGoouUgN
NmBA13VrNQLFkcfI74D+B9rcKQaRTCLwOMfGt9LOOlT3jJJL5G/Z9XmX8SU65v8W
Kez68QBiTFoX7V4JlS3h5AdYxg3lgUle6kEVmjoCO/8KAoAn1yY324gjnMx2kcFL
uyXQMsTtUk7cbLNoiiEcITcMYO+UceaO+9eWaYQ8P+mYMglhV6QD0fb2ifGO8jGA
OwkOfcBPOrKyL5+4ZXHY0ij+zYB/K+W74Mjv0NxVcFAw/LA3082QMHEGFNsaa9lO
bIuY8kc5/BtD5v78NFP2U3Lp2VZELPmlNLUHwyTV1HVuWmMaXvnH3jwEybYs351E
+Ma7ArBROnOAIV52YpQOueRYBrGwiJvg0lKBTrtmvdjQNkzHZN082q6sw10lTUr+
/AAG71heiTlZ11G57AppfWmHmZru7kQeVKA3jw9hW5tO9bNX7GKUccrng0BWl4bO
FpfGZqKESadepodeQTZf4DX5HwETJITq2ch0x6buIGye3DMPGzGM2O4HeOiYOckU
d0GBIXvLfA3Rg6aQWraVVhaB2HuTrp7pW6Y1ImGwPavL8cPWRpt7L+za6V+CYT4x
ILZZWGs6cCHK69h7HheFtQbpwFp935h7gyBTxN98YYlO1zp+zZwJgsI72G7O1jlo
92xTZ9bG0r0OKPkREC8aRi+uQhrSAlbfGlLvtGRfZ/rx8RsD677A4v5seyzG1Lg/
dMAPem2uXOCTstwhYnF2XdXyIvpLSS4pLRjUTezjV2u2q5QT2nhQr1kz0neijEVD
t6EvJXqERhakzxyZStHF8St/c40/8+wY37eTWjJGSDTeVsd/SpK/YDDpWW2pRnVn
QCr7DCG8QP0T8CzbSAuyfLntxxYOii8hFdx0NQPFalebmHSBJLmW5xRSTFGmuI4q
O6AeO9J8d+j8DpLMvDIyVt2a6ammfGqxLeUx8a2o3jul679mkilaibQKhsKzt9oH
S1GO3RBrWgSZy9NSmGdokQ3yYHWi+KbO1vO9Sira3HmorRVmrPbb4pa/Oy/hrhua
0tSdq0Xw+wUGy7lRt9ZEE5NacrjZ3TWaAqoOXFmgaL+XWTDbkBTehSxvUnkJpbJH
Hi4mgsYuGhmgs+raW26afgUVRrEonQlzSQGo68rQ3fJsoh7oIX7pziP/8StjjsPc
8We/LWeZgN1M2DhcPwRQLV86ycunYDfd5oxhJhQPKQ6pU5+ukrefDhO/W464ZMal
gBEwEJmnQ+/YAxLf6tOVXQEdkEZei9myg6GnwCS+OMl/wyapASh+OTTlgCaLa2qi
dav4SpIIY9nyFRr+SSCV5xvLttS80WsqX1+2h1bme40VF5vp6DWp4YKBaqXWiAGh
aKpXs5t8IX9fWlDEZXNiDl9qYiGMi4JsfLXgZ/ZMlbslr0CukfZ+vds94Ao4GUUF
a9RafosM2hOUcJDU0f0NclwhXDx23uqjnpGwhHsDPT4liYRvBGTdv0UbDWDUQmKP
NHHG0S/GG1a5WLnxK9voAIV4R/rvtiMl0HNjxodk55oBwnLtp0ZrdcXpsGa2SYxg
4rVwyYKMsGkuOXM97UaW0czL9s1YyLHh6m2lWmYuz/7rbaGZQEZUYonvBviyyVkh
TDkvAm60ww7jFt99d+8Wodb7797BS58uqHY9kpxnEOkkeKXeR7Ie3++Q+c8rSkAD
hnQBHxd8DrlmeM14Z9jwqOqhqpAHWh/XjWXxI+RTJc6IZk679epw+YX/Zij8bsf4
mDbOV3WF9k7VlwT+B0Rjx8RqoJnTD/bLvljOxo9a4GXeMJisoxhV8p29fbYKfl4g
zC6VdT3HLOc0Da8yzqSZYpn6PlwqUbV8eiulW0EArna/r7QFRm/cRQlxYyJovsJE
IwwKFsBhkjP2pn3dV5ijDk/af21lfdDZWXVAsOtV01QG2vtWJFLCrrJTWnZ7PJyh
BwiTnvMU4ECa764yHxwjF+ktrc4Ev3IlrjAG8ydyEJInvyXzvU4DWb/D3n13GfoY
Tb5kjS2ysCX3JdtT/QfvIvZMSOXJCumJutd3yHedSO8xcBsQutUlp9Ah5hbkyDjk
czkP5iDU4k/TwRSZUZTF1vZttcjyxhdANm1Sjmd2zGa2ORxF4T0FL+izzsi9O6Vl
3hX9ROHD18tzKjQuHtykF3Kn0Ld3aWuLK2NT6xp0gxnqhHNNr5unGRr4WGjlmh5y
w/up08PQVUFDjbZkKCdFB/qgTIq/ZcqWkxoWqebKNu44oqPOr89QAN5YFBdn6N+h
4te+DlLkCihjtgyfOj9aLuDBw069vW/62vF4C4U82//ICRZ6p0yQ32rCkCl5RBth
9VtfdS1ZRSO+J/ychBWveJNofzd8eAzuz/hKHkWsoK3UhEhkOS1q5GdpaJ7TzO32
oCOeE0hKzGEmvwyo1zgc57E7UQ8mo+1BDXFrAgJEV/+zwbI8wBCOK0b0Ovi3YbGt
bkYD//VxMJEmGDR7KLSSyQvnBcDIGX1PqFEhhGoHezOpJAEyZCcQDkO1YvPxB4n9
rUjJ5r23utKK0cbFaV7qbkQVKkqj1qIZhSSZNYNUw1a9gy/6przidvgwE3mYahj2
uvc0xl74qfpv5xeg5Bv4RRWMU9PyVJCVG0WjwLLJMKjD3nnvZcK+IxVYEya1G9TJ
4cU3JxGXP46cJquay4YxTel2GjpnIuc+Qsqgon6Fi6zYueVEjDavgQGwbk5mF/xD
ZuLxVtMnrOdNAhzjauizCTPGJZEjY2rIbPq5aCKZgksd5Iv/dqPnzEvkkOQsdztJ
/j7FS3p028t8bwpz0znclh1E530XW6G08hx+WFBzbaW1Tgme3T4XUdVxpKTe5Q5N
AdKhjP4c1taU5YH7sMUSRt8uOnOeba68X1MuYjD4s/mKBN3EDzhDv/MqjhzYOqcp
O8gMwzeNgd+kaKfghFTr6sHWo4BrSTHMjbrISFXop8THS+mLL6fer1/EDbTDAqa1
wxkDsjUpRvniGcbW+7zZbezE/+yUbaCHtAG16d9z22hQMdyC1cHL4JkU5dDjr9kt
Z08DY/Yg56vdBHBI/4+6gqbq20nBd6r67yPQkgG70G7Pj5N8JLPUVjN8ACzCtvMb
ugiPdbCjtp3fYfINm1AnwvFs2xTVqcuT9uFnbwXXDjZY3gtAWWOwPkHuyVqpwLyO
Lpx2fOiZvX4STcAdCGZXMbdgJDnMmv3HNzn/x+2pVnx7HQPLEv1rca+tHKmHi2p4
B/YG79dc2Aiu/ENagVj11WE6HJkEc1bqO4bEY34VQ9xUMn7cVfEf7yuv+ZjcySCZ
UW8qiWQFdUUcDLobXOldvkTpcuvTfOqhAeT1/sfjaA+Dc6iWI6hddIcPsLPxTKzA
cGotGTZKRlCHMqKaPrYpilD26sWMvwVcrVEljTo9sqje4J5RMSRY40S7bfYe/+he
ArBSmXaJzwI+VWMMe8caWaFPXG2GohwQ+x9Vw/D0yVyoEXV7QPwgw21lj47PEwky
xB4qRSHfaN6lFGr4Z1gijYtGKADDI8QcEPKFdtgjVedbg+Lm86mtC2zpLML6+8x7
UyLa3zY9op0hW20k5jaMkrxLaxEYBiPMOOiR/PZn9XAm69YDWO8+eGeFrDgJLkBW
ri7F4dz9bMJqBcvx+KK/6OYAil364QRozhkOaZNJ7+Brj4k1eAwgPRCFEeenTg1/
gTEaO8JFk45mfQPOhCy7tw0yJJdCRyZfqLabGpnY4DYGdCC5meG/F7A0u4oH+WJ6
5BsK2b+SIDGZPfSqvW0tRM0ndo8heER/MNBleQs6aZIHKXxN4ooVCEU60lT+auNc
T+//j3vPQbS9nzYb8GBmnI2IBeplsNCfiUZVA4mtETQQz8HuaNyNKahOs7yVq/lB
PrDmGi3JIcA+GJgBUD360xx0QQUS+cX3q+rsEakwv+0kg6LxUDo/W8qpb54eHEKw
VOx32/plWTe8cIcRoDXcsbGn+kXuiKN3DVpOFhuvFT0AnwiVy5DvtaOHMWzkSrpx
GoXW/EyVEMqh6J+8D/VZ2lZOWRuUsFA6GyODMi3PH9yxeBAl+q6sSZaGerOMpZoc
25XpYk4d7STGgjxbQBuj/+GE+GALe5Ps8rv4poEDsHxobEayej0fbm3Tu2AOM++2
sDzzGhCKe61zKAYiFN1n19WWWsKoZbSPbwzgaSN2HpaOV+2DP4uebMAZCq1XUIT+
Mq6mPJjJooGXqzNNahvHFQ8jxaYRUPB4Lw61LfMASJ3jFmr4L5JszuLwxmrvwIox
tJTETTXojoNuIDNZMt9v58At73qt7oW/SsLkZ6K4VhKC07DECrdHvzxCKlOecqTd
82ZoImQ6Q2hnhfsMsWKD5gqJIGs36Y/30q40DQfQi3dRPk8s41+UYi/ELB9yFR2V
`protect END_PROTECTED
