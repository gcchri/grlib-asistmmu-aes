`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZuhWrLAA1nnsIyAozkv+aUd82MHJt917xVbx40tqjAQNThf99z6OAwebvw9MPj6f
y3OnU4CkrLh9+QCePhPlRkXRp+vAcZbXjB9SA+xb22xbc+gR12GSivE8nXnJYFjK
XeCJmJlo/vdKEKiiQPuA7Qa4tgk8RC4ZqGRHbkHNAqbZsYMm7UerXkgqJDngjitV
A9JfLYAxaraDiCLH6EyLt1bHighzMmj7UUdW4kI5VqhJoSfijJxQxgzqouhj6p8X
ZYOolNPt59qT0U58nWDTI9asEml6P/VUPiVbFIk+7bRfs1Wvkfzdvq+yCooR0BqN
qqWjJyVXOMN3eBWwiNwsljfbHj5JjYMFrWkIgTalgl7TB3oKSh441G7JHvjomhBs
O3bGXOPLlkGaAeXMbcwovDn8Hipf7jgCoTrax6J+c06/rUBaGGtpQ+06jMMbxPfc
hsw8l7fieTUJtix59jEUtr9CjAK/MwqL4iqeTK37okgcAe8gJlFqRlqD10U8qgCi
7aH52s31lYe7W4crGpmsiW1q4/tl2QsnypvbBM7jT52QonoJdXMPrTeQQQJkOli2
PsPdkTTRfX7W7QFijHBt7UYmce4MFT1xPxvlVl2WpfIHH8OQdnmAEU/U29O1/VlO
yEcn2wHT1RgO5u94L5TU/CmhayRTiDF1V8fCGa9EYGnLfu852XK2ud6kLTa69+t5
`protect END_PROTECTED
