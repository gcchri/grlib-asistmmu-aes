`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/XJIO+KwAlPFx5Oo+eu5XGae8rvytXMMqz3LHKcZJRLkjekpzIVqduYjF+CY3mGh
HuOvnOkl2fpKzMr03mnlJ3bWcrCwlxUHopYrjo1pNZnVYSFWIuscc9wriwivx4zH
pdqSehAY8Fo8LLzwuAyBjp9JghAC6WkwkGbDpQP/duWLPuu57ATO7UhSYNSb6xJp
hRcM5Wmcfi8UKrRHJer+FX9z0p+os3vdqE1bG2DLKKALXpl4gatGT+tiYCK8p0Bj
EQXhdnJTjiLZ717i+53BGvYmNGEh0weHvDv/JyAX6icj9tPhI7pDOS0ANg+bILMB
`protect END_PROTECTED
