`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ek6r54MUEhNIqX2jTtS8n1OR69uXO+8n4szK+GdAJVpamVQRIsDi0E0oohPFf6GJ
obU5TjCwPVlb6nrT8IaKlf3nuoqncE4ddx5ZHmJoq5bcjGqhQMmTCkrTd4PuaiMu
d0BwOemU34onPRsOnfsS+vpoD2luDWwhQJ4x/rgMEDLjwjQnFcwQpg9vBEkMTVjP
VaG/i1IfPQKtIr4DxWm8palYTqmfvASPCBbhb1aYn07xdpz7RnoPtJqlstsgP+jO
TNCGj2saJyGclGOBSZwOz7Qrb6jugCePEEgewmtXsbH7okboSnh9QAYyxa0C2c/g
da031ssB33Uy6wiOrikSKJQaD6SmXe+0K/18j3uCOgaEo3aEEAJLAE2QzFTWeLzo
NxbHRWK98/9PxjqdqvWp+0bj0iPMKVIQBeJ30sPtwADKKyKUqVw2PYKaAIOh/xAZ
eu0HuLNYeQrhP84f21TqfSCR1VvRgHmuAMBrMJc3TJa4LY+BpplHlzTG1whn7Y/M
JhwzvtP1Metb6xBRaFQ03q2JnbdaQlpCZQ7mKM9r/lBI2obNbgpBAR19qhlhvo2V
f9jHenZx1Y4UEzu07V2z1Q/BvD7xjsDxqHjCTSmxz7qz14XbVtGzGjS2Hlus1UpS
Ruv78aBx+RFd1BglGqLL8FFSXjkneV0Fo/INKj//gQu0j29cGSwwhdNNPwiaeHSF
sd0A4jcnLV0qxLjTv87MF38dfOgliEka9PrT4+7AxRUs2IzyUrIpcZF5IovY3vuI
EeRd5RGpAywpfhJsvdaLcLH8u+svtfjsqpwN3GiuQ0hlvM2YqhNmzjDo8eqVkT6H
YeUz50mGX2aE0Cg/MLG50HB9FKJ4kVEaKmS1kTNHxe27NGq8/XXS4zKXa0fsqLo8
6NNL+NiwlE1wrwvpRlmMLBkUxUQ/mHN+s9KrmAkGRWy8ejutVzpUnxImuAa9xkiz
VyhJuM8cfnEg032/BO4kTDVMgmXvSeQ3mpzS83MpfeJUNZn17NufHWhQ+oGblVKN
ps+fqYkNTyMZo9vLmJDM1S55OxjrWCoT9OEYh66QI2+UOKczF5LaOAdS/F5Hsnj0
DxKW9dReAqdVhs25fqT3aYLJG7jXXvyHk9/Al4MW/FuWynMPABXok/doSXcERxl+
1V0HfJ7YHBfhhPEXSdhTPFt9m5YoIEMC92AK3fbOe0kanhhK/EXfbeLLdlQeKGWL
plNe20IOwBwkgUvdvGXbWv4SPKu8RRblY9+J2z42KepE4sEsIKi8G9qQpX8TV6no
`protect END_PROTECTED
