`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AcqrzwI9geKTVwO6Zm5GbbEMRVZG7bKnyk33rDcTULkiLs8VCDam8DiB9Gq8TyHQ
0Hktoi8biPcId5uxy8b2UBpmTxgqYlh8a4aiaHlNGM8g4l/3NrMyXVho6rYA+Vn4
f2bBRvAsV9r3bEW1TwMVtiDm961UMTuODHDNMuax3UDGQohmoQ6etLv8lNcNmtAh
/uTw7sI6MOuxtcUMTqAJ1M2jQ/toE9G7f5MEUhPoylpCFRfd2o9Mmi1TIFthz5lX
Xp/cBqfQD5Ave8ycDrRLOxMQcnzAGDPxr3d0c7rCZ7u7TrNj1qLN5aMObxocnrvS
usn9OyGdhr1QmuHoL8M6IQ==
`protect END_PROTECTED
