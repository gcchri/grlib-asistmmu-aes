`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UC9d6Hxz76P8ZbzWQAgbzEu6zeYSZcG4r1FVxm7DF+Oix7Kt7oOtCZJ5fcb4f4nH
PeWqp71HVpUo/F1uu8Dpxp4dnGMKH8LL5WFGP3Cee/K1rDI3EOyzHjZibOzblOGZ
OW2v2LX0e4AKXQb5e/Jx2rCU5s4ugnFqgeLDmxPn4xa62PytkzbEEMQhW/7vnr5P
miDSDyaKVvQrjcokCoiO2iTt0jbBTj9ZXiDfYNL+PnJNaBZre+ueEgY+nyiMBNtC
Yfgdjb7Qw8IJIkUWbGDQBvudo2ZeQSywEvL9FWW+0g3jaj2N5jihMbJFjrTIFYy6
3n8fHsCbi37paX8dJvwv0bXnhxUDexP3niZgQbrbl+aBhThKHU3CtMpoVWoNmL1K
zthV/vstlJewaY3IE65iemFs9rh/jwxycxiVbPfbNPv9iuWydcGFqfedhQuxxO4d
odrUsR0Hn/2VFgaDL9RPgepdPoNO5ZBrxreKJ+hVv1A2tR/GUWOLLRpjPTtimHh7
ykKCFFVJJEs6ZgR03+DdHRLOCZ3ptOy30gMGFMtpj0EeQcBzIYgOowLrEXOlj0M7
p+Cz+PlJTLliKr1w/CIdSaS6zKAiMEvbUqdxk4vT9hzTx5JRSIFaAqsLK0YX6Tn5
3YHP6mKlvFWWoXrzOIjJq92mEG3eeJsbn8nxzH4SHCVZ/ASNKdm5Oi+pJ2ZUnuJ2
5CVCw2/oFk57+RTGHko5DyIN8fI89Ow1TxNdtpNWw86x7U5twXdklzBdofParnoT
gJ3ZSxySG8JA3/+PLc/OZ/a8908mtlp69yWJX6b+TQS5kd6VGzNMdTrnwzutJWdt
bzO0y63o87tDqJ86U+Q4B67GMoJ8Ok3RmpTrykTrcfw7alhrlMMGK3YkR6dYD0wS
BFFStQG1/ikH9asaFH8dVFDokTsLPZBC47p6Zq4TUdkQ2Y1n8BB8p9xvnPlsLF8S
`protect END_PROTECTED
