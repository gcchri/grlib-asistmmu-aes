`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lU6Eycco6DMN7GxGWXE1mrhYyCJhH6B4ankb0Ovy4ZX3Fwdn82e6vi/LlaTbaOZM
Ebw6KYWvE85MouzHOWRRztnAuLH8eKmsJxm1FzqE70Nb2bDa8ENGm6B74MWuZjMu
uWvWAPUQ19fvnT/ufs0xjR6zTxzJOYdtqjqLjMfWN41+pFiaOy1/6qTKwe2IfUpK
/yRKHfaA5cIBVIzkYQPrA5phhPfUlKRlKtFY3/Opcva0Clfuxb+lZTO+0zltwsn3
HbEdxjCRhvR+f8IlFILRCDgwWCecNCNoU2IgvqUWCDNieptWSBwztwkCh3R0L8KP
/JawndM5gwdJr4K9oIxy/PQzAqFbb2R5akrpzwTTfEm5zydQkc1cAZPK9FzEN7+r
`protect END_PROTECTED
