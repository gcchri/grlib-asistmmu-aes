`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TtzlSTJvy+Ov2Y43FiVLzVsF8iCYdCHdB34ivJUW2N7q6tV/fXT5mJ0nD40DjMvG
SwjQ6fXpjn2NgntzTa24zV1AFISimxRWPCDIg40YOL7pCKLRUBlWd+6asQyOgBOG
D4DnBapCNK8mBizwKLrU1zpRf6DfMKkjmEKKDCf5/waBUqg3+aU9XKM9U1G4aOGu
MIG1AVaaYUy6yN2ng0vy5A7lxLs7ar+RMQt8G7rQG3tRJMesQHCfgI7EYjLjSyoC
H3TO4RABC11WjaWaswk+EzId1xWpVl2bFcsTSvKv0tRQVSiSKJqoQzzrOvnLXjSz
rA+7m+i71lYMI9jmv7wrBDrmaiUrqqQ2Ub7eV3ZIVVv3aGpyx2Ev1sdM8Elh8K6r
iCu8gbCEQvVPkurPocWWh2P8voHMYXIf54lD2+mZJg5i3CfjkOynZgNUZQMV4pN9
WuCm9JVGSlbPCR7Aow78RV3RrbHdPEgMKkgGYLLZuwBQOywb/eKX4Onc0RIv9LSt
M3KkAqsouA4bHJ6u22Z1cLkIk01YoIfd8TT0w8GObo1a2ZFKN68uRZXPOFXWPfx9
/Mq3yYDzqo7PrlsKKHR8VUaoR6rDsYrmTqDNGR2QNF0FylYkK6TRkuiW/UShCWkh
2jCM3x+BVABTT2cyWq/MD4BLh8Cf6gfWBHnuj30RuSC1gaMCRm5EwzH2xY28aG93
VR4gb69KcP2d87c4eglMGgH6J08hqjou/xNgXuShkvC2GpeWp/EHdwfxqJZtpcPR
jdlmGBSGMxJbWyDNaqV9bZZ8QCxHwhQ/to49yGyhdD/0rVTMxhT4p98YFY9AQDo7
/MhYagQcdB5Tuz/TqPEyzCJrYv532hF9Xibxtq1P8BU/DQDpFEuIQjp7G29uqIfh
FVDISNfe/NVngHJizbvaSybqOnu1kYzN3Pavs7i1ZJLRg4E60nKLN7EjHCqt7hhN
ghxI+TtCsBuU//FGpWEo18GBOG5x41wJV2jCPWdVM0ioxAzNAtXsozQ+1tMPoW59
rCijKY6J6WyY2RWhe0NqD9fU5kfi0XWb3FTAK+Rxh5xeGONkyKPqWFObAm1oC05L
LgJ/DdItutwvLG81s3mGmsNWziHbmuilFy6qjk8+GGUCmTgl0HgRPrj9sxiOyb6U
xmcLo1r+s5aXJAfnUiYGKGpXpKflHK7ZkiB8bp0r/8R18N9vu0JeOyoXy+6fXK8X
y35jhv66r2gcCCh8fkxHS8SkIgPYfwRanzEhz+ChmrUYAAWflmOlBw88mrUnY1s2
X/LRE3Ayhk5s/Ve0mIdnjKa7NzLSUehhp8ItwDsgQ3AYwstDUgyadUIlpTGNeUnt
M3xmCAf8Lv15O6i/g01fqMVzNuxI2n94ft66O/+qY4GJ/Anen5ElhIwrTo0OkdxF
X494zjjX6mF02CxnLJuXK8oc9fIeHufJ035YlL+wA6g52l6L5XF5L8nPCtMz04hM
DIfAA5gK9ERizY3lE1Vc1UR5mM4ROCXNY2jogfuRGuuGYcefA5qi0EhyujnO2pQX
bmPJITmBYoI+GcZiq0bzsZgVdk4lxwknjSuMK7a0sEea1Qb9HKhjPQb4BqE+aKVS
kTF1wnviiKPH44GJnOJycB7HdvxSxjh+gjqbpRf9X08psc+zG8cMsx8c0CCayRRi
yOAf4BOHIj0nuv7ghCer4TE3DNPLniqeSEdLWnKSGDviSiyD3dDhUMNZIfSpme26
JpA5joxr7rUdD5+74v3Bl/kthFjfWc8iJwILU4v68PIOJt6okTuvw9uf47XmCmvg
`protect END_PROTECTED
