`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bJXUYSTDDeg4KnFmIati4S6gVKtkSCaMsXW/xYaHjRyLuO149DmK0En3R3XN436b
qaLshJdrPgsT10axB10SoFkY9ayTXab7WfIdd9FPI4aUfqd53zvj/kJkQWPS4t4l
oejDKEf5Ypjh9bGMYhjm3+KhActJ7wVYhufznoeWcTdpKkEPkmd6+BPXRww4onw9
E7yBSBClnK/IFgnjIG0g55W5w9j3EHQtcCR/ydJ5DGlN0dvJmJ0DRVnk5Qnfaa+C
yZ8/gswdOdfy9VkF5QIb0O7y05idsMW5B8+tzABoweXsgws7qq1ELjGmF+ROjelm
J/JsG4MI1tNLp6mQX/Rrow==
`protect END_PROTECTED
