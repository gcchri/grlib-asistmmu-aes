`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pk0bH5vaLxjOqr8FyPs660iv0fMR1qR07Jar8ASfWITjUmPfxFQHoTGJRNgHoQ6b
A+6b1Ao/S0PhdjFDHOvMok+2LXmaLui7daTkNXRE2QHKdjtkwxQ9Ch6Q+rk0Nn6z
VPif/kB6rGYJw3M9nxbo62ZyOLWtAe57QnWpcMZcXfs1GRHWxvH0telScsFNvsTF
cL+F3jgS6zXpTK7CKFeXCt/k/sfzV9PPzOC+5q9aFlHjOfqCmWJCz2pKt44lv2Zl
W47v2uTOE3QvAxn1vjZ34j2+Ko0NMlDCbib9DTCtZRW2lQpkT8mu4LCGDXl0zaHj
l+X1mwde2kkVtR0IO+zACqjkjZUATXzdkffMav3iuwhJqOYW9Twtl+z5d7MG4eMa
EZ21Y/KTLb0pqM01p/URxw5UH/SwHv6GoXzz2+AlAoMVsIDzmzikBwwIZwFRMsLW
Ean5LPdw11lLR1Ap7yPUdziCd5KQmfKurY/Cw5JZMa7gaG3QUTk7dzCLoKlw9S1h
zaIQykssN7yAfGBv6c6b3Oa7W2VqwIZIZ3pgYH47A69muxkUx08YaWJim7Op6Tkp
54ebo1EGmAn5erQKSZkSwrU5vOvXEHceH9k/NsSI5v4=
`protect END_PROTECTED
