`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kLD5UN9VUk1aonOGsMQm7QjPRwQ9jZPUAN1tD5IcFeN0zWjRGcrK2vS5kq8PMad5
wAqjpqaqhMrglhEh2jzLaiciG0WcZCHa0D+2U0QeJwL1NPvIUh+3g0XfU5kFgHUl
WQF8HThmYfqc4LJQkA5P0GWoBiKOA4iKG+GJDdsmqiUHbAJDdpgr60PkWhGhY+pl
zAeaW0UV5xACcGfXAFY4ukEt2PmhGXFA/4/NGaLb+2IMDsgQcfWSVqqShToab0Ei
ha/obpfDO7lSQ7Fymy/+ipcPP1jHygonI56D1cc9P0Ix8I9iCtV9JzDu1JqHwmw+
LkxfGf5oKfe4YHO+4aT0VSUmKlZN37KnfI2XqBhCmE3rrDk9fI93YvTzA4kRBbYw
GZwyW7QwxNGq6BwonxYVndAfFOFLDmRD6hrVsBKpjkgmGBo9ZRM+L8mZ5pLEzXQl
Nu3IZpuG9NWGUWZ6mIEVoyPJhk6KIwEV5WFPqqovnIO2aLyZ4mMIJTQ5Hkg/V3Rj
VcyUUoWMMb7y/ohofUsXASex7XpAaDT34L7cANmzfZ7syQBAqmm/KfjMIyTVNgV9
kPK6L8KBMmRr0NzeSSpRdsWa+TqtuMIDlfvU6CF56ss8oxGRVrwvE+riWvtM0i42
hTvGx7anYmgzmFnDZ7CUqjnxshBQS5mXbw9eSeJ3HJvUWLg2dH4sCMzHt1oi7TKY
UZRYK0OznEjkobW9FJZMSYmZGKzD9uoA8AYtot9PXZrDZJLWl9fnMD9jx/SsfGcv
Ryrtf1f/EJgMjrgbWvnYGuPAC8e5BgfbHgvUWPgg0AFyqoh8C/39ztCHLtOQfN/S
6/viKvj62dbzVTVt7QhIzyX/JhOl/z7avFTgOmDU5/wHfeiMXXSjStq+z9j1twQL
RCs3pw4805JxjhUSpFJQzxRWGYrHYYrQdLgwX+qdQbW5OzWIvlRrlQDr8JsnG1H6
i4qcW6lym5qQTFwrCg+QrWxM4wmkb7XmpZbgvCBqYpyIr1gnWuVwXfduIXdYtUTd
uFuN4FxR9/L0FckFBrkz/yYJeRVXjEMT38/v5G4bP5ldKl2WOy45qpQNmsWof5VD
Ii6Fhv6kg/gyQdKM6IOqrYBKMg8T8rTSBlj8XvRZJ1bsFIU4/PyO+H3lKYntnPBt
LVre/m3Ryvwy6M7TGHWQ+0tY5Tlz+JHnXASn11NkvaKn9oTBwMNfcwPT2u8tdNoo
kHJPcdmX/hxIB+we3RwQEnh7o5xET685l/8088uDel/45t7ohnKz5ESEnw6ykQ6L
4M26CXBEMm/rbQP98EjpVCztXnjaTUZ/xQfpeZeopGWEp6wLLhGasksRJp/hjWVR
Sk7zxTHtZSrRvOyrY1cXgDBZPg0R7E3v08+ydZZ1Vrxn2hkz4hcAi80ufsUtA4F0
fpJGTmA8Pf8K/RGGrKCfZs1amtLX1YJc27QGqTkawyFcAv6iKOJDefkIT5IAtkHt
or3YdZlnPf/zbWsasXB8fj+Pt9gSbQvok80T79+I3D/ocw7FhyRiATBliaG3h764
MC5mXnQb1Hnls/pP1moFli4p60B4Hxw+tYkpkcdriMT+MGRSc2M1ULzBlSIRL8JB
Rc91XSQWw+bxblyZFqUNpf4tYgV78bzU8M+xYtAEB5zseFFW3vcvmgg76+VOvJ4G
OjuzPCzU3yfVqHbsdA8eYvz+04Ch9GgXdlZwpNGK9O6JODkFdMTCs7iHhSYfI4lD
QBwRaGbbSV+RPBUluY644RNmTTq1Djb0qjLM5aCMARj6sOyJHsIIzYGzBLAE29e6
zNV56I4R3ukEVZPmkRl5tAfO8RhhDE5GPymEfwHuXFMmJQDfDNQrKrdX0yTPKC/e
hHFHEEsCicEu56Kx+CcriaFW2gPQ4hg8OscURC8rBo7n7Oc5ZUNRUFmnutEMDQme
8hzRn9BvSKMOp37nGCIdopaSemXo/Zf7zzkMrYfkY3xWT3bn/zUke70dVQ6vy/oR
0nc9UDjsoPUrOLGMaoAbasdpCHXEv+MhzHg7lM95kn91LySFh4T9vZLECUxP/3ph
AQy1XVAA9v4XLP91BYWTOIAkl2o8RE8lwROqRcZMBFEursoXrrY/BhGbd7JNtWZF
Z4wtHReWc0aJ4D4RYCRBex4pg8YjstiAqyjN49VwyfkCKQGWpQpuSLU7ke+jgUJw
0UIDRGwoin3LpamK48ZoZb+rvJr1U9MacS/EmUm7yJXDDa09E+p2pTqadUmURLq6
kQbNo/uOCdzQaMDlsaVQQ8l3j0Xdxh465pBZfLCRq9ncRBpqeMnsV9n+JXvMwNd/
FknpGOivWcsJXWvVoX9PB0clne/es1Ad05UT6wY9HMb2+GhSBhJoALqnmfRZNmW6
AsQiCAy+IOXYq37/7H7IMuUeDFsE5NiXC/dghcBBQsEdQRHI21byNqlij8qJUh1+
gwxve5fny9JSF0eqX4S1/6ypGeQFzxkDD9vwlo4Z/AYStTfC4JpjN+NG3ttkBhon
GTyiPvQvW1cSDYa6ieuxt/5TNgt2mv/KkHzX4wdbBh8kqD2EUc2rJ873qWsWMWLu
18n7DpkPDP+pfnzR2wV6tUSnoAqfoGbTCAnb5tHeWJjDfLeIhgkMp1gVB4osc30J
kCGWLRxyEBCPfH0DxlmcP41SegzaVNb+ZbKXbQa5kIOASqz+cJv5OEHV4Vp8vGAJ
141O+G9M+FhMi4uj6JVku76vVi4H1bFTGk96Bk3H2E76Wcmu9tKsOctJu5FR8dzg
nZKsNJQl+rIvJplGNCD8HZkQzEZ6RgM5Ay8g/chxXCfkj9re0OQD+qcUKa3VOhDt
A+BhKpVzexqVxbXxj2Mr5oUeStGkcbpPdRQizq3oQwD5OHkQ9DULO+nm2kYaAXz8
MZ5+iUolJ1ve+uHOrqGPbbwc7Rp3LMQvYK9Ob+x1k5xPbpLA7asVTolFDMNOPBPd
cn8d0S4dSqUS9DPjGdtNKQ4G9e2+v7BPnIxCnI4fyf97hbAbz5XrSvLguaoZzjxv
c5NEKr4DRHJJRyrjIlaGGn3wfu0HDwaJU6lfHjrsA5Lx0pTKM2N3bPboBNcw9Iwk
Vw39qKqwjYXnWI5D2dxsrwrDOlM9OLNmIhJ32PzmRBKfl5LJPPBwDszWMjuAYmf1
weOPtB1aUvFEYGi1MbZpsJ0thFYZOmbtCwiMFTdrvw2W34V2APbPDwo/D7eVndKy
WqmImAFe7hQ0fqDPSBLN/S6VEOlqZSOLOGbAffbApYIbhQbL3hQ9VMrcX71ju7my
AGKsnJpL5CvNhmmTK3tLZy3dY3uRcWKW1SOfOkcI3NhTqY9rMV2oclTMAHeykdQf
HxXUOB+Y9/n9G3midakPSJ7uNtyqpKtunJjT0Qbwz+Ph529m3KXP/ooWQXZ999tM
UMVj3YEKNUZYtmF/V2CoI9tPAxiCqqiVpYqaWT+jU4QUqS+FjJFAfiVAf1+unK8F
OhumqbIRbMplPfsfkZnGXVB8mf8gh7903pNRbLQ0qJQ=
`protect END_PROTECTED
