`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z8BK9+7L3392Tf2CIlEtE3CfIHGH+83SHp/jS08I6FttEeR++O2ifKvb9bW6e/l+
4DcXCYGaNe+Dv0TJ0ij8Rk8QCgnbcUG7swps9aR4Rr+w+y9EPvppsuwontw9msOS
7BAwN0mLaLv/jL3t8ed2hyyt7Wksc9TFPZBqQHe/w+l4CAVsBjfmgHkreBVbWChZ
Id/mTEG07JrRul5/PkWdScz/oGAaseJjjVOUKsK0jkYjQs00FA4J97PLGKH7DVDg
WqXpKRHy1xUyfXSOZWKESiqQhgeDkcJlxTUnEgOjxyRWBDCGvHGJYrIOIcQ/fVgw
`protect END_PROTECTED
