`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2XpWbWM0eajZ+aocfYOAmNFZ7wFDWRQ4bV9ud9wdNEnf0WwzDN80Q1qBd0jq1eJi
NOa/KJ6wh20PugWcXr1TBAmpXExTEKtnFdfG/hklEdWibx+KrB5lKIYUNePkJCao
hPPvTyijfW/MY58Ce1q6+84RALKC+6c9Efx7/CCsPDf4IDeQTSF85kEVM8AP/yFH
XP/6sAbL9ZtwJPqg4pX+WBED3Y5GkO5hxgMfvRtLYsxBTVLsyo8KvOaDewEdsVfq
nM63/XVK852qsXoZpE8tUiw8rZrlar9iPm0stgjR1hVBO7Ai01psZsp0wjdrKnt5
JN6oggt/vzJISkMmghMrKQ==
`protect END_PROTECTED
