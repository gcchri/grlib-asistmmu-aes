`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cpd6ZG7Gq4geTG89W43C7G+Ikq8Sm6YfSorbUVq8RH3O7SMeMYSWVwy7b9mYrBK3
hkGpPnbHewezm2YNvwDia1+J2lvvVAgMfazlG2syKKLS0YaEiYgeSkqDBMoAh1VX
OMapk8iCdm8EP+I+E6ZSXWnyzF1ZAW31Rw2UgHAko+zkS69jtfHHfXR9WKPafHqe
HFlL6jkO65ldQyjTSbTwke7EtfPwpbaDJK0g3jUcbGcUGYwLFm2MKIp0vYdYUnQM
/XrykcdcCNVBoA1D/F7h8Vv6CK7qQ+bED6oUN3hJJIm6Kpi0meGsKGQZUP8YRV5h
Y41uJ0bn7WnljRhh/06II5HahDJmu5/0J7HfKyzkbKS4lapOTB8UZtjpS1MLLNWz
l8tszH3uDLCdzNlA0JHmWAxUzcx161bvGNBeJjdOGcCmpSxsrsODWiUhLNdfiYtO
2jQBJFOiEsg3P9tpvvF9bgnYbOAhdYBSqwPTsKS/gdUdbCoNR5S9jeROvYxiAhRe
ZzOXSEN18VvHd6bKT2te4BeQL2X1W+1Ks80IiBR+fBMhsLB6WetUuEKP+R+RbR39
T89KLtVSolluBBWR7+DZY6vBeL2tuOsDwx0GMH8oARnxircQqoa/56Bh0R+Zap7q
7TCYZR8Z5F9AJbANmfgol5QTcB2fcsNHtoF1Yg3kTood5dj1RIyWKhdU5tGYvAx0
XgKk0Ym+J4gfy6LqVdHiu9JZHJjxi3ujMGePP5eNg3GBA7gAe2RYPj0h58oYymKe
zTSKUe8tr2MUTGNL05rjfDfv4vpCzlzuh8mSLw+XCfQErMMfHXoeT+0ny6xgJqj9
s533NsrNUPJZSKDkSCUDW9/uIw25hgqWkHnxBW5WGjc/ov/E8FY8/FYmf9k7Phy9
x48oK7oiby5rPpScQdwJYSzZzUrkTCaxdbKEekKHU+w=
`protect END_PROTECTED
