`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Is2rig0P3oc0NCUluLWNRJ+PRHesMFSXjl+4nF26fZ262J5yD2YwB8SLAPg35aNy
QSVycDS9ppfAhpUxa4b9zwHpLg02AbexSiDUlngCjrEn7RL20tYMdoy2zNLkpeIj
NJC+aRF5VhdEm9NtJdiSUEyv+EW2r30dCOb89tNwRoOKa/esVurAVQFtjGo/P0Fy
fKry/OxYhx4SQViXJGknOmtOvArGErNY2rGfbGaQtR1MCqj9ypkapUg/TbpK1bdK
M8NFLE5EeSonJPRUax2ZELS0He88/+hSnmXvYM3324gF+sd07YtC5g5+I5hP0gDG
EdCb1JWg7mwmDBRHPnLfaQXprG8j4cWf6yt/6zmUr+Xj1zYeANQQrx0JD6oUH5OI
homdEGw+KsU5loc6B4KB+4ldBhkKJMIE4es4CElk9ieHI1X6LKdn3BPo4i1Lo1db
Ya6z10p6jwAd+A9kD4oDphZLomX9s9FXSjKADxaWqoHslAb5toEyT6fX9JL2tq3V
+eXdYuPTPK7UCQnoFFfEYG5EkAuPL6w3PY9X7l2c/rxNyQJOBUii3uRZWs21RFkE
4P6VSh7BqQbb8a9FT9a78S30I3btKmNXxtT2sFHvWs8SWxozps2Ze4HqXfHVcfpd
D2aKt9cS2L7Imqe0hqeuwCz9rYP3lJTTyVzhJ/sRct1ekq3j0n3xG6rMoyO8VhFO
fhKbIJpVh9PmYaZ9GHx1xpm/LJ4F2RntyQH2kPQHX3w=
`protect END_PROTECTED
