`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ygZRpbV7s1fSTidg4XUzTilx0J5nflUit7Mdqub0VkhLccDah5eLEWj0/gdnTklc
1+bARZK+lxxYMkbMeTeVeqR434noblOrVG5/qJWE5lybBeH4I/a2T2dEnKeCEbav
Mw9grBAjJGsaRPpw1efuFD8CQhSz3idUo6XqzyT71i6ri5mI/csMSB0AFkLYQR/9
ya2Etg/QWfpOyqwWGvzVnOWnq5XHSOdbSJInQ53z7kPmIiBsc+VlaW52wO5L8LLM
iUxByZ3OAGqJ3hL2/antGJG2YzKgPfc3c/l8ajYTzIS9P/hU1U8hRT84y4/S+22X
eCIcvsBsLIQ5wiykJSEuPhZFRZr3zhT2NtqXblenYm7qArFZ76OmF/POIq8ipnmL
glkNAkICk6+x18bEz4989Su5ePUMk+pEaui7C1K2bi0Tz7aqQzpVJHXrq6zBNgWi
mmGsyjCDQMt59vxH4IGd8VVFzXDDN3h3b8Q04Cqh9R5FA0haVryt7UGfWgIgQM/O
PtB/Nln1Q0IVgCa/aLt2AdXIKSwpKuI2ssR1KDl8nVyvnIPtmv8tYFN6utjSFPb7
Os+imRXHhw87N0k4KP+scV8zPHLurPCCcdB2EqgGKgC6yH7dTBXlcbe5AR29nlGh
I2bGewv9vbhIDeSUAvenWpHN3TCLR9Xa4zshmQ9eMK1sHp4lQlxa6zSrGXks5Hk9
`protect END_PROTECTED
