`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WKQHdvUtcRFeDaVDFbxc4WrRK5q8eK8x/aR9D3M8UJoOlt05Pri10o7qCa0WEBvo
03ou3m/NUr3ENJuSnzBXHPr70uTNqDlVLfNPj2iXIP1ogCJ3/1B3YhfZMmXaTJuK
HVuNCJvGLyA5/jVGWpbg0svQiviR7t42SdmWjO1lK1rRidPH79h5mYKwaUffHtyk
LAVQo4xL26bBI+tP1zXKaohdb0EnDH+rX6FCzcgG6i8vgBuSr3vaW1140aoH0S53
bsF7SADng08n4GlsKtUGKHBGQpGuGwo/eQaj3XmhLF7bSRdeyv6uhWtvVXHtfeUw
X5+edGdeF3egNgeO1GVLcajprOVcniiIXOeFKZyytJE4ikfbMyYgpiAGgELzcLmM
JOoMlVTZgAN8kzq3O2SwDjlu+YgUPS1u0F+jmd7nFTvAbqFAUQ53kmt3rpN2Pj8t
faTTuX8FkIQXvIwaW95iYQUkN/zW8Tz42ZRlWmQfcV0oeIqD0XgnmeF2Ik1+WcEy
y2QUWqsR+FtlkrevfI0ItyaMhb+hxkCf9LZ5PpgE98W48J4xwcS6JcITPF70i3o/
1uMsuAM7Fu+ovvx7NQSC7C15OQmv7ZkIeot0wRjCFnpOlSDp+gD40ix0EcNuQyTB
uLK+J/R/inVtrujajFrKG/6QlrohyxP86TTeeasaUibd62D/AAbP7q20z4Cpqvi/
LqBvkOti9OFHjED+SRF5FpQMePFEiuq2BR9RdPss3WC5/a26c3Y7P1JUlw4Lh+gq
ts02AgAat+sg5blElVxmiQ==
`protect END_PROTECTED
