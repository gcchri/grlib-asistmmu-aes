`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y6CEy8tkms76mGg3PAEta+D9bCcIRfgfwjv3qF8hVBRDQ14eZ7RHD/cSAnZyUB1/
vxDl4dsRFPuygR4TC4Fyxblr4teER1ruHqg2/ivFEZQ69RlrRUeB5KZEXStImHHK
/tZecoSMo58mbStKrCTQRJhdOyHlbhJS0sWVcIfmmVl+LF05geuz6L9okeoCPWgM
OAQgkogHBahjVcz6nqYOnNvhLVHOxQUz5oCoRACa4woeVZtPcAIfjbsfh2sHcUs5
rTApXL8wy+TqngvdcU9mPqHff673geNjtDwHmzeXEArnofH5CdCrdotR0BPth+Qm
BKUN7mCm9its4yw0KPkNeauOQ9YoXXOFmEadUodlOdvpT12LQQkm7myfcnXpqsn2
qif6nt8Od4baJMzuT93WnpqIQ6e68ZEqMtweAqrgktocKYxrltNGggUnHI7EP5DA
Cm03JPj4g85bhX9yrrbT0etNBVMXJlwRUicjpc953Lo=
`protect END_PROTECTED
