`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tFL1YRcCgOgFmqLfeZgupnYf2OUmsx2hp6T+b4hyklKrjWIWaGrofZ5K0JrDQP4s
86b8d2XQfrJ2zstEx/Li/Ljum/HesI/tD0GhIy01nAA8ci66atEuDSvp6Y+rb8HA
zas/KQ8JBWIA2H/l89NHkMX051JnPMASK8K1tuA/+WIs4BXhQocSRciTA0Jqwxam
LcGONHsy87EzBmwMQKTjCkGEvGGUmE5Z9iNgaqy11RKOhtjvcuWN10CBRLgQC7Az
BoluESQ7wTd4sbrXpyxBZkrdF1mWf+Yc8YbKsymlORF1zF+dwCNBdEYjaA/52uYP
oUDdCSf5LHGefPeCMqfWyvcn8hDTTOAxgmx/2JU0P9deg8JNrA8AeOhi98rTPzD8
ODRYbBX8MYpRQV4RWOWfyaydmtggXVe2emsBqC5YL4rd77SGur/w4TD2ZOtyS3CO
AeygCPx1EIoY5vTyv9Eouijn/eXMldTeoxG4fBoAGn7SZZ44mjb1ZN/xdF9SyzJL
xFGasJSbyHsZ6eRaTjm2qYRv+6noiVzoAVwt6G9O3drGLXA25gzvGYXGZwWwle4J
rm/xhzYWxVe+pvoVXOncwn92JH8xP1wXtOWrVlcPesF8C1NSzF31fcI88FAjZ6tq
JREFIYOg+t94yWBbPosj31qDVwhpzMZgeiFweq7/SRw=
`protect END_PROTECTED
