`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KMoInxnN9+FzRYoQb2SSOEx65fgnQOG8W5IwnOM4rLejebAYgoqQKa4yf3CY7wN8
qqfHUwTEaozTtX3PJSMabl5jnTtjQrx1Hb/qB2vSkzjs4ccA6MLh9klz02UTbwP8
5sxLB+ky1AYqH6fMdns8VZ7y26gDpT8g9S0rjkX9Aq5AEoDpytOxYMUM+lxZjcX4
3d3LAKVNIcMWBXD31zpW6cSjZLYQmGl5f8fZSCJoRfYQweuKDoBFfeOJq7kk1T39
Ihlmv95dmUYp4PvHU8GelbTL7V4lsuyAKfHbtNnYHFj2Tq+58AzJlhp14gL5/PLR
erkRrvCE4j25e6bkJ5oXcGLQ4VIvcj4kNAzXeW2v1i/C+HZCJywaZ+HTUO49M+d8
SWFfLPQAWaUijTCpAJbeRjrkOqvuDKTwVSGON7ARivY4cwYyxLT35Sin41JMh67o
MPFj9avl96vO/Vnd6fbLvRvY5RsPr/udG/dS7v0wpvi4/qbhiUacQN86CeNhikm2
meS98+oOvlZdzsETNM3Ei3htta61JC2G6gTJCNJ62WI6pjhh62zngdhtAr9Okanw
u56EbAIKQKeQ9tBpjcEqQICa8LX/IHpC/uyaYv7NsctVVNclQAqez5K43Nw0sWTf
YyEqtakyKRrbnCYpVByfgKknFzhYZCE/OyMxeahGEd7zjgAUTdxjeuI1RwTl2h9P
C/a04aSlssjeN+M1tmfiFNCzcdFupsDX8bvKrRLtoY6aKqhgAhbv+liydIGRp4st
r4/wntGI4kc4AiwRpHYh3oenBX3T91JP8RZK4PLuDLbTGWeWwNUHs58CuIGRsvFz
tBgboa+7qqr/UaJEJK9Wf6SExvBk5GpovggDDkkwLNOz3id9yvbHbSgi5zUjxO26
NOn6J4riqLUnD4OH5gOqVMkKkG2bVC1kxZb65JGgk1q9buXYJ9aveOaqUC362ess
8ZqfZCaIRO6Wxi63Nan8hezAP2+Oa64L7f90AdIe4LLLztw2ZRXazCkZ1MlqU/7o
`protect END_PROTECTED
