`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fxuwo0vhqGv7RrlvPAdEwBUWX3Ssup1xu1VbKhX3MQhJc/ROBEuj472DXQBoA9Y4
LbpKD0LSyqSByS6jx8JEWOYfomvc5FvUjjkpVf1OOCSr2o1uCH5tWuHIsJrTd05n
K9dtdg22H705NRa61sz0sEmFCAMwgh0d5CDvTELj3JW7gOtjZLFl7pk3x48RQ2Uv
itkbQtj5VXdt1/g+7Hdxp/niPhSQMIDD0cK5o4KPTaiR1C81XM4MKmWztm1FmAzD
O1XRd8VoJ1NhpOdzZFklloLPTaWnHIrcrDH24xtXNR/n5eQx9eRIS6THGKn6pE4u
8Q17kLYOvU1N/mfqKc+YPyV2kKddN/WRvJ2Y7PQzIGOZZeSxnqCZ//ctRrrHNK3j
dMs0joOcQBr3jqbKEocpMLqkWeJljQIGVt8UW/iO0Vwhb+rFDXu9Zno3zU9gWHs7
gdVpi3HLFlsSjUNDmrNswA5MRURlG1CGkb/aDzX2C6s=
`protect END_PROTECTED
