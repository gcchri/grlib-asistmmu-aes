`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rtcWU9Hi2gemyY5tOgHza5ohddGuyoB6eztvQBDm99Tp4SSClVaqLnsk96savliZ
NXLtMvxVqtsVEXRHDE9ML4/V2lAqPhUMXDJqRORMQX0+jm0bDZDpILVxCVkNOu/k
uU9nw6OtTzE5NllzJa3yhQsUQx2i3tZ0KdLHF7fSng9tBBmZ2/0RdSCNFnVufeJx
IsE7SZRu52z/ETaXnP7Y8V/xiV3sGH8JFXO2GDr4UmUd5eVYVFjdmBZVftsUlfyU
6oSaaMg87NcAIDDXWKmbQdcLUXQmlSzBFrZNZmS6yK5nwdoVdSf0bgM8qDRIs9BO
knaKbtO7gSqxX1bs1tJiPaoqx0K3YFGWsKeVnIdO6BCDa/CuMiJCVAFfSgvds2Gf
++pwAPtDpTorAbqkmkLKvkgqHSzCAuSQSFvwvJt4H6VI3IyiuTXIuPNvd+4BxRuv
q6VpLhJ56rmKxvWaGmqxUxz4aDuwrZk5yFjSO+pkFz02oPhS4KN2Q+QyTBNYCcH1
owp4Ia6pQQRWk/HcIeKc1WZDWwjXBb0HBaR4VbB3OTjQQsSWdOkJx3JNvtrt1hoT
8+6WJXc6kPJrxenH/2WDZrRDWzxwse1CqvgLhVwvZwT+2Svf9OHGNCMEZI2xbh4d
CtjGog7fCzC4FSsVdSVPBUjQBEjOQF/y2Op5vSDn1nwlUJ7c21ehUpu7Pm9CrRIb
Cxi11th3xYGDoQ0fI0pDOw==
`protect END_PROTECTED
