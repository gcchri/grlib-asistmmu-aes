`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3qmFrzQ1161iSsgB40qzAwt/g66FFgI5eC9i7Jqc69SUsDyEuWEuvjXBhUFD6JY6
M1E6pqF2r7fdi0VVlxCq80bGcZ36Doi+K+qgb+ps0oBG997iH3Np0B/jPCfMaCVL
bSxLNHVCMVf7EkjeMeIuuJNrIiUgsjuv/JntzdgV3itYrMG6eBK1BrDLG3fypuO4
mVDWAk7WTJ7jWLc1WIZ6vwMFlCNiqTN1t9ZBrO/Vejp1Lftzm0OBURkbGGuTEFub
0uBcu5P0W7+n7KndXZgM7+Fd9f9/A717tDDrG45A9ZCSD5FlviNjLaqCptT9izdL
1hxSHzIjzJhmrZyEdifIfqoXpzcNBHU4PWz7BJFFpOsIysVNOlOTf9hE3lLqaIka
`protect END_PROTECTED
