`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9driNG1wtMX6DbW+0GgEu6L2hH3MPgotLamUM0ehY888BuuYEb0/1PYDWaYSuMgV
5k6cRK27pL/jYKeOgpGQ2TKrxNd6/YTEZKq5Ita8rjWN+JNpN6iKJ72WQAn7bLIV
0uteOw3Dd3R6mRFfi3HdX8pDfuHms6Yd4bAWZiw7xnZCv/FhMl65WHGoEdgoDnSv
2Zcjd+NV/XeUoSqW1X4H7WPoprV3xZ6HLjCavUyLoKAKFF6wlFWn1fKKHG45UMd5
s13pLzj73D9UjJJxw5tx1veTmJ2jKj3T6g450gaxURkCl2fKxuOgkqqH3Ix9irf9
bkhWLqPbZ80z7pWTYPgnFa1QlXNoqlmhfRaTOFInqerluPT4GnzUBgDENgL9t0Kx
YBe1yblLqg88rh3E+qz40e0qJ6VmGBjoLLskaaE8WsdJ4RGWswHMyLN6VfwRH2Ve
FP1UH3lWATGNRet0HoNAD6YwxOhbi/PLKzkerfb8T+DwcBU5mi8BD9vsePZP/p24
wFYHJUUTVFXHwNCfn54xnFVNFclaNqCjNSDEo+OTz5nogAOmqvzXDrkkb0BXnKDy
Kn63WdNpxid2A9DuDAH7QqzcXHKBXz31Q3z/HiuCM2A=
`protect END_PROTECTED
