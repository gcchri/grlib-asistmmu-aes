`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
icjfFvCnFpmx2gqfhHKnorGbQT7XKGL8dDUQV+kOMJiwmeuxA+uWMPzHHjDuLnmx
592bWlHKgYFCWGuki39HrQ1cquFdr1ZDUl0dJNEkTjgklYk1va5TQ5aFWilW2PJl
6SGTPBTSMb8HT90EyuDUgadRJKAM7D3Cx0fuXrL4wRtHznD6x6vNlgAv9hObjyRF
dT1v0gKI9yOx5XdjB+QyfPSuBMgTomasz6jksSROKloIYt7uK+wiwWt5xIS4wWqz
STpV3rMG+1idYphukde7iMFIdF3A465fWIKeF4/4gUzxd07wHe39VInlGzKf3WnX
NY30nKZso1BZMWkp05UVroNgVZJLL3eVY491qUb6+EAzUTbgtPnECu0tEBv/JTiL
1pfOfZk/qs4nTnXk3fvqDDmA/3knvXXmp64vJ4yj3e9bAdSa9BqfTsiMTJSfEqIb
uRkMzxUg/8e2NFHctMmDhOsJamA85G/jLxV+W6Wm/FK3atrtNQHeGP8Wy/E9V/u6
JrN5HLkV1RAKQ0JEO4Tbsiy79WoWKpf0fjp/luk93VqR3vVMpofC61jDBrO5+myL
Kvgc6i9vImekkfc9Hr6AK5O6A7rMryF1x6xJXtg035Ljg01ESgQdclI+4JfaRUP5
81gMOa6lg+5D6EbBMQX/omknl7Noy8GXqeIkzCxzd0uta6I+FwFYm9etvZHUQmlG
4526ATbD0sF7O+XajcGh/ArDev91NQuBJtvyFUhDB6mLdKLm8L4oIIXPTJ8v9ZxZ
SU/wsey+AsTUi4kyno1RA5HU//FZAPd9Oawts/AOd9rc8+sKQ1KDT5SF1opgF3UT
D+G34k9exj+7N9oPkQK9F+0vAl5JeCYT3zNB/iFX/HG4+ZVW2+N1/6ZSEEGFhjGJ
hAwrXWUXY9/D2rwOE0VQN3sJhSqDdRvvqkuXbwHDZXE=
`protect END_PROTECTED
