`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rwUt5wwEFyj4HrSZ6Vij8VVT3hWkB+IYzdM+HeKMTuE14PgtXtovL75/Ox2u1xU0
K7XNvENjneddCePwsZkq58U4kunL/M06chKovLxLKmrNB1i7IyFFhB2Wexje4FGV
HziNE+j3lOdbeUt290WqfN4x5ClDUS+O9LUT43X3qfZZwMHbSfeprjWAllKsE7OA
qo4J9LaOloSxmeBIK2MtC/wXMW+hNnbn5rzTWIWxuaJes3wiJ7HJXpAIbAWSn08P
M3If2mkiQtqLuPwm9MHNVmOPprO2jhe8liamHDNDWDnOgocuCAF++TZkbfbrvaPn
vJ+ipTE9imMfz35RwXoA0Vz3fng/yJtfDZ8JjTu2OQBzOIZTntYdMgHAyu4atr2t
yZqQ7Lf+BfBI8xipHpJleNzgpMdUBHEDda3OMQqE4rRTo/ji+SIyDRc1pD+wJMjg
teFPsTmCitQXscEq7BdQoGBOmDFL+HnVRpuGvAeFcc7db3h4NElB6/dHvyD16Ptd
EO2eJitFpRqssUHy12k/KA==
`protect END_PROTECTED
