`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V8HXvXCwA64ItZiEY//fAK/LkLJZSeyFYtiFX0k0FEpB4A+4tlK+EmGNGR7l2BIN
HGwOeJrYmSQGj+2H05R8APrN082fhQ6YAGL57EG9OINMPs1RImDY+4Bi8FzTgvV6
cFrRmxyOdPa4KZM3BfAROOmvgwgQHQumKSb/XW0owIXVF/+6ATUkrFat2iwly4HF
KutAoGROJC8UZ9TlxZYgRzqXIHn8XQLPn1Z/81oSYsj1QjOvmrm9coSBTR+zkF0T
CRWuB6gbBjuK9DWwO+j87nKpjryxqspCI7MfCHFF5hdwyo/jX1ngk+tPYvof03OU
hlJEqg7C5KLvWpM08KkaX7FkDLABvHf9lNzjad4Pt9YopIvnKLXotOPnjFOSys74
CepJF8XZOYl5cdY1cudjSa0h9nBlZlY+amHOQJO0GMJyEt+4FAl2WWrtPvi1urv8
aWcjYcjCNJH4LlWvconO5nieiMwp/SWBgRfa15P8ususyhd6Sl32WSUao25lEKZx
2qwazgurhQya4Q49t3B+dPTVQtqceAqcgoRZMW7s8enDmThePsksNnNPGQTI0fOs
`protect END_PROTECTED
