`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GxL/UZmWiqazLF2IHeoWK0+kf+0qktRgY4xHdGmiM6NlnTwomneKllmBZ8nGmFue
ZvCXgHffzC5Ih8sCw/SPzfyl1jIKdW0E4ajrgH7BayWkFjfYch67LDriPewSV1kw
lhQH5ZI1tehM/oaND9zUna7nsedILtvsab+/WU6A7FB1HT+i0q/gZ6BJfsSddpvL
p4tUvqTZAd0Cmf5JBCmX/RAMuNjfekeZtmiWOgc8Z3d2PyvfTz0lh257cYW7r6L3
tV+4KUJNxi7bDWvZVNo0cK+jqFqmv+rIb5zmznWF0iHw2ZqWZNnc/mpy7qOPbW4t
ZwwVNpNON9flSfEvA1u8JNFdIsAOoBocgbkMiQu9KsIouwyZCMKGMVdvQBpH52kQ
tOgk46xH9BoBERCuTUuxkqkBEAKy0+N1+VLPPnfZTCX4ngEyWYqnmuA79tDn5Qjo
JOe2lFuEVFyuGmcmgpIDjMMmImhCmF62uxf5HUJ4iEQf8MIRFIBLp658iudRGmzz
H53mtgl1LoHoVanKPNsgy2+snuPJrD1JUI71/mEY/RPtfTvOZOxLq2VzX9wOzKmW
uT78ab12b7Qs7cA8Xu7+nhpWr5VeMKjHZE+S6a2qPhUVHDBGJFDQxLxUpEYmwMIb
KnEyxHOVqWJ/zl2vp5p+lVByEMeHIFpw5ef1rxU/kp5BFO/psazJH7FbGx1bbChR
YlnAdw2Vr70nsgeMRsVV5PMAU2K03XXtzKqW104FeeHYuZkHeK31SqN4lWy3Ss6p
4eIFa4ZKKxQbhTRwfgtuWcfRPiYI/a3kjdOVcDHtZvKq5a30kB4xme2P19R49jNf
DWt/QuD1tdf4QemgEWig7g8EpIa4T3DoqvbipATiJrG5ny/Dw/Q7ZmYEGmh5laai
SitakM+wo8MZA//xikaVhythfIqZTOUQ8Faybd1Yvis1eivTaMv/ef0sp/l+LhQj
h6WwONXW2AG7t+adFBuycw==
`protect END_PROTECTED
