`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vv9+uZflFstNzNn4OxqND/ZuOa37aVpXvD8pfqGEDfe/+muHS3wbjedimUNbefL7
fNOVQlf6xFUILJfOmrlZg1qIcE+US1lnwRtjWb4PbHz2XPGco8CE5N0hYAsTlZcC
jcpKmUZDZQZGZiBo+Xcfa/rbtui0dLpLVv8Yq9YfCpjefMG0Af7cwKcOqO3IgKBE
bwRJMNBnBosc7a9uc9BbpT2tBdxACbzf3YoumL2PkxRUHtT45KbIqHljFgaY90Lk
t6MBH1GL/sk79vFGwBQy/ZWmXKgY6/KwVq5sG7E2UwfDXG+s/oM3riQ1t6CoFolS
aYp0JAozmRxWfIvAhbWFtBWeq64TtVKKvnUoGY/o1DhcJvcZHkt1kWpUJN/gAJ7g
5t3m+dSs3LRAeM/ZsSXxJHdURBCVjScsv1GVPwdSwWhuh8mKgHQtJKDOUIr+UrED
QSrKwjv/WVgUdhCikQdOqZbamz1/oGzpyibfZg89uaJRnrtlqGmaVxDJgTIRn4Uu
bLTjHHY8Nmvu2KDmyaiWzjtDlGNHbVacQvzxVmuKaBIls1HLlfZ6bh/k7PdnpaQj
S0ODBZ3oQ3YMSbzftQhm14ykEg5oAfhkJjEJdYLxrZoWSbgcsVmaJ0hHwuLVJqc/
012SvLgAfaW7hP9O3NRzeJndr+yoG1mQD5N8PMmH1z1mL4g/tOMRdRTSLXXbTOHX
COVQm3Vs1A8fhOzgELV72WqGcpbnsfo2buOQEX8upPz9uGDfC7kPvHuOP3RGhpC2
Eu/0D/17x24rgmEXEy4bmAW+uliyjNLQT9uyoAsNkRaNxjiSO7QEkJmBYe4gl/Qz
7Su15lPpbqmShU83GmNoXtjuWz6ekM1KeQMT5V89q2Fp/OjA8unjSwC2JGVsz8Hp
bckOcEZPa5bzTecR0ewEv2z3tiVt4BiHcChVdh5TVfNEcsowKANnD8AmphazOG6e
Wf9CsQZ6C43OU+0emFHQjyFLe8I4uEqhUY+TBAf0VsidtZAhro0ppxTsM37zx9yI
TTw/EUCJGJKou/QSfJCsEa2TcbybvHtm/H0kbsnFU47/oIhQr8mPAt3i+PdKFNbz
z/bed8xa1hCE/l5+vJjkPzexCOPiORI49xM1Vwl26Bax1SMxP8OlHoNjRmEqkgz1
`protect END_PROTECTED
