`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sZGrKnZAdek/AlsTFopPTdBXnBAR83+F4v8tlWl5gFkgCyj3EEQgd7SMA2gQ0Rvs
0+dISAl9tcQFb6vwJjLPDXHnl2o+WuE4ky5kSIWG2N9CoGCTcriPs96UfJcqULbC
iUmHjoB7ls8i/lSsuGTRovRYUiaPvX90tQIV/2DOxrNhsH5ra1G/WnKAVyTdH1W2
K9RRYGojE/E20pgunPF40S3a27eEf2z84gdF0sYBDngMQ9ZirRcnJDFQ3EBhAcz8
h6IJ2qGWaE9RfA4tNm77jtL0npYUNqR9LQ+OOkIjamYUh8OTHPu/f3NeUUoYHfXy
4tSjJ7VQ/R91Q69rXcJ6VP0zJXBFeWe32faPCSumpJYGyTAVkzrzueMPdaiwtUVn
jXJtl7xZ76DGmGNV/RvxrdR8+8Rr3duc2Y4goyt814WQPO3G258zSWtdJViqjDQg
P1vdnHb7UZw2TbFuISnxCAAvEnS9buCVxU/FvRJUTFbb+0v4uQNjn3kkKyTr5bwx
ZPvtA6Nuz9C5YE8yXoBD4A==
`protect END_PROTECTED
