`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R6UDJxFiF2jWOkuJvNC0crMgbB/HRsdqat1o3+Uo7I3KqAbZrRVa3y3McIiWgq79
IE8F+N7lOUpToGvtUR4zHWmNc1vV9p4Z1JENo+BgNVm0a041XgmlqjFWIcYrKg8A
jd5l99+F1W8ChA2xSTN4wRgOcEF6ZoadxXYRWtd2PxQcNNVmJqOk+WkQXvpKkbhB
+apjMe0WEsmvrBzXVIl31z+WHenLUpXuIjR9dZ5q2ul0NcovswcOFkWBg1371hWi
yZER3y40uRou0GSi6Ll4ErUPUGm/CoeDOpVpiCrFSyjsoNYNaj/xEcZiFapnskkL
PESWGmN1at/gVqJUjFYGqZm4MXrHabX9BsUfkbsGOHuUd0iXatEMr9ugg/qg0qHs
J0nmkkcF4ef+/kk6TM+pk6t2KVln7ooTDydiXFLBAI4=
`protect END_PROTECTED
