`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YosYXRmy1GGi39ODlAIgtSyk7x4lS3iEL90hOhqxkkuZ0P2Fcd5TOYj0h+BddxqC
Pw4R+cgQhWuKIKQ9hWnveVG3C+LDwevtu1juwyXhv4y7MG77vpNuYRNXWqh9i9e7
hPSB+BaUeI5qCOI91Nnb0wtClIjlGyp4JMXF0ypqAc6onBNFnLE+xF60qXrcVHVd
8Ro3CR4mwvT82BwZFibhJQJeJO4wXB70NaV1X2ErU7ISbKBdjgWlm2FCFNMuMiB7
7XFyuFKLDGZnF2Zx03+iHVxRdUM8p06TM6aMgdZDPjR8o3a0uN1SpdP60rFalouW
wRzulXNWJiYZ62mdQNX+9vOXwLtkPdBMcVgu209jW/uNhnajbs8MXLLd1EUCgJUx
8BErAjY1rbuHeLTfby0Y0MzqXgmXHKNVmdz1HRIQXpvz6aXBOLPxeFCO/P9oxf+i
cErR7XIklroeQRsew6YHK6Otw/CbKCDjeYfJraJTE8YQmOoGbymFDaLh0cVQj1sy
7OBrFJpmwSncxbS5JegNuDDu2s5DSXxiUbaOxvynj8+AJNXVyPD3gN1Fho4jJXan
zqU+6ZpJTewb6hCzl9jyxjVUUSIlICum8l57HZb3WwNc6FU1kwlk4Ex9DpY7xvLI
bXNi5XsAQSYozDAQR/0e85lqyUAZaGZ0S7SKGYozm0yVo3g0l2RAuZyjZBYQ6J9X
95KltKfco6OE7QKrckD7QUJxanno9ihC5Q57c/L4BvqAvR+079cIGVqrUOsXKDpt
SEy/ZPqQXd67wSSGaBUpB8+eZnCgENW7QEbKcHCSATlf4b4o5G4f+y2zGtRuRQMb
IykG4MoKhniQwPIMhXTI6fy98pCxOQ8XZTd+kVg/EqQ=
`protect END_PROTECTED
