`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8aH1+JYoCcZjSmTiHOa7UpnesxxK3lZBn7Bquz/1Vb2yEPcl3kfsymhAM1Y1mwwb
jQVkMesJV6ZGcxNQPQx+tEqPgCXUKhthuXfSV54yfYRl4c3APyWvvEr3PIM2L8Uk
j0RLEbSYNBsg1+BJHJ2PgMA83rk9utiznojlqlURgrMo4n7HULh3oae4J6dUa48u
rMSOkjUpqm52qVX4g9cgtM0k1PegqML2k9awZyBnhKiE81d6544CaftgteV823kz
4qo1ThY6LZL0WGinqFTvRsUbbA5lOOgEevh8h3PWzEc=
`protect END_PROTECTED
