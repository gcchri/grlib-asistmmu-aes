`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ol0oNtXMxXi9qLAMAx4GDss4GzJ/iyAzqVwYuLL8zDCpf6Oommtk3IcBoRVburYW
26OYwTX9fMjk7SGZ84idd1wwuARUq+KTsWzQsLhvhqKAwtdgQyYeJbeILwvfljun
7TTaMdHcMdef/obQlYvO2OvtY0s8RWUO69g8BTEu681wgbmUpX65CIgesIEiXn3/
1ORJ+4SfY8zYsxYxuheao4VDrInNsRtgjackUBoNaFncXv/qwbgcRN5Q1+vh+U1w
j1WYFvIX+N9Xhm0efo8lt5McuNQbuOaEzxxJ4TsRraEdE1XM5GTbHzDjzG9wpp0M
fRdBd73jf6WoyUUMN+vrDksjW1ufZ9gpIRaqu+9M9D5eqKd40tpWiYQAqXQZxeid
WzIlJ2/vFLgZy34G+WHLnA==
`protect END_PROTECTED
