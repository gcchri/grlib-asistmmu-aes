`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vHUyGx5kCQPTztbnyRWy59m/bsyePe6iRR26V5S560zYC0GoqbJVRt9Xjfm71iGL
n7L54aAZouahF5jzk6CFmrwj1NhyhPVJROxCYPM+Vnxdcj8BlwZFJMJGdiGQO0cG
0WUdseBSCFHQBxgfoYGPfmh4Ar7JBt+Wst0544yEtSR4EMDn7AAG0sm9MroXOS+v
6zvWYDdE/UtYwNl0U0d0Ogfq6v7G1lRvW6vHltE3tOdpVWj2qB8xuyen2fqJ73+8
sN1901IuCuNxZ1aTx8PSiHpigqIJk/j4KXQIMOgH5upgQJyxwPfVxPrSV4Y7K+DI
3oeNdMNH+uT18USOZ5rZc2+kQ4wRL7bFEQWS2D6ec45fD1acgNvZZW0fCNQd4u1V
Kvx32JcRriJHi+BigMWa1BiWmrfWv990Vuc6RtkbrDlM/PZz7NcXSloYZqs8nGtx
AB1Dm0WeaJGFRmFKIdh7QRnSBHBYH5R5fNr+CkLEu90=
`protect END_PROTECTED
