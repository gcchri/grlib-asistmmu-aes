`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SuOQMfKY/Rsbs4FQXdgbp1aKr4HHBLJUpNDW6Cstyt4dxBEnND/DYs95h22sKWmL
5bni2Q1vLPrM/lextAuzJLufw4mROOCeJHaDfdVNMS+q1Pkldbk89NzoqDFH7vwH
WR+swDwE7++4KmLSRuLnBvP9G1n0/YrVG8+vz+Yq+U2Ci9Xc7T7MUNF6eaA7DKtu
0TNDIMoVSN6hppj9oTnY9NdIm0x7KbyeRCRQzKKJucDDbZDiD81EkMaxvImVUNMv
yF4iPj41Yt4VXg6q6EYaLCFyPTdWIpZAXiJ1Fl27q0iJA9+9HDdiYLLgRiSARMih
gHQzPcfhgaJaTQH+g0pTuiY9PDxc6Nq3UJlKJY5sZb2qGdAEeav8U3h0YEVl/dH7
oBxuGxx/bvADRQqlCk0w1CV3uGEdQu4fWjr4bvYd/5k5VPz5HGjVXF/6FsOYfDcX
0SxsWJHe0IFXzfMNlkk62IpVSUtNvuvJA/PkKU6P8PuQexcOOay5bnHDwzWU8U+R
`protect END_PROTECTED
