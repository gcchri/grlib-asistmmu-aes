`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FHj/m2b2Ofg+RsVEr9RF8BDaiLZrL2PJiP3SHw3IZFq/fbVbWZm4OlZ4YTIKxpqf
+nzjnL/1D95N+6QYZNyTjrgW2gw4sR1oEmATAgHJjvTTEUvyNFXtzCXl20mxddV5
3kpxv2xfcmFSXba++/xI7Pt7CjUyF13E6sUb7HRniAThaTlQ7UkC9yC6DN4otO1n
5BPJc0OC366LWINKNPGDJWTtPZSbKlNM4mRrpMtRPftgdg68tBtxZcmYYVxG3YJr
VB5pyjbRYnbTk9tPv+wcKwsTZUEibeTmVAytJQTnnVcBNQ72TAmZMvakHH/D0V4o
vlMW64Q+IHHJcZY6CQUxfySusmpe+6ryDAmW1PYGMJawRfhcgIxdQNVDfCgJsIih
WL2ziN+slGe62c3amzy5vapLs2b0zqu3WJ9m13WKTXxgwQvZ3LCX6HHFAOeXH8Us
PMhZyBp9MzgiH/xSF3I0HW9PhpHM7MnJgaINVe570njZHjd62K/uY7pCT01SPSoF
P7MFBV+vD92TwT8z+qKt9lLV8UzVdqWOEVSfkuX0GgoqyqAwrXWHBQPiCA6VAhLo
t0vKYiJz5eao4p7EBkMFZpHZj0pyfosClMCay8q9n0vgZlBinOLV+a7gjM8IukYc
2Rc3VAEy7LkphBe3eiEPsY8GierqdD/9pSKkkROnbuGLDKKz+ymhfjalQdkf/iza
Vx4SRpQ5/pvgHilX4thJFsN93ArvmTmaE99rHVBsrc9GQ/Os9FngQNhdGj/nPzue
XLGrb6MVJ34rrGyzLiftgaxTDm8vWSYdDTkJDpgJFGgOQhcllhP/ynVqg1lM3ipB
9v2QQxMoz8SyLRQn9NXXY13eKY/GHbC6LyG6k2jpJr2BpfPgHw03HJ2dWzykXvGr
N25TjrXIa1hEh7X6WQCkUARh4SNlfjqX2bHXLvxb99dXxa9vYZyAqmiSFEHChZU8
`protect END_PROTECTED
