`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
33g3b66wWY7UM9NYqPlRsPD7EkkXuh5PNa2m4UR1E7VmZCiHkCymx5CfbKIpeenk
FtyewR5lj8+wbe1oCJrPGl4IFm65cQdShjNn7e2EKnhlG6tg7rgXIy/BNA0WO6+t
n2/6zuKWdueyej6ijKZxR19TldjPKUOHc56SPdv/SHC0Nup/mqO5iZ+J0gkAwGWn
KngHeLKzEn1Zpl3lD26f4mNxGCS+Tg15hhmdECa5yo4kS7wla12nVoiYWJVKp8Xe
t+TQKK4qJuo9ODJO7dWXnA==
`protect END_PROTECTED
