`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aM9DLGBZxdkXC67NKd+/HacxPTTgY3KfRNbZdVPQzDcdlEESLCsPcvnMitOe/kqH
OxBWXabHH9zLAVA7CfEL7UiamOeKjBl1oU8VCIrsAoFszp2eCMyGGxZOpeNQX/aq
nW+38s6v9vjXiACaN+SsFAH8cJVcg1VZvrLQFXVoLbSNaLG2m1MHH/ZAa13fcD3P
lzAmJR8SoFK3QGw+rYR+J5lpPMSZde36nr9eiVTOhTEOaJtTthgnm/lwsPJKGwHe
aM9PzZq9YE8Vpms1yp/O4gI1cg2ff+bcSzbJm4kXOrJnuHHr6RRPB0IwY9jfitmk
EX4dx8QZQcfCGyEa0AFXkhHZ7sxvo5Po9mp8N4JtGjjuIGg1dQ4hdvgZZGucFb05
3R2V9LHj4siNBfjvQ779gdZN/nH+Y7s3MgdFv7lD6ust6hZHrD8lvDCAF1enIRaP
kGVhuqGXxMo6+GgFh10Wlw==
`protect END_PROTECTED
