`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d8HDbZzYk5bUYt6mHyEq6XzuKL0UE8WF3wgcufOqhDsrgal/igLmBUAs0f7Mp/gA
bs5CQ93jn/SULXo9hzPFw+y6629OPs58unIHNKwWGyg2KQ3pMCSvJ4vPMB/wZ5uD
AVUxUAlacTYEAOZgZaVp29r8Dt6UHXY9hTXwpHyoGDemLAGZZGtFX74tdJ/S3rd5
82BgKXMrGv1M4JApl/ccUF9BX/nQdwXd1TMmSCHAxR8Ust7GQg9vQumwHzvh5j9u
2eAsWj5+5IdzrkqKy55u41ysy+M2u8ExY3vDiHbO6RlQlUoS1YeJ1mkEp9ddsTeO
`protect END_PROTECTED
