`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
89ZZS3Sz7jNtG7h5SJObdXBPUecI+koR+6B9TRe4/uWU+f9etibJFI9hznZLR3wZ
p+12z3pq6bKLpT8bXwhEpdknqiM1U+mRH601kpWTLRO31kza2FE/Bjfq5ujrush4
kTxLBALGZ2kertBFvsZm0C8d8XGvuUADLTSd2z2XscWVUgQe4X/usdkLEv9WQtkY
YHUWqqGfIXwUxtO3V1JRK6XGqV8agVApO0qT6/kq9ihmhCIE4PLHAWAtbwMY+qFT
rPhPcSbsGs/RYBLmi2pAE/zKfYP/h6gQy8rq2yOKB5Ute9QqPOJqgnBmy98Q3ZKv
GjSfh20rTWU5/YfvlGS3s4MhcOVLc8ext+ug6b8T73K+HkukL0uz9jjS43JMY6jq
64GeqE8eKZAAmRevkY+EvaqhBpZql17UuJy7IWE73NqyJdn1A0aqnOyLxEIoNIDl
xnibg1u3842flS9yhS/vgqoxgqV3EiYsxDrQoEdP2yERy8SNcwPqWsLdHXSe7Sh6
pFVk94eopCDFs+sFVWXZq/hGlCP8I1X55wCdcwaS6S1JnFrGyH4M8tS/O7aHSJg0
DuSUX7tI0R4GBfGUx0N9YW3+VsadDDneNTaet9P2exlsIHFY7aW7yB79Wwme30g7
H26HsiW7+AQIRc/ftaxJop65fLpX78diV/wpcpSHwXOni1+tZ8Ef/Eb5tgT1FnaD
v/BlNijuUXww71YekgvUpfFhkLRJiQnXCsneC+b66F0GTqIlLM7pVHS/muGeLcn3
SaC7UqPDLtVqCNPaZw1VTqebKQTIrFrk4pCHwjOva8yp45OykduEH9oJWwOr4yDy
fPECozlEnulh3QN7LDW8q1ElvQ9FbyBBWu/9PFnxFG9ArUHKPdkCxmPjWeLnvojM
47jlno08Ek8s3MlEaXOowjCmFRBDmMw4TcUGrm/Fx7G9+1zPGrpZmnBNNOP7JFLd
5Sjrav5EUsYOS6R8NUhVBMRAqYF2YYn7NhRWGkEKjVEf5z3kgCOe1Iy8+1O5Y881
zlLIaGGEJvlwCo+JSzJjJT3gyDDgSKV4HFmBRKe0v+QQPFKaNByPhd7hik/z5af/
TjNDIUkEZVQXsQDjayOmgna25ggM6bJrpNI3SroFaPjpmPGlWbtHu/H1TCG5RoIl
mPdWIQWmveURXheT/wpcShSBpbrYFjj4UMOP0eE4l9eAJXu6DPvln9XmchUrajEX
6BOJi7YxiApVvULDww970Jit+O+nM7HQdpAFdPbq2W0fj6lJqbOOdGR7aY1UFGjb
BNEtxCkj37Heex9MdMKTzwcRiuOWCp/CD4VlH2pEL+P4CvnAb0iJIQRRXLq+vcz4
hbZsMrWvfeq2bfReCUhAqjG/xXs+bgCYYdAwkDNQJKGP9fUcCMbFp/u1Pj+zTwY9
CTNKL3C2CB5XUIs+UnAHOL3e33+55VEbB5LPdw1Lxi0kbWAppTJk5b7ABuaC+s/Q
ltYLfSVOYCixnRovfiu7CfR/l2Ov1nTZz21iy1V2QlKJEQZhZY6ShkcGGGp8ACcO
PFKuQbdbtQRGFTsPURPUGG+dR9B1oPKZPHIqZtU1mDaukW9sUtfVrEVVm97ICEnX
Z+vUdSVmFwgJVppCtsM/eJxAWK/Y5C+e6xkShDkOV7BPOZ855SMsjx2CpR4PKYXJ
IE2P/3lSq7fpSf0r3E2gQ61JJTGehDBcxx+/nLudJ092dBRx/H1eqq+BLkyQ/mVc
KAxF14WScRamaH+C+PYKd0K7mNApRsz1LS7e7rcuVTABmD1hDND0FBd024bn6qjN
xHWUNQcKVULGZBZyBWr9uKBESdd3umJ0xi53Emq7lwpzYCG8krWuoTHLyw94kO9I
6FAWm1bKv48n9kLgFcEloNKAyC0gE7KqrY+pMitRMVblZ3/ca0dvX8l+daLSDYxb
81I118HmNxuDzDEw/N3PXgbimYVvxHxC1dGAbhqh0lklLgpyj+GT7FAx8XgZaPJI
XaD5Z7l+igaNaV0IH5oIX1DrKYTT3wXzJdRV5D0mjFfGDHWSslXH21nFBTlmEJV+
VIeEzyjBkMc2V0sw/tQyCb7ACr2KzvuC783bMoOTMQXNtRjWYabdUsf4OTPpIP8w
d72HZwWufQDy8TC+g7P4Gc8xxGDCADhG4ExSkVF59XXVlGjsxvbWkTVYMdxc2Qu7
gYUmk8p9iY6uNop+hzD5Z/JCCqr+YC9HT/VN7+wNL+RgiZMsepyePf+1nyxb9tmG
SfjiGVJm2obie2fsBLsBf5JHzVeGGs1zxgd+KswXFn20F05Grki7XJSze8YPqZQ+
mzpkmSZN08VZ0bP42SIqgKCWKRtcMsXBVHYa900HP1u4u7B18h/pW76y5EWovORi
Rmq2KgsBunMX1pimMbnr+7Z/3HM4OzSXZNrndRifz0o93MVhHTQcFYtgiw8oY5hB
ECIC718agu4BiYTCNtkZvwhFnTEDIMrKreYfMs5j4MWIbh8ia/kktAgPzYtpjJO7
HFg2me1geoqvFkdDcy26Lj/6zk2Rn+TlE3SrMxKf1cXj2yJBM2DjNxXvf5emZTcf
wjF28lH3vY3L89O2oz9yQ19bE6K8whsSdwWBHz5yZRWfT6PTMWe1ap4ESelG1n0V
AvU5oKYxPqgrngSMevIgwrKTc9ATcUXQZ+nL5FupH3hnb8qXoqKCwHReg+MihtFw
c2vod5wm38ZrEms7ZI1n9IdN5rjhVSIuZRx/oLm7zw8h6JJGL6+WZnhaB4zF/yac
cYVeYB+2jpe6ci36UWrGKlXmMGKpcBjylqyptcVWBzMok1gH5gnJAZesX5PGf9Dv
qlJEQDnlSJolbFWliR1L+werzIhgJ9f0LxRaqOxeEkFBtl0FnAx5pgVASR6dXu3m
6DHcp5xeLDWNkLKhHVwyYI4mt8lscpAipXkS5NlG4SVmr3G9VYyWvjqTGNhPbX+K
ctSEeOvKTZSHr2WIM0tmM6Fj/FPHJFqRift99AE2IEavZYLQ+j4+Zlcy/no34VZ3
TPPRjRVbkwGkRpJxVBWR9o47YnFHfwioAL+eG7h/ebSfKwTK1RG53V9NGknBGlx6
L/DPjuFZUx8hqMeqp+XWda5xyyf0ZxMtqIPcrv9hQA4KDmmTgwsY+0AJhe++h9/G
tqcHUTAkVJudEs6A9hnSDYTmBJgAL1XakjSBM7PAGlgIJxjJwYl82aBVHk5/vRDQ
eZxJVltYOVVDjXBngT5s/ZWuxXNrh6rx/HDzndaUiXGHJl6xEpoJTNMgA7dZQhQT
KtYGwclhguHhCLybk+VbWWN1GCqW4IfXEbNoaJFikRA=
`protect END_PROTECTED
