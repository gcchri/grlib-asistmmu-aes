`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
09lPKLI7A2g0yDJ4EyPusASD5w7y3UNBRXMxNgKK/gmfgWYLQOsDl1VEz+24QRJL
4V33IGu5sI/IZUqtpIUMGxRIuHQbYuUp/EV2vtXQ4+DiOoRyKdFROVBoBsperCeW
+95ZAD/oLgi1oz+PD04cNAQkcXyDVm7tMp3TU13LJ3TUYIHaS2gaaeXYVzBP62aD
H4g15arbl+SdNh8Y9rs/EdLsF/jHaH3iYTb3cXZU+IIwYxRfBEblwOvQTyr57wEO
h0V8Hj8IwhfxgPHgbSCz+8lLq0RFCww/3yq0MA0mwydGjJqXqU69aOb5f3Sf+lay
SzL1kFDAxw+cM13r9x3an8krP5TheJu68CCIV9RcJ6FBt0+DFh2tT/zy3XIhW6Oi
He9k6tySF8gL45K7erY6OrQwK7bZZvNzAhYkmONaLAd8ELL7Z3t6SMrQpcMpHrdh
hQyLCxeEiR7iNgzHcvkpbz3O7kqnKfXeKCeH2nBnwsE5/SCQzYdgQf8hK7JUYqQQ
GkT82qNj3XSF2/FHojrih5X8oRIU1bbEQrIu3IcfvC2rVN5+7I+z95vPherXkUPH
yyPuinWyu7q/1D6/ohhYSw==
`protect END_PROTECTED
