`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qO7sKk1wQXdWUngw5sZ/LUI/Rm9kFKVN/Qjbwu+Q9E7ukSKcJSE/uIW7v7Kps0wo
r34yoMr/dhut7xZMm+mkQdhqHkOxu2SddbcSB39w40SJNBNwUGudWS0JL1Qofk5P
9fm4rYxXobpI/MqCkiLyqnaoN0erK0iwxQ1StGhlwjOtZbbEIQo2T/vxxkpc8JPL
0MH3xZpylUjvCb/aOudbbYXYXfuxfEVWwTqlFv+Po9Kl2eWjbRKe7mvPDzB/pHyq
sZHC8s31USm56/Zy/6zWX9zDQ/HZKPslbb4RMnxHqKNy/YBaHblz+7XTrUfEhw/r
/nHtyTY7B8G0xywr0RV3sPIA6bAH5d91tjQxeYA250XYqe+gVD688TLWql/0Ngrt
9HIid9w88HBklf0AAbFrUN+OWOY87Y/yB65FqVlZnndaMlY31dYzBDEzSEf98i8z
w2OWx62vXD30PmS7oYQ9mBFzxXU0AxH0adVVwglLr6ePRmLxzdZWdvAJ8cLz3Mqe
wIRXokhkPw3CfOX8BZL1OwYm+Rf8vKgzC290uuUhKg0YZCiYygFlMxtGdIvfwvTB
XQvpKZzu225IkrqBQP2OLhAbfkl6evuwDbPBkfTK/CwtQT5oHrmUBSf3u3XJ4gb2
0dydzM82Nb77K5q7DSsnU6//6RpZpJBBskVU5mNIoRo0zxKg+1S8HarlOg+eBMWg
SGJql/XJgR575dg7sXmnQQ==
`protect END_PROTECTED
