`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hAfXCD7sGiyvZ63xPDVIKoJi19vCnmcoC1twWKUvQb9LGj2d48q1hf54TVaIv8Ui
spvLbcplckKS+vxWT8eeUmnCa4xWJ87F5HaqWqXT4oIJe9ssj1NZlCKcB0t75oRA
5TVtGVFFJpgJfjo5YfGr8vtmYd7GOxSqszFkQRt7MgUUVQbI+k/hVGHzFzlh2bQR
hp7oBnZnKJYqLS7YmygadlTOQn1iX1Sg7D4CCXof7ojQk2jL/UOw7XXOeZXW3/Pv
54N3TSFuH9ygi0kFi2ZGOAfhGcQ+AgJSfbB/jTRo38MZEDr3f0c8pEmxAINsLwcs
GlL3PWPBvgGPcQlFYk3MG2obOOysVJDg9dkTdiu5bW1xhFrfBkS5C82D4R+yD/vm
h1FfJG14YIFfRRg2efab1A==
`protect END_PROTECTED
