`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BX6dB6x5jqRT84yZBO05prt1f/aAjAxoLTQuodMdjH60nQKZQjqiZUM6Wj2IkggP
plSqV2Y+8HHjmv9yXb7qiEe5IsZFt07wzNw5VQTcALzyzMkPudTrsxY3oiqgrVml
WCs1mXUEYMf1G3J2GVvu5h2hmgUkiYT9FOqus1wlyeMQjkckzxQ1MqWaO/nYVgoy
6m1CguIdif6cOZwRIyLL5ZTTfq2zvGX4zgDyfFijhrqlyjIv3m5e69xs7kwiubni
uI669DG3CSCaE04lgYtu8RrT0/GPpkJiGjBq3u66XZB655dWNTwXj05nsY3MXpCs
GgxwHKQuXqpyKZnULoTaG/ZA3Qk30E57VP0/zjzPA80c7dxRjonpWcPXe7eEiOpt
ZFukTVPnfKZiB4Arergii41gaGMcmjoacx2Eo+5vy52MA9tJQ/R2g6xlT25/l9ha
ow8VC9g/z93kAT3GBRWMSt4BbeYCYp8oRsH62HnKg2N4BizZBtxnKLMSkRrAzaUB
kSX7lPMS2ACco3KdKc2RFCZ/FIIi2SJmBma5qCQgNNiTuhyooE70fZpcIPEw/X7S
fh+BNJ8wAL9y1LVkfuq3+q39gCBASj81V7T4HPw6G5wSmswgNgy3nX7EK2d23kNH
s+8x99agtk5S+IFoa4CUE19ZGmqT2Ss1mwbj26jZySeRqx3wvr7YvxYq+9u/TwL9
tHCI9Y/dLaOr3AHxJkNRJx7OlxPnAOjS0MwOBvSI8e/W0Fb6jRrLtVKDRx4+ki5j
Kz6M/GH5tz0d4CUnYl8Ld6YqiLwejuOWgCtHvZvkHxSMcvIfBHAXiHdy8gCtlk9M
9vD89zLTwjwvBB3VhtnMW/L4qxviBE6PytiFhiTpBpYz7h9bUkoQeBMHfv92eZYW
ROloOvVE4UmdMc7sOgmGFilWWVVlm+hR4oKfj9DYqkSOiLUWLPStUVojisyMgNYD
kgiV0LLct4qTs+S/oBlfytbxeyS2zXTHrb3t/mFpmQPIufvWpAsaQrXePKPqkBj/
QtWKqT2KljIQCzRczl+ckDjalmsiWdKHgcPwDuI+yA8zumwHsIrrYfaX6ppQqOcG
k3th6Jwom2y26AY0rBkTZglsHI36PLbt/1Yl9ny1fvyyyRcH0qMyjoxXK3fqnzp2
JpVBfEKzbm+vNeR0/s+VJ9Kh2AirFYpdjIDHZgglDDhZZbVjVXSWNHOY0GxZfd0z
sExt0CnMMAsmxPCsOVC4v9QxXGX6vnF4gr/pI5lR+dcfxC5f5iTV6pcXBT8q0G+p
C8dEaezbZTB9+Q0eB2BXVlyY8a1q1JsgKF7GUwHDyNEv7GBn3xO+PGYeu49VaUs0
mR0ScHEGku4Qjy1zgac80tJmfwcxs532Wr83CAHldh5wrPDij1LZd7A44iQGiJ1Y
RYhcvPGiAeKiQAmvId3Fa4tU4+uE2drmZGyeKfmpjexu7yP4UYFy0ERV0vxjoGUT
1PRhdNojSpWKsxchDf0RecJtEzloeocWks/ClpPov9b+jt08hY+qg9Pmgc8f8wHD
E7VEf97TuI0C8dQ4MoyvZAmO3Dc6GwR3dNs+oINxOIBOMd+WR8TotgkBEheBLYii
RYKWSn5BxEM5ZQes4Nm17rsxGUmawRcwt3D6AfcwlSup89s3DUB81zuuNYToBzE2
BtPjzppvxRFK79gc/cbEJKTlsyRXGnQrM+Xcj1Ee5gdNPxSJVEb/1QiFi13gRz2v
2wVWjWJ7bLzYdvYgl6T+33pGUzri/JuQkzcqPWZEqeY=
`protect END_PROTECTED
