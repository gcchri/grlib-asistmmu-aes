`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QVVe+RaI+fomYo2pnL4lLZJMxVCznS5OtmrHjxWfwyUsLNUjfxNmTy2agWaPAIWi
TapcR7wSNNWPbcvIq8MJk+fh1ysxVGGRSgh5lePjWCq5RN40wXz+cQksM2iqIFD8
WKy4p+fc0Kwb9/AIkrcqjuvO9uBzRsuA6rXombpQTT2/LdCVbcW21n+SlAawl73B
OsrNTXVTEgWQJWaJmxe4/egXJ2AJ9NgnG3AxD649QbIwW5luUWePgRhpJajBeC5c
11YJxuK+mgS978SVFmFI/kYi+pkKb8mRWprjCcn5JK4vGftft5kuu6ptQ9D7hvdw
+8MJW5BfxZ/B/Y4y9d70Gn9dpXWDktR4BBFYs9GEav+9kKV1gy758cgq/ys4UTJp
fJh3Ro4fmd3XtuXy0ULeU0ekAffEs/RuQ8+U3pMLasnlHplEUd6w7E5r/PeyL99E
JUGdu6z5FsLfWL8JakM+1QsLm7PMgelsutYqfQJuveFgYHwM1kIrT+4JqaYClcfJ
kvROm6su0SEe1AAoUvcHpF0JSR3nVqodIAU0FKghtMqHazwAKI7LpHroGAeXDOcJ
ZzlkpIQsQDc/OX3GEMD+R/F8t415UMf7Ro13DldmQyaDyBBu7lKxREsqvrl3pUP6
i5A/JY/ZRqarA21nrkpGbRgO/8RtwUoAXUGMWonzv8OGyl0UWEtXiNOZ8g5fa6xv
p0KUKo9YCKfscxwz5YMBWwtvhonlf02biHQOMbwD4oyFmKeKjB/5syitcngdw9eI
AL8iQTj0kAcwKOb3bnOrTpK63ujoVnx7NHCxu4oPCy8o8xhvp+TixP9KwYlIOvhi
j+ARzUckf+ZPfGALJwEzW1+x5ORtM5wsvOONqPuborIjYVoQNXjwkMgxv93Td/nV
UhDGy6YWDE5sKDRFSXSyEDtkbnli/fxSk36iod5ux3beUP36/mnxQWglwRIpCTH+
xGL6KfMkCvBXYu4M+W/lx4nFxGFIsHKVZl023V0+9vGG2Zke1R0ISjalLxmkTHSu
m7TMMsFJqcumuE6ha/ifl1/nBlf0YETzdwwdsg+qLGSSFzt+4I+PWDJCnn3p9yCr
yHmMadBDdKXnrKlqkTc8KO2Q4eg/KOkz7k2DQKP+hnJ9SJsvmvP2r3Qx9hI3Iaz2
Ot/y7Y6HtgCIOQfrJQfb2BIlABODJJsdfgo3QvbmWsUg3sg7UHzISOBzZd5gQKX9
qv1c0LNnJp4scttYeqmrUfeZK2Ea7Gj3161piqSDBD7SRQoQsCEUdO54YYPgcU5E
GEOA7uBXgZWlLNqd5tZXbCLMLxggCHa21a6w5gnxjUB/LQpD4Ij5kzTr+Js9eXKu
eVPg6heUGVlJh8opPMmmhEmSjscLbTnmAP+U4adqKFMQCeONG2+IC53MdxmfCmWF
bl8wOV9sHOfB9o/Jb3NIyqDt8f01bBcIYt3duBEXK7x4wpTJEPTd7nqlMy4ArNXI
Je2O+zxVXmewwrWqz/6li2raHCKWHFzD5hDAb2eRlJecYRVXhy+Z3SCAPmS+CupS
YG/8VHLR2A57CmavFDJqZUil3Ce0QwWHkAMfLejDOJMb8AT29IBkuhl4Kq/oPbfo
hPBKXyg7PPQ4NetjrHKpcDpR1xHq8DwhRYOkjNWG4YWx+iAxvmHuiOiHLj39qXpk
fDkMTwu5xAig8MAtGcYqOXyc3uixsNojw5XGqcVI9rBpTo7hXAGYPK1ljiZ5cCbw
HI7u6Yfec4OVakfCOEXeaj+bi2wVdI11G3u/Y7edBtV3dnLbNlvKVKYzpZBVBg4j
Gr7WDUgp4W7IeqAw8/1tbCbclTzEup7V5WJPU0JFPNyOMjz4ly7ftWshAjHOIH84
i9TpTDH80JKYEg7CBEBhQIyTeoKHloNgiYpc5Hz+H5FdD61yfuAAD6DpaWtr7XwC
9YWDtkecEZuJqUJpDDPX3k7Npzd6vM46cG4Wp3eSSWxP3xb9s5hjHkXzoO2P/Anq
FCRVK60SUrl5Ag+aPWdSh45ChF14nzXTICo7e6mJGsuvVM94lzsrKFIz6orKBzoX
Rz9iBU6hQoB8Y5309jOKKF7NToRvOqidNaU3RC1pa9FV4X/3M9f1MaPOmUZOnQUU
/qNqjws5pqIHWMpC71g6471BlUMJCNliVHrEquCtq1uc276WrOFH/anPE4i88dFf
WZPCKEcGClIWmo0j5VOg54RJQyv3ah6+FpuhEeGnpvzwQ5deBQJEmgAFT+3oWPK1
6wyqOGYp9YSsty7WEVGoYwBeoiLaRJ9h+IwMrPHVammY/ssMLbwJS7UeFMP065Sn
GHWS5k2vQAiodSuAVfVauFUAUtusl4r7LXWJ577k4xxamZXPjEn8Hb2uFxQ2b3fz
TEvDp/zT4AkIRVAvOf+XljCc1ZXBTAzdVsVmcZiaHDp3bPpareGh38u7RWOS83VW
r87q9blG0ssp9vBhyCUHGqJFTzJEHwZvGEWetUIdFRGNakjkDXceM2ttFB7VcEub
VWneZGlcnVaw6ek1qJid+ZWGuIXzQp73lsmr3u5pfv0B1FkGXoqrNCc9doBvNw9U
9/lfU3x0nEeTs5h9i9x7mcMUAAO1wAxQvQpRx9Owm0mvPTmn260phXEbCQk9LBBt
FZaXbTaAFLO8pFmEipony3hEpkdE7YHkUMott9MIeUi3l4GcySM/Cl/BMIyMq+Ty
KB8lwJL2BIxCUnIOEVT9zK6+0wJ7ekArTiVj4WV4M0oNHTtH5U245Ylb9SAoGl9J
iv/4fxL9Z5M3ygnmeP98V2NDjEoMJTKg3+zkQUUQeVnUqFDuD+5IfO7E4RUmOtU7
acjwwyFeYjZnEpe8XzkQiyGn01M+MWNAI+ANhzyNwK0cGa8bNGlGH+wnGRiiZmxB
JCSuWhwfDGw2OZR4+5bzbDXRNtAIbLh0AH/ktTJrqFRQiUsgXyv+un+aysoxeOAm
Y99GRIoPkLFOsvgGxLT2gY+8MGfQ4T/wrZCqLFlfgFCEffQbMSQxAZ4szfrwJa41
BppW9Y+wIHew2AqAJfTBkFQDEr3doBV/eHF/rKKXvNo52cm153JvivwKKuhBmqhB
gCAUdmPaTdAFCngU+esh1k9S7aaO3VBTlHhK1ZmYPPmSU4/6pLgluX/F+W+zlwfM
ncHLRoijoHXpvuM/GD/SuZkI9kOhppQLDLhq0O6dzQuXoTrMHrBbfuzj3dktAwRm
Li6B3GoN2JZQLyJW7iXFC/18UMTO1T1FwU/uqNEF3xSUaqxuukbcQ4AQhV8SFKBM
Dbqqp1Aeqea/eVnVFSPVcDe/4WMw6lrGzidQa1h4ZjcPg1mC9ZsRbu1tsdwvUezI
AKocBNy+FW5tb8RSGV/pmC8KoJHi6n9Bc1RhE1MtQVEoGQzApzFuB5XA+xbf772k
Qx8zJenexBXtvCf9mFh12qTrvW84h2Hq9+4t4mRFpt5b6StHYtYxPnsxgkrCrzoq
ZzpBp697lbi4E5+3vgI8dCRJpS1hJc8FvCC7+xpAPnjiC66Fjs0ebf/KrD+I4rvy
qO4Dp5wZA0+ghaFHG8FVnfQw+/ng9SVVIZtc+BfjckJd90Jt2asWZMmM1nEI7UKE
PGfpvM7an4hq+2jqnLF/llfuy63ncUGQ/bezpd0HDV11HuevkyvT0pgKw6S6DnqL
CJ6/AfGjyhLTD3GJMmOe5+Jyh1MQsDv3zQ+F0zUk5EJkgFCAY8mEUbBGuibDH/st
CPlmvdj31zdiD6nT6Pl3oIgsrcVdMSItkp1UYS/hIR24+yK6wuCgFPDUa4pMweRU
2k1zTW95Ku45D7JUB37aIxAoidG31D1BLGGDGwJWumOftUn+r7i7ZzQREdpYEWMV
4Hn1Z3H/dfSiX3qvUl6gNjNJFT+zTAz1Q2YIW8bTizh073Tnn3siiP++WE0OO4Id
MhwZnL/eT9+TX4zSbqoNnTnl/Gzi+Cw7Zcizyz5y2lIruM+QigrsoK6R5nGXU4HT
E/o3y3/mrZuRKnWoNJLC1Rx/ITMlnI7FAb7BNqofNmlZ29gwkbiYWVOnsFw2Q5Wt
OiNkO50/8xbM/GEPLf0vghNYXgsEBtOGnw35WNCcftN9kVEflIfDL/JmNYA7KxKq
GblNDNzdN4Vi+N3hxh78kU5v3o3CXRyyAZU/oi5MoEjMnUbD4U7u8GW6GKfZcyVE
bK6O1+2eZQw96qEyWJB25nfsirko0UZc2qoqNsmCLIuqyp2GD2J0Na+xB3IbKyek
twyCT/fhIScs2Gs2j52qaE0ucuhGZrKAcQK/BCodvqDQ62YeOgLfbSxkF4B+M50b
/5A61HwMmTueRBDXHM/cdDeYW8qFa6O9WaEPTSh2vr21em0bFoJlVxvfPLfi/ZrE
hdo2FVHAFnigP/kdfSBF5TMoKZNePU5NoxvyoooRG9VL9wOnYAyk8pNgjP6KuX2y
WDzmm34r3EtM/03AIvrmju2PYdVxcbzkW6v5XlV5PGxkZbw9Y8AzdeB/tQ7rXNYT
6zgCRPYBfhkBp8rfGh4A9OVaxaDviQxc9vaICAx8yXaJLOoQqdAICDmvt+VjzCo1
wqM4Mha/HC9DzJE2qxdNn7Dl3L72U5M7wo8/h7N1qwVB49Gbgi7fJAr0PTVRbSEp
uDsXD9n9/nLDYb1QRZsSj78AKDyZ+ksOPSMj+0ygssNcKzNGan4bYMcm8jWCQ2NY
5CQRmGFOt7v4EYuEiSO6UyZ4pLIr+u8r1ADmhFUu0Oldn3H77jMgQpd1j3s+LMN+
fxsinLW55TQwnK2EUusMCduOv2M8veiSdJufMl72amDhK8CInoeAPvgm0HMhD9CH
EwaklZxhHjqyikY1yn5YI3+SG9ZQ2mgwAFo9Z2a2tjXnozD6M+fqNMVV53avKs/Y
3icIIaysBM8bWADtJ1OHKTeFBNSd4m8c1rauq9vyqVvZIbhGeAHcaIwWDOb+5vjJ
5RObW6inj7ALlBhePaqdplX5bIXe2PAudyKdwm5l0gwhtXhPEkVVD2wTjdg5G4G8
E/NJVoIh6A5AMd3nJltLQXjD+su4e8LGqWn8AZG/EuzzcDhcoorpinoTpQTlSAWg
nUlxd1u0ExEASGk2kzSr6yTLNKHh0Ovt6hl5yd28PrMPNLKYKhwarG+/jzJwDEB0
Fy99Mpis8HQsvkg7H8Ugsee3axMHvPQHQR9oK6EePFtbQBDBXHx14KUeXoP3fSZc
rcy7j3XXg59Gx/0A71wBl3he5w9xuJovYW3gvO/ZTSpc6OWR8QTcE16ro5fQqHFO
L5a+4aPc6JC54TZHuyTR6vKNG7fG4CUyupSyxpUOIhI9PCehY9KWyZaSw1TbNW7U
ST6qZOfFo0G6ZR1IxD8ivauAcOYgVnFLEj3oDwayVq3+rFtCqP79Z1rmHrTsud8y
jier+qaLgQm2iCYtvOYVJhImbbahVSLaiNtbPZ+Tp+eAf2FydwRx4Wtwli7Zw5UD
BDHFau4H16uK0BN1m69BnO/9YVZiwIH9GUojwuTuq0qiKE6UbUcIPp6qD3qdXnIx
YLk5tHLWhKscT0nG496EFPOqniPM5P5rNhNlZDIz/GWag6XyIxJIPxVKaiCwxBqw
dwuOgjn1kmHtBdbCVITVrPbU4o26WasNqpCiEaUcNsTim9xsUrxacDCQvnTv6Fqr
tjlZUaTEIcDChwhL2jGLCmQMBeoe+d0S00w5KJ6y2DeHZsKyWCpr5c+5/v5RnD3j
Vsh0upKxMLq67FWcdxvNm0QTTh7SWwJgFmGgZom2azvQJqI6Ow1AP2lDKWCk2KwE
LdhaPmapBNscGS8t/RnQ/ZLSVJBwOBow+T2hM/LgT1mqrqswfpSfCYCao2x+dh1g
byno4+/VcZF0BiyPy5nVz6nqL+TaE4Vll7Hn9DuHESlcJyfEtlemlpWwL1hSLVI+
2y81xHvIiRSjeEtiqGeqVsOHk76owFp9DDRsjNDHwdaPL9NZehJK4K/F+ITk4cov
pwE3JXF/bsPnyFZAiEIyrKvRsdug0QcPyfUBP8g+G0ligczautWkLSeXcvyDsPMR
QQBmZzyT7M5f2xhvdMLK4gpDzejrXPIueQITgQwPIyHJuYDlka5gAlLalF9cOJtq
VLmmK9Yfwe3quHJHcEfpGZuVpPPcNITlR3pJMilab3g5vJvYV04xkhbx13uT9Ga1
1UMhdtN/5E1aD9voYNzwhrPDr/VqiAh/oT2rJHYNmXIw3/WKdUtOfRkgFbwlkD7G
G4e7VSQwmYHA053wEbo+fbRWkgaGc5Fnr5OGiL+77yeNcX9VGwJyKFxL+kpMnsNV
m4S2FV2ZEip5RxBrk0ceTnK0M0yOfgYWp4vCgvl/kzU2zjhiXJUL6zRjrmg9tgsi
BXjJwTuQFTX2Z3gxIY6o2rLCOOaKtj4cI3WOjrzDaTysEagRw7PvanREHi3bulKn
bXk9DA8qVO3W2Pemz82Pe/O+aUYHJWNCIIW0vtSIC8e7BhLd6Wl6E64Ut9CUDG/k
CGgrlwUMxy/m4JvcDK6JINeqcXZrzjIoExGph1rcVdcd2OhnL1IuyBelZO9dQZYQ
HysGyYZEUWPK5iEJqDvIsDTDd5EaoGDDr5fwOkevAvjpk4apyx0JPn1y07KADRIm
uLyPVxrzYtjKPkwUUgS2RuWTbVTzQKh+OhTUBdTFkCQYTBLovWORmOJulqnfEHUf
sSldkpmdTHnVbCApbaY35EXGu850SR70S9ySzD5qiR+RzUkCJGttrudp0qPrOCEV
6s3TeY2Lr4XGd5cezERUTscvG32whwHYhk23U0YmpFN2cOTRIzfaEhRF5NjBYGh/
+pOtGfZz7cE7o4D0hQbR+Qj0HpLSRud3uwpvK9O6IZHlwflJKjEtPu/GLGUfBGMV
gpCxndpz9DEw9VBJinI6NyD/MO6NduK0nfJq1+sN0Nls0QgEJi/QmITO0Plq73zf
ztZ9dYDm4QeX98aSNpmFX9fBEW1i6zZGQ/ugpfo3CqXA/o9xaxAd/qkMoonWmd6n
U7K9a7Yz4w8E9m6Kh/IlpsHAZCIQWqxW4NOdjfXPQtZKnD+sGGvkWbgBZ9Zj3chK
CiNLGHMApOays+HoHGVivnv/ylDAVLNwndODR2c8SZvigpB5x1hTFfNUU9IPqea/
F10Tt8wEZgiP8nLBCjabqfQaZaFohw9d/ye3gJD8GrC+jzbkis5kZrijX9tNRNx7
zaLlx/SSDdHdmneeUgs9TGNBRSC1GcICWBBH8iUbvCm3Xm8myS3YZZaEvaECJ1vB
EWZP3mcUM3yetB1lqxSQaa/WPotYcV5TwwX94ONvk+XdBSy9YGM0O/hgwUtMJXUN
MP2+u8o8zhv5eBT4Ltnv84kSMBaTJLRI7Gad4Cxya0dfOrMlMfFGxvEWsUJhF47N
X7CqtZBjlU3IZ7gRFQlSQHCUgj4zn39BumRYvPd7A4KRPdYw+dYDfZK+81QgX/fD
iH1WemZ0EFkrKYCQWQOi9g3ctUr0fEJIO6LN+67+Pe8OPB4gcURNTDOJsE3nbXJr
5/cPOU5DWPAoBfPjZ4Tx/LeC9JfkgYsV65sIN6kljdOEJkE5RWD/+oU6JixEbIxo
hi7TUKnazb1O5Bf5q15SobF+IIx8dkWNQDsu/kZ/heDFC9axFSYyiZ3oxUWhoF74
uMt0vFohyxn5tY88pBX4N7x9uhQ3iZ0p4XTUflao29cOhQD/mqRx3Lni9T9V5An0
zb5JHAvuKn9GrzZb06nf9azV/JylNfKjDs3vuQP1c3p+S7kRPbfaehAgqj3HCAdW
IHwvieJz8UDHRbC8o/QtKxLmavVQNGDcscyWHp1MIgwTHqo3kLNyJA4WJQkD2SuJ
O2xt3koPgZ1HnkXHCNo1YASWn4c9GLXne610O0r36qyKkOawevXeztJVwSUGPKVu
dNUZ9hFcAbv53V62WzwiqNybKwFau2n3nXJ9Dq2Y/FdmfW6+SMSD3OHAFi0BTTys
GS/5z0RmGru6rtpaoUPaMKHdVSXvr+TwHmaUeAzsbyYQDfJRBkNBRcdDyikgsuxL
nTn8G2J0/N3BOreDxvhgs4qijTqy83fLD/T9FVi6ApKCMOJx65c2ojdiG0JYU8+9
7c/dd+uaRIFCLqhZ+3UpToPkEtPBhaPNNj+Ha/A9Y62i6EHy6haMqSWCmXwg6hu7
KhO0nKK500XHLgDzvDhKZatICwwZgRXIOgWhTRV72OFCPsRDhGLh5jcvy3Xo9iMt
EDzV98H7wKhsUYtUjY795JHyRy6IaosEsbDPzv5L0iGlYNeZsaZxHBlNYHOdC2du
B7G/TgSwrF4EXm6WzZrSt3SkRmX3db3Q6lTRYw9b9rJ9nUXAFAJpyznts2FP2HvY
YQYI5XxIFS5WnanzOiqn6kq13ef8HLKYZsk1dAcNv9UpPLKhw0Xpx5yDFy1ycAZQ
DK8oEXCPApVJG3KyC6fmTlrbJWpD7uZEXj5Bd5CzMR2hII74cNvovclwzHDrFTDN
NZPBAuX8JITQrA/fNTocXzObPc0mwiH9QNYeyvcFMP/0fGA36Liu1AZe5fSMlI5X
T/6S9GQJfbDvaZMT6gWcZ1P4SSUwG214y0cIm1H5c5M8gJu4+/N/PhDPIaEU+hfd
+Kz5XDKrIjtLgvg8/WIwopkN8WnfVG3OpfAWI+UuooYe7OW1/AhwqBKXaj40Lr1E
SWhPRe0UnQs/CXsyaYR/m/A2TjF4Qkfd1wOLlellkxQAVHPoBLwxFr83Ob2ZmuzO
o4KWc7Ki93V11uEE71UOJK5YsaeSqFdd0EbT41YvDfjMwzhCbot6JiHp4JwIOvhM
M3n8S3zgADuXrRSY+Yf+LRRJpLr6Ml0FiL1Bal1AZ/2uZ/JFIUE/+qAsGIkgZOX7
UGqAEou/cLIqqw0FXyPwwkTBDyNv+kpb1CvcX+AkEzWQZUbfkHGg/bX3IMv+XlHo
rDIuB6ucVrYRdNEFCAirQEA3cGoJL06uQQFsBdHnre++3HWuEIJOnV2ZqnhbEYXL
TxF7LwC9yURbDpw6eJf00r8C3ZGO3qeDjIBDngaQGqb5+8p+qNWrunA8tXlWkGQd
m98XJ7FznauzGckfgaxrBQghYE6tZJSF5QnJaupYASAXVZL8LUCQrzHDbYMNsbt5
oYOXR0w8FfuRATD3YYrzQWff2SEFHZk2qCgKRWwvd5Fo2Xv+Ke82EtN9kfrYOby7
EJm15l5qwhKjeTScifutEIOv22UFg3rCNUiz0K4q6+lkfLrKsT8OSBBW1HjFRTxy
VTzYnrhcclOK5qzNCIb8k5YOlfRFPegkoovPNrPWQST1/jtsoZP/TAPHWQ6mXTa2
6l1ogS02M6mWclrS/h//dT2bXlUzHnrJiGjVJWWQWnxuyAPU7DW/tqkmvjv/ZMWT
bCwf5QiM2FwtZ0tMeuIqYJ10CdhCOK2OC/IGg5jxtHwlymR8wGhVnoyDjn83FqN9
gcwGKnTEchJBhmQ/2DOyc4ybY+yfjzaGggzxzjLZEJ0woOKxUZSm662g41nc2H8I
98h6d8DTrivjo78qCOrrc9UQ6z6AvmhAJKhyKaDpgpTnGaXQT+y/eU5BgQYKOThg
/QqIq3ERY2/XhQM3l0kHEs0Uwc12dKMDTqNgjZWldDX16QgaUd9+Xu+WMOy6uJiQ
YJiOb8VR0FFo+bT2GRxXy7lS/lpac2+FNsJTYNr3ZoAeLSmGs20jtyNC60X5RH5Q
k9/e3dZ1qvGsEbzS9Lnvw58L44UVols6gqUBMHyWQzdLixrIIORV7fgpX1KqGt5D
48ty2fQzkMbbrS57r9DZ1TgyA0ibmbUorq3K1JHA9kAaWRjqjMsaHwFeTpqtGi62
GR+A3YJxKM4WDyOJBXO+tqPzjchPGXcOENrYg+dN7+hvWsmrwwG5fEH4p8wok0rx
VvDqNTN7DE/ZCRMkwjacvbZmolK/VgVmP3Rm02FHdkDGdDoKeukmB3cTLKM6UB1D
RyeVrdlxNKWyKbvhkyey4fEWuOO8wvgtvTwpUg+8CtC2749M+Hk7vz06HLSJ32Bm
hziJBuru6BwfqWNSB6Xc3itQVfs8762HYZycDe10mBk6r4+EKeuUNBiw/KzVcFba
o2GO36z1N01yfUN+5AF6U1g6aedJv9JO+WSVG5w3q1OzqNmh8gO3Q/yQiYzH0DSL
4uGm60Z7KJVWE8E3RF2pY7D6NeSMkLKN0lcbeRCu/k9TiN83d+sJZ8x4nV3aXi26
gLsalDc4ndOwCnmQqRmBp126wGjehOWCmmbpUFmmNkzoFawD3oGE+jLF79llmlKT
Ojf5JaqBTkyI4LzWC4UMndkMwCKAXIVd68t9/CokvbubekkJiBaooycRi1jnAw5h
r7ka5FLd+0AxzQJ7sn/4cN+lYTSAHX6hhMCdgTQi1MBwr/8eBRd+BHGFhDF3DSmZ
k7NR3u+9E7H7CwPu0HVI3UFA1GkXvpasuRNOko+m3W50PLSL8RxTkgKncCI+eoXr
awxNXJ0J8xfvB7nNwZgerO4qGrUIYeXqpHENk4xYEC9Sd4C9IMYM//2XmJiREz6I
E7GJN7ZtZtyAcg4DOi5aK5g4bU17LDMibtG82eZvV7fvztOogUuVA0+0fwxm0g5f
5SyHuPlDLPqyjfB4S7G91UwbYtd6hsjCc17KLcJoCyc5GFJ05aWCRnMe11z5q4NU
HYG0sYYr+eEKmjhWS+jxMrxBWLOP3rRkebJC2wnazm5ft0nZSu8JR/ZJtcCzu6i2
FBAKLQgpOGM0nTo/hk7p5Dgf6xIaB98mgsJrBlj32djDzqI5wzfYXt6MRR0cLST/
ZtvcSnVCZXGcB/4G/uHsdVvqVC4AyFOFaCr8Ep/NdKYPJtN3EbM/1VEAKmNAOVLK
PLDuVDQ5NzhWOm1USEDY4bPVqZUmUi3sSMxr5U0o9TDz7y8w9wFstGx7zdpsIcQU
oFVH2gA4OMK2lIAM3aq4ooyTs9TvGR7TF8VHScISLJuPksTkoFwVne/pHYMbhtVC
U2IK9Hf5/5UFfCwtVKPLA2OhWghsoMwaHYFhM5Zkni38CkUJNfCrPn6lvHTBDmTM
8isS9YBV0RqvAtkRweWUAcO+kgVXWnz5V4jP6iIK4KMrpi3/8SY8fDEV058fHn+w
dxbqtCCv9jfAWcUQzD/ThHqf1HM1OAbuwZd3e2l+u44ruf0VLo4Wb0d+pE9ZZsq9
FrU4QIlvdKGHZ5j2fPEMJdjzte30Je0cE3WTLfRwKb+r6gS36bVDDRXQDvcM9d9L
uKa+gv4ke0oSdsgLcYTQT9EmkneX2uPNN4f+XBNnbHfYT2yX1oBWmv/3TgdZ/pOK
PC3qdyxL4yzMI22yDwqE7bKTamcAjc8jSDujMCziAW0cVkKX8l/WnacLeiHmsLjB
Hq94MgdpsOGSnkR72LuHscoo9s8WgggCzwWgDARqIDmGqx/DGTyOYKjjjSDbkmwF
Wnl7zcJqNAfXyjXMYOXlKRqMFOPomvBpWNPUG2HtLAKPXe3LEjeZyDPHca7uWjQH
5iiYeQb6QMxUpWCy7wSEKBpTKWAbUWx/lqVYm1Aulkmn9qY96v3Km/igYwBS+D2C
O1ERB8l6hVam+pdUXkLO4LDtpLiAcNqCyIKYRqGizH8u1h437nN3foGCiQP6/FK4
I0EItnWzO2OYR94dWHgWHDaNXJjsb91mugkzXXB0uAJ6Ge7AmKAyneW73sOUf1z8
yJKOOLzW311Xa4qPSOV+PgfaC21K/VGJZG0h/J0J/lKpMGhPknuce8Ozkfrd/b0H
e9CLtz4PyvzmvBabdWScrRNc8fNp30wJ63D5hZPtb9nNAB8sVuINWDsHgEfX5vqO
YY35z3ICde6rMBnDxnYp6jaCWmV0Z12dsiOlbomiAqFpK1sCnZ73ZtFXyaM10KDN
hF70AeSqd3YAOFM1X0cUm5t/bQh/8iwGiaXGJtdxuYzhYmndYklL31h5nJ7pctoi
2Q+7OQ+6TSxWYYDuyu+HjaSUnDkzheyheyEKtJa4YmwiVttMQqroWq3PrWWItydq
RpLl6PRJnXS+hYh6ie8RIeSS5jRu4/ZdV9KwTYky1YdbhzKjFsAxvvUNattcX1vF
Hwre5LpovydyeXwEmx2JIWsVWHHXBZbI5p+DkerWQSzf4RjChQDhILJJeAF7ai5B
2FqCi7EZDpFNfU5z5BJSnVk1UXr45ETiS2lG3Y2ik5pX+dmsd368mWFZ0bvgnh4I
4o8oB/k7/ik//K7QmnATjSBebD+JiUhMp8qn8wRQhp2l1b52b4818MLiRl2XA86u
SAS1pEOoFojWTLr8wb+oU6CZr4QLV7y0+RXM2/5NdP/N/VgXxNb0+h3vVdisxWYt
2i1yplUk6M8WAqNa1FzUVpUnrj3OZxwghsDB2UDIQ/lQ8Maq7mRcny5dZBb3kOWe
kBDrHschEvDAl5kjWOElEi6ba0rplU7u3N9FxwzfCaejQiItSb4w7JIl6ewYkEgm
hA3v/fFfyHB14aLD/AiLQOTwsalX8mxiyDBGKpbR4qH+CK5BurNiR2996hehgQB1
AHKwM3Reb4Migha0iHoCVHqZfnPiN4Laa2z6R0iQasB28P+fAGQ3kTxBWWup5VGH
LPEstfvLmM9BH/E1RVhbk9gYQupxcfjNB3J8madFmvaF1CUFC/OfXIgwHTndBy/5
LvX+gF/RadmHELrcY9G2xT6A438pErmKBxuOVp1qZtZH/ff+JDV8zitZTGlGBd61
T2XRhJF7/5Dyiv383lFeYbyF+PzAJTzjQCcC1RVyhxO3fTNkGzYQ3DCEHFfseX8t
uMI6HZDrMaPlJ3CCAPQtDnoaU4fCjOUql5rW1ryuP/XwwhWFEVRyiU9D2e0D9jzc
6sPto9zu4FaTN95PnWXfOC+BqE10K3MwbAeFR4Y54zabqCZAsogQHU8CoqNrfjse
lJPaSpWpydaajhGxdbywMoOjGdRPqQQFHD7H0rJMOWD6E1yXqraI10mQnArjrA7A
NzBO0EZ4BsCVfN4BVb0fELIo99bAuZh8MOb0qvBLWQT4onEGBIB9w5IfqOc7t+x/
F2R0itFBg+EHShL8uSy8Tikgqtr1UE4PUoSRbz2PoTkUH6f1FzgSX1X6PbJ0YAn2
pvBVtFlfplB28OCoMUUkSXxKYnOt/za/bZ/WhFR7IpiyK6BqOK18JSUouYYl9/01
i6OVicNlepVWHC892fHxyl2cblyyZFG/nFN17McNAmqX82OYdUf47FWDpXAmYhG0
2DQ0YkmuoZgmfAx6QkTXBmKcjFamwTO8IDDVyMcNJWcznIjVuJrZaDSeD6oWmLnw
+Scc3pnjgd93/wgz022rCbnHEFoW+C2zFQ+YCNEGRILgwXhTKs1NeuXW3qiwDORa
MwIf854QcLlCyWpvgU84PS9/1ENUP5pCl9/q6KMbkU+fH3DOolgup4WQBpszvnBE
GeWQWnXETQFvjRVLG88COkbWpR7YxRm7rds+BlWa7F2Nh53uAG2QSn/tQCNM44hb
4am0Az9T1tQy/25ye2A8ujMR/BDpwP8kmspN1MvJfKeHZA7xFChQYEqpuvRlfLkc
clAbcR7tZjroJ1dlVqcOaIObwJDFD6IWDhKigKrFBMHV0+Zm/5aZXUzsP8zRlfEo
lWygS+iuyxZY1CX9QGyn0pCm6NKzHX0f7yNa9D1t4VCWuIz8gNwCZfS6KhJXQ87U
AqecJ8uHqA+drjRIs/znfUdKVV2hnmLSRlFAq5Cf/CNtcyWTiKtoFs94D+10bU/m
qQWq+LpUPFbUJ/WnqWYkVVzJ582IOaNuaX2VztMHVwjBCynOt62hwG3wBmGIeamb
YriIhGS1Ft1+MxZ2irf7sVmdmSmGhNoM1FB9S3zsKsDRPh5fZxY4XlGIkyFCbV1A
Z6qrzwM6lJxunhbNKzvC8kJyDcyuVvEV1u49NSwaENNCMUclHOoOXq1Hkl3n2n+Q
DhrD3eThx+u54/NyDbQ+Po1UJJHdRaZIT7s5PlO0hGxerIXZn83+G4Dhswtfg0NF
+UV0HAmGP8vgdW5ka4nelAGhjv/2Y4joUwtTVkc3gn5mrBbIhx7LnKUf2QBqwUEW
ko15rcNwag8xkX1/8ZNtrrALoaU+jloGzEBWy4iYei4yycxdlqbw2pLo8nfcdV/0
NRLw0XMMsBWGe/kE9+VYaO8LExwnH1XufaGK6oM/zv1dnKw1JuEdSXSQSdSBLli/
XnA6EsmiGCnifHsT9bxLJEDDNYTy+kQQFfw8iwt8AxGufsUFfjJv3QGnnpzfxYqX
WOT0WqX8skfNC++XOw/GEhVeos+pQ5xcaI+Mt2rNATX2NJ1sTXbekGbw2AZGxfuR
pZUCLQtrlz6T6UpB3Rz+siYKTsw913ZLNIx1LN00LuK+k7FxSIc4jlZ58+Qk+gRp
yxAYEyNdamr9GsZwL8WYIRYqCKOpWpQqoIoYkxZ61l3eXyo8cdqwwRhd+Pd4rwqj
w8yCeXbUFcY+fiSGAJ4zy3o7P0ldcCMhnMmXwXsER1zNyN3toAU7xcUE+inFW0nr
W2Zespq0WWf0zj1zwI2cW0ruOgm7+IiofoLZ4g30RfZC1yC8cy3XvukBDL+i9Q/E
sa9WshaJO6kCYJQ4XpiR4xZSHapBrPyEEC3nX86LTRUvNj02htsmLH4HnGXaneGz
ONu7LvHfVH/wBbcdSyq/yOznmDZCdanLQO10vC/nBelKpu3aQo49ER7Qh4yxr/ht
hIUMlnlY019q9yc3fifpgR4h13blVndvzKFF4Kpw1DUyR6coZts8xa3MtnjXWyeo
bbi5YVgvV6q+k2i2z0rXNxOR9UAQjix1HNz8bL+GzoocEmur7oQeEKO1RnkQg4Eb
31YWLpRI/YDymbGPN2qzig459pkudLOEhRzLochNjQAggIcKWKe8EVrAkaJCrUMk
NdCCwtRknp60XrsrOo9k7uEOBsMbMZKjeIv0Kc5eflTU0Gs0xqQ2Jbt06dm9CETR
8S+ltp08zT5tg1hXKPh8x6dXzMDFkxLxgcpWKJpoc1Jw/dYStXye0bQ4Jwf7Ew5I
oF+k/Ut69cGj6hJCebIeyKasJJTXZrt1aHS7hzkgiBWqYzmLJ9oyviOQUMlynk3O
HPOBjzOPHeXiXHr+g47AyAAgSd9k1lJXkoTOljR+JnCLyaOmY3g2UNJG+VJ4H8OB
nuAgcaVcySxcOPXZzJ4yD8wMCCRDJw1hdUADLhPg6oE0NfvKLBqOgDYkeXsRrHcU
E8ojbOtiiGD/PKgxMwOyT5sI4e6jfIiA19WzS1iAtpmF+oM/mWx5WCFiTwYdMOSb
fGz+JwAMp2PafpuSEMbfzOMG4WHifFPoabhmt8yhAS756Et15fzFqS3OiaqRnQvn
MIgNxdIujKsrgrKDZtFZFHDUr6faIlaECY3Gd2VhqXO/f6Pizs8CZsg9LW5mLGk4
PYun9A8nSxOr4AEWx9iW7eo+G0ZIsdurKZk+CuZ67LKPbLkFl+EVzloN8cBhR+V0
U/c6sc6d78f7d55Y4fl80WVw46sQKSRbIkpHt82DdTq6wW3eUYlCu4Uf/EewIIEq
hWdNiLp4P6XLWdJ6VQY9WVWFf/pUKGt9dOreNXPIO7yHFCu8TSPTUMBa3AUjBnvh
55pboXwVI5JV+jPhZtmGbYAXR9w5LSc/NpLeobdD8iWMIYJWdVwBWyvMq6rZhpxW
v08aGaeGwQrTt/DojUS40rW2owr26+mE3gEKfkIAU37JbTt0HsUH84S9Bj/Y81Sv
d8MSOYDAh1aR5C416Edpzky41Vt8ehl3HaR2UGHgAgpb1npSODpXMX14yag4/1Yc
47tpxBgegElSB/SaS9Aef91O4GE5aeAnxYV732+4pBRpaFmT6bWlOwFSlsXSaa7G
peNrbNDKhBfckBUEwSjNdt+gnnvXWmPG59wP3CxND3kzs05AtvCVfQj43gBOQ2H/
t26LCs2hNm02QQXyDBGzToGHYFw/dJvq4e0kTZkCbG5AUcbKCKvCFIloaOx3eGrj
Cj5vx7FGQlcqlxAyj++JvWBWi54WXmJGXHnlTlC8vA0Geiq0qiPEMbpZIX/7X8GW
eeFOh6EU3V8C3IdCsDsTDlBEKftFXh/RgSjFEsvdnVScYAj1d5gm0RrrZxq7Wvzw
AzePGQqJzX5NTyPnYNXgb7/ccs4zAkeVwwyl4zriojNOT4qTFOL+COgItwIfT1oT
Us60i1RuOBiqNF8yyGUjfbcqqVUVleDzbqLhNAY5zaSJRGYR4L4OQJ10BD1C92iw
Es5X0jXm6zdd8q4PnVTka20qe4RZCcQmxfjq84KuKn7NBlFdCIabgLMCtboCY8px
7X0tyw+2sSoI2WYtMUNBhNwuGleu64vqm2FQ0MF/mz2+Y65fvwAB6jwMs7O0IM1V
7qqXfiGtNUkJv5AidMX1yPWeuK8YtjJlgAPTcGgMWnis6cQwIOyzeylWynZzTdm3
VpmzcqJ9m3+/v3O064ohs2GlQyk8PI0RhsAHd/h24HH4wBBp+wf0DubD9sEsgDN5
yxMkCWy2Rx5DKrwSdoV5xbkzJj3dPf3VsQD3kNOrQV/b2l3qWTUgNclvJpyw4tgM
tqSl95jncbTttMthqcSunB5U9aHQ2sw62mZXZiPJhxaS6jfF9shtaxBUX5Sni72K
+scTizE8W9pkLG1QK4g+KirBa/cd+pbRoL3sEUVoGNh1cBk5ngbDKicHdLWkKkdu
ToPZwwDc/aHflEB8BhvkhPqTO2T1+kRQnrzLiZaTdRGRDV/XHqwYQ7PVmUu1JsXA
3f4nyYp4AWtMwY97njxq/NQhN3M9xQyhpOEQFiY7cdtWE3CSLml07h6j7/+29+Y7
2jqyzIgxZg+hSG5yrZ/BGbtfqOBOJ8LKRPK9EVpSrxDgQvOfQbJIPSPkBlKEG1Th
IaX4jzG162Yt1Gerc4fOqdYNAp9/nKmm9zvI+R31n5eFgJER02XUEIYtVHMlh7Fk
aqyRzhSzIhZ7jd2Yjmk2aGuDsW6PfMV7PBfTy+pODHvXX1nUjP87JWQl2M+JAKCM
JypJBJeLyU8nhOr73bh9vDQ6dibdnY3Wd7wEbHN6nDg1d2wV/FoA+M6i46MoaSke
VAoOHZmU7tRgBzkxT9/s9UblyBHWp3f0OWIr4WM5CbnZ3BHEzGrMBldSAYnc5oM5
BA45eB9VCeVnELgZOdrPtWiQIFv5XnKlV2gXTXTI3DG8bQwQJUEj+ueRdx4uSrJR
PPr5jyicOA1zmzPQV/aB0AA2CKxCqNpCtU6aNjYxGksxCGH6eW/fOaKD2w+U7vvA
nq+LznzCvbvQ7tsPMxvAWlNtg9+IVdVv/3mK4num8orgcCwnlB2netrTn5+yJGCn
7T7bQkUycziUoAWifUKQvBNAsBakP1hDZGme4Bc+n7uLlzvAK8yYIgpwNt5WlPpW
lj1QqQS4WGwFdIIqxwJy09YcREeh4SrCdJxa4ukGDvI8N7ajvTrfFyKr0qfeZqQU
/aN4QKmyGddAAKW3dxzFlGctJuitILzO+ry/jC0ykDNZvvKSqUmbp7NybgPjI1xG
ZHxk1hDjkIJioyMvBnIxO/w5c4XHBo+TjI4GNQcORWUYvHj73hAcY1YMBUm45PaQ
1lhfMSSvPLgAHXIjP9pLFLoflYiOCI5tXBwsb2+CxB+ONFe/aRW8OHcHbm5cF+VV
J09CnvqHM8xd51nImH5RPYc5LFmnvI74e1+uF/s5kfFqqaLnzuiYlcZ2KwQWxT+/
30LK9AOSuWyqzrx3Pj6Fejha6tJhggJn521BJz6ui9PHaNcdrM1I0djMy2xFi7DN
MQV7bZgd5IVlIl65G0at88KzNcEGabiUf1vaVbHMCF5aO8+4RA/0TxkREbSBdIV/
jbS7si7R9Zee/QQmDJXCgpaSd6/qHf21JUV61G5/f+OFnXUjicNEOTJ6Z9m4pktp
COnWBgPVWGyP4HxLPJmUuRpHY8EFsqGCw9JWgEq6wPoe1iCtVZyjK1hHeXhfIgMB
XsWl4rg6bH+w+n9Ln2eGYBpeaWk/LmOvziBNsOu55p2GbJshO6fKmyGyGmV0AJ/2
m6LmPygFr4t2IM3v/sa8qSWKwv3gMW3tlfuU9SNWw0MO37uTGmhcU57u0drkqQm6
LZ5TLf3WsmBCKKb2nleMxjCjtJ1Ed6xX9q0tFKDe8BjvignOsp4JvXOGfzJFvnbj
IGDI9ZmvLGWdxBJg+o93kjKFx4a9w48t/Ho56LxEiFd6Goq7TzxRIJJx2eYGhSX0
M+tqd+qSt5F2k/Zhk0+A1LTplGYBMlEJAmAb3uRkUp1nBAnMRi4AKydkn4sD3Cw1
LL/xk1NovaxXHqr/HSibe1/AkDotXv5XaqkqCtYBT2In71SLw7w4zL1Ucl1xRzJY
6m4NpJTvgYn+YR7MJld/VrbMLt3VIsdLiqcfNLv+NDljESLFdjgrVgyXgCvJd2sP
yFb6QZhcL/ZNPn5vwBPDoUvIkgZVu0rdzboscgrQrg8KwKdzJEK4xPOtcntNdX1u
caxQ0AOvekole5bmS1RVCFX/3dMiFoMKyFQyl5mVPqlYhOYy+hNujtERCH6yIQtw
j/QGXFrU8Z3s50+rGwEEu9jHVxFFC3533+oVapNdTaDJnegu40h8FL5mcoGu1Lq+
EoHDHGiYt78cLLDygqUyuCBHzuoFkbain7AuDvPH+RxAMQgumGdhW4a2exgsCKiu
qr9RDDj+h1XN/360E6VktWZ/l4RY3jb7sR13eI8nHgPOrnUb2BQ1QoGKXw4abtMd
jdsgfIg6sk6C7diwkmWC9gDKjml2pFNdqbwFWZqKKwEPUwWZme24/nwpXIVZ1R42
eOA0rZeSYoCfcSNSFm3Qxm+DcpZcBDMYTOayeHtOImqguDgxu/zmYUmc1kqj/ZgG
nSXMaZrs27O5RKtk9YEB1JRiJjJYVdp3HHE9RFbdDIQxqxBjxKR2fDVqnTW0mjwV
5a4UYjK3D6VdrY8uYlt203DRnoBKbJdVQK2RYIVe/jHNkuSfS1v5UUvOHu6RIDud
wvYwi7rvAHSGoAEvjvwei+Uhi5J5T/lMM88fbchPtUhhqONkJUx9g7kx3Mbggc+1
1ZQr+UaQqHvRQsjYTo7XJ+Y8HKh2F1T4iaU29zPZzd7vrgqA0byp9GjPwK5xgc8k
Z6fqW4EG5QtfpOXUx6VEqAUJw82gr1dABWbVt+/ytBiR5cB8XBBFfDvxm6IAO4MS
LVxCr5XM7RejKthlXM7iwjUYcyMIrCC5Wl2yUePKmHSLaGVcRL9dKFby/y9K57Ky
OHwiHVbiBacZgGUOVnexkkKEegSIDwIWoBx7Jdk/MtL94KTTBmvdY5O5XBnrSLpW
VSMbHjiA7cHP6nD+kU6sHpKGRjyxyxDVvvOV+FzF/qKGLGKWb3hXRrNrSH713FLW
WmPF63ndTKaLU1GWjKWZJBTu2L2opAvBiMakwlX4f46u4mBI/8wh+YA/go3dWOGz
LKAnQqVovVBcuQ2/bjloFkd9ixthHCB1UhI5OHmJaVC1bwh5nc08oKQOw9lMPxSs
tToKm3n40t3aiyArfX2KKQ4eCznSTBVfEeqMgCpiUsHNm1a1T7A5hD6HGXsxYWNj
vx65tYu8m8gK4EkMzK4Kd9RoGb/R29a4eljsmAZdKRyr494RyZoyKt8ff4Z1PPcq
AoDSpHXGJPn8ypzPx1XyZepw7wSDV72orRGKM1Ixy+si7lxdfrWGcfjTop56DuuA
9AheS8COSe37loirMUdsUpuYpgXg7inEu9c4L6kqDv+s0nY7uYEGpu+iRLv81kkq
tWoEObOlPBFn8hwebk+Y8svlW+VmBHVTLMoEpcAnQ/KmE2f7gqG/KzlwY5ic9JEE
YpSqdoIwhFwQxGi9Ml9PQQhJ2y1jyKI/UUq9H1FBjs90Z/bjpIvY418JN/VkT4F9
tlGRs3oOTsvy/144AlJIB5bencX0nsCGeOOo+z5vZrugssMcfMSZTIy6lT8b2C0x
eNHONek6Uv309QLVqslmLP+73ghknZ41Ge4VtKLDHQ4zjkypTeBWqeezwKmVyOzd
7IuajDhh8R8XMg0ryjQqqWydBpbP+M2h5dRBZERgaUMiaL9bPCo96AxdyZ3cm9Fs
L6aeMNqPknwpp+miBZ1ehBsnspcRBGmLjVamybYYK199F1k8HdTGKCE/7ADbIifg
WZDjkk8ZirKEpcRAb4spgk/lCsYgxkPpUwondiZrl7JPjLCZpJRq3g/6iCmqelnH
m7YNLC5m3jtOCPLdhnF0squ3UWCoGGYCmrKXC+RuKFCVVxLWqN9QdCQGT3kc6Nc0
bkv5UNk3p7I00CjBoqenvTYHpoWqaMKU8YG9iYKbGj2+l7vv23sf64YGabBU93y0
mywkAUmQmZUyDjHz+TpooSzya4Rti78nzk4DY5a1TkiA12i95DYGRfYQXfKM5CIl
FrE511qWrgMeSKHcF6QkeK1pY5PpG7uAjZ20ZonKzL/Elf5piDRXJbo10qSbDW+Y
xU68fz/cFavjBaXdUYzkkZT0vUQdvCiv/iwwpo50mdatC+Ib+k2wEtW2j0XFSXdc
O8iiirmpvDDSVNef3R8XRrjI6cZdCYrm3/pCdA2TXqMZV49ADhUxLXIoeJjuCSn3
o+gjuKXZzmdjO4Y2YaeeLJd8xjfQ6iKHveHVjzoiZBYJuruZqIfGZhM2cT4Ic8/h
7JumAASTC2McLs2jU3FF8EiZQBQNqXpaeI1aBvGL2NEHkoQgHd3OBfDdDzVwuCrc
0rgVL/hIUueScDiM3ki+6+Xct7f59AWHLnpM9pBaODmot4NML/wnKTUQjU3lGxa7
6+ixAMSgkYxGy8ebpzCgabEYwIN2WLIohjf9VGC9lDqdYqpcwdXk53gM44PxM4Ek
7kk68PS2he/TzIjvp3XW6SSPRIgZ3tiPfhSWDcouB/WLGMHrX3l2risaOo39mAx6
FJ0Ho1MTmLlbAkJBC8bBHN3k+FYu4H/SS94E8MA1jJWfydnbMecPoqPY2XpIl4um
DeUCWBTU5LGEF+5jkCeuvS+LNjU91OUMUHwwyCXE4XK/h+mBm4TL6qPrqxIj4Cd7
SETo80KIGR+WgNi+e2fNcBV59RnmSWKymp2uRZlhxnp2fOmeWypBnr7I/RKVdEC6
Q5/SBqovfLyR1dehCRm9SV5P7CVqam+PcI6x2VMlibnVEELGjscPP1hwlJDPZ+uY
TcGMtxqqHVJ+HoM/M+iylhQJEG+vC7nnddqjsMN71V8Zy7wIBBIqv6aLqPmB8Dm3
m3J5ts+HxhbW/7rzGIXaQ0zoJ1TRhO5Q51QA9ius5F1JCeViJCr4KYmm5Lff4FZT
YsleFviMbdWZRyZ/Hu+wmmeBjRHqC9lSM1PGDosgdFG71rwzOMbsYiaVi6HVf7gz
zmhNNz0jc50qbY/VaDvw3q9IfZFommDXacnAbvW0Z1iNYYA14SZd0V0HYaIcG+14
ee9N567oA5nSOblhoFIbbQKIvqRioBvaieUNkvTUZzzhP47Jv1S+lFKqImhJJQ2F
g6z2pYKnlV2qCgYn0LkVhE0wNUaYERkDDj1T4cp8VqPwnoEATKfEpjiZic4NdeAN
vnebXVgbJO6DTMf3V6+oM7xstHEa2KGPMhCj45FU8lM/tPTVvyKRxfRsI7uc2bMG
EXc3KIQcDNnh/E3s5QujbN5RehInqUc7Z+/kfSYPMYjzqxRjBVwSjpqVGNVMk9u3
7/grK1Y74da0ep3bebFWH7Z2q+If3T5ULIsQM0wpO6VRbb95eh3rWTxe+Q5v/nCw
XdDFGs/uURLfAd0/8eZO1dGDDlD3G0yA3Z/LRN4VyrCear23fvJvytxWNuslOfbL
4YfhVg/LFRzYdnN6sq7txaYMul7kpuV9GSRhRMwI5Bed3jcxm8GYmGIrkO2NLlnL
wMAplLXSiT58q25inXP2dbMuXMOYdxNaVRXvFyK9b/IUMSfXXYEXyQ7/+xxyZmnB
GudvI6LiJt6VkWvPhk6R6Es7unjJkKZV2ek5/f1DUVuVl9caLAI89wqNR6rohk5r
e9ygXOyjGCebAU32AUDceXrZ4Be8V8fmrrwGnyONmtqRBw7qJCSz16obBmVMYsET
ZBbNOcPGPIBS3RScCPMxjP73/pWPf54X9E0V2y6cMiaNUR1evkjs6ySKeRvLrT/A
9IyrLz+VwgSsZP6gbOAdPuqnHM3kCoSNlhdX5TsbnS2fhzUwjg92fIcCcgy9BiGr
RPslDDuL4mZSJe2tXfO45HUA+LGREACWStJL8h5rMGJ44BdyGPQZVDXqMTVg24sT
d6VKDHRj2l0BS5orkna2gcL3SBq2WXnVSIjREke7NWSBpXs6zycHfJ5qFDGuWn+N
jzO7kTsTA4TFVxC0XeP0XvJ+ItFRlunx2OHTwvB9DKw119K/yZXuGnOhL9YETBL6
oB5h2TtMYj2AndFNaHZg7aOFJPmb4XpUlq6lhRq0/JuOFuooFouAU5FeJkWOrDa8
L8odVPeRwrdw7K+hGj7M45TITOASfiS9ycVLsBEx/x4rwHhvQwOLRiSwzZvraLWC
1+8c012tKp6eMPS8qMQjvvg4hhTYS/zjX57RJdUg/9IIrqjV4xeLmiSKvD4O7i8x
9L/IBqtHpwldjVi3sI2OaMoGnHIJWqmVagZzt8iNig5z4MijG45vwqZE0ouJhzAL
NoeXcPRSjma6pfpTw08kOdvVeEwsiru3nbfqKyytwcMvKZMOHZZPhlUlaN6KFyFo
C3aJRqw/4WwOOxZ7JzNzfktMAp44gUxffZAS9/6mSPz0iDXK+kKky66PR5iZj2A8
ihasc2bjdEDRpYLT6wQWxBNeOXgGaRqqa9o9t0k2sSWCd5Ds4YJ+7qy2bfZustls
62+zzi4UXiRcI1O/BLkqLZ8ZCc8TxDG6haEUiwLq5oKLp4svzALZLAHoHtX93JrI
3fMY5AdxwxgKk349ggE2oHHBGU2XFXd/v+TwldTJQ3lgCimEL0q3YlQmJpmYPTxW
uOAORR7hk+BCNii0FdOs9p7CNxEht9enXcexABZNOJvUZOXpnhvvNekojSVod5ly
GR/u+JIV9ilSUhSQyyvcdUbHk2bIOK+geDCdh5MoG7xrcr7n6L4X9CnlQNY5me4f
d305xMotbd7JLC4lnIiTdpRoXfQBpLF1Wg2kWUxXNDPNC0/QhuSpvsJ/pv9Sd3eJ
Gu/ho2mS+RrpbxkH2aQZZM3+6lY3PR1CjeXiLf0gNaoJqlObofcWPJ2+dqCkgjVS
zcvOyX1I/iMvvhVJcbvLCzMUxxs0KNdrViJO0w+WujmBccARFpTvafZ+x2vQ6gza
V43GCF3sNheoHM9EuQkQ4tLSySJ5xGp/HPioeJnUWEWkXTPj9RJsXupCYg/CNZxk
JiNsFIAxC4uIpAmzVMQEZwDKsur1yh+U86jVRqgAZ8enqghWNMFkIfB31yZCWqhA
IDylWGuG2xaixttbb61OI15vRiPW56WC1qWlZyzp0kFb+Ruyfk78SYgBG43tN5qC
PkfuQ7Mhou1ZIPri5FWW3CxnKh3hE131OnZOjCKvSThclcosMHUnK2xfqjk7Y5va
eGIQjmtI99ScfcTgxeMwjGNQw2rOO4lWkyLca1fjJK4Utk/JGlqygnXrakhdhOBq
5X/OcIzMD1a2jic/BwDoiU9GD6Sq47dIVoURzkYxaZmdxtP/IYU4O1Jkt8ZfXL7c
tw4QhqXMJ8/oVatXcslBBYpO6ZFkEnaewRSqxPF2DkDVpuCJXi3wiYcHsUF/gUXD
SL9ExrAVz0p7X1cddCMewlWPmO0ixbhZHOnVw4cimN5RKVRDmS0ya24X20taGEh6
YQdUemlL7Y2IkC08KZ5jCQejSIy6RSSreVxOgGVfpoOVPkAe8dsDAu0wHwXBevEF
wsff3FSBueJ6hWrQeDH2HZ+m294tZ43/qBr0bu6SQemc+Clc9b/fqyuLSuL0P2+Z
NqdNpPYCLh4MSWCYXBbxQAqxpge1rdzr5dsbIGkWvZC6BfVyIkeZ4AHtnqfus1LU
FXB2Bzm2JS+7lD9URFpbJG03e8AWxtmPzqa/OZWBR1sk+gz0RuArxdBTvtCsiC5E
hLum9cKImY4yKe5RExCzJ0keWeRIEz/IkcCWytdZ/7Pn1wnhQ7kCnui7DGn/hc4v
MHGNGGmpusPrRvJ/EjviVfmVXGyymaLj4qMFOMJVzim2VTrhd8kgeLcdtq0qsAOR
1/qbuyDhkV4+qROgqmPEGgzuJavssRiv57beQ7PRm7xdL6jk5javVqjbH7jkrk70
4i1uf83ikO/XajdwdJZjUXeN8NboGKnKTtH32jepNVm/Q3vam2NyXEoW2YXbhVpc
jrG81XyLUmuZCCT8/HiwuB24Q+PhoZ0zkpSoZ8MgpdkOOkdFZ7HM4HDwsPJF5ZVs
SZMW25TtnlEiiQIC7rXSLEhOmYcOmLbGc5KRGrBW3btH6pR+FJpOI47r7cAKelhb
dxkuLyNgnMdYU4ipoMcuGhq/qdcwi3BeoY765VQpRfgvywcd1C8rFjY3GMJdjeQA
WyJXiO6xl4G/EDDOHJ0Ar05r3zZllLlWu/ahUy4CCuPo10Teq8uEAFryPnN1iXro
ckiPAj/rGmnS3eoloNTtiyqr9EjkBTBcLVGPDjhwpXF+WV0qf78SDVQiXpwKKrMi
+r5Xpb3KO5ZsJf1fzmV8b6PSO3DYtubT3IgOuZVun5trk8FchKuJv0J6MZ7CgckP
b106SnoD/8MaH1w1P5F8LXE3Ye1M4zVFw1OFCa95N8h3epb0/7EJaUhlDPXsDnjw
7BuwD2XpuSPOVAsceGfH364AoZkhtCXU05fi6au19x1W1QNi+igYU8/M2Qf6WpDE
AC9MvmDrqYcqr9U36sMKQKpsWuNPGNWiJ6mLPl4OaQOKYuFAzPYk3aj0DWbpceYG
XsgFv2YOTh4+8moesHJWIqfm4ejnqyG/ASRC378j2p4qwx1Zk1yaGGzWo5fjKz6Y
ugkJObHpL+WYHW11FLQ7z/ffz6UYomRaIFZv+Z8fp0Mx0FA3X42RerZwwbUwTVwP
T1bzizxOB+qVuRUxDG0tVrtt1QJfVNq3z5XTa+BpXJrte2+fasdQkXkZ1ECma1G5
KebaFDuE7oRkLb5GepoyM9jwYzlzhs9kzUIzabxQrta71NVnfNJLj7nMA2o/TP98
zPFRhTUhE5mt3/Olc0Zq9JGNFIT4HQGAa5Zf75MIfMiw6CRXPSduKXgvfPUrzYNk
BrI5Cuc/VQfK0BPVO/LylIMna76pQz6o6mKV5tn1dRzGLL3kJRb/SGUEjHLKPDOj
bM2R2LYOaR413/7oILFU29tsqpwlVgUJv0IcUTUncMPejLBi2lhH4PIN51n/3USJ
MI8GescrU/LtGVHK922fC65pSs+s+hHlvHH+ceQm/mTKTMZvy1ABdBQFXYvj6RR/
1cejQzjLfGbQRmQDsEmJ3N8ovmRWqJKgpbhYA3lRE/7o3QDg41Y3zd66ApGSmp3W
cmvydqFMxY8lRTQHeHF2KtXmisWAs6td4Q4AtjxFitNqIvUxJ0e4wD0sOJYp8llh
jsOkJ6NXwjssHdwt97ev4fknozwqO90P01qYY3cJsURVQmQ8BJ3PLJmh6Swk+cHK
rWvjui1cQI/fC3AJ7r+wHU25BC6Wt71tTnPo05ncOlkC0nBS+AZNCgP3YRPw9y62
pdiT5N1R1Fc6ODMCzVgIquFW3gzbzHN6QArp02Wh+kWxrQDpvJpchSxn1CS/8ksG
xevyKfTedDu+8HnXaIinb9NowbWnSV+lQrH5kQMmO9jAIWou4rhQh4kSaiIXYel3
RcUF5vJE7ClMzIAksZZsQkVzjZvksxE9UhZuRjXcdellIDzafUNWN6o+a8nbiLI+
ownL3iv8Utxs2vRhIdLWtoK++E7dtG5L5bTcLObX1VoaWvlv/Dt5pMQ8bdiEQMd/
pvxshZOjff0Ah38GymZg9Vr9PhCSY+tWm51XiBnpbeOSdeXm3A4Y5mJ9D79f6QX6
Is8H4Xe2ez4hXxppGViwD+3tKRpOKz1QxcgD75EjAsMHr7RSQjrgJOejSpiL0zoQ
5j226sxExOCY/Tr3pAeyE+LNNGeVRBZtWQWT0mwoztSRnta/W3Wus+8U7e6aJs7o
AdrqNiib+WLgIa4oI6Q/JbSL6sqYeHYxgC4nYYO0n7VtZGqRN4Sv/k79LK/Dytvv
E4d+siRp/AXiZiqbShXi+qNCwjCiR0zNF6baHY/N7u5U37O8RsXLIcChc5HnK6kE
glmEkrzVRHzaQfC2/V3f52M+057VmDMMpIblpGbC7ffMuTN9YNe609OtGhfuPwal
b4puVnLgQSgr57mfELiGJsWrymQCf945M6g2LbdIRHxuSy9AM2zF2QYoQ4gYjol/
3QKA1B4BXwmfQQxUZErPfKq9IueAr3dGyw1OQfuRaTqxVqJPLhjmP/NNy2Avk+ro
VyGulLu2hTILQZcYvo4hoO7TUOYlpWtpMQ0tpKU0cvQQR0e3mvLcpRO5xmEAzZpQ
IC4arLHns7vSjGTkN79UBUm9CsybjI6OqaNO3RD9yHKket9ZEIgZbIP/OLCJwCSW
2G9A0lbGdy8qJ5mNpubsLrwSWMzj2iv0MH+vaJSdMXOLXQUV2gxcPkK+Sf8F/S+X
0Km4ZXJNViWqtMvkLl8tFq1K/DXoA9o+Q2gjkh7goDLmcNSXmc6wgNzth24EfC+F
6cDoUP+vqBlpjEcPCw61W3K5ia2iEcbMiQod994yASQT4nXVoXybh8GXFWD0NB9L
qfC1p3WQ4wrHe7BvnDChTvyqKmRQ7llN53VsXozSbS5F2wUZV4FRdGl8iDWM7Uus
2a9DnzO+BzbiEiuRRgtGsAPgdgHGxNlAapj053G/evpmdOD0r+yRnNoY8DDBPIST
/NIqqqP9RgTxNolxa9AY1s5iLRoAzBRib8iTVQBRacC4u7Nss/NMshha1Rcw1WPY
h60jNcJQreU3eAShslXIo895mNz8EITSAbYXDzgT91ErrevFyS9j+PTaCBBCs0Z/
El11NizLPfJih9SNxq7cIF8uS0bW+Nn1tRloTcq5itJG+LfqzUS6SY7pt2yvAQL/
lMnziCfjsVx+5lUykpNg93XnrnT6i3/YIOaqIngOgX0WxsHPpXOVuOqLjJAbeGoB
77HiWOSWrR6rFL02aEkP/7PNnIoCjISKqqSfLXiNJrJsYfs1x5HV7A+TWECprudB
Cbx6I7VT0VQjHWQL0ruEbB0o0GgY0+OS4ckVpgAxa35CPz+wjbbif5+p+OqV8/HI
qtRuzxpN/djW7KiMb8BCWV9sPi29GW22+ygrT7ZrO5lyQrBciyHZZeyHwtdYA0fC
YqSOXYNLuq0NEJnddjRf+FcntWhxveVKUoeafUldLKONevXFj1pb02N3GWPuKEmb
NdJvGOw5gX42MqIBQP8XZd6tE8DrXFQjMaBcjx1ehWdd5X53mmNR+X+NsiRp5Axn
LZBY0vt0TX/+8KBDflgc49mFKQNEhvzAtbFN7fEjswoth3c4O8Gk/61aOILqsaHS
c7v+vfm2jWbtM6r0CkPcCe14Y1cZ2Y8skhJStQ+a20rD10l1UEFSFUiSv1MACnSP
zafm10/oWnqbMgoeHRnjidwkW7206Z6eFUjLLbKxni3pUg3m58XQvGrzEnJoBrlr
xdZR5TjlYmpYVQHG1cvwAz6d062iiN7hXmnqEyc9v13C5J9ifrXl0kaFQAap9vfK
tNkP89Yp3iaF3RnXlmV6pRkwBk2rwMFPhxtVMLw+zLfadZUDwmxKCHY1oT9faByu
4GEaXdnkAcYWBWYg3ZRQHnu6P37RsiMd54bfb7T5N1mZJuyU2qn2MJ1w5bSegnnw
ZE3mjna7MrEvArO32b8GxY6iG73R23pXc48JZp6HliwG/UbdWymYk3RVcP4BYxCF
hHAsL0TPkUtsAL8D5hE4/Vi5O8r6k4qIgPWqRalTFLcbS1+PhFbcaRVruW2gQEnv
ElPAuN9zt51S3CHItbr7taSocmXx8mM0KtU+lOUgEIa5KOG72jZ4lij/G8OqjX+K
FeuosjGZp1XCAOjZxDy/GnpKGMrNSf33xiL5gjhstKPeZ72U3VKI8q0PdrWBlJIC
WDzbsL6QsPFEIgsMqOCzzqChu0lmrdIyJkl0bdiA7Gj0gE+Gik9/IXVaqCIJm8y2
uJpFDEcbvSxKj5nEvrMgz9Sk8SLktj+FsrwonO0cPKwSg3RU0T3yxk6TVFWsH9KO
RloNGbK/vVVVcST9PsgIDDfqPikCU9ZxXx6XGep+r0LqoSh7zQaxpq0hnFUFvFa0
EPRgSwLh1eJr5DLoZGnGTAqh6OcD1XSET9D0xDpdrhCq+pWz0+s2gIU27d7XwpgP
WR+vbkN1Uxfda+vuRCSd8qvy5rYBum9ER8gCkYp6DQ1zfuqcvjOoFdpaezA2u2T3
tJ2ybfg1xuEumevZXC+CIN3auLoRWR5v65DxiNeDgF/BY6vMnIeyTsI5BM86yu/G
yu4UHnWoJ3gbT2II01JISHO6dv0Wop6VMdsQa85eyuQ=
`protect END_PROTECTED
