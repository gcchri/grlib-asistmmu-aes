`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jiYJXsVylcYvCcYt6N6lS6VdKdkClRtE0wlhhBCpx3+tDfclQ+QX7tAOESwVP6Xw
+kDq4VPmrva7vcMKfiwXYeg/Q20Op39K7rTIMHzwzVqwbhfSTkkK9TuWZqwpTldH
DL8ZJ1IsVrJiqdKr65gLy6QDMLezi3fFDnJQkqT4uqd9O0ERHfogaTeXoA4g6S0A
UmwcIymtgX4pbu/2PqmNsUUn1KlPeQBKXd9V491Wtppvro9oZ2AMHki8EF3fYrhG
zUadGgyZSy/mh++dtFWn6zzDovt42mD77NqL0Yb4w6dJd2il/FRQc4I7xyktsFfW
SUw4gY261ZjR+TDuiM/0FJCcRZW2gu5SVco+ssVgOM3WqwbQtiG4Skx5Q9CMsTvJ
M/uuag9gA+oTNlNGJzSB0O2uX9OKsn81QIjPY0M3aMbK28tQO56MAtu51EX0ppV/
`protect END_PROTECTED
