`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
js8sdEd4r2Ms3rcb2O4g7ikDY/exeE0R5Zs5aJpJI1h4l+NkRVh88i6sIDr66TDt
cWVDzrwah+8sm11GsAMOXua0Ndwk5ClXLVC/GGlEeFL3yRNeHt1bQ/YQPcDC9lTG
m+RykrlItc+GMg30OyOaDFJlVUafKQvJt7eOsOOk727JxWpfne8EcLLSqetwb5UL
pY8t70igua0CIIQreNgpQDiY+KkYIs0Jfc7mdtg/KSChsENQl8yAwnAS0m7Zyc+q
MQ8xmJxO0tJ/WZfMEO2tFYrZ89Rnoha+XQkSshK+I+frM28ql/CZRDNpSwvkQFl1
AlVIXn/U0+gChZ8IYR15IWWnAO6WhGaPfPko/EWB3rhOIKCtHqzjVHaVKlTbsLmd
W9zmOrbrC4/Nw2yG/ZOvDvtPA4KJ1Ef07mptuhe/JjJqc0hUqwtJ8m9C2pSaEkcm
CGI/Bpq05E0J+Coxo8z49OMrhxFyzRBzO1zz5T9BvTrV6NN6t0NrZyygUge5WXzK
vKnmI6Hydf1jgdMPNYkGM+pgG8A8YmRhGsYw5T2L69P+G1au+3xI+dCJmdojqKqS
rSYnoItk37KaiNqF/faGeUgt9ANxbFeV8heiOIHFBl1TBtFjKGHLYQEDGjYi1IOA
LvjKIjZNOwoosmvEqOC9IMghJ1opCd/wzodm0TrQ59um9LpuoCbTCwLPh7lYKRlm
FO5p8ej+krzrPO+vehdph1OF/7o1BNjHir93CYAtxy30C5RSb7P/aBIwLRbSxdtp
N61uCbTWZzxgmHKeVf0tfCjRZjUbXiHLAr02CHn/MvsueBg7XqIzdCGaifZrndLs
E7dspSF17cFc2aqGfMEe3Z+on38Ynuhg1EUI+MR2s66m4WgytnsFci1h0smABJYS
qMeNatM9tWy4ATVOmB9ZdEGGBqg8oygITqBPtGVdL4znLzwkkQXJcX1EXGNjsWzI
2aD0HL8sKYGSu3aL3VcDJ4syy+iTbDfvZj+Be24WCzg=
`protect END_PROTECTED
