`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iH6kXHwkM6eleFy2/KJtSrwg+3UmwRe8me2rXpk/JxmT5Bjuz308ls96G1EVaF76
yF5dwMJndXnF08L8ZVYkZ5X7NcLAVHlZZTY1r1D1ML9X2WT0zE4jLaDGFIuLc4t4
/TV63f6xlZOSMLyWB045ThYwerezgJpQeiIqD+dAzAa55tHXNWh1ofbII8yyN98g
2oQhqVChNhlBgAjz3r0UdKpUzXVsUKtYH/rvMX79zGJN+pBX+uOy8BvJO9hePMBP
VwA9NwbrL7Miv7v1XaQQw1Z0bEPyEdf6mznc3GD7L63dTjoZhFz5TkN8gVI7dV4T
4F4tl/yGrvEAJ8n2K1OSIcLosrcCG9NAIRuvOn3uU0f5gLAoRIyuGvuuoXNbH0Nm
9qYvfVcifYNJK2bWgmFc++EXZmm45V8vcFWfLksW/cpX9lq4SNhuMxDV5uHVkZ8g
tRglW0s/2V1U+XG8SBOh1M4oXJm1PtDoaUptOoIPXTM0QicssiQUpWzkWvhAronB
jYvXj4dIpTWRA7hwfNSXZrTcE76ksBKnwRnjq0WqwqCtLA61vdnMrGxF2+ueE6DZ
/iwYXtT4ueZYVJy7RfNXLhB4//PryqQDi2K59ehywCZXgtVAmnev25blcZ+K++sE
6Tr6w1KjQnV8dER5/Mpc+67dRfpLO3v3xhZGiN90b4Y0XSRR6rxzE53O3oBtNAP4
+P9ZqmmA+WO/LyqbfCxFjNqEqCgqsURF516y+idvWmzpzluRUeOzzW9kHor1/NCq
O2fPb4djEAE8H+OF262SDA==
`protect END_PROTECTED
