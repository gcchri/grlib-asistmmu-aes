`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z2n/yUGnd+zoO3jNgbm/r2e5v5cT8QweWgBVpWfKIuzlAdJL2jENckqfFHsqvpRh
q4o9wTZLR5dNis29zvzg32+WNpRNPBF2TIelu+Vo8Wg5VHtD96W4aom+olhPHbkI
MqQZ/sfieP4WOlym1+acsOvdiGeHVOa4sNubJ5Z2iJxJsHIH/CsGm5UFVY22DmL5
CWFXiFHIN0pdaOzPKDRXgDTQUusprVXgWUeBCezX7scu9F2G6DTHdAAAFD8jiUTP
W2dVt2p+7oBiWwfPuL+Cssc+f6dcylOAKP3ctIK/KyRoWr62+bmIjFGaVgRLOkQT
zou9NzKANLTP0D7hSdpvq+gnHADMqjTtNZWQMhI3O77uhEkolRZJeTFrVsEyU+qK
L70ahe/4Oa9LecxL28UkQr2bWTZdp7JWbVafED+PZWM=
`protect END_PROTECTED
