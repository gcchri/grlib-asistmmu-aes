`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
899AfywKg6s2CX6LwzYiEmg2FMiEKoWlXg3TQfSb/lWjHMcH/u87ytnOoK96bwjY
WaAizjyVPZdREaSPuuptiazNNIU7Xo3/+8qF7bOAt3ogz/uxx+YqkJZaoglgvTVQ
xLoZ98DzDmGVMo152drU6X/EWpEqvZJoKxGLZ/3+MqwZNmrSwB/b+Pvf/Q4XK6HC
QVX4lj0BVzy+WEhHyQ1IwKgm7vU2XwdoXV24yvxd+F05AD0dIRcA/j0SNLg9bYkO
wcTY3KoEGOimgGaRcj8LhQ815ffIHx3w25dEdDOztXiIPqa1cmfZuIXtc0DeJoZZ
zsavKJKYbx8Li/mjDwQDQ6BRow6qD0kD9ObuLqfg1RB/Oq1puNhW8jML/WMar6cr
ZWsTY4lnzAHl9BgJgAXqUNa33ZgjmqNKUW9U0uQeHvpyTpZUsKXqDwP9CqSpp2Np
BZfZdKIUREPe/eHxjgfFUxgzRaX6nSmzMVIC3ISbvSghpc/p34c54Pz6HO/gXfFf
Sgjqot/GTMKdiysOOU/GD09+znidZkf0X7AsmFUA+npD2mXl16A+GV+Ks9nFBJGt
RwcXXnmwxaIji/TznaE6yOEY6x9pTHQlq+mzTSzKfyod247eqtD1V4hnVhu2FFsO
MMq9qEPmyuxVRcEMxuLNslZFlmGDUc0vae5IdPXoi8htjDdOtot+EY01udN/DKnH
q4zJk9jw4wkUFDj8vmO6XSO0N/A5jggl0aBCTTfKPQRYtBVA3+5A4E/+sA3VIqGZ
g3PgD/uEV4CI0BEOG5eGa6shTAhH5kzgTjxSAtXgGA3qATI9YsCnfiKzjzlQv5tL
GgUaf+cCLZivy0T1tabb6wTgSP/Bhti8tNRiIqfsCDhjlJJM4HHbPlLP1NoPutm2
WEA3KNoezIDlaJGyz6ykQnNJ4Q449+oiRy/GiFMoFQoKTU3SRNAZnqy4i5wxoK/W
Qh9r1ki4F56DLFRBLAgCyQlB3q/uJaiIGIKz7qtbCPY=
`protect END_PROTECTED
