`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7dBO+Wp4RgddAhIfDwKXbzrdbXdyO9H/1To/Pmx6WNDJ0hXKPfSXmMFTf93zK6I/
H4ztxqEgWSAfRgdD/wv34t2zx6u8h8TXbuwzWz90ckjPPhAK+678SnVkgy2sBHb5
eHdofo7FOnZIe22X1RWThAh5Aftgx0t+XyM4evjCiMHOFd9D3eGs4LlI4i8wVSm+
FZY+93kgREFt0nxYad7/81R7AQiGqMkekkH4PiryP3Pu7NDg+n55VX7HQWDF2CyQ
9ULBY4F69qbo8OBFc7cZCcUFeu7LwArJeMIMD9U1uiQFRLv6A+SOB6pOEq3WFzh+
KloxYbyFKequwgVSFhzsi18Fn2XOQjl9liNJd6hxU0xkMai8wSGrbs01cnyQlE8G
nElCYWJ4WOXTSoCc3rpI7eo9LjfWRE4mey1yQaiWmi2m3oJO9xj4PtRSOKF4buma
FuyVDIIhqAuyTb9gG26iyt6me3Pxr2AC7UoFUYHyL01Q0YV5W8kxvzZJ74a/laNe
Q9YShFaV0WSRwrLQQgeAoYMf9mzAuNV+xvGGsToJX5Th26zkJRYmOYepRxeW0IbD
NBb/T0GofEFBAPdnVs34KCewvMOXwao8UzTc1ntqXYJVTyHFJedd3kbbETlbHMHH
yDtEEeCfNK2zY2R7D12Y+mAhEGj4If/0O2IEQ6zWzz0YV2xxkFTKXQo//tFArgLe
VCUUrLV4Zce9yWtKp7e/SQ==
`protect END_PROTECTED
