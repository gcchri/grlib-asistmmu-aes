`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fIFMckUSNlpCoK8ksEUgV9WkNZFggp00WKz0bF2dS2RdBmiu9+kupgbAIwpf5ymc
M3RDpYvHIilPiBUkYsuKi+JemnM9tA2K/1JqKfuu005F0k15eLDKy2mimbPgGlIK
6mo9LXcRO0PloSXLDYMI0B/G+nYOWsUC/yJKhdSik0qb7euObuy2vLEgPpaU5zQX
6RqAeYKx1Tkc0wO5V89/QlvtL+rgAwOou382BmmYGtA5CzttobjMjHZAojHAgtwB
e18s883IkyOwp3kBVqhAz2bHYRtmd/LkjlnFvszyVX7yhOU/Dl35GmUtyrOnuGNC
zSmOtK230xk5i/L3C9Zg+/Ckz400bgLS9kMEk6vYq7mOeW3zHeJtoOVJU7u1IfnP
yVtQGuaGSiiw05L6ObV51euPEYq7RKb0qsPLL+LCJCUoH/DFa9WnwaCT5qe+xyZD
2rnAIIhkwTzvMSpJDkYpHjER5ZJXfxW8ezZFB0UlZc1OwOHN5giX30fnW1kPmcrL
tnsQqxnK/96mVTTfG45TXrdaOoeohPopRn3iEN81xXZ8LQK+BFk9iKG4K9LHYRrG
NT4+IKuwbaUpnzkB8/xMBWfJNddnGGEZhsst34bZBd8PNXY4w/eNQ9NETvs9Bt/l
E4Q7/Oo3peMAwR+amqapZqDU4ZpDZLqDfyiWIvvXsDB1uvskIXz/5kXV5NZKapa2
hv6NGFRGQulHBOtmdwv0hzJUj8UZr3P9r8ygH7njJr09dgAHaZDqEVkMGB6X95gK
tbYNAp+jiQ160yP3evfB2cLO+4BH0gG0gn5u5fXdL+OsVbU5voDZWSE0YZazdHIl
Xzj0FKM8JhknV3/w2w3l1QGfkYVCvAumMefrCRFabc/Aqi8rOf/0l4teTtKhtd90
78xZBphaUozYtUhyCE1qRo48M6dUZGeVYZ1xAShInHyKtXMDprE9QxBPZ8ajlTbG
EzNA+KOARABiG4Z1uv+A8UPsqRucTkS3HaoEVQypKPxgEQrmb+0Qs2dRiWWwIWHd
hB2DXNSvdyIMVtTz+c8w97LsCO0Xd5K3aWHLIiX3SZNTs6usnv43cT0/YO1iByhG
MDfd8MaRMJKAViukifMBlChy0sMWJMjQ4b/DgsAsDeHmeHgiPEv7q72xaYfH8kjK
VZl3RL9H7swTMswnFlkunz+YABvbEun7KoXrayw/UO53iZRYO148dLjhOr8TpTpS
+3XgpGr2MB3mi7v2TGWhX0NzMLV4JM5bgnRYFdC05eFyS1b8K3iclRChH9UKa17q
GvxQ+BlnGr1GRALcQg6whrGxb7Yc3P7vDp5DMqeKyi8NjUt2cYygMVVB71GKCzNZ
HQE7AMce83A8KkvOxebBsLTAzPj6moVM/G6ouIFvJVjHL4tAQzylC5keO9qQpnRx
ZDNr05OkAPJdXl6ybEqYvb7bU66ICIwjryCGBnbzkb3h93zha1b4ymxZv3Rqn4R0
pA58RNuYstl0k/CGVoDq2LhxdMWgVTz0PJastninmnlMTT/H/vl38KKtrwHNmO1z
Va6sYVyR+sD6+vX1198jXnlxe0769rOr/ve5DKwqeXMldkHA3Cmh5RA57jZJY5uv
1Lu+KtLC8vqdZ+rISCV3D6Fur+zKUFdJPNRhAok1noErNg0fCDFjnbDY8gK9KeSQ
jZHMLwX+Z6ORo1sKA+sBhRi1mfXv4do0AhTs4DN8RIlnVPFY0gJSsqxWfuYFq1Ri
iUMXfh6TNqDsr+DyqNchE4BBGk8Wd9IKE1L+d2ArwT+W7lvuh7evUOfSlh1gJbXL
/dP5gOwc0ArrL2hsbgD6PHDAyh0mErMMsmB0sUhSRn0=
`protect END_PROTECTED
