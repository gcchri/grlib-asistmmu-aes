`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZOU4vDGzWXp1UXcBh5/5uBvbEZBQKKDqBJA9zACeI4hgGY7ccs7TORdippflkMRq
pTt7cme3TOigxBhX5IlMQaPPRBuR3mUiprR6Bjy/Bl9MDWt9zRBEIHFCNaTKnvlk
1O35hWNAW/XmZvM6EvGZ1oBinEhQQR7Ra8io02pPu0IWc3JzBz9QyYXIflgI+PRO
79i8gBmPS3EgG2CXV7YS6gav9jwn8ivCKd8juD2qUEvEfDZ/qguBd1lr2iUKWHqC
tDtR1SU9BAlp/X0mkBz0KpYLIPzfqhRIgFnkMUswgsmAgjek9Pvok93ot5sXg2zA
D2TGhrlwLUd1AMTFqM2cbacyFVCR7tYPFVqioViR3wdvMS1+aahKU2K2pj5eEYVu
RyYGF/YhPRu/AMsB8movsletN06sBY8Uc4fu0IjmIDxh6k5/2QJmAYefUTnoQu+p
`protect END_PROTECTED
