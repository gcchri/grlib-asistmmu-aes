`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7tuc5pfpN25DPa2hBNC1K5dX0EalThYYFMKL6TUgzhqJYdyINFoWzCAeJZwLwTwk
izjcytV60Hw4VOEsN500/l71SsO2eJ3BzbAqDAKRlcy4VxYNL+LRdeLuKzsax7jH
Q/od2VhZ5vyvQJhkzTyw4ZVlWoAgno5VCY8iGqpPdXg0GNUxp8T5tSBaXnZwkEfG
ptD+GnZZTC+7o4n4mY7rdG/b1hgKDPJ4Qz8bXnd/fvc71u8Ali2OPELxsdt5YQPW
`protect END_PROTECTED
