`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r0JZ/NsgvJQA9rKk0nYKYHDGBVe4wOROIcvoskGn9RA1mvrryOGi8oLwk4tcSowY
abwwr6XGgVJ9mZmBMsL1DvADPuByB0ND6nglXol3UPOhNV8F7DIzmmWS14+MomB9
5yYE4kgzMzCfS7YoxJMq0GylhO12qTL2q27EjJ4heTLVuENi139VMmGMetq56G2f
zqFWIxGP8P2BFkILPXhpG88SLM+mj4IPRZhPuyo+Z+BPqW0TZ+GzcCNO5YBKDkBs
gNK0RHSciwUQxm4OTBladY2PNlwVgsDPSbJmyQp/idQ6NeJkmi19gvAJdCZCUu3R
ROp9MKHVB1orWmlFg23O0EMFp+jSose8IMiMuM8IcD7aiC6P7DO0uyBXYAeAQAON
nS1ymBgHNS0iatlrFQbmBhPw8bgA0mpqJtc6mnZo+I+tj3N720N4haNyHRSVi08D
KKx/sHeoZyzmAR8Yw0T38a3DgIgmtDo57qr4GqacKj1MQTGneCoCNTQH6VgDSTXv
vowWaLvZQxWy5GhJ8wEyAa2UyA5zg/yLmN8Y1AOgSoE=
`protect END_PROTECTED
