`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zcx6ltYM8t/3jjezKhanJTGlqBi6P5sqpUgHxe5w0qgwyUJOdEGVfNK5WIQPf5CM
yqOPoHUzCKsKe148ojFS599lhuSBbtBcw36hUA08+sQVFSAUD2D9jjHEmYkOYFve
OFq18n7fQhPV2RpIAvoVwST/L/VsEA4Ra127gbWX2n1ekIpz4kxCC7qT08naf24s
jusIyhwwX7hgLd4i8NYLX/TZG6EZQEpn2liP8CAjFmo0mHuS5A657Pt6L9zcFUtC
QYW+GXXg9K+XXGYrIVzaXjHNw7bs/rd+kSWlqA0vLUQSn9T1uSN5mEKSYHgnO5tf
raes0+LTXXd8anmvWNFuYoU/80bfEibgaVefiKNZ5Q0uCjE5Wx8hgK7M+SBFeifQ
wHtOIIZutpyMAqmCn78kC7UreXcnj+ZiPkOkrITU/OQmmFaLPVvjljzWHzpxoWMf
+ELi7nUGqSrMqkytC8e3U32tN++/W165EoBD8fDK2vRWAAU+L3sGiXb4NrSuTlcE
99LmH+j9xSWMdzVtJxhCuEi/oCMOwgrjbaua1fE4el/bV0scAqeJJYi5aYChDzdX
Us0ipnR+W9SXBkfwp+6kJFITywN4r0AoqUEhy96G6sdX4W6qcGf/N6fg91ABCqi2
Eu/zNOl/So8nHMY0tgG4nfe3OPWfN0kwvhzykNahHH1KGbr8d+c9/4juDRjNpaRZ
RbwFVKXdm6bYb6BmDTC0wVvgSPKpbqS79PxIylBHHLaXaBjjW/Qbue4hNc5ItpT4
j35skLN82/fTgwt69MI2HnCtlLOi5v5+x8OabMe2VH4WJQsWzsE5gI6TyJwTJ4pQ
uA7qPtjGvSyLbeoywsOR6x192upHczHyQJbKtNhUQ8NI4lV4Q6Xclk9V86smurYX
3Unx92fwmXILLfxSD96jIK8JLTy/I5PywUFuheqh5B8CZ4u53nkDYELiUPQZJIWL
SdSOC2xu7eFBgfDJOxo6mlppzaVKeUgxgG2lG4EcLpztS14Jy/6fSEGk5XPjEwye
7U5wSIotoaZeiZVO2uPk7fxmT30iUWqa7twmbKhe/MfJL6KzlYzfeVcRA5kNU6zZ
4MaWuw8MKVgT/pbGxPO3LKpN1tpVXAbxObMzqNt0aUMySM88X04rfkkrkbk9YCG8
sHqFTdvMRuPPUsfEMc+uz88olOmyChuniYiqVNk3Q8lWSMUwRYUMLowtShOWHcfl
mVo/Wx1OfeKAEKUV7SWSNuoOQtax5KESohPpeeBDHkRCPvV2wAx48xmPHpVicDJp
7MB5MzUSoJoN/WjO3MvuVrntaJBh0pNi4tjmEH5dE9DQRiVz1Hmp3FC7CQeMFq6o
UwUf3xh01UN7UACGZXOzmscGu/h0SIvozehR0Bc3+8EfvdKpsCE4nl1NDJJKN4Ui
uSceSRtip1u1mpeatJwljShYROu4/fOBwNrBops2VfMDuB44zIhN84M2iUgZl1C4
biCwEvqgifO2i0eIrqtdoZdNOl9r4F9PSiVJqZ4iHrrpoMZMjKUBXY8rWDBLNfJg
YhxgHnZmtE3OrVsRCsY3LpM+7uVCjn4ywF/okPrhChCsHD8Qc5xfTPW3C2Xau1pL
y9PNQVBKfZkY3BZFWIhmg1yqEC4viLLWFkGoUfIPmenK6ipU6t7HqcqhZtHnY188
5AAbFwsS7uU5Rhbrh6/1RjTGVMuY6nz4nLoEsRf1q9w8tC5ZgdeqiyAKNtALvQZ4
ZqkrmTvHwjqVk3mgGSCYoGzhS2dw04CmOpgup8WRK4FKuZmMykRqmDtux7VzBRun
Jc8zBsoGRsiKZro6nEuQnCZrR7MAaZZiMgzxwAYkbNQxNYL+mX/JUGRayNIxliiC
Rd2QzCOcmfLKXY2lL2h4YPze7TezbVDg0XhHePHeauxK3tlTiNJThuexBgslEeD/
oWQ6R72xVVaX14t4RMkpDddaunmSzGFtbm1AEJ6S54cv4/dVYOJfmzbKxohsegW7
Oa0Hf3scuP+zMjKeL95wVir2Ha0/P0uW/vZLAC20jOTBbMFV210CqHQJgtour8Vq
yxxSz7+XexrxRkRf0uwZ2se610vatSS2V5TiWSnLDDz/8yBYfzdN8gVHakUL5yzy
ZbpAh0ryGZ4dzmq/jU/F7aajPxlC59c0ytawp7AtzgCQ7QJJoxEdXJvDQEMbItjX
rpes1LKXu021+0zIhB0P7BFxQH30jLMFtFnxuzleRTB6Y3MSlpG2qrMt2dPSL/Qf
Cq+xxP9hWJcCCJfVWqfJ7UB/+HiVIXNFbBpaCcmS86/x3tjxNP8JiPDqA2HecEll
PWjSSVszWRsWtSCehSGMc9YKDhQpij9/mRxa9WeCg/mPnyrL1WVvDmHIzOVudn+v
VDaPh98BfAvgFEwPO+0X9F634UBNOTPnVZMfT3GMyqGKAi6Wo1P3tW9noTMXEEPZ
2zaV/h/Hy4cr3iw0H6sJSTGJDu2s+EDEYt2t5v+USBXLZdIr0w+ZgQyogTy2ahVB
LVZLYQH7bIRTyTCerdRKzMAFfqBRhLlLV/AtcKsfLPjRwYb6hx/6DEKYrh2RhPSk
qP1F0S9ZQgMwQroZJJ4LjjhF+PUC0BXnZCI72mh6e6+8S9m7aK7yRD10aKgtN0eO
ocm4e2bhmX9DPR/xSVAlUpLos52J8RZG+7fz1qCAEfPA6sQXeV8tyHGu4aQZGqCL
Ht1fxQMvsV4RlpQ9ozuSmKGlzqaqcGvhaeiG0t0pklfDf0LRhEl/dJ2t6g38v1A4
ImShudJyWn2kn3S4LZi8+Pzwa6mxvkabyk/mC3O14/S8GovSuLLh/8whrqyIjSIq
w+Y+S71RToiVuLf8MldABwGOKbmMZqVMp/KKC0hRlpHZyc5JI04o6LuwU7mpqD7u
rjgLl9l4J3goDzT/0Bwjv3QKN5IqfsMEn7Uk881NFieaYoAUketLLZGxW+30rviE
q0JXN3wFD0NfbbdCq4SK9AVIwjknmHNGfCOIrHEhUhPKR1ib7jzzrJwu/l8J4Nc7
IVOGcqVlUdCcmLfw4S1IcGo5TjxYM5MDiuBrNrtYCwDbAWoNZEL5ZSvKOe5vcvwT
36G8E+o3/Ur6+rh/8lr1ZsSwNCB4FCM1YJDg34OZ7rZaFtdv3cCh/+voFnxeI8UC
ivNcU/LFNCdZ5Xf9Ixa7DEe9ey3otsjhLW5HP2+mePKSTzCKedlvv/d8bL0adMR0
dLqym2+ht2GxsiRNOlbSHujMd3uqm4mw0nhXrxOHHuuepNDGnjewuDUKnV2Hqhmy
HKNn+ribzYBD3ck4JSfBjSBwB+vrYCdJg0+uC71h0mw1DkWPqcxabDyqC8Ifuods
g2ZW4JjB8h6F0dThIGSILpW9p5nMhNxWex05xet003vEQuaM7iXaFyvyIdr2RRWB
4PXZF9nTstarJAWGPml/iEqGSbfdZ+LboPPTZzNpjggotSQuUUfX0+1Xrt5nT2kU
ef0jnDcBKoAEtobH5xszCyz64IDalLqrx5Fjrs4CBHak3wXlvGrYue10uZ65Tpkg
70zNVFHgc1oq8GoxUJpWvEqtbcTKiTkK6Dh+pxJBCVVgr+hViWz3Cx8k74GDE4po
VcblN+D2jRprSBdLUCJ3VAJd86I+6zwYGTCPWUSeczOMwUvlvINq5swIUjXgI5/w
b1jcKVb0wEZD+WwhGNRLOnAyDBgJUYOXueMMXSmyoh27MLB+c0TNgs28L7oh0b6X
dxaSyYunHQd+t3F7Y7G7F8yNB6MY8ftLiAsbuuFk+OxcVw24WM4laPqAnSFVk69F
K+Kml21+WVYdjLpyiVRXbbI8FANrjmOrhxNZYLLFplAog8YMUuxgbXYwt6B1CVTE
UAgIgnHWdZxYzWKpQokx1KF4yfNXFvYdnitCuuQUHVKL7znatmC9cp7zTyXBQI8M
qVoR0UjpuoYzAFUFGutYak2wXtIInhUf/q57A+p5bUaWwfj13R6VhMbzJ7qOCdHh
9RFZIHCoR1RwwJUkdAMsxEckE3NWt84+TY+P4q2kT6nmD9uzufz001Ajq1KVmwZr
H84KFfAE+mdO4n6P7Isx4YVm2GmMyaHySmOl9evkPCWCv3sr6rZLSuX4AYT2rqDp
GqbE+AHzwDXXMzcdXuGdd13Srn8S6b7SWeu8h8s9t8d/IeHMvzQepNuJROqOKvvM
fA9zLCbpWfHUaklzlLtW8cilgmdt9vDUxhzie4B8med3VE7lsAWvDh9J43WuysGI
dukKksgYs+MaRgy78Pqwzf81aryQHDShBk/PR3SIPjTeFJzyHT6gWdl56NK+PhS4
G12414Tn6fAqPiR3XRSoquWGe74us00Cr6Xkmtzu0ozq3r+x4d2cZeiu+L0T6n4k
OIZmq2fRWg3C7rOOK7Z9EpYdgQuRh6zInx9RmCss8SHrUmmi640AGh8O8LN4XjVU
2Rbs7bDyTgZa5z45wlkrjWnWm5rcoWwRuXkm4E7HRPhG8w3MIA3NL3m6O9SdRd2S
xP97Bs+kWSzdaR1k0v5rZeQefsCDHWAR+EMqp6aBsglvnYRO5l1yDZGBIFHHMkDT
8pwLrpCHlvZF1VMJOf8zEbyOak5fb9x0Hyp6iLf6fJ/Ef8zouArU7Gk1fxia+vjv
arKpyWtyjUsyCeycaQENGmSZH9R/oCOfU6bw+cRjOdxqWt05lsz4WofS5QqPhwvY
A2RZI9tlEP7DE24KzqfBMU0omfZOyMA2qiu8soq9Dr3jYglphngwe2mzGw6IOeea
8Vz2uCmBeti56+43w5rY9v6QMYYm7+9VZTVcSer+EvXIFv8jBLBJUD3bwqAgwJ1E
U/cTWuXtncYDu21vs6WuSoIhTxO0tp6iOI9AtV0EY2YVoxBvoXsBW14ylxPJphav
ldZOhLDIXu06DLtDIBqYf3J8zJDiSrCY3KrA+o9UmvdIAGOIBeYh77Yi2IXGJt6o
c4neGoCROmoaTEfgK/xeB5JYod0NxScU962UJvh92iLwg8N1LNaA9ORpNP1EBOKU
iUmDZnMTHLUnK79Z1xK51bxIHzNVpPvgf1s3242Dsi0TW8EobsdxYyhvc6vt0bN8
vbP/byx2QQqLlviu+wBMD2Dmt7e1kkSSjFXGLfb/F+e7Jd/gj0vyfn//G8fheY2V
A+qa0hjn/igUVZsLtTTptEoDEVRyIE9SxaHie4a/kCEp+UeCVv/P+5YhZJPo2L+/
NjPigQaqpZ4Ue4iEF2h+EYKrmvjcTbKRtEoy7hOer5YRRnImnYRSSKXOnUwBJLxV
F/xceEt4qFSbY5+0sjOwWjZnddgFFZIpfptURoJFkIsv2ks3eAb7EcwMtnpK+kzu
rc823ZF0UCXtOr1BfGUcPVZqsYyC391KIGuxipiCgYNoONlPYKLEfP1iwTRc7Shs
PJHZW2UEJOzvOYAjVDsq1nItln/WXAGHg10Lwgczsl5N57qqz66YNl56yfa2HEso
lIZePQK+aWjX5wX/JcHAir5EN1kIoTz6a9sMCM+GgI8EcKhXqCPZGBhXW2arCJzI
TLs2NRkcDzYxOaWrIjGOX+6y15NOYknqDzpWrSqHf4srTJjxbUXf3OlbRkJS95tZ
qvFl2h6k0W5TzoKDvP81RsgftegIxKBgw/Of2FZYeK+79Cl/1clBoM7ea2gpulgr
8eGXG+mWBoPpT4O9uSMHKlquDYwKhYpKV0VecpdCbbHhkcxMqKxNfWPvqnyAWaCw
smx8QidyEKPfBoHF1N9qh8M9nGM5/ZSXAbL2EOxeu1YXJZXE+wHv5EFjsXTr41Fs
vKl5qsMcWz8yFOH/NN8+hhb7wIQ7g0Jp88GeTm6kufS8hLJY3nHAjgD/z6+IFvBQ
V5/tuGob7klOSXo3wIh5pLoxFPQM8sOU2KngKDW8GG38Xhkj6YpuvPGNIu0m7pmk
IiiX01vFQcPEaOgPg9YQbEvHhw+mIFfAVWdCkxaBslvCthfdsxDdVXIV0/jZN7wb
C+4cxCDZDobL8pwTWQhiaQKMP6f5OSBau+0x+BUEBtnluQmDf0KJsJLBPVazHWnw
e1dRrCtGC7Q0x/2bUSjLOZdVoOppTYCYgjP6Uvn9WpkIfmOy8hgWwXGU53z65Klh
/rMzKmkXcgEHG5Qzx40GdlaX25TcbQFnQFmN04lQOMe+vVcffX9EkvlHOpo/jc6+
kjicB6gTyUnk6my2ymkUIvJkQV3pVka7niK6xU1Nu9QaabCnDmqKQmTrGfOcDR/E
FO0i7BbFd62xzkbYlOybCYCbqfG/uKeWWANeuflsMxfgYGEnmlOj4b/NxbkAmz9U
2fu7wMlVujYofLwf06PrtBqppChG4GHEOpZvjcvJp/LFG+OPW16C1E/ZGqNtKNbO
K2sTVRSjM8MUDBkjwOe25pwpzNbqoouaNVmW9QtMZcVPtmIDtYkxohLrZxBIVpxw
EY6xUNppS9ftiLphb27azn53RmOTrLytJw9sKPVAsgRZx4MIXKRNS3/644HHQXxm
P8yTwXAh6VT7cMhVGIpF6eutpUOT4NfDY3ZSIQyzqrwbh4Mlsw9rnol6XQ3Qvqw0
tHVPdzNNdcso72PR9L7igT9PsSMayu9E7gvBh0BxoenEDNNDagMp0fU1judDflZk
T+XjT0Zq5Q0wxUycfPz7oRiwlhM2zy0sYvADIFlkeaKNBtDM7nqXY3IzmIspt39L
p0ZZ3lH0B9+aBTqvc7W+wJVDwCgoCZfrLbpCpdZOpsAJrLt5RqIGj9CcnVv1v6SH
RG1GTI2fI9gDJ/Yycc9qMagVVVq8WYkg4j9o5URxa3/tJKifot5/+QYpoqgKYkba
7B6we3ebGs5/Tl6Y5pTF2ssHigGTjPdpEnEekzJ5147/WqB2oWpy3WCeF/HO9uqr
9XMvo675RWgPOE6wviefJBzpaZ4ohZ7ch7CbLwYs4jZ1yuYy2HFicVjKyPnFBvaD
9qFhAo4Dbw/aIzVsEMq7NtBOTHWOm4PyLm+16SuVbMgMJSP9IadDj6cvSbNK3EjQ
AExMukb6GK6iEfIrYW1l6Gjn9E1yL83ksKlSlnJK9Oqqmy4SBEJLtQSCkUv7FdEN
ZTlDXkWrEwDwplg9+PvMJ6Y6H9I8eHfFofR8vFVKbLg+oKf+qmQOSm9QYNpLhpbx
/DfWJxHUfcKQdBFC7SBQNXdrPkl2e9vvEMcpikxLoGfQQZka8C+4Pi1tg74Pj+CN
bdAykVMMFi5Uvv3y82sRTXhp1YwxWzj+aPu5AP+cR+Vnc8oQid+gFeCMiJoXnF1m
ryxJBH98+Yqze4Ijj1ijtNg/TXGVymzlpnK2q8Ofav1UapcSbJSuPhycKv+zAJQd
quuzfVjS5UbuOc3ITTcn7R0YFfiPAKmAi32gpBCmwqWKolxEhP/W2Z8yw1Lx2QXT
YIMgHXGctJjfS896hNV6tJ7dh20cUIE1v5fDFB8qohcJD8RacnztViDdUMMYWS2z
A/+jC5FReCbYJSySzNxD4uM8mGdiuROSfI7GO3xF1KuyPRV3auCTMcQVRjbHCvVh
CN4KEGEFlLiJh+1H1yaqPiGHLJ7ly8kYc/ZFP8X5G32XENRVhkraK+oREVWi0r0l
ADYWGP3mcxmARpzlmE9h1RzxyTHwZBP6wvT21RZ8oumYc6V/CFC4da5xME6UKRpc
wbx5C9p0katmDbX0blUREfGYrP1dVBK0/21K2KflILzKGNFdcjhYo0/uj+fAMcsI
A7h6uxVGv83eJfhGB4HVaE0ByCt2i+N7Qp3L0n34X4G5dg5Sb3UOtesNGPMCGYXS
EQaNPQPq4O+coqiKVJ1OMVnd0RywuVqgKJ5jwBYc9NEUwXCOJLeKAJCztNyRJ/zf
4cAsVtJazvAN0CFpjM3oWhqY/AOlIxV670TB4KCCpkNqPVEzJmYW3fhb6xmP9n6t
XbeobC/HaQ+OWl50PJLWug7sAyTRnTw/Q0FT2J8yQMQKnmOsmWvZVnqVZC5b4XYM
opO5aV6xVa0yxQLUEX4wNDrdOaPStH+5N4zpNgxgZOEsErGgUTKPs3PU0tD2ZO1j
kvvfwAKQy0oqSbi7tPldFvqTMducOnQbYzTsWvCUwVesuwSkkUwbdFSbdhQnW0+y
1+HuYIfxNxDv6j3uor8DL8P2G46u6m20XxOkVLvcsQOYi6YtCbfecODJ7gqrq1mN
4BQiyGI8N2tiJXxTmxXdLAUN9AX8/ajVETXIEaHIzUScasxcPswEeuchbYcilUcS
urLjxM0eFEMnMYqBdqD89/13Z7avqq9z/SCbTQOmAd4YX0eG833EpbfpHH0oU3OR
PkI0DV8I6Ro022sl5XfNvrhiwBfo7uNkECSwYYqKLql6a4BpnRvk+Hk3GcBaqfYX
QtGOLQe401pcEJ7yutXTFA5dz6UbYi+XNh4yI76uqS1rh/j+61Zmqkb+nvI2je2C
I1MlCbv/4SRGRydh5cb4szBkayknx7GrPuGi5bFWjEAMvmoXZpCCmxzUli+MNaCE
xEobQK1GJ7hWKhjEPNHHG9F3OVVhFpuMQmr25ZXOCm6Oul8tR14l+c+74o5RbM/0
85ozQKVDQstUFoeK/js8sqGG4Ejv9bIXUF2RWFKs4f0ocYfsGMDRQw/+nNV85zE5
VBN89oytsACmpPtASp9a0sY4jsQ4KmI4DlxMgjc2FgRsltW+BuYOviT/y7gNjolv
sg7i4E3arOkIeOGz6Nbu0iSpGdDw+eYVPDKCWGOGVNUxueFjXmPUsI4mw5tcfT2V
ojM1rLt4Uetop9tK6e1X+rjbwn4ry7xjD0FzdDW2wQlPyo/M8B0zA4z+rCDV0cd6
aqQec4UzcQgvsWd8gYo3/ByS7au/r1kFhC9gGPCCTY2A215+DdXoj+H7COQwTlJN
EzkSxryAzwDNb2m9zPnDgmfuFvqtUeWqRlcVQjjsS5po6jHuV/D58vDrzXbgBkq+
zBbGJaISXkPvv9wTj/53TbU7AdBIN7RM5V0aQvgUyukPNvA/Bjn039XxcJsMc6Sy
ut5fLZ52U6OodHnR7nJ41zG5UuaahUYYMEX6c3PNEcOid3Zzu2LmzOaQwUNLkLD0
M0gYR/+nAYQEnOBtXvk7voAeg4p3PLxVzZktu161/drTXeJKCQcA4SkFh6Ilh/tG
9k2jyRrVTlu75QX6auU9GgmtTML1ozPC7t1u4XI2hGxdpfBO6EDR3xxbacCYRkRa
Uup+czOusS+WWiKajFc8uZekfR6fyV15OlNHBsjo5kg82u/onL/8luVfm1R3hj04
3FbMjlKi5us0kppXLC8kS+IYY6dkVm3DfGvH9A4bP/KNj6hBY5DQMeBcYRi/Ybwv
rygwT0CIWpUyv4OItnEaZRHJHOhWZ1aTiHLnkOpJ5Xmhxg3PI4X5Z2XdKvJIljFL
q8OSLwDL/ATdKKyKzxexeCX+tPQF5bO4Mpi5qSkpd0G4bNEs/0ADlPMG+K+HtECS
kTumh4E4NujmU+DkWUuYmEVK0hjMSzioqsvtWqtrWXJOCQ9ej61gk1hLni37X3wa
SVD9tKLotfoN4A21wOCr/gqNE3R3UYhm574iVZ2hgMhcAI16TNFpkzhelzxT8H2i
m4b0ogz78brTonMoDIsvYUY6yYXTNkbxqce22um3k/hSD6wwDdq+jSqbqonA5FQh
QxaU1lEQDWi+GKSC5hMXM3OJfEaIsbU37/Vbh1/fpRO8yknK0D6HVZN2SrswPfCs
cJAj/qHZYYKhECn/Y+Px5sDUroFnPNHW/ndoBVePgwNCXflF2/UX//Dogn43fit9
o1J5Pphu31mcQQZyuhE7jSMEQu0i+8JCGE+tBW+3B4VqmdOHoSbJhiZ/eUQtry5f
ZZKsqeTdUKdT5VU2ztrLNnCcGjG9S4vUZr7IIojDWFbOc5ZFuKq3q3j6Z+qitPOz
PAUo7EewTWWD6MRp0zOvQWAKpm2JsJ5h7W7r4vm5ZJmg3bFO7JDjldJ46Ucl+0q8
u6rdSx1J9Herh5OuTCXTrK5NGaPf7Oi7nuNjjXBXlqIDKjF71f7Ac1NDuPTf+P0F
mc8Pxt8DX9T8mZ+wkAfTgeZ47MP8B/9xWcr9u21ZCb/IX2wkLmg7Tsbvi5pLq/Ta
oNm1FhktM8p5BGPLxI32DKEDohL4jNMueRaIKv/YuBN6DkR7D70LB2Z9nyN+V2TF
B89P+JzJlsPIL8QqDKqhrtd2qHAHJyVHLxC39BaPfS0Rll580RHsx7zGbsNv9WbY
1NvcThoWRP/Q9s5QKprh+nCv27IgHklSg5Av9jyvJOOcoP5Ju1l5rXFu5+v95Wc1
YTDdC7nvIfYz6zOeu9/BhHcoiFVYBJ6BQJ779BfaKu81QwL+L0jhv4dI3cIZ4lTY
MwQReEWcDdJkN09SqzUpixZYqdlkoui/v178rgWCPdT0Mw3+VH/XgsMuWFikUW0I
NvpgDIOiQB/c/qFR1+3UyMTE7c8Z0g9CGI19qKn/3ddJrXR89DroH1O0DRykq6mp
wXjPQQfvbmToVqZ6V+0QWE+Ki+XIUdq/JkR9G6u4UNDbJu5S0X+mfJAhvFILFsB6
JPgHgypOsWTMIK0Q1SqSN3T1NnocEWAlrbDvVxynWwLyvU+x6eggpYoRFTCDweL+
KumXWz+PcTkfCCEMSPpwkLyWsWHOr911c9C3p2tcT5tJMSZQ8dzFyoXP+W6y0OzN
mznUM+VWnfB8SqqtqVSwNgaMu59POP1K5xnhIzIKGrhR7Xd0R85zSJZB+KQTlfyt
FJfZbqHjdMk6GrOFc0m04Rq8TUPpDino3Cr6fwkoMvNUjI1o0zD5dRnR35G+Mak9
9aWbAfcKTo5/gqDg34e4bLXc5t6Fg7lvggYMd72msAS/8up37NU9WU1ii4XjCc7m
f16NOY3tSN7yr+p81U4KW4CEwQj+NTUuzVJe+rEeQc7uLjFIRQo7aDP0bn7FsdYN
P1wsVxC+Z1pE7Lv71dzLot/04hEbPcMFrspZA6j7mLaP+rLkYUvKpUQVaPx6mjiK
oofF5O0lfWTbd3vCaIEJ+4lSCLJyIKfwpy/BgXlXB8MCxbCRfd78jsefu/PAoEp9
/OBG9OwNZ7VSxU+T/NjBZJOyN6aYSntik+ROdQB92OMiT/D+OBwTDyoiTt28YmkY
hJfHQD4MjFiKxGAvCFbuAOOiwBX3u0evi4ui9NDKjT705Ti3FRSqbzWLVYLHUoOl
/zJRUO/dDsnBPbQCg1mx2E9GLLQBID2R1KKGa1zy1YDWSw9jUUxUfBxHnWq+z8Gd
XoDGhPwAWwNoDTHjOsNhvdnm2WP2NQo6mr3q6POXyJYYvuFRnjpJ/ZmBn5URkpDr
F2xH1EXbC++8C1K9l9+vS+Wuv9GINAcifBQyZCHrCYmfbCnmwS+vpL0GBhknK0Xg
wL+sMuIDSY5+D873Aw17uusSrwffhG9+Hc/olbsiIz2/SFeFZs2Odxyq+hbFv343
e7IuDn6M/xFFgKIg5DGEMPpMzbeYcSV3GW3RGdIk65FmRv4JoPcMkLKnVNe8FsVJ
hO+6m7ZTdUe8dhtiRelos8fZ7nLal6//gaeC9ZPwr14cWsIfdXrpTcE9tsrUctwh
BpD7lBDoyDtqXFDBHCR2n0gejDjGppiXSiwQX+FWlv5p3YDOjOgUwLAoEWOJsvuP
gtq3DZs2Wj1slRn2wT5nRnK/qhpeH+gExaRfFDZNy2nw9p9dgfys00HFG9GH7pD8
zgqLK6vXvG5tSy7kUawF+ny4rjXZSurgrmmpm1s/14WonY4HmPm68TfDHKixHcvP
vXXLDgBo7LHByF9J3AUHhROVWH0ZhV4k2FAsFw0Ytq5hh6NTlEJUhrfTu+zNKiNj
kJwa9zWJsqrYcKjcSiZqjduomRsSeYk1C/V5m7exWiRfSJCV04ohs78qMW/XcrLZ
FoK3l/PY6NfNKaQiSseDTnNydR6SDDfIpWKw+xmm1rNItMyTOPhaamTTF6QPFMvC
BMecsVcpC2eIFvGPPVvx6JNwVT0RAJmURC1LbX+E9kWBDycBBDYwcAp9QQk2cPgf
yt7P0lcQqPh0HEXNTwlpgkK+qJso9DBtBVh4gpkXg52n6hEvUfOO/IbjnjnYCap7
A1FHi2tiYJPkcEi4YBG+9VE55+L0SxOOSTqqveDtVoe3FTbRbWqeLhz3X8Lp1eqL
y6/3+ltCaUMgbhZSlT06qH11+M9Cc6+dw8h9c7xgvQWQ+fO7yHVvq+DN9zR4laxb
sCMNEHhgWTb1YeO/1hM4lDkfiNgAfdwASNlyRsuxfSJJ30OsDFHyVYNYrgfXmhml
Yb04jBi3HQfOwosOxWRgQZffHTYEvqcrlbjVGAQ0jh9Ipl0tPkq7Q5I5gBKRSFvz
RcjtHsYZG8CkabIIO4wL2HC9i1c+SGHzRPjhpdGHK15VLWFMVCTvr/qqDZnaWu2k
x9tOWrEQq3b6NctkpEzaB1vOYt6GzHL7/jNAktU8UWwcWiDZHpNAjkrIEejrNu/1
mCC5CRM25sOlC7jffHLPYQTOlg3BvHQE0XEKXmxYoKYRfBvlqkwD+c5AHy9z7vnS
Ho9x6WMN93OwNw+8MqOR3Ww7Y1kMxf3tloUPKf2Y96E8IJQD080PHhKtX57RO+V3
1RerVZNto13qxwHM1xL05np3UH+eEfaDDizGYUP9OEPq7s032LWdfvZBNtkH1DIY
pydmnYvuxLyA70fKuUXaGYlI0oYctS/Q6rjcIfr5P25B9/Y/E0UNY5D7e/MjBLkW
8eOtM9X/6IJViA1poZ2sCpp0K0aFKisOJ0Gcch8I89L9qVoQwLYcP32NO/pqrJIH
fCnWdPSoOliF0fNA+8LFqid0TFOlIiWtBL+vRANlt9Mi2D1r3aELObztq4tq+2vc
VZ7bpWTW7nbOQSa3BBxWrtXwLhMqKleTnJQ3Dj1wLHjZPzAKmWDhnd2ykPcLPfw6
uz430rlpHooeIIb/Q0pA1Jmn8w2/S5pop4TgDe++uKmsd5JO3pZ5Lc9LflSlDynh
ci3ZUmeufAJZ14wH0lprrNP2vv2eGqa8xqNyKmIjzdSRQmXVtcjM9O0b9TG/Umcw
vNj6QNFYs2HMEFJpIZRTY16/+IElE82F5Vj1FO6Dp9TL3jUWHNhiKF3jopq/qvaf
xH5+8T3Lr28RDNaCCImP6VE63QVI+ft6Um8gN1Q3FfPph9BSMlX2LLO6GX/bQpSC
txqtqYKLe/rKw5C+7aX8XvEauCIUqSmrLiwNHV+1X7kNFBiy48hj5lfY/Tuys83i
eFR8ManvjGMWiFF7wvrqOhQQfUOj5zpXBsr6FahJJQGoBl92TneOpjQHu+xnHK/j
WZKAsysRMjNmupM146+VvutS5zi0Q7JyfvxEDl1rradFxlimv3XBifTijkPFk1hD
yfCSD7Jy+wDv2yKUNFoNWMi9oiAOZNM8jsaLOEmbeUIYS2xL468hvzDj2FbkryTA
NM5M1ZFvs1QxaXSghEGz4QLZaJESgZ4+AdZNUhps2O2vCdjJDshhsZ+pCggJmyQh
t4O1XeSDsdtzal2hKdkoFzRbye19f9uoxMmOcWb+L91nvFZS+Q0KlhVMW2dhNCQC
f8g4HuvhqUL9rjdFj0Q/R8DIzO00B3MjQUtaXBfqmeOwCiNz/ArDwl1/kzVRQwa5
0pO8UZ9vo0VIW5x5N4+vWaG5oNorSCETJWO7JY8kPn1odFwLWJXy8nsL892qRlE7
8qKXAr/lgy+eaqN7Ad9I/xRY0Gg9QYwvqismrK+WpieOLAhGqBqjxRrwhumk9K5A
hzO0xb+0Ojicii2iFtyo5jjdsO5UlgpN9e/CoJtyRzhXWE3GZaasPVLHW6jEkkZq
c9QOjtiA26Xz4iks1MCWIDxjnmW9WdXKCnE+Y1sAy/PVu7d/5WwmMevr9tMrjmkw
7Uts0n2OASFYK049pnCtTby5mv079OI8jEIQHQSF7fu3w5OY04PbqpEzuyUrlQVN
/ByTmJkc8pCj7Dn6A9rYAO/IsuQpkNIiWUtcAoAZJLfJ6szjUmVIbXs2XZN8h9LR
GBen/fd4pd08Ew3tJJ5I/G0yvNpm3btsW9tKS+ZJJBQe85vWoTfE6F5XO2kWlII5
DMm6KGksu3qS0ZpeuBjoS0qTdGMMbi5u7EAaf/Wa2yckD2xLrGefhvpoeEZPEyOe
T0oZ3+bTm51S2TYHFYhZCWNG/jXBzgo7wsO6ydWJ38CQzpveDCaTACNnZXCFkdV9
vHDmPl3S30fUs/mvRia2bCYQhHp6At51BoUNQxjMzHTGQH/wkelD2sj1ceRAZc4d
U9INBc3UHfgeW9WWxufT+OcgOhMOeACUpiaBNULc//KDhI2XmQKyY0MpVePGTF/l
RR4ddqswRAFUnlQfLtc/R/5zFnwDRg9YXMItOm25WJRX1z0If6dP4TWLVnhkYnyu
KsGgTUTVF13zDciXyGTq6IMZxEE+gk4ek1Rn1LQeA9bc+0XobKt1XvKTMNdoz0Fk
hFi9A7fMc6n2N+YYjFYvbEKui+y2T6G6nas8aQSqJ3lcyCxan//ILxJcRjFNwsOW
aeZTzYFqYuXH74QGq5MLaKVnt/8Yzu4w0p/eBPJ0CsbY6Xp4ZJZfBQacY3WmPgAZ
8I3dteuhRsoyrdY3WigWtDLywvI7gYfYmgsV/YeJgFc7jSicGrd/f4cJHerv3dIG
EGAZ7DKTDdg4xE9tH7JEQbAgoQ8V+FL6Zavgm8gJz66V1gGtBxS3j/y37qOTK3yd
bqowU8xALhwZzmKowFXpC9GddTmwX2yMB0TJUDZh7Ot9+vFGHWIImWrHm1VAO/47
V35OwzsQ3Un30vZ7fDSJRoNvj1k3YB38AVIriRqOSVT5cIgz5/Z/7PLkndsvQ5Aj
TMR4ZU89leQB96I78BZd0I4I8uK0XlZKXGePfezi0eYW96boRSibhdzvKL5Vs1PO
/e6GXygXrRDJof2awwKSeN+qpVnJzXxS9hlg9Do07nJXHBMaypLGbRvyb5kQHzo6
s7Su0spwg1FvWKDVIFv+oTnEFrr37rVbFU6oubShGUgSKDqy+Lnid07RjuydarmM
UEbQKQyknNVPHwB2OIzh4ECyfKUOvy43ykBYP196sGWpp4PEmZLtJH/nO/luxi8l
v07lbDtgKeEaWTo9f4wtJgciQW74I5OhGsP2TDuKv7O9olawVzoA/qXB1yhwyeH7
VrcxEhEzs49VrDrLq+dcn2wV/7mO04nbC/P4C0QPJKI1qtfSv6YLdyWNVamvbjIp
cuwcNo2CHkWk1f4XSn9ei2Q/Pn4Sn4LPoKEdBkkD92BOgttIKm4MzTv445A1PRJN
ne6aY5SRFZAXFxAiCSwwEKwiE1qaWdnm0Zd2bJN9TZLtvmcbcBKCSqHyBETDqpBX
3vlZURg3j6TZnk+BZ5SsSQhwT0sKo/mjl3g2cMjEZUj6yM3dHkExK4GY5PP7UJRP
g6Xz4qn6pYmqDUkYHUkwlfKLIEBRQUQdoaCxRFxek7Hc032JG/zKBWgMTmta0KWs
aWYHkz/YKPLDGCM+V4Ij7L3HiEsI4joUV8RJZIT6XNs5rNaL1eLYbxSYEr4aeBD1
o4Ow/G4KsEMELLwSEgTRpN6AXNcmszWYiXsLNWC3CNozVpyEC3rEHEUeT+5w7ggo
UfzB4Ks9z1SqCoe5AMVw/1SJ0b6xgPleE01EgX7fr9tOnqQdHfCxibA3L8aBoEVe
NvtyjuB2TzSBPXItYXEB9Je9TIiOFOMtbKg5jDtPsCIC8e5Vy8AlASu5q2rumcR7
ETV2tk9ALB5Tk//L33n6r2to5Ebew1O+QvZ0EB8kfP+g77T6pbm6AYdIkhCB4zC4
TYa+1rUdUuk/2bVlxTGeo5h6NOltCTimeaPfHgyqC5FVLqsr+bHIPLrnQ1RyuY5e
HscyxB1VwdAKXmAJzvjwjeZkbg7G8aJX3Gza40BYkkRcevC9vdJFWzoCssbWZO/Y
XacTfV6EqrMFWNQSTwrj6xaRyFT+AMSgZSj2pzVFMuAkMyDRxxpnTD7/aKvXc1Br
viua5fXq5Ewr3IbL/msbGBI/grS4Vzb1SCamupLGr3tc5kBENP6kk/SdhAJZGRow
ZnSrmh/gnhdSgqhTF9GgdAXv8jFuGYCTns5GqyTyb08nK3XWI+nL25wiQ3+/efro
tOMRvZQTGnsjuAl/iD9qaISYbUqyxj6wA5YHcb5rN8m9WXoJIBoaSbr3hWABPnkL
NnUHbH/mCEZUZtZCWLq2YTrpXLiigsvUVXAXbAfjpj3j1CAj6HR+e5xtPbKW20VL
EZwBdYEregfrdX97QGRBvsuGrqkAFCNaj0719uxg7cSA5YdeaZScxGjOh+FoHHWa
obA3viaW0+GcjQGFGHTnqLyxX1loGaK1i68HXfT9JBz0fh2PlnHP49Z1O2SsqXnQ
ELiUvq4LxNQoNR6GbXpIBCb0ONp2K/2dnYdLwyPsXs5U/MpkydvY/+dfgfRfVINW
OYATkBbMAU773YY/KMN6/4l/FyCu7TziZ1vJ3oJRyFvz2hhgd7TY1FzxEwSFRSxm
uxQeXzTCsoUBm9krwLKwj8HKnSRaxyVORlCm/igqa2Zm0zzw4+wi2cxZAN9LLiJc
dcell/taE0P7k9XEqlxAjziAFuryi9VSFIHkuNS2Pf3AybJ05gu8tXtWDHLk78lH
sbt6xdk2cPDuk0sVXBZgJG8xSFMrQtpKEP+hOGJ9Mi0ULcJTbTDk14mTSwfzkp47
h+SXbqQoDHsU4KwRKwGOV/jgEGWkW/lO7C9eRsrZ+V93dsMkOPxOqkKMdZ3f2YwD
iocpU8b4RbsbFvwPfij8Ih+olMv85VpsO8jqxeNAYIoZUayR9VtI0P/2SmpZrmb5
cFNKJu1Hqbu8F9NVHcTV0OBSvx2xlbzbMRIGa37yMC5GRvtbYIG5IeLvhlVL89bp
o46lxYg/Wj2KOgKcUVt6C0Vxgceccd95DMuG0aDxRJT7ODpriI7nP6uan3WBkRQe
XxeUd0auFG3veZVY1ZmfiOLYOjOKQ3fYzj3oupNMMzo6rH1VkQ00mxY0x7cc1vUe
iQgk0IN4/69pWqKdwRHbgTtf10aEbqorBN3GcwLiUmzZd+GPg2h6+UGWmzaJPge9
0R+KJRTBugzEYN/i9tJ404699TG5eLfXXobUr9C1SnuLdeIq8oSvMOfv2411wY+p
u4rATKp+DEy9ElGNlQRqkt/5nkTgsv/IIeRheoA2IT8QNObGEWVBTQqRr85zI2OI
rV2Jf0CrSBtI/Fm8rotEkzbPB59SFN55hAQ4Vww+b5PIaQu6qksAF+6f2QScCt5v
9gBCrP+YFFGH184UzJwv83hhZaJBhy4VGLCyohnlsLSgwP+MPObDB80W9uMLjFm+
WJxhpGGyna3ptovpadfss57dirM4wFO0GJqMCTJx4pU6MCkq2biGclvcuUb6UddP
Qwn1LTI5o433fq/cUnJtH4k8uY79h9MnWPbJmIPK/p3bfxHda/VWOvm2jR/BCTBx
u2q9zB0GPRyiRfV5aiY3tKaTOKKA5QVbswcG0uCDW2lxISeWpSHGwbWZo5Mp9bLj
Vp3yXekIHRII3W3O1IJKDwElO3OEvSQTRKbowFPuAxY72+lWGwspGFJUnPTFnCOt
pouELpvvVgZzcbD2539a+F0vx25P2qALtaUWOS3xOrSZ2RGUuUb5UD4KFQkH2Zy0
3aiYafiWaX2Ed20MYA5nk8HdV2feUZcxwlfpPQfGnXAaxNs7PcMNi0L67+IOw+O4
wjT3+Q1l1Zkp735vMZGA/YQyyIp2F1rYdx2m3zOGCfdhDAOjJUt1YN1IfQupUEcA
PyRRN6qqiJauI3WiQ1mj6xyGMo3c+WY+jkiB1fnOZB84iWT1k3/SEW6rwCGrQgUj
jAG6ixJlDhjRhWezmGPO3WOX2FHKYa87tsE2ZtQcyhb4q9rbA6+zpN1bRu5e8M3S
ueuNYGLqVUH2ZJnkN4hTBwiTYU/9IEHlb+RAKGSUd0aI8Hpawtv4t5KF24EtjXiv
AULw7Yl5nFF/35m9UN8sx8tPN0xQffDAK41IpGow2rDdhVRj4ScjfjHkhHgtKnDh
IO97Vx54JOkRAqP6vU7tFD0Q4Snk0eVNTeNXSrlznHi0r2uwDGckkELvZ7L49wFW
OVl7hLWoV1EFpiOqGOEilnFgUX/ZRLL/KR4ArPz2yqAjVj9VsHHmc5gicFeRwtKA
pokHlWCFtCxOrINmabj2uyVpULsQ+3vLxCkY8FFVz79q4PAZXElVgxBa+4u3ehYg
rWJQ/vnBwk0fXBDAigankV5216CVvQsAJVdjwetRNNhD2HvKVssiPtZdqYYDndY3
sm5apVOt1zlVnVpwaXAHP9ftIR0tWpTIyEzUYqOMEdJdAhWPrZLvXkN88Bno14X8
+UcEkNalRdXFafxyif0mnY6wTaZH0eWgW9CkjsJFTYxPsjJaHKSCIDKZON19q1B+
mZt+mvmTV/sgHiRkFPLOdTXFTes6OA7qJG6Wh5sRDWzOWdOzNwdQYV8rpxvpoc9L
hYF7JpkS/7OEDyfYG0a2KUWQ3+mm2snzs65f/MZl/I1Qtcwm+2HWvKv68NtzC+HE
rJ0DUFKHfyIw2DiJsQEusd+mbY+0InFjGNXvtazAIf+iv6XDx3my2Vox+nAqoj4k
AmI8w+McAhZTNP7Xtscy/Uy23UxjaDWloq3vbl97+2CT1fagX6ZeVIrxw5qb2Hm8
F5qCjpqg8jIvl6OzKCD80rZ+2IIxhbn5nJwegfCFUW80ROuQia9Mu1Pu7IQdX97f
j3Zg3vNNYWngQ5QFqn6Kg0kt/r3ANMCAk3W+R9h6Z0UBTu8apx9cJ9qtqZ7akKjE
VDdhT0efnLxc4NNiy79ax0OqM9JEFtGhYLH64IwYIaH9AjvZgqe4v+0RayqUPbDw
6b9stQmb2UNCXpAMTXTjCamcI/WO5kAh11lxM0pMS7wfx+AQhjLMR6BJnmU8kcn9
WBuTmkIPvp7jfXzZxEvV9VNdys4CL0CWXNT0MEjdblDjbrDUcf1CkDweneKL3CFi
DnulbuVShh4TbvAqU6Ua6np9p6B5e9uBEoeeCcOkL8o/OJybFi/5VYoUOiPlGDMS
9tNmlQkylj3sTWgVr+QLSlVW3hfhY2gjOPcCfRP0JCb6I/FBA7H4YAB9AxiZbnIt
Epm6qPPMOTBs75Gqhp4FELgbxG9j56aULjA6XjPHr5Qs2GGXjZttOpw7DA/tLfE6
hyHFL2XmU6gvUZ/0GCar22T9sIYgFtqvDHUkucLtflONIo7u89giNihgO4OsWphh
kYWfmoz4/aO5n0um0JNdAuIrKwOL3/sHpNAJpyc8KOOLZTDUrYfFXHnBEngKuRho
qb8how00gQIQea6DF3S5U/wyljLzCD+UlS8VZbhEvS5C0pCGoJFQyVjH4cSnYqmw
b61+qOtY/OVEtfzzEWRiCnUpYVxYvSYNoehBfW4Fk6McyAh+LHcHDK4r8x8i87m2
ZVkPaYa7hkWWU8hwkvbQnC2dfzAoeZB8zr7cvkQrFBrtv7PloltIem3Ur4GulGcV
H0x22RBGA52G5n6iO7dmpxKcUdRwsSjtkVxH8lBHsDFj0+hzykOv6OekuzkKX8DU
mtJWZnmETcO8T1iUx7B4OtHL17Plc10Gb+4dti9Q8pQew56wnfM/2xrqxDKVhJ/s
O5ZadcLKFZIhL495kzLnOdAdDNlKX4tlsbFMf9VAJfzutjiEP0Rtig9uadHXJyF1
anXipvmgGlaonEgS+L30b8+CL4GXNp70rbfMk9n1wUd4A+apLIZlDZKBFmuxcHq7
`protect END_PROTECTED
