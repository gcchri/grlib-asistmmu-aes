`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f+LvQimzSj8VREzKVPzRcBe3plS4swCP9lT5OXtNv03bfhUkaMnmCphO0iCpoonM
hOiF4Az8v3qGXrA+K9PhU2qVZddjaXvTaq23kAYuaEzQH1RHrbiGLKngczl2+5Sh
o3gH6vUoqcL6prGADExLGAL7F6HB85m11Fy6ryUINrzhYxULe7/RdY/FeoN0uUte
tCbFhstrKIDnVDvvIMTUMvstG7TBZsmABiBpmt6jCtR3W9/HOQJo2/TBjK2HShvH
siXkVRIrvexzaAXheNhAag==
`protect END_PROTECTED
