`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yQq6yP3nTW9UFyexYVcr5/jRXAA4tEgSr9qQ+kbnlql+BL6tXw1P7q/EJ33mg7lo
ncqvOnEJc3F45kU0voWv6rJhq9Tm0scnmR9izf6SzJIB7vbpzA87G2ujqONMvtwe
ltuds/gTmrhBiN5NGBhc7/u2uzhLVQ7envA0HoQwNcmEANip6fnoZd5UKIS+P0jV
Ir065H+n8AO07GAP1nvInofY/JlUc8BQ8y2yIRZtSrGrP9adtVR5CVevBWTs57Gu
GCJ1vzxYJNPoKAKQavBEGjDFNxcJxdgGQeG70WKZihZaag+B0PdQXgmscrB2v1E3
UTOxubdqC6gMhFEdf+7W183jo34lY0CPfio6r0o4Xfnc1MbuidKMTWACAKgEgNfy
dJfT8WhsSBsLLKO87lgueLo1t/4swUPv7KQsh5QPwFiFgDk8LfDPboruR8EVj9Xw
BU1Vmy5+MoB5W9NDwSPPhZn1o+bjE7eNFuJw8Lf+RoiFSKxo49SBoJRf2P5L+tDg
UwQiMT6ZcfGP+AWfWG/TUPD34lMVeaVI3DEFbcrXXXRF282CJgb7tWloZ0Pgoy+V
p32U7KfkpGdho+YWupuQMY6qVzhAKNtXS+0vYCaAgvijsOle1rh1uWtK/eERVsPK
tnFtd+xkxd8QHGasLeI0MpyfSItTF05ivt6oERRLJrXnuJmFMxeyIJifqbTV1gCd
ewkK9DJwOTemQLJwR+WEbWK5PaFROr2linXVnaxO4B7MId2NIMOfZIYJtqPPweRL
LOnr3gvcgL0N1YXEZqGpPzt7x4IghCNkeyvMaj3jMqayga9PCmQtYoFes4niLdnx
wa3lBignyTpiP7zvF+smkhAXdOktbg9TcadwpkP/z+rYMkR60wrTOo26JHD69RH4
GYAOeO/6/qnMIbErCKhIuaQBkZGrePHUY3eUcb8A11f91ckvisQ0NRWjjRAfdIRg
CFyHZYgbEXODM34UAPBhthQ+CG7IvBJTKxBztk88pfqA5hcxK8aEFJUDQZRPqA7q
AuzVgsjkwz1qvk4aqPgOrZmG50Ablidi+kPN1Q3a4RsxoJk52RQkaM0+I/ehBpm4
iLkOXg+tgLxWCNKKJVPfYA==
`protect END_PROTECTED
