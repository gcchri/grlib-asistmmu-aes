`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AJSlqvG+lRLZNmI8QAj7UbX28FhEP1/qtr5g7Z7gxp9v1WqroEjbdmcWSGtOyubp
dhxdn6tAZatSoilUFB0JBqPQTNEvwmwcHEIhKpcNtEvWT/ADwR4cy6Ukx/T80eq3
b7FpuX2A2KHbvAWEvARPpvdMXzl8gYJoQZtoYdc2KawYPU++znTDWF/IZZ2UsrJH
II2CSLXzBtNBrlFkJpgpuW5DYyE0rM6AiCwLSHRDhCvLInsZVvKGq76f8QN6oxKc
kdgIm1I4mTYIZTDres2OptWmqGdsBQrfGBRU7jnGnEQe4xHBnl0bF9eSUkpZ/994
6UJ4wXIzP+v43axvhdHMcENBaMrDMEoQw5QDC5+FmzufgBZWNl/taLvJqhumZpAb
xpb3+Wb9Nzoh3aBnb9Lx1AXphDHOQhKrHpC+j0lA6o7MfuLU8zb2VYr1h+ymX8EE
5RS6b4zOouB3faPfg0yFQc+F7Ou1UAvAB2Pd5ZEHQ+QSpMYlQhinGK6r3e8dmOYk
VSyDQ1Pd2TTehsJIBem2VXVi/NRjLMe5SEI/V7Ku/H4g7DmSp04f8LEdg6s+SF+E
IrNEPvFss8l3h/5bd+xgt6hNmrauN9wfYCPI4vyIa/2JYYHMfXxLPn2yCQFjAmOX
bckm9XZq6DIl77coE0KsjZ6NR1QklgnjUuaaul40S/Bw7hJ1MJJzJNJQvEMBmx8D
0pQC59LTl9H7FAr7Zx5jZWSOrifGVB6MDNpIzjelGsLaiqpz3lUQjYHonExeJOWY
JLNpWNjCARKbAjvy7xskGjgLY13XeetHULJTRQ3wwCNuXrVOQ6a9+nLlKGLMG1kC
zMcl8Q59qvBrl71wttk0Y4WXGuj2lpJdDH5mIIazuumMnL8v+htzZrPm2oUml+Eb
slj0lhp+dJ2spL7LawVKaxobV6/WK+JcUkIjcXXEPGEx/WZt/+3XmwewOQBGQv2Y
AGA4DpDdpEjGYaksO3Tgt9nZ211PbC4fYDecnKLTzdTcNbI4KIf4hs80PLA5VMtX
ZeK1HG6ZEJPcRngsEBGopsVJES5KigyM8adafNNmJSc=
`protect END_PROTECTED
