`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CTr4Aq643pSk2FRC9+axymMSauNTUR8rbU17GMf4w8lykV6YFiqovRsGuQX28k5x
0r99glHoacvndY+hCeGpenn7Y+u0LHYSqdvDeIMn0T6+s20O5+DiqFdbpXHrAw56
IIpZvvRZYKOyF6dgrhHDH/qcAYdgPMZfrpNncJbOblMnjQ2BG7ZRbAGkW2pC1S0y
WnKPC9Tx9GGmHgG+K3bSzY/EI/p6hY0xhL+gS4ZfF2zenlcirGBLwwqEDa3+tnTW
7cy7V46oW7CyCPjIBIGT5yqWsedHNomYn4CjlKu0M5I85OA69kDtwCeK6ucc2eXD
AmOZsr9fLTDkWWW9gOKPRg==
`protect END_PROTECTED
