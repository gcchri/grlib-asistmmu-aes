`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kW2Gb5zcqjAuvkkUJbrhkmH4vctCnjgnSsuFGeZ7K6CuvkYzQSk1Xq0vws4+qVLc
fPgpG+Gtv8ZA3sz6neFh9xABR/NpFnh1uoI8h1Kdk/rKatD8jBQq7rGOzZ09yrkW
ecEp4Bzku9M3WA7s6DtfoMHas/gy1RxkLd8rkpCj8pezm0B1aXh7WPnSDM3q1S9Y
NWXVAwRgclPdaxooSyliEj1nPzrUkTcmwaAAN2EeiErmTSIawTlma5N0Q5SA9gJ6
K00NPREbqvuu5Gon6RMa5P8buDIc5lLGKhlTtS5tLxdAahtoDrZxlUZGXOA7s5ed
nYZ4sO1rxaw8YOPpcGP7uTVX/Aoj2mUu6UKmwet7XOhP4c9bx8I5TGjS1mh+nK2G
zbLaxol76YwlkZs0qDt2Ek4hlcuBZSO+I9F7lSG+K1oxGxrAE/E8aHEx0uH5n9BX
Gedhi8B02WucsHMJtMN3lf2/mQdizKQCZCG9W1/YMRxkDL8Oio11nF9eDuT57JEu
LQ5OFdF/u1QqAYB1k2OaLOP/yMozGAsWRRQFMl+E6dSbud8S1ur/RYX7MRZMJlNf
3Zyjfj4jk20NsQ+KBByxDCSeHHUdEibdSUYatZ36seMYpWocSPlMD7TnS1qlV7WC
fbrASzp7XpnPW4SWnLoDU5F4dZR+gt1v2dcLjXRlBb73+HtNHVzFvhCZ+eXIGj/i
bdp1WgaMrGVIWSd3hOQjkMRkAYRqY1f0Vuc6zOtPt/x5W7YuOnBUAJ46u+DV+Irb
NZcp2L68rZf3PUuqxrmHcAAs9zHH/C2KclFsIN0BSkFixDRxYgAdoU6VskQdR6ys
BHCRyr8ywZQvqYuvJkOtMHasEX6OJX12ST8MP584k8QMenwSYb02w4+F+AKDtjVY
omnCFv1HUV4szZIhmu2ruAM7e6cNMEqFKUm8hj9CLAk2SGVm+xFjiv+3Qt98njgz
aYi9MBfmcfdd0fjOYk/mmFS+1059jrvIGnDnWCEQp9HtrjcmYsU7/8vixVc1vYlS
AEzxPZZDTeTyTXdJLy/uVdY+3eDBbCEoeCH38tDpDkp/GJE2s3EhK904v0W+TOfY
gR2wSuVsvsO9iGDdpDYQY7SiUk3XdyBq2vmL0OLJcj5eg46e0yrHUizaMoY6C5E8
NMgX/AWU5d8ZlZ0PbegHgEtdsrvl3GdpCx5gLu2lrKeDlGUzdsa5jZcq0gW4vrx8
S9YKBxhqrFkNawPsIst69RV5lJ9uphFHfDsQDVGegkSw1/MPg/eDEIZeGInJ+bMI
vBBPH5oW2cTEi5D/h+dFQP8HFnL+LjTM8LQQh3UpvTIVwhSL5EyG/MylXGOUdhs6
OL1n/UVQlvKfssmvWMhM17KRyoDEiepY2Cge6nSxuHQY2fEu6tlQrOZOQQ/ddtDf
4lVF2+lxOGTqSTc5M/3DeryjE0g+CihnisW9fWu4yF4uHwUFDPxJllvDPapCRbzB
ssZZnic/zr1RhdOzNKQW5YGEZRFr958VRgIJdY8K2sY3829jIr4exrLRmOrnE/s3
Y+qt6F9L/5xN7cP7ohwK15hN+DzJ/2WlmEqoNeR6PJdkTbuFxmkIFD3F4s9KEoSq
gOoumcIgjIpOQNGIc6S9mgNfBZXodH8DOgD/VhgJaMEo8oLy0iR6L7VOo2aEIqrH
JUB2PPlho3wYG1R4APz31aZQRSmlYIzhrvwKOlj6CRyPLB6vVB96H7h6gPMXmimR
N7OKymhdOWZUY09yfl8oJu1YzTjMACCBFx9r8opahT5Rz3hCdc1ofwpc4v50gpej
uQ/m4UhDq+Fs1Ye8/fLdeWcj/cUi/fL7qkdb3E/sWfkQwjqAaMCrztxsTT1Pe45T
hYnlEZVlHYeM17P2bmmEejvgD03rMORRzrmGSZ8lQSWUb0rdNC2hzzey0ynUENae
vLnC9DAfy8mqXU9CID7o/q6Yojfxw75saZNnn8NG4Ku2bAyB0RnyzTSakk86f80y
MIgPAl548mknXx+DInpOqEwp6Rs7WH/tC5K+fFjAgSHmBl+aoREjfVB0le90Sx07
7poWml6a2Vshg/uF6KJovT+JYaHXkTxFaONb3/GnhaUNIncrzPF3mxcLnwFEbOR5
CJyQevHrsGw9jR8Z+lL+x3gPBHzgoDwaQHGgEaaCm69gwAxlzLTpTrKsJIQTuYNP
hiVYbfF3k10YSztSni08ItwFy1bOGDooXVhuuRAeLsYXetWxQRaJ82n2TCMy58/N
2nkvwMyP86NuoxsUX+DxZJ+Enxeu/RFJRqSe0bJ5HOyuLveNq2jWDdPRRZjMy0Ez
2pKJ+ETmrZ4XX29cwxm+EkR0esbe8EMNgPWpE/bmOviUVALT4XwVfNMtdn+lyuE5
UeIgMLlYn7aqTXLLI6mFc5x7evGDbLsdsH1cRVb/CyvVF5+qGt3Srjcu7k13+p9b
ii/H8nXujZUVe4npGtXhSDSNT8SzNZbTN27IaDjGa7xjLrijmF/8oVwxFk41kmWK
KHVXbdS8j61BVR1+zJZaCqPp1mbdqGfx9WHPleQ54zDg1B1uTgPQW97L9krsyOdc
VlM+M7FqF+R0UwC+tJFaTsddltFWO4DqjOrgu8tzVi88G3u2kP6PM9SWMHVgXfUn
aC4RNAMHkMy3tgiFJXGLyyYF+IkZq8JxIgYUJvZhuKk/FTNYKuGlx5eDdejYuNOe
dURP1q6fBU6YRqqUEf5+oKMPRypkZk+YqagB2xw4ob5youte67guuiBkcpOZCTkH
3VYgkfLdTKzfDXCXZgRD4X/O/QNJyegJqQA82jZx+MBZssWYLUkZGYERNsZlHUkg
j1Ag+LcoFzD94YaWGm3tewnnUsLjiWU30CPFexo52OszKWcWSxBRk1P/gXKVFtVC
S2vxTB/uVKui15HcCpUa7p5/02FbBmN43z3Z7f6hwS7tE2h44l6i+rnJ22D+rxQ/
fbnmN7lpmeUcI2TkxrkkoZdbhEjpTuG08/E10KIWIMprCRAA0D6HHaiGj4XMk5lQ
UbNh/CmKyvc9LljCCuF65YUn+eV5DzAqsitWXQcLF5ewOE/k9Hqqt3S0Hj1mIW5m
GQaxU/nK9FBhwXlPjcRSBQxsYAyMJIu6qUrHpjK0HUWPJsdFWLTHDHvW8RFnZ2G9
ra7CejLsBybu9T9pfFCzRIrquIcZlR2uNNX260C+EGpMl+geZzoTzMCmUI8VqQ+S
MWZXRnm3aBJ1TO/n4r0aG222B/30XLqYx5cXV+oi9EIltIiU3a+ncwe1wU3vzK/y
I1XZyJRlPijjDYDQkc+VQYPf8xHVck5hnN/ZE8rw4e7N+CLI/Ndx/SrFwFZjJxzs
uLJmFhK48lqjmEGrUPlLnKZSO3YeJDfrlzTV9NDQ8o9udFzBtjSK2HNGypsboIeA
qXTwib0SnJxTkorNgCPY8Whr14PGuHFrvGlXepHCkjuPHx3qiFT+9StK6Y2e2m3e
lxLutig3p3jZKMg912o1V57Uurr0TNFink7vsMGa8zTAUQHoXZtfp9x9pllSYUyB
hPEVckVdNYsMzojyXOZrP6ehh5WN4dw3So6Ec4RPpujss10qwm2BIJDks6QdQ3Pa
ARgEnrmRuh673iYpGTNxD0VLBeDYjIhgH6z7fseM10S8MHBOmGNQGbwg2dOeaJMw
rwD6OjNl8X+y5Q6eDKnU9Tnmg4t4K9tcEM9v1bv5nSaXMVMlfF4TaMng3lz7CcsJ
aF81RsdJJ5z6Xaaz+fgMR3skHQ8dkoX3L0DXmA+BthMxbIbyBgw7AmF18NeCxDOS
Hm8s3iauub8VaNbZpqshRoo1NOaji5bPfqvBRmZVBQA0kl/dPn1zAqnf6rq4J4SZ
vmHrL82BlNdz4y5I7xig0DyEpqyUU9jxpp0HTXskJmZ9a6x704mC1yEpgmUhIX4S
QB91pDc0jpHsbhOanyYUqSdVwBLJgt6euDTKnlVTReTzwJG+1VFQN0Cr04zeZ24X
D80N0ZHuINFCQsnBVOlJY0MEFXxV2a9WvgIM7M5xTBP38pFN4XSQylj6aM91jciy
5X7fHCq1zExhfhkuf0zKUJY22BtMQZLS5DagQJ2tuAvFeV660f5bhQQ359jVzIl7
IrSKald556jhcKEawfay4bMFwQQmRRQpLoP7g3yxxtN2QDhz9PgDrkWt5MUSNK8t
qgRF2Qn9xt//iIHXS3XN9jY79ZFuaw2CMOqRxcNSI52atMb2A8tv25IvkzIy149Q
HuOsP6rQ4w7lFbnRLo8+Xsy3+Y7uw+XP/jO5LBcbdZEi18YggfSsnD9k7XLyBPrm
LcUovp8jJ+rIGW/oevXz9/KrHXGNRhzShPD2lLetYadukjNJA5XPolvk0uCYYatL
8Wy382+zieeMwwSFdL0pmkzr4IaKkz1L4b0jcL9m7DOkkSmorkk0B1RvsXiaiYhk
7PzxgUMYTkSqbdhzijPasb94UoEXYKIFF+0gGSKyTb7S1Q/nv1dtkJ361fYoNDKY
W68AwE7owUFLTRC0PItW7s3t416tgAFsjYiy8Fk0Jt6SzhnLpuC/6WeyJwLykHc0
lB7q983OmA9lEe2rHZ/m2Bx9gxwOs4lb/17HMD4ir2JxV8IZ4bGHkcVpRTe18zEp
sFlMeHchMBB6TVjvoBbyXlTT5wc7Ew575iVaoBaXcRHIu8JbkHaYPX7mqfFfJ5eD
NttaAjO8JcG2vJeIiDu0SLbEGtz+YNSbfYoKYMXVlraGABPe5GCH4ewV4qoiAyPC
PlLTf5Bc96pkgZdCpIgqaGT6NPId3Va8ayONZvG/9soZCWsmRYM01LAUNoErf1Xy
Utw7Kg5Ir4522jo9Z6YQrDfUcepOKu//mOwtv4HZCVp9hXDn3d9Uz5pmNAEnVjVp
iLdwZ1pNjew4euFuFFQ1t1dcUO6+Yz1zuf/dXpRoLdlx9i6QE4PaoNuEy8sfPrVZ
mEWtts0iTe+RLDtEyhIgBwZfpszYLVzPARtZJcR9RQxZqpBYkciSaaO717uorh6N
/ZI8lg35yMWeGDF+BtAY43qVPh2khc2ovpptUkJxnqe00j4OP0nquD3UZtQmFjpv
olRz0Zhetq9PVfA+BaTdxaGOn5rp81ysf5CLE4xnv57mIDK4tDgZUzb3D/IKf/K+
fQO7mOykn4UXV/Ino8F3Q5b/6tJC6it9ZKO/HfSrcrcF1SHD+1DrjtiT3RiwIRbO
AKkqMPqX1qwKnNcHhE7/OF7nMs9gUa0Ia2kBmr8S05NTA3H5XCkcV2dwTKv5eP0X
9oSKsZ6AVk430aEmlOLBUG0XPneG27VU24rdH28u5IlSbIsw0W/aw5bUwULi8NHT
VxFRODXQxs0lRIsI02ZrMT1sABQRqCBYkIdKj6Oex4SCCkiNfIIYdKOsTTb1wvKk
4c8lvZ6mhUWp8SWm0NxkKVWQEYTkAkzw3Cf1j3HMfgDzujVRtrb0B1ZW+4BtgPUh
qE8Ly5VcSU9JnsGOGVLuly4iI+e5IKRz6rGWz3BTNw8dALhn3YiDBPKWH3myRGqU
1jeOqHplfgg+JFuaI+XnvnhWTAKc7HFU4b2ocZU+Mo5rXqroRAMXVpl040dPeseP
OpV7i/GTvs9/YZ++fWJqImkonJp3IuwlvRdqW8I+hnzIFQJf73P6OpLem6E5zoil
ShMfQ2r+f+h7SFwFUHu0A5SeMOm2my0SmQpUI61abOf0bKicMPHb9sO8hMWNvJPq
srLypB82XNV/Ea7MKyBza5ktmcSzAPtvK2SAl9GT55JM84xX7BHALlvlF0qgN0wf
DedPsG3OQymwqGP2cuMC04mTdeyzWgfKDlhPT9XMvshV4ISLuVB8x7yxbU4l4P6B
7TzqXavbsN+/JCiSzGPzujXpLDQ5M2xqeaRu7Os8CoCtVSajcaI5KxnDV+nrmY04
L8UxYmWj8dvI7nzgq8vZ8bimayWzjRwIZ0gqTr2s6DvccRrrI12Um9g+wBC/ieyC
G+dFnqdeySxmO9SiD1S3KQSOjqFlAKimM521uWIR8s/AH81tClexKFMK5su7WWPH
9l6y2XQ+ThIJM59BnPsiOls86TojoR+A+3h0zPZPynT3rnr1FhDudsscJGMM3jQI
WFBaBk4CGhERPuc7liy3cTBYlIYNfJY4mIpHFnZP9uUPU8eKacl4De55bBHG6mx/
asNOhPu+IxZ2zq9FBArf4SOy5+xndJQRrpD+gYkx5v8qZ/ZPNPeYSNVyLVdpsZj7
toA+p169y3hRhc5Rq56/NrF+bzR4fz3ZiNJB0mIVwKd/t5wX3X9RMIe9+h9Spi0S
FiJkJcCwuRShzarm8+cXD3GCD6Ch1f3ynCS/yvpEc5kDyTOP9BAQOsAhHnxvFw6j
Pb3kCQMZQ015uP96z4f+ZefENXPVV38nE2zD9/hIjuIr9ciKm3tS13be3R1O8+Ln
IjJRy/vFOvF8AymkpEziykc3cMxHL2QOoSCtrcufYFgJC/R6XJoOF7da8jyZICIp
xVdFQpvtlOnaZ4zO9V18q2iOhorWJVoUgTOqX8iNMe6GkpvJ7ndQux77SSzLntJA
Uyk9O/USp9SNzVFlLPqYsbtVyBZkTUwlGAKXCUJ60nYG7Gju5IZ2J7dIkisecIwn
aHk8a9u5Dh+OfVtIzLo7Co1a+C1haK0MCWmpl2WN0crgy2QiMCS6pH40nAGTOYYX
lg6Cx+yvzmagrpT+kToTt/YmLCfr6n8qdui3BUGMfVZ/u4U8Np9aR9gmCwinY42I
DBkddo330iP7CPWI+udlLSOA9m6aXeK8w+rRLwBKPD3X09zNwyv/kiI/3TGTrMOf
wgywFLzBajFkCWYJl9cYmCTbMbj3hQQ3rp/a8h3VLNlomDnkF6e5Vhqgid8cymqk
rS5wM3uDbRPdXtYf19bKS4gGgPl27FvhjuaamoPI7UwHI0ToLajq+5xbBooXsKks
SMYSrTGzm9HcyS/I7If1lNJG/t6oEsPHILD6Tg7E6mYjrkIdc4UHdrtbQ01xnQSh
9dLwT0N/9n8L7DeUJkutDdZuD5J74Kflj8mEij4sjKgftcsj7AVswD2p+fxhCb2Y
uL4l8OGQAYuXGNypD39o2oJ4wVg0+ba7qLYltMwoZoij38bCS4204AHZXq2UAx0Z
CVy94I0YR9CILBlY+1h+N0F7i3KKJhaJUa+aC00bRI5QRstafHh784W3vxT8Lweq
0/pis1oj49BYjGReLJunk2h6Dx9DGliuhscR9lwT1ts6gerK6Yhfc9qCpihBn5GC
lxh1Y9Zjyzul7zth7sHyVxcyi3fmxk+P8qzXTXM56365vCqX0uQPqnDa7taPUxx7
xLTGy6KtUltwIlp3xE7aa0D/SUqsrcuZF4+8YPRTsy9mNpaRexRwa5Pc/vwA2bMN
GG67Cv8cfYed+Pi1yEAONCanTMNUThuq2nS6MTo1IsknxQ2uu72Kh+2CVn2EAFbP
ZS8GLsHQTcTXBbxv55EkvM7Hh2hEpwyC5CzYebv8YYzpgQysskn71OcJgZs8XIIk
YrdPHjPVVwbpHIa5jQLvmaKNfh9luJcg5eVZVxWtIswpGBRfjVoKjujotK2j1pLa
krN82Mye7lnRCG5DCYhpDwRIUmKM7qsLq3jYtlLfBkPcWA2/7rh0wQmG2GRwEf9A
imGAMwS1GtQ/yXrfol5sj1yGY+/70wA0dkDVSpGnroGpW7fnQzh0hyj7DB5LW+M+
Uv7arvJ0EThQPoDHhGL2VSbJbbfaQiVccxiiPPt9PiFVa0R0bJmR64dPeZGyejah
vPH8wxI/rMXdylhxKw6znubWrTKikSUAzjYVsrwOVq32RQ3+db2WBfUiXp3ecHN2
s6c46nNWS9KxQU/6rrI1GgHZO2ijrZXkpDsWL0HsWRQKzOG3u54qqTSsyYQ7/sRl
1tE9QW4kd/GjHaCiad9ct8IQOHqNIvIz/jNyXjTb2I59Zay0ig1mbKdPVgW7dE9w
qOOqlKiUJ6jycJy9odFwq7j3OVnB4vJLu2IFhvnp/DOO8ukSwUOcwgWmpOzwgJXL
cplifO9sv+zJXNQhWG9Ce4+g0yZLZXbI7Th9HHQNNdgrT7lQpCYg6dddM7wI8INz
bZqYZhQN9pt9pN3CpDYmNrbm0Rq/+mhsvciv/n+AXrbwQqBEQm988qlI0RMsCG9J
Np3qgIoMlJmxjTs9EF9oBGdGQenjNHZfxRN1sodgjZadWA2xYtkh1lzxBga3nZvx
PCQdJ6oFitkw4OFBQnnz7L+drOJZ7R4gfL6Eut7mFEQD5KpnZwUZ8L9w/pch4EMk
0EsuC/dWLqb9r4cJ3XLAkuNRxaI4zyNASospinVa68uexQi94Gm2EZreMMGSRyHU
G9+8bWw3n+LvrJzbxfPWQP/gHbRqwR4Qr36pkhE6/QUBvy3335rWfVQRoIatCdsO
pCeDuJbBgyLyM4XYnlbPqp9gu6ZecHnFNL17kkeDDVBSh0WmcTQG/GidK9WlFkKA
fZ8YFV77JPgo0gD8kou26nhZSCYpoqlOQn0KFnZYekIIPGsV2AXOXjvpiQ8aPRMH
q+nkBcnIGoPjO2LmiNXEhH/hn45EJhdmtsAjwsiVapoJWCmrm0GtK2Cnm3tKPefE
KwkfPV0vy9NtUadE641OzLKG/bt3JdIUdSOs9Y28ABc1K7Tyu6YGptjPzzzkD9xj
mJzY5/kX/hmt3QHiSKFzeovNNO3BjO6ZjEKQzc47NoBPrJIPV3qp9dBAxurE0n6m
FjwAH8dg2wjDJlZp9G6hvSdMF1QDbL+6aLVi1bCLLLadfdgDwwlQSgFNDnC5MBaY
wm4n89U9HvA6SZNqXneJOHTuAzSSxqOELAEoZGkoJWb7MRFKecvMrQGKBVRZpcvD
TEAfTC72ZiUnBytMt4wrJKQ/Ejq/9X6Q+Ms7O8WpghuLZY7SSsnOBglE3Vi5rDXE
0VxOVBVFDlqrXGPKj1/HlN0gc6Qz5iSF5LYJW/bjEWswXHEgUIYxSTlmGPtshEwe
zkuiOyUKIdp66emDVfkf7wSERg0+tL6M4DrTeATaNHf1quyoGSGs2bSgA7jAgdms
XTPZD3FmV/2lf2ww+sb+V7MBaG9h0sN7bigTEzWZWg3HeNuc97+btLBd8mGV2zgX
/W6ycJOlZ4kjohJNxoxgpVIqpRj8of5o3j/4gd4sPwrxOOBDrfGNwKnTOr+T8tkG
hycnr4V5dicJbWASLeYiP5IfcGCu3ndP3LBGCR3xkVp90bGKytP9h12ZbIojE6cm
aRsst9WHrCdHC4EP5VoLgllqJ1shwsraxWM+P4t6YCHDa3AfKYkb5kXU2ZPijDxw
oHJukWKz2Dtg58rHHqBYLA9horR1aNLdKu6UUGVEewUDGMAMQDgeKz2SqrPb567r
xxrx8/ntuNfXTeX5qr5EdfIMT5Cw7agz5AJmbmQcJ8cnsMVL5dPTGLtD16+L+bCF
jsgUL48DexfSBY+Jd7GAZ5SbF2DouLGkzOTtsZt1hEvVG/W4PwTjXUtA0SM5sXou
ZopcGcc9wX/ezXlQPYMv6e0USQWzqy6mXK84hO8hy/8NUVjjxkF14kIY+dyfFM8L
fnhSxZpNNluSKsow2O+/65x4elv2sdVEjv5rM2RdygIYNIZv1H2ErqeqENrnXteE
lSY5e932ZdALVwuSBCSRNakfeLILxkapeOLAoN0s28IVMAbcbw0pg50J22Smytvk
LGGKvh8AGpKrVERmR8oupgneWoKY1l++gPFKo0+zkNHkCrS9IUx2+jpre3O8XdIF
BMf2OPatDHmEwo7ca6U6hgUzun3OBr6SSbLsRu/LLAAVl4WMjH05/2Uumr90R2aS
s3LGgYN+w46vL2k9tWQevTAIExt4XvMq93nU4Pucmbf+m2E2C2ZznnDAupvLCPJM
rzNG1yIbCbue7Dh9ctnALJdvHRMrCa9aTy1B3opH2FfTKmu8oiqP50QDlWAlmoj7
0APLXhE38WbgHWEm+L1IdPKRoKWQOe9LTMzBclKEPVo3MUFLb8m4F5Z4qjVPAhJT
hHNRf2bH36epWc+hITQvdZjF4qyRE/1/I+bHoySZMlCdXBh2iTRwJsgFBa3ywhcN
FXImKCP0PjB/FbLh5yWTPW77zePk0tiqkMI/xzkva3BHVatfGkeVg95gKYSnqQVO
9YP1mUXjItqdAczg0xldxV4b7wJUjKIwcT4L7PoLolkwJOjoS+4ANj8HANOy/eXw
HG5H8pgLKLJ1jIO0ULNysHrh+3c0QElbvRTSo57Tvx6HMt57WeGwCIhNCf7rIZ+2
nsOiolQJ8NR6L8Cwu4FSSE+KKMkao5JS710pEekhq6kLMfRYvZilcmzXgsdPp5FE
rm6lnWTSukupECpMROr9gIxK9Raivx3pHP28gxeAs8tkoytDPjo4lDuGzW/Q+pqw
BlpNTRv6/5ofywt6FtAVzly2exzEK4HvsEXvQyKgz6KuzbrJoxj6ga6ruJ3Hn1N5
gaijlrvEiGRyE6dxyI9ALbLygQWo+chAlNjPC2w/okqX7QRnfPwjXb5V+x99W3az
c5bCambPYP32Vpox1jVLUZDCvjM68DlxqFkH5T+Xoi0X3LXc2lA2duFWRqsUW7Qf
qiS/dmEqEDlKgBmmviQht+SC4bLt0a7pjg8kiSw4LWdBRTl9a+Jost7w2oNIUr51
tg8tTsSdGoyR/1rqmvb3YmioFqiEjJTTW3wq752uy0TtiriPFfFvSqp8Bw99RW2R
c3fzZmxF0lxwnzs6JMXBVty0ak8yu2l4blxRp/6GDB84ttbgs6iceWyMjiVTYieM
jwvSzQLiLBG+xbXeq0fPAamWtXGweAKu5Ud1tVRLV7XcmEtItT5y0UW82+r0RoR5
2dfW8Wpnj2RqxBv0xRu1BEOcVnTjl4I6GilzNuH6XRw1ITGXWFRjSn55FUGfpAPG
`protect END_PROTECTED
