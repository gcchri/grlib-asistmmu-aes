`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9QCMdRCuceBmCjY3T2PaYfV2HmQQTW7IcTqOfLv1D1bGbubtiid2Pg0ElAsZHh+/
BsXNKLr1KAx037rnxpackWIllO0hiEmf4OOj7HbnznioZgaVDSIQ7+4t4agvgu23
i8QHlsdNylO/bdepasDeYVbfT8VUS+vnyz9HnVEgxx4yK+5QCyTo4jFPtUgqPXwL
UCIUzL7RJ1XHOy70JHXNlGYIr4UGM1LLtdU9sXG0+z/Szz76NNaTc1w7oJgW64aa
/dv5br6Lu9390ccpSebUn9Sm7amUeIdlT12vtg9ZMMGpnAwm10D1FTZSwSUOMF8O
4+1YbZLkcnxfsdskAu3CNw==
`protect END_PROTECTED
