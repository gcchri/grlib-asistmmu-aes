`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gtWKI9mXff3nc8KvDVMfPqa3lXq29iQicocUvCg27VI6h0KOLqgtSbdzjLJ+NDRb
03Xd3cs8r8qHBeMb+a1akRP64/NuMPDs9XP6EpDZdLmdXi9Lhdc4ebXdLWXM28qY
kgwsFV9zpG2hYUuM3DHUf5hNh/Jzh0M1M26mNBqtNs/wS+dbEu9S+x/7tfGfBoPB
rkV+JlEBZRyF6gZMdoFmAs7tlseaHp9zK9CdVW331KrLwVinncxSX5h3v129Ja1c
FLRKoJz+Vk8w4NMpw30dF5rP8hhdrJWnOPG47goeZr4m/Jgp3EQ8+GmN5pRpiFZx
cYHsrHou4b0IQHdyedGS0ny4LTXTsvcaIBy4tx8HN7/p1fO6FuAlVkufCiMZEO36
HqYGXEpCL/G72ZKA1zURGjfmVaK6tfQuTyDTCOQGESOV2gq45xVF4vy41VUhANHI
4Y0EkW5baTffncIBjTvf1TYr83YJgo8aVxtY9e7zoUwMLANb/VmeBkts1uJK8NUE
EsIronPVqszNtas/pCd388tgWPxTMI8w3smxaeh8w/1KGvLVnkyvHGiCz9M1XaAq
IuG6I7G5qpTGMybXWGWWX51vDTBPpmUkC6uV1lowKthTvagrx5SYLpG2jcgCyBDD
JpdvRr6Et0AAJ+6BD+/uFx87YCfrBGsMd+Sg7tnBX7RwwLsKWWc5tAbxOjv54PRb
3pG5DryZbtVihY5WwvIFeA==
`protect END_PROTECTED
