`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EkSWUW4m/lIYZDTaQTEt/aAc8HhOnmQZt/er8ObsHURn3R4j9OpsxErhoN+rZ8cT
Xuy1oPreVuAe4pWn6V3uvrFNbtzczFKsmkYwWbTBChzA8IpRouziB+U6JsSlUB86
xcTyO/rOYsKj1nQXO9SaZoA42bmFtQH1HLxEMAM2/IaNNeANnTOfR+P6uww4HcnF
D/X0hB4EhtdIKeeHaAz9EzhUYGGZ/n1Tjw01AH0Hfb9U/qWPoqWUY2A+w7tTu/Vt
FguRUhyDbNmF6MswOtpERn//iTWaGuYY9dhGnzjwBe33UrXZCs5qHNhESQeE7Mgi
BzNWltzz2AhNWbqiHzE8YGoXIQN0qgzv6ylNguX6GhPE90fFv8P96wCOHtclZUJy
GcN4SUfI/qoZ0dSUYtO2EBSPKoAyEpzbScFMISJCskI=
`protect END_PROTECTED
