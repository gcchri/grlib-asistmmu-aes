`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TZC7H3BoU59VC1YjX5Gm3Q8oRsyZFSnPwltuBuJP/w0vszkrwkcZWS23Tfgy5lJ4
W5au72bj43BN+V5ZhlR56P2xMlVZOGJebBvHT2Lt8HIhE2QMwKfEuuNidFWHZ5Ig
MnZWieXzEIFQ9apSDiK5SwILVsS9G74Ms9tgGBwQOv7MCmo+8Uql3mgeQBgkZMN3
TYb3SGutmkC9TQ1Lz9RNzr0wWe+Hmy+CL6agEpSJWLKpGsbP7OHf9AtOF8+AxNFC
lRvLbkXBaNqwNwwu3cnmfzMvsP0kNbxGBaClmGfxbuhwyLiBS2b7xwhM8Md5RnL5
ZaCGlZcCgGTtkelQfBKPqUTHKikKEZHEH/6wjcvmyEyNk3jHU7NpnyCWnU0I38oQ
PHc8OaiCGObd7zt1vMmGoQ==
`protect END_PROTECTED
