`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4msW6oaF5L8EahBQK0qZ1bvEvzeh0na/T/03p+TKoo8HN3A7q4kZBoFEyuXZOqtu
g00jGxA5NnVGAHx3C7R5Zq/S9Rx2GPbOTU7IDHb8+TJBeN4nsoKDraR8EAiX5vCG
rk+tbQcuRHySzFgl3S+dqRgAK/plMlF4WU6RMb6Uts5k6owTFWE8AfciMcW045Pl
MZe3JacbFXjLT02F+2XcmmYKR4Vfuz/EGWIjUAUQsoqNMKvbjB1rFAPvCHhk6zJy
U9pf4GjLrPtQRBCW6mNdTOSkbnh83ynV8oyO1PvkWczzJhW7RjnIeGliqI98/bVG
Y3BpiD/JlH57amhRnUrLeQ==
`protect END_PROTECTED
