`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qx0hCn2e17Gm9SCsbiP4d/0XFqV+fgR/AaXlHzcWHP/WAbaG+m9zU6cy4m5sCc7O
dyVdMlC9iNPJ7TiQ5OZZeMMfVD7ArkxDtUMc2nfAVS/32x8jjaqptX7HDKIVGZ7E
6W7XoecWXys0KIc9gE20gbRHjxJJdG1fOdc8XEQHmdz3lbiIDcCML2rD7ZyfIHHx
typ/hzAdRZa3z1qnONjTqL6vwGjW2u1UTAfAiGIqC5i/qutpDcXB/71zJojb/7jA
psCCT8BxBxQgJiSfvlBAFw==
`protect END_PROTECTED
