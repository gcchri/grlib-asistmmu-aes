`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hU+m7CihEO0E2ArsXjTt6PwD/3n5PC/PozM9DYilCdiAhwecFSYpcdxmEFn6TGpZ
GDFmWWcLVMKLX/yGMkvHa/51Mr1iYvyyFgFaT4TZagAqEORRuQZ8lR9B3TElBfL/
kQgXBzljC/eOtSy2YpcyEq+1VVSFVmO9BIzWEA0CrfOnDh+HOYOCd9qX9wLrE9nA
Oc3Ke69R1fDZtBr8ctR0TH0UxRH0UAOdrh4MzQXs/iLo34VQ8quIQXsWjXP9kqeJ
aJ7feKK8qhW2vcpdBBWCSMlE9ylD3x+EkNXd+/d9EfjGxZzGDYQcZX7BZo8VonMw
aedHeQ3h/2sqF6PZi3TKZ6GJfHu0cNkWQfOC9HqeL+2sxOSsvjFCBb+NhW/xSNfY
lyob2Kb4X80Ne4e7OTjDI7b8MsFGAeTFs+49ezX5Fp9IUGEgu7oSCsqCsucXCZNV
g3BOxBevhAVxLjEhDe066w8rolv4WeGLP+62V9Kq9JGHs5zl83GxupOkyA/niR2N
ah/nl93ZzKilLDwtYgS7AqQuD79phNkzkXiwh3gR7s43MisxXqG2dVh+4VuIbI0o
TqL9UB/Nirf4Ze7xU0zy7do2xzd7FJL0yPcO8PrqiVhctAkEzgjE3YqnJnmWttiS
AZsSfU7dXgsnorGtIKXhCGy3cDznVPhH9Pam22pYflNFk0/TjZs8Vcgu/HOhDSJ5
/BNG+AMT/PhQ5F5jpbPed5rGRxqe8Cj6oFzoBQmgjVyS/ZGnUZoUjr0cwWAzR3dd
PkuK3OMZSfE8AqCUWocb6WAfXFQbVGtSIUM1rvLhaEjx9REKKZ+iZ4KVnIM2hX0k
neBMg8vAeXQBAYizje5rkZLHzy4+KXX6Fp/sxhMaSjoNsFtRwwJN2qUujYwGhwnU
MlTqUOuhRSINEEjGIzXLg159w4E382wS52bAv3+qP/T+AT+FiW72cWSEpfiTt8Qv
SZC0esRTpqMkA6eTblmTqXLLX68ndWwA6wX2CLeRXTWBZpdfc82Y7uiWmYu2MLwq
iU6B3eMh/BceXvuiDI2KiOHry2QZdosWgFJ04merixV3Zo+L3ngnuPhTlH1hpIMr
1zKM49l+OjcygzvAiF9T7JFp9UMDUZi1lF3HLo1Nj8QEq96qV0NoBmpAS0ooPv30
kJGvBWQpuYugZYfIw/kf9afRcM9LeG62AYSDVY+gwupJdjXz6K2eeRLuVBKY6NEC
6aYoudLoqsNsVjH4jz8VnzRz9Npo1/qyVZbpKuxOtRphwQVMwpKKGJ1fxUy1Zf/u
jbLoKmEjQLad8/ivgkSSeJg53pFWnu/XxkqGfHPQlYd8KoEL0t9oadcxJP5LjLYV
rRlw1/byOQB7Bcp1EyPGEuVbgoAoAMneUrctdo5W0JLl/cIVcBEtxVPfILAl6eWZ
U1emddpowsdM11K9PolMMUdiZgNxcWpmjWj2UjUxKVyj07Ac/N1jHm3gPfnotf95
l0+ntX5PU6HtLbzz0JirjKrU71PzTDL68lgX4sT1YI8+o0YbFLOeYxYMEZIs5CI+
tnv77Mxp47sCl4YOnI02SnBJhc4fu+eL6vgR7IIal2SOKoo8g70UcxeVSqoCQs6u
/z8QqELWkqm0sQJN36fmrbsZR8amTnjzCktcQTxSmwahNq7S3FjX6GXDiMjkxPtZ
FLHC7QmPPuC/NECG4nmCB/SjR+LsySVYQjOMbCeQFZSnkOZeoQuwIv3bCx9wtSZ5
lTTIDl07G0WIAPrNfN5nP7IMFfzhGpfeqTdZ47LL1kaQF5GA/P/RfM3kgGtlMSbO
YWs4wr/xdvOpSYLBgIda+zi+DdXGqiuiMboXDkjw6nprW5ZDxsrzhPUwh1F//XrH
`protect END_PROTECTED
