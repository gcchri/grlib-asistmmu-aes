`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xxzWljU8yCONkALN67OzGqUIBbNjDQ6reibTuuhrW5LCbvb6Xkggb4l2CKvYxU0/
CPYz/csHcvp22oViDBZYiDljbXQgNs0unfLYVb4pcEvyepRp7MI6UEme6Y3LUsca
cSzRdXCEAG9exaB3K2yVXHzKDuavBnHWQzfde5h2vTdkukjoqsT/5xzRAykIZpJ6
EYte90BrUxbFxQMQl+2BMZjPeuT+am/hF+3OjDB8mRaI5lrvCBA55c1wfV5JuFiJ
lmUmGOFIMQW8vlFDmfEnhdlkCkwEUxuSz/29iInhc+IvQkmeKiXAWXohbqkwc9Yn
Xs/0Leu5Zgr4ADMVJp89mVpM7v5WJBaOI7Ru0itpSmIvkvtiGPnLU4j1rKpPLbwd
qhYWlKK5Yi5FDbxdPKGabJLPktHry/5l+2Q900BCUNAZeWL24tWPDkXe4rLTXD9+
GEnicS5AGtA5Qjd3tFGmTsGOXGe1Ai+VC79R5IyP++cWZV5mFhyFax39qRZyyz1F
`protect END_PROTECTED
