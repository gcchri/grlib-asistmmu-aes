`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XY8/6OJMNVWd3PCnBmWJgYOxoipeNsaru/WpYh1i+53WN9fwlQSbAN6mBDo9dtRB
u09vSV+kVTQoEkcHiwNMqA87gzNlhzhO3HbxZk7NBoga5OtLWDyfxLbOrKkv1sgo
Cy7sgXlYft9k1jGF8fcHslnmBKDRb4vPk4Xm4r1IEtjmS+3EnxOwK/RVvPUbqj7y
t1Z9Juf1SlqwEcHMwJDlWudfINiOfo50Icip7xlYNQ1HmvC7D4ieZK6dx+vUpLBy
PfO2uIFvp1W4kXmX3lQ2SJHX4VS2+faDoa4zkcffUIqTVbUQ7eOdyQ1n1FrtxY5H
5nNl5/EK1L9VT5U6OaVZxSgVDxgG0sQZ+/o5NzPwK84=
`protect END_PROTECTED
