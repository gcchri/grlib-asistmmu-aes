`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h9DQ5snnfugEGE545Cg31UOk/RfEHKEE6V/EQptAREpi6g/2jNiGtTH3h4s643xM
OVphLi0wQj9P0MO2R5EclakgJENm5CQXnrW7e4aw46I7WvTGCcW+qdH78eKMpt9G
eyPO9PqbnB4VTjwz0uwCm00hb5kIysi93qgmTYtFuMlgkBoEXTqkIzXiE26hDFnL
2Wjo2Vy8zxzaEEB+27aV4BFaFaLvvn4e0HC1Fyc5CdpABmRba1iMqwLysHxR7HJb
iH3W/KjWPB2t2V3UX1+59WI70+BMP8TbXE4KeSnk0LA=
`protect END_PROTECTED
