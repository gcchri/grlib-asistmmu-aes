`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VeG5QSDOauUmKwPdTKf01njZbc+hiP3EYpMlxHxzxlyR/cdehSNOzOzp7jbBTHzu
0N+O7u/gqnJnMrjgI9l5X2aucSinSNXBqCqNxVnTl4rYP+S9pMjl/dpgEOWikrky
p3eyPLCiJx9XVvfkcRO+0HBd9W5ZSWTqKYgW9tiaXLIYPeMfYfZbdo+HqZhioAvA
icAY+lFspLNpoIdj1ThQ8DWFrJVVJMVwBvToHxi92AWJpWXutc/j142+hwZ243H7
Cf1/uGlTkYFGneBUHsSlanV0j/7K34fgpkRDKjEOMHDvuQunpbQwHGFUM8iehlyJ
SMTo8qW2eQo5oXdF1pR0LocCHRtYaDzkuNonC5MFjfTaQqKSGye550T1VltbQ97Q
JM90hzam6ZPAyQkIcmKs3hrF58RRwoICvbAhOPUSArM=
`protect END_PROTECTED
