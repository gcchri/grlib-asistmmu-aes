`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XH3TUFEyIY34skhOBwuCofIW7BKUlTlD7Agb6t4IkNq6q+gSLkiMyoUn+LXAZ08+
DAJTuW9sHUrQXmURb7S4SJ8ed0lhmnPpujdup4sa0/UstFKEpuKhjixZ7pYfMFs/
R5xawratTxZHjY5agNMwBwHDAY0b6GKtJfkHwtfIYSzNPRQDImFlUpkMg8A/gsYj
njAJAA78wqimvfcE8EdNLQ2Ze+L/hTyqbyuyrzMKbcfQk4qc4RDVyOWkDBJqBvbx
g7+dtMhicYBKeilIIB4MIA==
`protect END_PROTECTED
