`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
deU8MwJNFeV6OxN+J4DOeL0ccABj9BpQcZII22wvsEDD7rGo7U3zCmGEjAqqIrRf
CV+F5rffbNwt/OwUwYz6cMX+5lyEmceF9Fvbv3keVV17zo8GhHoaU1HVkl69ZJRO
ILlGdxd0ZdkcG77MkqVtaP1ihvq2fJKNI/smrMR3XDr7Cxz2pCXpO70pPl/rlW/i
Ke0nU1FIqGRDVD7TAMl7fE+Tqy71Zl0It5cYO9i7MkSBHQdSccK7tbVE/NGL20st
jHgX5bKVwH0OFuW10GHyrvCfeukn9yQzSPVdSrv2INA/9k4f7vDIekFY0VQeUBuN
bsEKCDrjgsxYprEtbxpl5AFBLHxxiNNh434N2bbqVRDAVO2jt1F8a3Uhs099oBOY
AyviTiKOUJtIDoG+2ShKPA==
`protect END_PROTECTED
