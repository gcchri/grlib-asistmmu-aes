`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dB1XufEPzIrL+k25Ebw5mgIb8NRe1qv48gJ1Ali+6o7UNJmQ3moHQ6dlrTDDsmwe
7UZvMlr7kmki4l56e0M4sXS5nSt6gTXf+vnsHQrJpSSplpDWp08syagSIjDQDEfi
M4ClEOzE/+i83oOQmRUFPIn4eCJbXUHBYViJjbdRn3J6ArqKmuR3j0XKHJHT9W5a
Lq7rGmI+QS9i6oXBmz0HxKnZ03xGF2KAKgQfWGGK9K4DfxShX+Yvvp+uYeGcLu1X
Vop5KiMvV8ehQVOXIacBJhiZiDO9FODRtvgSTnSYz5xqL/jBPKODL7JDsAQBjg0U
EEvFElJqo/Lb6dsoVOVzHfWwBOa+C3TCqPt/ZulbySPjbnX7JixnsEqyS17n1ICu
HVw8bvS2evFTd8vgmaIui7pHtU7wQSs0nZX4ZCTKn6VsLi6KquKHgiKgpuBYP91x
nuEWG7Mp2nit5Pt/h1U77us1Ds7TcDA5mFY4tJx9C71fzBzSSSz4MYiYeDvEUBD4
+07T1C5PCMdDr4P6NvTe2KmAxiasEHc2+QXcMoAgnRxQBLodeWor0rM04+sBZrve
hz8Bw648++9IitByb0MvPoovojITqxQ5JNap63cY9MRrUTiX081+ke09xpWQxkti
2P+zikecD92iOeeEhEkIqq3Ne67+QLC5faW2/gCgvKf+9yjQh1TS9RjAuPp6St/v
Og6Ul2e9qeW8VWer0yrU7hN6wy6l0E4Y9CK7Ydxwiz4GS66vIjV+je0zEAKrdb6C
8kLszfyKaRluOqJNXmbqIGIfErKtGvolvis8iOhtQHfqCCIXalTbM3VY5Rmyoy5F
jZiUHRovr96oNyH5SH5GBgI1vtmp79AGFzdi6miDQWGHvIya1ID6hlMaHl22VcbG
1So2ilac4yK46k88LZj0bxh470p1pgXX4wP9gutf1LNMGw4Qf4qlUt1rVOBJ6ZlM
WPmHxNsOF1jRMLICymE9V7UawrtsMiCZKnx3iJ4USb9INtiO4RpyOur/dCgm2d/X
nDMs0P0u+3AvIuslYQSlfNCjw+Juit4XirFzeEWLc43cK76faaxnpERWXU90D1Wj
PcUM9Z1rk/wrTt12aEf9rNbsY8Gmkk2dCobD5aKDRIMXehqkJgQWkokkPt3leP1b
x0pJs0QSHaF+t5mrtX0xDmTLOKsd0a8qZu8rhMk1ZiF0A8Y5n753O750Ke6yzlCn
0lx73C32az2DVyAPhg15x2yPME4ssvzKzQSDNbB7jTbectOYO193qJ6pgV4nb9Ob
`protect END_PROTECTED
