`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RTkCQK09Jn62cX2+uBBsyUeYO4uz/sJdbxNbTrkiuEHOTJa390MG7tpbOS418y4z
OtQGrMdiJEaeStsIPjicwok4KTOfNrhZSDNrr4sO2q8KsONZ/ZRbAuFvhCGo/fIS
EY4IHFdrG/WGorXk7nqt9+G6MY4erbsCepRTly+IwBZDQN/0w0Be1a1fUq/FB6AF
Apw1S2en6rRYWE66M/rI8A0mY5suLm1ubukzZBrjcZtd/BX4tw3H8KU40NMxwnki
kyJ2tZ4ghSo+1dvm11y5rl1VL4eWurGPTDQx+7V18HtmBDBH9XNrK73jvKAMV+5d
vMIagCA4H2EwcvTVi/pEQfFHofv89hN+4+B9CGWa+SRO7M+IMGASoXC4zsLivEKD
hpkpA9fCZ4MedK9e3NQeuTL+/YUPHIJMvFTaZ6J7fwg=
`protect END_PROTECTED
