`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gCPvlogGAqpNHTEEXTQFWai2rr6D60fBXweauwkp/ZAIKCJLeupq2hpQ38K8DClp
yzuqeIxWRazsOzWSspG3Ui87pRAjvy+ds4kI4NZD549VrZ4fM3VZJ9IVBPtYJLn2
JkTBORV5XbZKWJ8R3H7vnZG99hMuiXEhbwj8Dza00kcJS7qUkZT79l556Uf7VYma
CL22W1Yab9vl/nrSOHUVAc5QE9AC3mbfcbrQShAOx+PKeojh7Jbs6UYFnpcs91Kg
wuxUk5BPULO1H6Y4zeXh2vUZlOEgfhUgkF572njs89cKlMe4r/5vxVqQ5SgOsd9d
N0zgYTiWHPANKT/ofHs08Vk/uROxiKjWcatdZ/XDwWmh80FeYchxZCnof3CbyZ/V
MUKDUGPEPuEICJFEaDu7wHmTzLbb+oA6aDdC1wZOgXU8oOFlOLooNJTFqV5lUl9l
I2xm2FRjgdGudhVDbTf++mon6Jqy2ltV/sAVYkWuIpnzy0ga9jQWDoZxM/AUPSMf
`protect END_PROTECTED
