`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VcEAm5ZREL2MWXitk0FrGf4iRMCw7XIptrFYHum1wvMn5aljuOTalSTjZTx4VXId
tCYkhiGa5mSviyjw/GpFpjtyERjryajPOyn8H8+K1ZpUhTdZcCYhk+LwDLll/lY2
lu4TbZKU7wvqblr0fRlujo/oHdMoTpL3kY+x+Wl4eKKlbiYUaHkRuBaWOraAMPxD
4/Wx4r6jK+pRUhOsPIm2PwgzjvH1xPibSUdsXhz3DIPOk51VaHtn/GhCgtih6e6F
`protect END_PROTECTED
