`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TLweNJhN91EPtlcTAuvYFwVfRQwkoEsQKJr0PDfI0m1hopz8OO1Anwu1lhBdeP97
bA9McX3L21eVphig6CDXP/68KLR7BHVDIehOEm6UjNkXKTLCFqHd1VFFHNTqIsjq
uAvum9pGFGYL51rAyasjHBln1MMxno7mx6NUA3pjQixOEK567O8CJrnc3nTs5BRp
Th3ZUS++fFvmJBs1VkQNSuOa1G76jkEzTCYSz+Ph9K8TbmfFxPb5N0FEsvdM1nHB
k9mCM0r7xmPdgWYQ2DaXX7QyDiHMtNhenZnve08cPvo9DCpGTmArwg24LmYVUjPO
kgETTp243kCidkxOHTuBHImsCh1UcZ/Knm/KOJ9O6i0nnY9o4UYLfZRmUtDJqfz/
OrH2s7QRnjWYuV/RYf7qyqit9Th4W93uSTBR0NCl9hDyq2vOeO1zvoDWIH9vFGyi
nOqUWtMWMDlXnUf+5fogXjygkxRXSF6N/eS6IEFOfABpENLVv6Ilub3EhAhbNaOm
aUz0TuqaEhzeY9BNEVcHL/ByhPZvxa8u4Drr3zhjDerujZVrRpDF+gYZn4zskviH
xO/q8c/HPQqDOH5qVekTHp31yMmdT27d7D0giARAoiHJbLzUQqq5KJGGUfoEmlMh
mzQH1g++snMW5S4pDioLYO5KE0m94/LOIDci9J//gI/o8rBpj74dtFOOzLU8uRxL
k1X0+FfsRR8KfxfAYGXtIjc3gs9KGviheeDflwE2Klc=
`protect END_PROTECTED
