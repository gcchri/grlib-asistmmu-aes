`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SkYFwWHgsoP2mqWhJcn1+BAM/A8nkUaE3kR+79YxdV51/3tZ6YMiezoGkDUB/+C1
WaZ+TE6/UJ1LjrQ+MnafzQYkONgTFOhq1Uq6azbqFt7pt6W7CVDXkgWQPGimsvjW
uP/9yaLoPvNdRiYDWX+pvuWTEXyE+tFHTgJViQ2z/wMcXUzcM9zkEGRTiKv//5Ib
5iX3TfOE8cJlP0dNnkQ/b6tK4mDOCfz4fmnCgZU/0AVT0/onbY7fNS36YQFuSowx
ogUewxSbfg/q7rggCdvUUQRrLwkTM67tnQt1gSKNS8hmJoY17iSNzt3oZSe+zlIt
x13TMRko2vNat0OiFyb35AxFR+oPWJ8BtROXeaja+log8lpHWBmRcJ4iKINeoL3o
q7TqUuGkUG3v0ogMEYrgfg8ov9x5m+sZDn2vaCrbBNUx2f1Ym3Z/dIzRPYlPV1ct
2Y/o37o5oyBnATLgbb8ZVMWrFe84BCc7ytdN/U9WMKDVeLSIPy/956R/Hfbsekcz
BburENNF52geN/LblkqsmhxN3gBoMuGJ0J1etSR7f8TdLEYIB7NRFpIiSLUcIBNO
pKjPQp+FKfba81f1fgOlDmJ7X4NNrgGbHM5T52L12BLztJUGGClYWXirbXVtlsSe
lI7WvNe6SVblbb2J2tKSpPsi7/ndHq3Xd2Zqebb/9iJHHUv/5DVo/E5yeU1eGAFW
F5lmTx2MdoOMjYKkXIuxnHbjIKQklTT7t0y/1UO1X0EH5lk6Gd7UmCMs9c6gVrZK
zZesejd8zrgRFLshEXxV9XXCMXAgpbK5tOW7xsQuHyhK9mU8rTImNRQDJaz93uJ/
o4v+vfclGDBgALGaTlz/8Y14t1kBVHOIbMIAQk+EEjBcn4P1W1TwsFW53RltlK6t
+yZ4TCutQOUQMwrqXLVl2n6GG7GrlnXc8aInRq45P5HGZ4dqpfsPxsW8ELyf81mc
ieOihWGBy2WHErI13/oHUQPtSjkwtSARlBVSnGaN8uMFha+K4fwSOKE3c100Z7cU
bJbWpXnAjG6xgruVF8iWCYjxHE2IrWF88C8XFCEGbHcXK9RzT3calb3/WOooGjQL
KUuSxfg576IXoHOJSNqh3x8VxH8DV/fYA/fiziOxNZcLkvhNeOyTKQwED0XIRDVw
CC1xKhchDnHAXMJQPzO2IIjCNwJC05Wr77UBWQRwX9QdmcKhCnHUrHjukrLPKb+3
Wg9QF3DloNdSeMpYZxsy1PGI8e0Xhpl/zam6qGXH5Zh/Fp9H/HIbltoRv9z+VFT7
oxLlM8346Q8H5VrHes33lodK/iSkNL81aekPGWEoYFLArhceL2H+OEb87NlGzvKw
9A/6p9KcwCJQznCfn0xtD8Hrk6mZttLecKUpIF6JaKFEhDFJj+gWReNMqrnGZa4+
ihok0F01ytZzjTjLrkaQhM2TrR44TOToYBkQvCavdCgNixPo7WszTWliCuA6+hlQ
aIYoj+jFfU38IPMb6Soe03VoK7Gvv64TnHMzB50Gr3mESE0kjXRAz+T8Msy113l4
kxMuOjkonafqIIWmP+DquSpNBRYSKZn69xEy2WsRwiLokY6/GBUcG1UNklYn/ZSx
DI5OTYsp74S4urdav3YR44kZHhRdiV6MzJAuGruj2c4JSENb4MXUtCWa1MF2Chhc
kljFYZRmdNGS6mEvElosKrDmELqaP9o2T6zzGqY9AoyxkEvAenk/iW9jzfSRRH0s
+IJuYcyOcRthrSStGrciAQ80NTstkPLNTWIhHufLefOW03lcAnFfwzyIvztSpXYm
f7Bp9eVKZ33KgOA+YlFZHQkbpDOCrJc8Chh+V+tKJ8VSUynyifvd3/VRYNqSULGS
ss0PO5SMu/P6pFGN/fnkmYVbDWaswqh+5anHjJfDU2t5rs6GMjlcSPK73atgmiCP
ETXJo8wDfNGk0jssbZ9y5IXV4/gWMPd7McPdYswzfItXv+lXVs+ZTK/FwW4NcQ0J
bpjehjqPcanRcVmUPXDzcQqRWULeIAwZIKq3wiQAG8NNI9WqM0Q0RHQo7ePEYcmC
vIyJ4NFJGT/5vU0K0iEdZkxh7lh9pe1wxj6wUwVyQwXIaxUySoyIPu0/AklVCMAQ
LEkH0I2xF3jSeukA/4WGAXfnpDntFA1A12EJ2QUfwDGAdTeqLsvTZB2u1msO6uOi
6sJk+0jy5WZVvdR6UtUC4KlvSd/YbVNvPqO7OAM5lMUzO3r3EK9GBOIXyxsXQgAz
GExgcYnI1qkTB+7TjEYIQQHzM4k0JwQskgmUUzTyfHaN03JBq4Q0Psq0M4oQwmeM
08snSLTo+Bk2urThKb6hI/LvZaJSxE1TcyNCVIZZUN6qJPy1jDqqps1rDzkaaLE0
IU9wXDNPyn01ge06tUjumhaHDaJpgxz+aOzkh2bYDIOJ6alqsPrN252u/ZtAYev9
B7CDGLVK9SdbW67PaFZGFMeaY5LL/ZwfhFuNMSuoC1Sgnnib1+FXALAjqGnKbyu0
ezU4fijfNVh61rsQn/FQScqryqcxvvhsH51evoxJDvxzxA60nTYwK6ZJGzcgwupC
8hHEcozo6qAg3wMNL6KG2PlCh6lvBARnTjwW6eGQPNfdrLiBmS1RrQr0QAmo3p5O
s9otG9mBq8FYLmWWx8zjr+cyZ/NGQgXuimczQOxoufbaEc+6y6FoF475xkC+IZbL
OrkbNEozxSH/dqVEIugdfRdsXWECC1YRipqpyXjZv/W8ILNaxN4mAYi/zPi2FLt1
Wbb66MiEWyzrth8G3TPBdEBQc2X8I//yyy2eANNaBLQcHx754IFcGy4a4u/ztIC0
T52pcli3/uBWvWKYBeLjTHI6G/q4whLgyIXuAWiXTrsEUltV2vyBrqaaU+6zWpls
mCdbIbo7IiYl3HHAAG2U/Tp1HWTOeuCu3nwjgnp8ZGWRHq/rVGmiWXITOmIEthuE
MEU9VBR36jhMTG12YTe8bInG1gYfM3IjP/aHAiSVYacXOdSJg3jTIylXtVlUbH6x
z9xWq8nGws5sFd8PLgJlgVRaZ4wPSXaMKxOkQsyT0vQ7BweCOIqX79D53HNlUqcg
VcL9GSijF4XDurmfFFsSVLFoI1ZUkfy/ZU+BFw7IgmZXgJt9xzbiji9bkI32VEz+
F5uB+ZGwi647AGY1C2Xpzd3WMixqb6l/6N71eS2QbcWIb7JnX17SIUtlBuO3Q9rq
U7gbkczz3IGdL/0sd3jp8HtYzThCOnRxK6+F2evjON5NNUw71W8bWVj1/byBRVsN
DOLKFMaZI74gGg6GTRzIFFpqsi2hmDXBLcpt7Q0N3Ea8deJp0YDjeidNFUkzWFCw
hm5VG7rp0HqN63cx+PnVBM1/Rje6n0uCoyCS+sLxwbp1GU0k3ACcfpy+kd+TGdaR
c7SyL2CfRE/Lb2EC5qnARQYTfkIfy7gPuXeL0QyNRJ6YpF5zV1iqwiiRwoVaVUY7
TqS1SUX9e9qEDeF/0Q1Rh8Lcf2R/67Ug3R+PUiZDdFwfhWB7KiqlxrcZs8LvhebE
a/R7hOKAAciSspoEfJuJ01crCIdQoPOse62PVK4PP41LEiJDNBnaWUfcOvxlLO1i
2Sv86eEZRxISi1V7tr10cvOW2HWm6x14ciU1GgkO3T3xgSfxoRuCqWV9QU+3/qo6
wf5zg8SFnSbIaMxPCp8JhR1rRfHzv+F1X5lSm9yo0H8oLgzjV6YGG2RTIz7BNaM5
QlQKOEGs67xVbDwkxgmHlMHB4rwXqOO5FwTnZ8CLsXqz4Ii5PNDCCvbdTxFsNAAL
Bq3+6R+vxYZR4rNkrzvC293p+oN8CvybvnbJnNmNh3Hky7hrAvoRi2/IpuHicoAu
D5MXEZb/Mek0DPUv3/GlyxDdDmKMbzsxcfKboRhGJyEVCCaIuxFZzqUYiU9UXAW2
vfTYXIN5vvOl8w9CYH98uXmZ0eYV/F3DUUCNawq6qQOHTQdyXotrXSRKbyEasyje
kKMpfsUklelbvmYBSidWXkqbmciMmhh2mLNP1LZqcxV0c9uJKdfUKMI2ogV98/Zj
oanAGL82Ec0BrVKyX/0/EhGukDu+61PEGwfYpteBiR3VYX3ICFaWIyRB6Dxj8EvD
IyqEIUvfjlTOuk+p90uvLJ5zW85a/GzY0ZV9otW4hLZQmjE1zAXbnlhXofRhKBqD
tvVL4zFAfjTUSs+2tITE7Ifew0DjHGC7/kve1tVe448Vp2//XLdvX78J/cgoKPky
/ffZ8BwRtXrTtz92rtFNu3dNM4osKF3e0UP16X9Xum/mAWXo1cBE0vIKy32dlzKA
E3bTcJmhYLLI54bydgasIzqkoY2FLX9fsRPjdZa+JAEK3EEy0hpWJUY1Kl1DE8fc
DpEGkW35GM/MBwmAk73XSHdXGZo/No6k7ThH3I1h+ZA0U5vShmL491fvc4t3WbKD
MGT3BgVXlOyO9lBD2KUL93Y7ZAMPcWJEoVpKl35urU43GHh40jyheq0arI/G7IiJ
bLsQnBicWSJnD2S4kUcIwkiq0mspOmddWwmKtM/Apk3TL5EKAlB8ogTCBJrGEq52
7VC91bRzJH61lGXfyVEFatnWVeEQyg1//y7hoIq1Ny06bLBWBeryOoegDd/48W3/
ONrOXSAGtiGv975kakx370Wt5+YkSSEH1y0lf35CFl+lPIOnUeTvnhtTQWepJTZW
NdWnv454wH2yp0ACXnbZ/9N7hmXW7L7XFDSsvQfAo028Gf15Do/R65wOcmw/GyTP
96y/88k0hEoxBXulu5LtCDobob9vwo0TpNyin1uXX/rh7tvBDJQml3ZGwNBL7Ecs
/NiqE9lIZ/SiZrzEMP2FYG1Ku8yuJr1vgiuQq9a7SsKMHWRVPX/c4dgOVy1XFM+P
SKYWbvAYY8/Yt8VojSsG3rJWDtV6RK64KUh/cjP384UHaPICQYdx7SwtFaBo+KBG
rX8lwA5T+7wVJSJEgID1bivqatZUK7VNr+KoZNGJd5bo+CLkxsiAVknqeGItyhAR
o0aWaKJ6ubtNh4/doAN+8tui8T/TrEEPHEnT2v+zEkdoKzMYqeNrCasQdfX41HSH
uC5q5KmUJhd4LaQMhU3rdhNc5t0C2X1cJ2LCrdHOny7jH3dh5apXphUEjf8zXvtu
hSgfSjKZt8IheIenrEw15R+t3iJASqOudAZ6p1LaIJmspFvCkZEb8V778VCVW9fI
Y0MfDhfYFQsmrtzu74ril78esiydPbg+ZxjaSWKEFWjmMEk9dahGMvuyLKc+LFcl
vOjTi1lBk+/7ZuSMl2EBJ29vxmEqbc08uBHZH4/Sz90Mm1TjjH+0OxZGHEjhoy2a
hrz4ioaCLRtfKX5fcNotVnKcJ3lDDgp6kMaarO8BY79FRXnI9L+s3RG+wUZzavkV
xvogGKUr67fEnz6e0drhYpERtpqRyF/gXCTdWxX+fTSSmPvS8zjbj5oz3VpMqR4H
pRIQAf0SGRUf/1mIgTjnesJmcBuxzmZlRg9no5HxYhilSj2mnq8KJ5HScjxEDYfh
VXjryXNut7gwTuCOA+XMvMQVgYCWDcOvnY0Km9pGuIEOvZx+QXIB1hMH3B3x+nXj
4VDK9KRvrholG1DBieE43j2ykHIKL9DopXp35ou0f/IFJ6A959tMJRpvvPs/O96L
cQgF2yeI8yiacLbR+mmEMiUK4H03Xo6p0K1bfxod/qBbzcl9cfNSayzES7ptmmFs
I8ssppUQeUF/dLlFscHh52JnKv7wyNHwdpFNUtmEV+ET1akmOX77xZcn8cfbDhUM
IQRKDZZiZoXvfpJUlilpXjdiL9jZYmE/WyZIC/DyyFdDAHuUGPoCmB0Tf1pkhoJJ
p8S/ZLqHAGor4rA7mKSi5fv5p6tKhXBChpoOO9INMSeGTosVZhCP/+5ulzh3MKPm
N8YchUO85bQKcdQt9ZvXYnITvG1xVAQIJ0Z3I1AmMPRvsnU2Lxqh3C1bg/ZPV4t7
bw00jZa6A/qMefWljAz4+W6PGUpXI8O4uSvVp+GYPF6pT3TPEV/koI7t/ZqPCqvZ
APrJIe5d+/ah1e4Y8KHP3eQpTeE+LIg90wH/v8l/7UY2CTgB/oD4lmHttUG15/bx
/R8MSuJavfl9rZMScokGzPioxFRdA5gc/0gLcfwBksQyMz678L8sQ5S6Q7PUkCTD
OlDivvLxFxxIt28un3se4AJZLWGPNSXeIfQOJSb9RhBvE1YwUWDoeRjSGVyMB8CK
/7vgx0w7M9SfTFpeOZ1NNjQrtYMsjG9qK9ef60ZFBBUg+FMVK3WiKN7vq17u30iB
nTXM4b5AOcdnwXgES5IWsCdsQlSHLW32XyugKtgTHJT+tSdb8HSR8dvuj+NJBKzj
RY0/JNKN/u20/ZKe8v/+Rt9vN0pqSccFvhlfS7wwEUWQXfWnGAUzt6unaQYXeEbF
E3S2aF/zBFRCNnAdyYV1fwNm3QyHfftsfTzN6bH32P1zWauKJCHieQYgm7jlb3ax
X4rxdVg3d+YBbv1sZGUtTur1+CZe99mOOj1PIks0aMY4WJv9edjXK82bEODNy0Fh
RZYXgQ3SE9r4tdMF/CcxQBrmeAw07LLo2CUdoSoIdpT5M7H2Gu0hq5FKL+yhOi9k
MKfLuaaItZPG9XLNpU6ENrW9FRKtzDWAOhn8zmfXZzqWxT0VfwgJBkCtSPwMgRmD
MD/OeJCL3Iv0n387yAU0MMV7m2IU10iSJwCszHAOurtlwFPStrEaKtX8OaGOrw5f
zGYMiU0jKpes17MWoRmdUAwCaiwX5aS8gqZ3o+dxsyVG4oqqvz04aOsIpclQmngH
RXje27sDjd43H6MKS+/24wXsf0ITMuOOfI/XbwF2/HJdvb4PH3uyHElmVsVEuCE+
muCY1KykoT2fVZaQrCMtQUhJxgbav9WSpb4h/jB48CNDVPPgonOR1bs3/HwNadn0
2vWIe1VMVIXW1xk5oFGa4jNB72xftg1MefeeFO/NF97LKO7HPeMTZErMriJgIQnA
5bPZXcTHpX/kUwafGJHQTs2s5dU9WtF0Y2WHn4pMgIkctkk3caFQGBkBrvHEGiYe
xHvkDiWNcrDTMbvscaB0R8X2B3uAbmx0moWHEfoMcb7f24pN+pKtiCZpzDNiF77c
4m0myQEf71vPxyugcH7EDcmZgc0pvPEizgbyNs2E2Y/ORG7eJCFxwVdKWZhovOTt
dk+9YrBJbEyHUb0CIuxL+iU3q72W846/LG9Oisu6kzlnZHhvaWZ6Ca6yuY6vt9w0
xWYzhP+rUvWGv0Ye3LAK/6xSvGGFJNIMrHcu6YPkWW2su0+QJcuKW7BHLi0Ea4/x
La3aHflUhNz01be7eefiQbOeOAlJ+k+TRswkf65PcsJFVOJWmUlcnDvyIdhXYlPJ
197k86dt5xEAbcLRWSiCgJXZrJtlWx2vEDtryCd8FfC27+pRuXNrwxnnM9ofnHvD
I/Tdm8hB3tlgwEg1pykQ9zBmKt88/Ojw/qd0NrIeYftLFORYotFjpyKzbXwnbjtT
1JgdQc9GlA1VMBS2G3h+KLQSG/jjaBCiP2Re/wz/JDyNlcNrel4gJMMhu5vAQ6/u
LauWE1bELjjZ3s/IizTqjur9vyu1f8vvfIDzMRqUbOIRGECFk6Sxb2+qqQgHTmhy
JuvWJ5KrmN5jq65FPtxIqaZKFrTp120PZL5aXZeIRPqmhr3BNPTLATnWoOiEmBXO
AZA1XcSHUPyfiA7IJnFE5j94UmxOX5a7C7GYSoVAo9KJ2gHuws52IECFR0xwTOST
Cwdr8p/RJJsO6IVBmSx8NupTzKdhhE/TfrKwTgYeNauAKoBSEHo3UeCEsn5g90kl
1TMbZBFJIhk8QpUMXWHqiQ5W3TBjsm+yPYEsgU5RPa3N/bO6sYAvPGlYRfL2aH8k
udC2qCEFh3N0gOlSp6duR6MwINaVaxLw1SbFj9/feOb5+55zDkLYoUS1gn4QSqu0
VN/0ilHvyOBnZBbfUF7JGalpHJm9fkubDzxod1QFn/CEFK3pUfeFB3aqDoBajiMJ
0FEDSmL/6oU1WtyG6JJSqK6bdcEiTUY3AHtg1IuZSmQ5+rTVECNwBtM1lo6rMfqk
V4FF6lxaMmeTebDYqfM8N0vYc/byOkDQHaKieSOVg0pypweDUjuArutBkqknOr1R
EnJ8pTz1pVmmI4UxY9uU1qislMXBkV4mejqUVDSu5M0Pm0/r0x20POEA17pdmuRP
mzcE4lOogXC4icR7tZIKMSIHxEowR5enFaEBjSWxK6zzkiZo8hTat4pedwRUHAT+
ogd/SFVyH1WMOCTs6V3wSHXF8JUbMYe+KOrKqFoo840kbX7eCza7XW2xzHxRP2y5
dkPTL9wPoKFnJ4EBAU5HdktXJRVDc0ED1p2hVByGeGy2Nfhg1EVhXLUN4rKSZLF2
a8dDxPuTAUsZ2ziZ9HRqClyyE65NeommTYw5pZXHYlTRVVzbXLkryKaCQyY1HYVd
KA76CdaY9Af1k2YspHCkuLT+IFV4D77FDlRjXzuqHoakuBb2ZjDHU9dvef+frjbv
w3POONlpAYXduYDfBSIsybeJRVyppBReqRHtPJo17/e44kLH0wcQgM7BhEuXyuMS
8bU3E0H2wU7pvf+jzpj509XUmdJjmTbd5OZWErByea6jOW0hE05x01VkKTV/9gG5
rg2mJkK+nImRWZ/eJSCuJ8ibW5AEnESThKx3J4dAdIOJtpg8mF/QD+xleezJy6ns
BdmMCBIGtDJsmyG/jsRHjJSkJY7Q1EsUlRt/9Cwt2DfAbeqb6wj7YOMmlYQykXmd
htQlzBI7WaUDzIsvvHeHp3mHeboUagLDwT5B7hdlGHJSXmZ3Uo7yK5C80COk0lOd
MVAaMBBkbjaiE68pQr9JJ5b7fq4G2peI+t48Nnfu9IGhzFotJTMPmT6+YSqjVNyq
6Xc8UV8reIIlOwRLJVxANmYr97nrhvEdMazZftwIGqoo/tWb9SQXdpashRPicZt/
3r/Xt1sQyu479Ld8zaAn0OvQkfACnrGRZ68O3yWjOgpP3lXJzWee8pXJoxVa2+wU
ZNf7t8E0gGez4Kr1eaRdHVaZq6gfLlxQ+AvEgmy+ZacRrVDYUCKg/YmRL6y/dEIl
C/Wwe9qjXhkc1ZUTXDuK1saskdjF5bi3bcuNObeY5clyRS0GdC/M4b+ZKyPZQpTr
SSOldq01LTW8NqSkp+CNt5l+dtNHrAL9+g8rEMvuFXAcyUYrVPrGACp2AqEq5qkX
mtVREwgMVnSreHZ40dFLVsvlYUQYyKm+AGuEcMJ5Q8wbQjj8N0oE5+WZ2Q4Lcs+q
y55nLbdEoXcJMtwccodMDqN3xeFVEWaS6O16aSOMgJNJtl1N6KTDrdX56fyJ4rhL
qDxsMhmp+nkQbbm9Q2yq3T8hItVwmhzBRbNnHNHtUDeoIa9p69+ExzIza0+ddVEP
FDSxp8HhXSEPsxP8cUuCidNnmAbm5TGe6Nf8/Ne/5z+CyRElfW7TVd01/ou4Pase
vJLmAZn+cDNSlHm1sapBg+8IqEpNn0hRutTiEK8V0Lbb/ZzU6l6UelZGchSnmrAK
M9YvzIbi0C+SKvpiZUvTJOc2ZWOv7xcsrGEW2ip8Q8zvL/aJNKkZDkUQU7wBmEbF
iq+qPnM/MSyJNco6ZXrjwKt/PsLoP9A6kgaDWD2CNBJ9mRSdKCPrz0pvCO5hfskY
yHA8FAR1bkUN1TM/LZJvInHPRAemZnW7H51PJKN70PM+0xp3wt7+ShdxRQpzkJrq
pZCarMZYQabJQDk1daOHKPV6rNft6ufjTenjWrPxLHXKF/ebQFHCA4iKiy7x/zbx
OlXQc7mvqdFDslR0WFbDiNluucg0anhKQeroTeEnpzDcl8RkKCFt+e37T8RaNKT6
sruwPqY7l5i1dAY9gDY9UNMcyCJOHp/+z9rBjDkpOxhjSyRRBxiYi3ocT3NyCvj3
w1r9dgsoomSo3BtMEIvYq0bJ1Qo2EFJl/btuxU6Usr1lOdgG/nk0vLB6c5KNMe/6
jH4/nBYbwgq0lGdtDkwr9cb412AC/gTuYFADQJl1BvrjtKNynaIq07dY5XLouOvV
8zX7Cxfph+RtIlpyeVN4ehibM3abtuQZ88owk8S5xGxbEdQ29g2CDuZIU8QRcG79
eZmEDzZq2+LeWUN86wq62W+ZysVAnqDL7v067+efsmbEIko4Tm2efpootcTJlTVG
aU4Q2f46k5oEeGrp1vPNYLorHnjWpCf8oUAVW2OkrFdsHeddhe1AFLi2nbru2LYJ
3r7V01hZvvlfNlWQBbD42rn3Kr+p25w11uCHl4EFKGXMyNyiykSsGeNvNRBKueiO
njLdP+pwVBgItHMe0ZgG7pHoYL37jRzHv0y31m5H11puP65bc4C/24Yf9IhOhHmw
dDo/WTDj9eV7GHOVnIQBNql5Axh6S/JK48EuSh74zDHK1UPbdozgXbLshAK3PVH8
I0eEKrBm23z6ViEWBl1UcKxlecF6kI8LJhnaX45F3PNmS5qhf5n3Oej9avZMW2O0
+CZi1+4MzFG+cu2dtfOcm1tixDAPSvpF2pQFge0g9+zpK3zgStUhIHvVdRS2Twnu
oD90HjZw3ShITCo9armLcNl+Wf9BD4ZxYO6r/1M3yRlYBILwymbg0FRAe/kt//gi
WPL0YpAyAJjLGyWTG16StpvHrQz+GYPbP75sHYvES8fkfuRJLP1+0cOuUxQ9bJ3J
mWFCRf//Xb4Y/0R1mn0Y73Y2yNA6w8DnR02Ss4zfpl3nhK4Kgvox+KvVjDONCsBb
12M3EF1EX3IQqiPfdPkU0KOFX95Ao6krOyXwVWkao/2Sy5J93gFU5ANLXB8RKOgl
EjShchgRAcVc7dtGhAJSThxD4PQKhpg01l78H5WlHRGkJaDRTEiIx8bfMZb4yW8q
Zr9KywE4v1MZqQ23kf6G+0rMWygoEapwaKsRjjodLo2ZS6wafiys/VlIsOEJOWUO
bsWJc5DbSXe8riZqPBimHwu1u7x7LdlTcV0ejnqeiTsZ1VLojPpkvf+c/nD3MnaR
4UTNpx9bGFW7hE85SFrivs3LOk+xBDMUoFO/+IMDCb6qLvlynxuPoXZt0fXn3XT4
eOpd9qkA81b1Me5Wu5qHnhytw1z8ZMrJNTzPZvF7xihpulQ/eWYV76jsD/h7YmTH
aTuVBcKoutg01r5h3cKlluLkYn8Qlos6hq0Jo9Z79r9LYQ1gO3rIIQUfrztKwbR5
5jFnZAKeBXYdf7AW6Yzj/VsG7pAV2c6IhcDi7jlXyQjP5Bnsa19onDSHJVGDPBhh
TIJb9qkVZ23Vpvz9QTxMf3coxYdqtw0SDIJqaTP/9h1ZrJgjUoIE/tef24x2a8lL
1BMlWivGLKOgkucaTwwJjHzYIZDs+SgtxEshxDh14NeC9QAhs3oh5jgV5b85ohI6
FdUTUOl83DW3t5MHr28wE79phpVpbOLPa/sAHysth0FFKHNOsTJlN4lYj+niOqsP
RBKksEf0ZNdSeyqIJKqxYr4ccVtwHlhjD1eQj8bDOWkc8Zg+2w/NyEaVcGtoTQQo
dUmCvna9vaKEzIUlFw7OGmBJbxvMQZbx6oeaGdHstrEtHShareK1LF4M66XffBxT
FPcm6Su75SV6Ss2g2iS+jsYMnI59Ba3GXt2Zw9z8DMyMF0rMnIRjrpyu+dqR3Hik
U+Fqcnw2FKUiTxrz+Y5mT5cOEximpuuFgQ1z6D7v+kstbSNAHxeNuBXRn8dYL1Mg
+fFrobH39l0OCJajoSrT+xNUefzTUfF3vz3UFDlFMlIoo1Lw9iC175fTgO5HoElj
nQC5H3GKVHopXNFy6BRFVGjJCzTeR0y5Ecoa8NFzjz6qvE1bvL8lK4DUKJLwwiez
ugHKhGgCuknYCFBiWt5jVcqbe+7yjwwwvxgh4CIYBPJ6ZjR8czQbbvj71sDEUuzg
ZmFnaOSRS5cRgjbmEFWt2ed+jrNhkdAqFMx6o08qhKyi9SoUhgwnv9rVcC01Q+4d
mN2+devbAxxrlvSbPDTIPmfZlXwT3x/GaedilSdgqY+PnMm2hE/wZBR8WF6bIx+S
kfMyHCWMA3RbPj9uXI1/Jn8GAsEEZXsOSHv4H40VttOdVjeCo4pc/iAigIHiJ9rt
9+pk4G1Rb+XlCcIrj4JxAIM6gy+DnnXBGCBptWmNuht7JvN24Dr3ecSsWvDL4dUG
gPoXA4RVHZHwV3eoed1TZXjyZRQnvzbzWayrZLiPnY3Mof0pDMrX4FR3NxpWfUBM
XqLJmXj6R6yfGMEvpRWulg8NCZSMHzmWpv1fPjYfSrNLzo1BRltBeZv7CW65vwNn
U01ZsJtOQf0YKz3jqBG+4cmci55c0QTBklS6l1KhcfUaaF++KAP88X/okUu+ixSX
Yb4YcFeLvDNOQwde74ohZUIjMFrZZYutoQITKjdlRxAoGxVQnQNE30Jqdy09dF+N
IwKZVhjYx8dUQ44tbrkmeN5I6n89/N5EnBQsEuTuaEYQ311f3lfJSVGlnnagNKP2
lqqHhmzFFeCtoFzBsQTZxwoitIZPdthq/SkAyO2Pi2Ay7tKPFmY6biutdCPa8SyY
CLQ2k7DqqSWBEzRH+Etk6EZKe7D1MNjVAAeYLhVuk8xJoZdaqpz3JFFDGwk3NgD8
/fkEIRu1PFduzdK2jREtfw5l5iWtutJ8RtDLeke7yzTctTtse8xqnZekOYem/o+D
vypWY1XLYfke4/VvfmVG4Vsb9xV66LiWiGQnjBk35nM7F1lZ8QUVXPOvbkLxzwe2
QIpoCF1iqe7sLi8Kv+ajvjgTnuHgnKeO9l74OdtipvMd3j8g19cyYzbV/c7nLxBY
eNXnniTTub73FsEAjJT50vkz2g2wF8bNjJFVvQGXpGnjn/kqsN0Q++oNSf4DCGeR
jFdnZ12VZFcbBi2HV7VKJ49LtfTE9GfvTxKaSS/WAUsqhmYz5PkbJHKIZxL1kLX5
CDuU7/bQyQRn+iAEtNBc11pDDK+xGr9uroOpMX84mbXqy4cA5lo78oj/hM4/CZoM
xuurAYhzojyweoCZF7VMRz/X3xmlb6wRf53qzUpZOybaP/sW96zguYcNdMdfXKpd
lHHH0xYitJI5BlcOBJBPfAT3B2FQXz/vRicKjG2WYQI7y5hloYlOhw+Lcy5ON+IT
7NG0URLNZRhu5b8fuO8ykEv7HZkJ61QSadeprCzbCqrWtX/9xlrEwOlEA18eI+HD
hulx1rT16OkYTpC50hAGDYntjct6F/jKMIRw3/89H2jZE51VL7XHYmTB87JUyG2+
LXs5Of2xQ1IcpgnEgR5ysGvpSkEUrW+5iD6fAdO64mumTcXbPsgjdBxO1J4QACgB
LSigE+fewkITJxMYggSAYxnlw7XYgzZcaNRbPvZcGUwuzQDsw+Lp2Ca6BR+KaNb+
E3uzpV2IL2qSp8k9dDbVyTLQ3b5VpEyuuq+UTWinanDVp1fqwLzvvGpRnZTeZrzP
81pExUc+epenVv+c2qLViJ9+uS005CyAHGodaDkx+pp0GJUIB2D0Xj7HRCwme9DC
EytfX9na68NleGxJ5fZHV1XUy42+d2qcd57Z66njTqjG9GyfsEvAAOAJcM7QAtgh
dSVwlAzXikiGL3ejzJB6wqelfPVrFKI/HYrZJW3sN7y6RM63UoAFSLbeak5gCROq
FZCvkkVSZBehywDoD9/QwXIcLQGuAO4fvyvnRpCJLgdKuzvCc9iwSiFIr5AGJJrm
FDzpz47Gzs/xux53nhZIgpUFrvweI6x0ecfJ45uRQ06YUeFzCoktm0+x4M0xhbHQ
nljWiF28OiZKgI+yG9LaaZ+W2Tdyje9Bj/6ogBgDPbvDFpPjZ+XVU8RaObn3WPeZ
Yz/u1KOMOfkJUGrjGqNddpYup5KX49wMU08E4EzojbF5eJ95c9vGi0wmrKtHP94S
xvZMHkkP9fsN0b1Q8ZU96i4BqYY6+OGmSYHDLeLMfRdsIgaT2pJS/d0s9O0jv3QI
laUNWt+mXJyvPJPLhQ3SePeekuyhW8dzFpY2ZI/Lzqxb76r+tzgRynWAyKFvI5Ut
gtsIMo2DSK1yw7UnX0R8VUD32+FsmU+240ceRc7tM0PZ1Pes1SfzLEjZoN/ovL2k
mv5e7Z69V8hVKkB8tyfcpgKsK4JSZU3kZ46TseP32VUjZLw599PjM2oiUrxgCr4o
VsBTOfafiXDc/jxV8bGsZkfZzDofmVmRi3W32Opmw9I/DYX0IQMp7bP8pH3O7YNX
tg0eogQOm6a4/zFjaFaJomue4S6zYHetp6ypsJSuDsgvR51a5TIvl7xz45eUdcdY
FqZYqv4BHLYZmSzOALGOnAO0Bo4Iu3QZclFdkirT7D+dYHmNlPp3zxatDxLUDfWU
+JXbg9WQWUfDyGMA8PrSAD/P0zJVeAnFmq5EL8Gh6AvUrq0PN+V0VIImqhm2kPqP
lNuhxayjsUgmPakwKW6J4Xp7QFwzVANlxpGcdidJlT2z+k/sfy/s/xCRsF6UgOqa
EN2gAiDuetBPYwcT8XolnTXsyTy1pNcKDWj/bYnTayvrRMY+oNyj5V3ydnG2UwqX
mJvq8aF4ejFg5XNqRL9KHlpBW59awfgWCZFFHI04AF/B2K8yk5O8k6rowZFLhpl4
BbpvZUXq7dPSBD9NGeLf4KAZQv9K/dpFbsus6qwRjYLt+fARfmUKIC3LJbub4er9
BBayBAoeYgrTdmvmtQp6Ly2oPL2lsHB2wWbWRdFBQx7Y1ELaqgfCZ9z0XqH4/ba/
pBj9+2Dux74rlz8W+tIcYSxsjuc8rEJkQ1AT+H7qvRwrLShKdU5vCZwsG5DTeMeH
WArXDS9lFCwZw1Sgw0R4FdF9aOi6NeVkBJ+MOm1aEKPsUjdCsH7BHQMVztYR/39f
GsAtQ2YSwx/Ywb8NxD5ThDud+dvdZLBYCT1I4ykZESQuWOODr9RSLUAEEGuYe/Mn
nCWMOyQoBeZ30mQiEd+e8WtJJNYjJd3sjslTOcb4IxSLJL3j4d+QFETrkVFuoowU
iwTp4Ke8zhRQK8lBJVb1VazH+oFZ89LaPuqwW3s2Wb7iLD/uNuQhIt5XdlDFMh56
lwxoLfeVFc6AttTDWRtVQLkfSft9slRZl2TDbkrFOvnrjrYJ7EhDb4dhzntdWrgd
i4ZJ4P7fIANjderuGpVKAsbrY19UpJPlm047AC8hj+SGftK8OOYx7oLLOCVblzIx
IMejIyra9ezrneu2VpBm4TXoDl1os/pe+h1rONUn6itQniYuSZPiBa1x/OSPyJhp
JCYPRL+NZ5rVpAn4gNPd2vHecxkgi3Najq0RnFkdD5Xy1e+6YhIYcMgTkyxeG8ws
HeFF6qLNdhHZ6w4xCZzJ5m0Fh09U1kk1ylR89hFuu5AvjRDDsogJmLxQiwJmyRki
R677TQDGFxMxHn4FWSaKaUk+I2A4vP69NsuRT1MQZ/qu+XkJ2sjJHYQ9b57ZjRLj
q/qterHaKCiZgB1Ikq7zg4WrvIyxmQpIXDI9XaH5eBEg3gWFfZcPltwLrfFkmy6S
PySAmVCzHjSjA0ZsocuK0bHWUIdW5Widt8zB8Q3R0yQct5UJYTz94ywe83Yxbvi5
/F26N9bxKhLraKZR39/ZQNa3yEna+pnbDn2BvtpxS0Qv+8ymvyb1UBOierlytvbh
D7IhTDlEGCIhDGlhMmQg7KzdfpqKOBD0s7tyWGeHyZKaYrccHBzubS3vYJGFBAu7
LGWFNebfHMozexxMQSz1OIIqxHsmPPqNMG+5SSWMeMlZ9TQP5bwwjoxPQc9syFCy
Q7uVPwJtSZuwQwIIx2m1XMjdTodzRn1Q8nwoak2w70JyM8Wgsr7GJhxC2YiF4GoL
g7RZh0aENFqAbH4jxzHJsgynxSMXty9ll6JcL17EVMbgGI88+vyZe5qBAriAHjTR
aP3YGEmHdC3L131Jh2gZoSZ7BahNYAegF3SylM2Ob5mG7AoNfCGTYeectiWHwHCs
uimr8WxlVk7+QiMR/JF86xHIW+++yCML8l/KCkjHAjMtjglm+mC06sOcYzDZXQq5
IjtKgSh1dRDZywITdXJ4idFwoVpMO4Xti+orxfXRzZK3B9E0djKkB2NtCc5f1YD7
pBWqjL3G1/Zo9egv1P+NFLqLNXMdfl6+603cFYoKWrQ4k+34ooyipz12Zil3BaF6
7svKC4+amkARINSfNjW2T+fPnxPuwbE5zVDpLx69n1kUpanivX7uvVc4oI9aMYjA
4HSo1aPuh/zbkRuGUcdePVWdo5pN7idecLl3GZQzyLkdGEw1JdRRH0msviOwTxfV
u8VUsEK9qt6+sd2XS6ESp4zyhc5GYL+i5kbhi2y0HBA/h6Cz45d1V1RIBsl418Pw
CsKrbUsoX975wxo60velBm1RdeXDIuTBVRU/bCOTEiZb2xedY/dKldWr0TOBhZNt
qqDgzGSvBKE4YZTClMcFdJsad76Ibyxp95jBtD6iaLFzGE/fUkGuoJ9zl+Z0EcrC
9rKg6KrGLuByU/ydYGJ7rwClLAMAaMCg9mxIsKJ81MevLIWbIwCGnuIrWfDlsfTf
XUaLXmNjBDDSeRlVzwzUD+ee8fzvqr3l3PvqeIP37hEFEGzp/7dA+XnvPO3SbNoK
PK3ftLSiQorJwcEP9rxZ6bBU6az1xuzGvLzP4LgvtlBRfSAeh+7lWxo7AboR/hOs
fn/2uxTU2YGR1IBRxe44Th4do8CJiSkO+gvgTF7T7CA5060lxEy7tB2GPBqvHaeG
zKzgsrm+UvEzT3VL1UvdaXLn8wfZRHp7LSLHjr4RSgioQ9vkYQjVZxEEkYEQBaSC
QsBhBJzsr8W3yZEvMVpm7vu/dEpPxZFuGsIrzn8ZHxfaJPGDV7YvFGb6RPXBKWAn
LZfXpCD5l2cxRPPqo8LjU9lLZXJyJQBudubcOG7WNAJ87mjBMfWh/Z50r6TCr8eN
Kbbt+1+8kuXmD+zeDHRjt7lM8hL711cO0ivEmO94W5fi4bV3oergfhuF2BfIY5tQ
Uo+Wru14Cf4N5RCSGZMsyQdaisxthfpBBMD8zY4GO4hq0FoIfC1wPN9+LjE8tkD1
tf5zXuugEL61YwbsCe4j8RJMrVnc118WB0F0Hj8HjbHt42sFoy7fq535zIRy4R/F
5CJyFKXk5K2QgtVaR071wXivhCHSIrJw9VFIw0BRdViHtPircWr04vCdAuQiaxeH
OijT3+1eRUiAP6ExOEVo/ayGpWV7UqcbN7JSiGJcZJSTftvl2axS0pCuHVrs4cTG
QIn4rzqj5975TWk9QrYE+7KAuPywgetQE2E2V8KEsXWOrcq5ohI+hG/rUURf787W
ketBepwJZ1eE3DUzmQxRT4QSy4suI6R0f1DWYY9jrzkAtsy4/4jAHvVayo9QBWZE
yvX/oUpqkNmD+NNunVvfWUXRXxKPcRg3v4f/pYpuyp6BJA++ybVa62osflxjW/5D
ar/xTsobwZaXd1OO5wWjDn8sIwmJNbOQy5W/5TcwcIfivQrsAIcA3oqjzgrRlUCx
OYyzazAWi5+I24XO7cXCfZjJ8OnzQMo45WbQXI5CtA7dnD9/TmpxokY5LA1wEnBI
r8ntYVM4sR2yN9H+3ImsuOTdUx8gKtf31tZqGB54GkiVMN5ZQxTZfBLL3QbymoLm
m1kJL8YT0FqkmblByWpiyJxTk9WH17W2mZu2412d64mWxZNA3G1ANc7fZZNn3D7D
bagvzQ7Lwe9/cmE2dPFb2AZVCdY8tGvcndrmUJ2nFp0FajfL1ubSYW91tLLlu8Fx
e70r9lMsekwROczrWCos9/UHlAwA/zfMR6u2vDOIMk4sFKWZnX7K8MC4GuJR+L8y
pc7vMhw3vbDtZ2Lf7m08SrBKFBploKiYW/M9W1Dwc1iB8jL9k53ZIlcrBEaga0gp
xNFbzpXBm14+UNFTqFoHTt0aIXkHkx2/v0iEBBXjw9Rkp46wpHZXj6w8B1YRLilL
5evy1aYpHbY2HsAqT2EkpLLnIq0LQKD99nLKb2ovdlDB4MJAS+vr3KEJJicGywu8
TQep0h/PbTXVLivSPM2/ZiGWmsIJDtFKmXDLDuzdo53pMvEtyyP2wqJilp9yEdK3
T2Sbzuira7qGPQhqFHVh7DBNEVinjDiKDmIdHuyi6HkNi0p/dR/pclghB5ntYoaG
WL6B9MFhyYXls16Fyipq5ZrM/wu/v9a5azNvCpq+Rihlj0Wm6ZYOJUh5j/bdZ+sn
iMldGPKXac95+Xy7gcdCqhjDtS4MrlrxKi+gw1Y3O7bbv8Lgk4VzuPTlr6jHyPLo
oEVLP57nIm53LL19C4iYtuw0ZLTAc5I+PgDyloeZ+5o/dVWWXGeFt60wxEw4wGdV
T138JotN5VmHFjDODbL3O9R2juTq/oKpaPWJAZ4zQZ1pcbbtO0hnXmlqJUZ6lntz
RYlw1kMdLaEV5vljpgeS2OiPkALdfHdgwlLtib9nlQcwxidW6sKj6xDMA7eQxBdQ
qPV0IBNlAni9EFp/c9GxF5GuJXj3HwcD6eWO/txlKWx3iiGoumqmN2F7Ko+skJP0
QnhJSBGAIuG7gZm9yLOpgnqc/+9BtONTTkQZu9Y+oDX/ADpijMl0TB3wfjoOBDiO
DcWZZs6EuUmV9Wi9s0bGjWLIwM7bdCe13KbCytrkanPwwOn8HUYgrjDWjfdldDaw
dl8dNhn1YGHly/10nn54F8wxKKOu27Q4yfs8yc9m5BAuymQ7TkMCBW9vsT4WWp9p
YSayfdQdlx1wmLfrUiSkggQFYixZ0vXTsIAnQVKnwCwwpIV4eH2lGcmOjL3vXrxp
0HyU58ORNyEtUod5Rk/HqcubmtylY2qTGGzuvFyUha8Qo6yieS/jDUZO07mOF6js
XOtzBPgaoJLiZ3TViuVVKHnynmqed2iZpoVdLksend6bXkZXjokDbRetxQ7Dccch
hjtmfsLQzcBZN6AGl6S2CZ+RWRAzKhE+0q26/iXe84+1JW5RG1ylv+2E6P+a3VGB
A+POtBEAkDQ0EVfQ5IynnDyS8uOvAiu4BwlvQTvdoxCJVk28PMKwNapzYDvVMTT4
DBJyHRKkkYEKXUbonEZRzCvbM8YQhguIXaYQUGqv4HbPPP1V8ewtjaCErfg6+mwV
HZ4qDFtt4rOeEYvg7XvNwtI/lj/SmezdipHuN+6Mp1q+UPWIk+s5jbQV/92s1kvc
7irBwr/q01F4BhwBqW5eWMbfouz8eSlR6jwj2Kzf31DTF773vyclRc0UjEYwK4of
Lkv8W437vtheu5KTs3ql5aFDiHNvUZErmvzUVGTtNWFuB9cE1Ung8+wowUAeYbW5
FpIOx8iNUr770XEdhZ+s+SYklRGP1E4rkIrVMo22l8BQAOH2MYlHqMvUbdENRfap
4kVqwMtxQpgzuX/vAmI37oYV9dmO1CXwGr8TYpB/5U1VN2xlVZkzGybYDIynsisg
N2PsuPvOMlthqyuk5rm9GtqNCgKmd9YhMGo45x6M8J5KGp5y77sGr1NilIm11fWK
8OhEmLAOm3aiT+yQ+nB0R7yyjHbc+73AARJ3IcK5EI+WeEVYvKgbyBfSq1hyYlod
BYH+fuCecHEQHHWGm5m5/Xc7CqwhWRO6EKVimnDWpH0PZfbRmbpVy34h8pYaed+z
7XtVyth0PGxe5W+geyDnqR0P4gqFK2LxCWnse3BKWfbAJ4S+w/5IYgppTUduWd0O
Msb1hZHhfyk/2SzTIKWJA51jcn9fGMuI0Mstz0DK1JMKt56XP6IXmIpHdtDlr/GH
fPpEMiwi4xCh5b9AWHj9RlG3TfGph6dVRa/MhVUuq9DrTbsBh/hHeLELLy/sfsBn
XsduE5hI8mwcFWwBEKmfWAuX9GGP/uC2VsitlSzAoLoEwBodczi9smS83egYt5A6
3TcPqDKebTbrMyHE3ka8mcr/HbThKiQzJHK/5zQMtPgkk60fLYYyfSE+xfLDmOol
NMPw3qejkuGwllu2r6MN9Wrjvjf5v5FPTp+ne8wwdtfbqz3Uv+kPTvw8A3b5vgkR
KtDhU3e7cILCEDUsqgeNxWjj6b4m24Fdpl54b7YXIJSpNiXX2xlv0oX1QIFw4qSj
x3TF47Za974NxJAH6bhmKX10AfucYrNDP00WpT9ljl2MNmzNqhoTza+7knS/fz0V
RZ64Jlp4FdPfHArZ4qGeHnCO/ryLBhFoP88rncKiJQ53oIFWT2m3o1to5CVava7T
ZH/f5yPX1bhgw93GNmkXR3m6IBhmBX5Jv4CAHeOGa/miEpSM3zVtNEAsbbwEx70M
6yvQPe+FeexJ/DAzvCo8J5ZTMNWsyd/v6Xq2pzoqq5hs77chwpJ2jJZ6hGxLcuxI
FFa3EZfFc0QPnT7kIRKEl+gr62FQa2hv80xlqlQCrajAI5CcusjS8/2HuZ3VmP+Q
CIXZvUG7oUxYGT/PktivwId89gUrhKcQDLC28GXVsfg9fqgi/UEw0+mz88kuJxWU
y2WyCSZzHMm1Hw2nLWV2rCIUr4gODs8uM1y38kgfHXJZ6a6hUoS15KTEfmdNFBHU
SGOuYMB4Q0pZZQ5dyAnGAlWkg/JXM8laeh3iEoZIRyUa0TF8TVaS0BmbL/KxlPvo
Yc7sOPB9Dsjl5aIX3VgBSCQ8tlBqHJmnviqigRCnHTkau0r//jBeRFxI7FIgNyhl
kaCQWqHVU9l5f5G6DqtC4EA2cHnEx9k7Lt010++AdDSVzSx06yrkhsldswkStK2F
ZHYkKfDUTkz9NynNafPRew+Cl47t2Lv18vXzQuyTT2o3f3we70xtxn781z2LbTdV
5DIpw7/s2UhVnnKHA96iMt6xo9eQsTgeiKc7as5Kglr7ifuaPppVocGEJYYri99w
yxU6OJeNoFDMtGUfU5J+DSyOBqCj6cg9UKTyXinXepWSHh9fqkf034TdSeDtPp24
9xVGQ/8rtlw7s+kewEVaLHQUXouwi/T2heaEIUK3FkM9BWlx5CGjjtwhedh+/6iC
fpTd2xlnMJMy4PTMQM9FIhKadIPzpjx/wTzyE/9kxvQtUDysxLQ1ApFo1XBZF/u6
g4Gr9sqxwry7220f+yrvgizaDHWjtPTObDUA+QqTIEShH5yiu+AuHQjlc/KEAWTa
nMMgWAn+9Lp3PKWYqKaA8v1hvJk0zC7P9bCcwHrMDsG29EtfnEkuOQ2OSKTnXP7r
OO9UC+djSRyczychdHZeu8VyGCleYYO7BoIkI6qm61hrodft5Y04xg4sd0IdcInT
EWaLXfGPDzJ8SE2V9atdMZ1GHeJzJ5wLvqq8Mag0tRA1yPCMNbSNB6VPSFZA6/kE
z9VI0fqEixN7w6LRU8sBASEzyhBCovZWsqo3bXhmapjEH4KDstZBaHuNax+WFCH2
gKikCCSnQd8UIcrqQKzaFfHmc8n/0PCcEYJ0ntExHMv3GbpLXdwbSF6/4xMGdyxE
t8HTPE59P8QehScHWJVCYmRVWnUSLNbl8y1thcr8NeP+hnFTTuVgEAv1j63Kct9p
HJJQ7NRAa+qjwH2sWpsi8LcUq0auwmndXnaKGhsJZKMJUecCK0RoBlcoz8AfTlvx
PgqFZL0j6M8glOifAwckn0oD8ONLUygn0tqicQl/ewVasJn06vJzQ1exP65+yQLX
fw+js9a/6VMw4QGybB0ZSLBUh7Ol4AHA2N2H+BIdiZG5SfQn2bllTN70QMEMHEKD
BEbhml2chUoFb56HIeXJpZgO/2jHceIjps0t/HppNh8wv1M0mPlyLRrz73HwQUoP
RePGXwomrU+xqIxGoaV5Hq3BqSQmLnF0f5LybXwf+65VkXj2vppYTtl0DT+V8MT3
x0buhtSu8Nvw9MFvNSnwX90D9o/i2RQ8zqI1b+AkN7MPHdANHHvW9GkQ/DheTI2N
+yvqieGAVnzxpBypKJ1BdJiPeOCobTR/nXHhC4UwmClMxZgf3L1cFGhyGsZ0nPHN
F70q6iInDyVp2eRlwAt9MuR+0Ixje3m+OciUC5oKlFeHL8BzOIZ/j40UUWDyVLsz
temI8wO2OX81f9YmjRKDhuHDVtbGXsFz9NV5r+et3MHOS2dPYQir6OwdyqGQ330i
SwduHLwH1zVQo55cXy9Y9HCfy4aUCepR3IxxtypF/S5pLf0K02szJsMoTSDpCdEp
AkGZzKTzwGRc4vBs6tP0KGp2VyLpzKdBSLp/3I/CRR+6Q76IBWVd8YALA/vy4I3p
gh9lr9eg/Qkuo8umE/+QxRREok7vhC2WNStOav6j0r5ulntvXFHnCo42eGrU2zZP
Zf+54hPh41+3Bp+rfHs6uLtsD8JKXNqg88qXWZDJ2RmbSK1u4hHy/aqyTJry6Rc2
GO8pmhjgoRSyZRFlCh6fXMUhrzbvA6Qga6X1zvWzyKdIJuaZJPJTcioM/IGINe/w
7DgyF7BMEi9BNE9YGzVwgdekhClHr7vd2r6YuwGInjniESMM4nP/0smMXv9H45Se
xLObmX6RXbsHHzffc2xsXl/5hAvKTzoAmdZQg2ljggHb1FE9Fn4LXkPJICAeYQw6
5/DCNoL35uplpVJQazPpdTVOR3lwry6xBH8tbLtu3cDb7RWoHgbsv50JgGDzsdTE
F74zDpGbMXNuKagRm2j/HbFm1GakzQZDnVQlAndAtDUzXxTaCcB41KqBjd6DAkvw
/XjK0NDWcFTJy04lAfeAlz7nB5L+BVoR4+JRydBWj1h9zSI9upN6rP2cS6odhuWt
H/nVgJY1vdIzgVjerj6aqIn20Ha+HPYaSZsVupvI8Hx/3D9hhQMIJSenQMov1LX9
M+jSUDHx3sNvIW8h7tY1V18TO4FeDNvG4bC+P6LBCxEicsvU8T44uWBgw6gTC8Vu
ugckYjkvEx4L5nZ3GUxO1yZ7gZG/D/Uy62YOE5WdoRl3m2MuODTFVVmkL7m7YvTV
myvVh04KisogrrwhvTYs8CCeKrMWS5/UZIAhVhoQmxAKhWf5WEzeBfGysxeZxw9B
Ad69rGSpY5XJ+MzdHfBcR+4dyTjWFo+XNJeHj4sVrlMnYFaRZlc4oipm1HrsjaRo
8yJmpRVtksUGJmmbCSUNfEjtj2D0sZ/L3zZQ+4pSliwtJnwZXnKbcIkxhP+v22KL
kuolyBI2CWLutrmavV5t3qx1ZOo+f9rCCfQxyDOH8XIV7waGcpYskNF/1TJi8FzF
3nEcWo+bXM3k30X9YHclCFn1/XbZXu0WfREqG0EFMYsmTsFXfB26xmfn+1TeAE6o
LOgaH4zuLrjFbUI33VJXEinUIkNIlqLiX7sSxnXRpDQRNiEuuZBjW4Ow3nbA80K1
4QXJ12A+/HQRyvNhWhh7dbkmvmaTM3vylfyfUhYF69b/A1cfsl4iMN8Zcrma6//g
EAPjRlnTwwWiQMyncBYLzESEI7HN2wbwtNoMMiC5FEeQM4tpnc8Iku5bmphaZ+SK
3VTNQ45mJmgve0oCQ1OW4wRO01wVu7fnv791NLRCaET+iRwFfaC/Lqh6UwjA6iAv
7zt747mosFbEAECRJcv5Zd+vyhqOTW8Lh1zsUdLg++fvrdBbrpKUMAReCLDt0898
rzMeVbCwwtxkGwRajep+T5UmGtB++8AurtvRKee2SMlJJUb+IRA00d7AU1zN6jUD
nNIP+2BY0n2fSmonRVL7+w1X8gqU5O4LdxAGp5WVfvf/koemNICxAGrKZF7Enras
n1TJN7PUCDEs7jAqbX3ZfEJDqW9JNGX8r+ic7N3a5QHcxDKWcmHgSmTEOgVtKRao
yn09fQdp2JaijRkjLwlczDR9i65C1uZWdyOOrJL1itEZZp+Vy+VFjfLKu+IHPDKS
FKSZZLzJOnHqKAQTkCn3xIUVX+zSpFbwkL9b1dJFOYyobo77ddz+1vKn0I4Mw6UI
MZQmDSIEexF6s7T2/fo2f7f/4DXla10PlZey3DlN/u+Srz5YhhQ6oLwEkHEwdjlr
uTyDD5y3moZuaPXKImAqPGKF1TfO8nn616ChE562IDxO6PPyUCaOS9AcBuIj3KCZ
5XgMDZprlt0DCnWKEtT09XFnzEhgn9a0o2NqqnO2cskam42sh99MejmIdmEBja/r
l6LvocDWB3ifRQaIF89U0NNcAgmcfip6i2CZKgktCbGzufIXACepG+Go2JMVr7L5
Ah2NsvTHoduU20izXZeye7+cvd/UdTV1ARcrfH0JZZcuKVWMvyqn1kX0s/0TUxgQ
XgJ8uAq9+E4OnNJZgAfMN2RdN60xOTKDa4Fuu1a2/Iov6en+1qLlLkyvbfGRL4T+
tiaVe9o2A5Un5V/NTEdipLt067CThDjQQN15PX1qkTs=
`protect END_PROTECTED
