`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Mty3aR7pLtpFb054zpSSVInTPK4fjVLUyRZSooQY4sbjxr7BIbGrtdMjh5M65qp
iErANCz9jULPsNB32wILD/9dLB5aOS5g6hkR9mLhTv7l7lHLmRwrAcL08PLIoGzt
+0VDQHkBU7vw4SApzGxIWChlb7p3EwuZXVxv8DkQmV7QnnG62nXh+wC3Smi12N5e
XlLOmCqQM90in3/wdT/8Bi2E5QP5PLBWNwqU1gbfIjPITX2FSA2f8TubLwh1kYVB
2aGWYgM2eubCBgzYfqs/eFcQ4B3ax6BlV5E+kVD+/WTHwqZ6liGgBz5SCxhvnDhj
mxiDvQlgGCG/8R763i9/51HU/YcTZzvkQPT0sOf+G177SsWe9P5L0QfYplZRh852
oEB+l7DGqsZWgOnFcuD/iHmgX91YToz5RGFIz+QKPgefZt5ISzCfnVbVYZrSv5xq
kxpLl0GYqFqcplMXmLus5Al7VMUmQt+LUWCQKjrTeZlCGKpy/dVfu0pqei994SRG
HzCAt1zWCV4o7o4wWhHOEvdl+InabMm9OMgzBRk4kVYMqP6HVTUmH39fIfed6Hc6
ML5lQPMDMQilwKwK/NPji4boDzhPi/FZcXayCXVAUV+ogoa6ADx5VMOYnCzBLGoW
s2KoHkT5PtZW6SsO8Elq68V9CUvU8/Rm5ed9D2MaOvwtkp4rkwwG5w5SjGg767a2
7yAw7urDr9xwpYypNa3sE785t66uT6CVcr/HWBA+yoRpNYOSSAfTv4rEUJGdfivF
9XjTTEl6s/LzErjW0jlia+qTGkSYh3n2lUDtbK+xOy6LadywdTkLhKW6oddhmoQt
NifeXai9vsIW1gudvfRJ3+V31rF0KypX3OY/rXg1414Hk3ArVhyDpkYdKpOJGGIw
/WqyKB2xGal6TEy1lVlQGOEfgcu6ipj0Mv3oAGaMy6//AJRCgtdzYZK7reuD989x
`protect END_PROTECTED
