`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b8qGN6FK5v6CNVvisvZuHMatIwKbzlpECBub2RErLeQD8C6WBUMx/ceZhP+aUzxv
7Fn75RBVFLwr1q4rcxwdgck/51wl+CFtlArgjg7otzcjioSHFIWL5ZsbsmYipwRJ
cGyqtoGAnS4Nseo5nBG57rn+GeGvmDg7KoQxQ35LnNRQIA1cGD4Af3TLWrZ34SMB
ZzdJcOpjt8D2249dUQDIKn0bYBlKFl6AeSkhyTtScOnMvURwnK1rPJ/Fb82tUMj3
0hbUFvSxGwcGaRRGmdEGfULhFLRTPvDdahrvHxae7yU=
`protect END_PROTECTED
