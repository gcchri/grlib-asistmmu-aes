`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PoenmVCMGAHWxlEETExcTkc2mzmgRfWz822UZAmQAETb9U+aifgzC8FxAhFyRp62
YC2QL7X8k8bR6xq7L0p3aDB+xDVn0Hw60D4ZoxJvmLDNDjw2c3RkX1aB0FXNw22I
aJXFtrb0F3Fr/7HdjWltlDugezMQpXxdYC23WRmwFhEY0RHjUzs0d2tmtfP7LTdQ
S2gsQH7C2AIBCTjrwv2UWkZbL3GE0isMAeiH7u/0Ds89s4sx7xcGriiy1G6KDQcn
91KG2mFuoWlqYWpLBDKCPFu72ZA43B8zhoO9+po0qXL5PYy6aWXEI6Zyp6GXlriw
ZKiyvVajLiUJPpjTfNkhCNThjY0F9RiT++UpPvoWqAgzKEF4BSkWS7DoFzBKimV5
Ti8vCip3wsgDpIIm8lK8+AIpmrBZAl/T4NnWVPXNS+g5ZF/KGALOXYsbP55u+n79
Ro0gwRXsBomkACKu+ewhEg==
`protect END_PROTECTED
