`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4yLpZKxNqtSx1K0jleDHhK8vWeP0TvJ2cl6/A+7G11rLSrNgDHqsydr5TdR3H4AP
iGH99fbbzGiXxHM9YNVzWni+7Pzi5ujwZsVVZ4aDr7IwMGkE/bt05JgM2T0SCD6I
ZPyl4WTJvx3Umx9cAzqzhJyu05W011ylRqi9prPsQkH1UOzA2TXdk1pfs7NtvELJ
W2GpYZRdYMu8TPgsHZPgpIj+TxRNsPuinFsAPXllNXWsQgPmjH370t3VTg9sO7Mi
HKKOZtIkuswdceXBoxQeteHHk3/BkgCaBwcOEZVxRRx1P9ygYNW4hM7UfVyqqjI3
fweSabB2JzRZDsnZKQVAkT+0PNZItA9TUEi0DVyyrzdgqmxQF8RuA9EoelE1TeHK
dsXNWg4dPvGX6xNSzgrRuj1tiUX4x1rquHOf7ZPP8zs=
`protect END_PROTECTED
