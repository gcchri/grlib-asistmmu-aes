`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/e2IdA8ZioHHdXhfIVhHKcV6UvIBz+TZrUH+4JMl6YsyDncc6tSUcuiTT8+XHvG2
aJ49RHmhbfTZPPe1nGPfM9vnAPf3e4dnHvv5M0tXKx+HoLJKKVKpEPU7SmvfWD+s
EkRw84phMSf8AKyzyESYTTEhIQtT8rbqIRAGLEf7x3+RgiHAY6rwV5SnC1lNdiXI
0cfRFf39X6k3Ft86CVvJP2Drm+5K32P9K0DnwSIKtGi8S2aj1G7NaAkFOp0wKTBs
pBZw37drtPyTCLuwYU4gRFVd2Op9wIBmofki3mpnQow=
`protect END_PROTECTED
