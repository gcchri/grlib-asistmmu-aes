`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fOoXCreJYXclDLLmORChnFotT9y/o2dmhtzy/m9K6F9G0eLP9fN/2zUPJDVXvQTV
vsOpRh9NQs2IdhlpWE+lbfHwhU44KsuLBMWOiKj8oM4pXmUi4jwIXXV0QIrhfKtE
el2CCE13/MwXpfhJGFa7JVGOMTOc/PwNTSmgbLiyUbUCIXay52UBnuIeO+FKZYjY
EB/N3S8eg3atqzZpc6gACt5crtlaEPgus119nUtATbawzIxDPBNWOlYxRajC+JD0
+OJirS31SR4hzR+nIwNaluYweCpyH8tsCNFHy6PxT01mSGUkdUJ16W+6MgMHJyDp
bCWoi6nPvfZOoTb0VIQQP1j+bOw+RDRiRyXtKlNLduNlJ8IQfwkmhS9f3USSkkuK
`protect END_PROTECTED
