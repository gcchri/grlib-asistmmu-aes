`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rOUJGtZms0fJtZb9PhpSdXv/o8ZZ7Njb7VHiE7UTK4F4i52nsrOddmt48KF6gzNt
8WYj/W3/7H0XQqsYPfsPHwurkXiv5xRY1JXI/5iTtgKU5135YqzcuWu2di25mLnU
xJyRU1u/VwyXOUBi8ya+2x5HZfoP4fQOTYN95j9TgipIdh3OYkGwkhp89ERlKZll
5vFFsfac48KR+/S6+NgoTALNI8fHpsqAuGwppNYVTNvrX+GZNJjawy+ia78Gt5BC
iASPXVoQ+or0WTrwA0VUXkWyLO7w+kATrH3K/mh4/f/MJOUCcYy/A7PUDfrpYZq6
lf4CsFq0vwn80EShIySgLSUmDk5NmWqxacJykM9qGTPcieAghj/u8LOhOdKxzLxY
FnL35HEy/4otrWZjJX2dmiNtpx23xZh4zgbdne4alZMOCbagg/Y1vCTSrQobHKpA
UH6pCY7jzVGxzM6qwDT1icz3SrfYQq4ISRG+nDh31NE17ibE2X+c2H+iGuJ0htwR
vSNQ2QNUg7Rhml/uSeF7iKczGfQdt19htnUpVnfVNXJ30kWk7j5+/L5/Rwthv7g+
irHwb85Q/LCxq9erXm8DRGYf7yUWX0n6VxBFicSkTsRloxgjt/eePBjv/+hEQsxu
aIap3/vuOwoohW3XEtjGxs8GtG3ptjlkM2ujexjQJotmfVD8e0+5vpWFFPnPBQz3
Y8rBWzMmkVs1nBEjhCYtaTFSNZfIlO9Ty637ZtrVKPCQvWYFUXlgcbGk3Kugyxgp
SVzFm6ll4ZlUlabIJP5NNEm4XQGfsAwaV7h8hGobQbFnp6psYf503cuFnrn9ygWO
64Xgd+z/DxBnU8aFxdeMtf26v2kepS3kJqRTyMN5kqhYX998tt8QBzWhFxrV57B2
`protect END_PROTECTED
