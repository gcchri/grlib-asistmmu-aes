`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DHDPBCIz4PM6G24CcyCsZ0jrHkFP4GNAj11Mq6Ae9LVvJtql1WArI0KIOP8mAMQA
ezpQMlj8I/gKMvlvWz8e0d+lzRJPdcvREvWs13vtPHBD5xjTCAK90YEP0iVNtsyI
0SNqe0U08MJDukCCCSyqFAfHgnk9cNJpxgb8Ki9io16apXLH9O6eBhPblRj3bvOU
QZ8KgdW7wSc86BmDkPjkpwbGUTJjaDJJt/ycPq2ktfzbdRHF8BLH4rzyKXE9txkD
PujQE9wSu9tZDB+G//d1jtgzSLJp95PaVoR/YXejyCX4kHJid8uetxAgi+xswxYZ
natqWbQtfHgV9vsdXHD24hNskDlHWVUk75uWMHAsMBBv01S337uTA7dRlXRzWCu/
JCdxXwkhBsJYYE2E4XJIUSSusXdfhXVU8zjc+AXAeVRCULDx+BzONSeKIVxJOBVk
y6ICyFx70eCY6BlAGDQ8+dWiCJBzxEfodvV90ygtjgThu8W++WyTu1j0TprvqKKJ
vXngDY5SL7wOwaRvOz9fQZhTmvBOgpKV5AsnjMQ6D3hn0t1PwTYe4L/uHNfWMgdK
d+8A7T1ZlnTZPdfKGUsK+vYo/n7jsfpPXV4PLe1EoffLYd0AA1NRt0ERYnHo1hnT
`protect END_PROTECTED
