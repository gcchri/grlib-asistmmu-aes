`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MB6SE8ybYXwaFluZLjHJFFErcP1YPO7XgWkc6sCnou8lJG4m8pYdz6WWNuVPUPIe
ojrBoHLcPgcLURXzoWsgnUXdrkszEUpbL4FJSknoA4oATV2sOksXlXnp6nBmBa6Y
vET1ysyGraFwgJzYIKklag+Mi7EXYzwN3CSlKddGy0o9hd/RpUSZ0aybJNWox8xE
Vze7HlE//mnC6tN6uY7bg2NC8GYgkUdExwYzEungaVNlgV53znmUz3avqtsbfRSC
/vZ6MxlzrZ94dSwMInjlpk7nw7ul0m+4SMh4eGah6qZeWZgLp13J0e6ktNUBF7Pl
pUy7aneDShQk+7a74RctLg==
`protect END_PROTECTED
