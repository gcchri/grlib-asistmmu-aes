`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2hZXZuamYsWr0Mih2DMW8ypDByJM9sUqvLCHMbKzd4b/Tfk1LcIPpOqdFWUgjIFo
KlE3sU/h5cdbgBaRZlzDdLEV4RLxHMro/4gk6BCBSWe+ks9z57SpG+8SWe0NeX9q
aI5lOX1sVuQPMQjkDAFoIE2m5V5IXe7DJAQtTYpZhmz8STof9RXF55QBaJK1PJRh
CIDo+Xz1GhR5XoDnNhQY/EWBhVDMDlyNG4U+2ijlFtQ6A712awtYKuqwizOcbVpt
YXohE+0n7OY7lQ6tGGPISmiH3No1mhQkDgsjcuuKp2BColFOHKgXFReMa7YJ0pYN
NbdCcQR6JKLixPP1KdcQwOYIZ4nR0+tH/FmUkLJ2nVYC5JgnN8RcbCbSK8kGP41c
5NHkmu0OdQgkuI5m+QdBM5DEW379F4g7N9dtW0r1GaOBp8+jZYzTimgM/6DL+xMx
pQt1Xn+eI0DpnEb13UqxKZE1x/EIVvnQ1bH8xuWSKmTeaHmRyKIgx5CFivAKUpid
h+4oHCylmDIiQ7qeNPdyhDirKwNGUcA1IgUZ9ziOpt9e5V0Jj2/4BSViE0TSLM6Q
d96xhuwyccqnMUNu6IcmC3T6dhEZbfYmj9jwXOe1znNKiifVVNDCrxzZMcaLaT0H
sJWf3UXXx62eSvrFAahJIMLOD/myE9cc+dQeUYXs25ZHWdJ4RPuD1d1huTVEfcqP
8qTqCCjOsGO3207LFzTuxKPSr8vP17LhhZVyGRSiyxQykvDqtBGfAdpYsQYCx2Vz
19Ln3cNzWo5B+36W9iTaD9TcDk0ud4fxMFjzZ7VFw1uosXUUP5jYlysPtPnDWs+K
wOdO3POQ8GaCoswZRq/u8yNAAXaOcMOHfR9VA+aRwSu/4CG/3OXpXDiHYYcIowE5
ILw71PG7s9KsVMRW4oCqC+jUiE2ELTQftjkHzX3IHucbdWqs+5YbRDbtetF9wuzT
n0x7p/jXI6EpxfrDmqMbg0Se9i0vEVgPFJguUbHPUZH1bNdqNKZQCUPVIgaEreR3
zSO2jig15aMomRvLrHHi1mQkwEDnyp87E7IjsSaAdW9A6tcWvEBLVea6EOPJA+os
/rM4nFGo6kT5dQ7z8yyIjlUpjyMWZoVQA5Nw1xHYE4taL3j6a9Yra2IegaXRBxvg
PLN0A22tYx9WcUdcdKjTgXaqHXgiU4L6PZljDAWw/fUrlLUb4VUmGQrlyErzF7jp
itlZDe+0c5raltJ8kRi80AJEJ1GgqV0g9rjGmAzWXh+lWAn/2O4oDc/VwtMk4DL3
R/mnyBZmeEkXtonCGGSEV0c95Pb6R9aanEosBFhSbOqOp7ry/WxnfiGPOH0EDC5b
gmoA335EH2VHQlFetBqEHGL3jYXXr9lEEEb5TzPeFNVjER1L93MXHMEapbaJP5kp
wqWOJhpxqXXIHzMuqTDWgqJnyjjVrBXhkxE3QCrKGpSTh0Uwx7Sc+OEZmnVX65Hh
tN3LBlWX/oyIOm20GZGY3+9Z6VkU6GMtkdV16bBDOpfb3O4WGu+LW5ZM0CQJRq8L
TuXjFGseibe/AtFQnPUH7aMc0+3Qxveb6g7PX4IlqgTHi47iRLL8XpkZ+o6VTliD
7Rh9eo3Az3xJceCzUg9yLyT2xUbzEtCDBOOsS0Vqd+x6LyySookX1bgyZLuCHQJH
r96dNMaIh2Q/QIU8FkKDDxUa7NOLfR4jfm3XmjLz7kGgFfC5lYErX9sF4MBHGZqn
8Ig/IFpJpzNNR2BWMiTFPt210M2P+5sIAZC/oiY15jmy26WwRUX2IKQG/Hw2naWr
emb6A5RY2XzugoTXdCbwOuiVdeTFvk7CyIQKiCsfNV0L7ZbqRZCYXmrZxh765EEm
MKc1MU/KT+yKXxkBlllU1DGirdZ6m97SYTI7CzxvbZZXhPLViRrMK0nAzEueNUph
yBkwNf4b8qzKBG36uFsPQTFJfx72hT8FhlO9SbOpsky5HmowYs6HSSZImxeT2c1T
z4NOItWwt/Qf0xqh19fMW48KdEMIK76uNCszsNCTG3JXbTnT6JzjoKXrG1FtpuWn
/Uq012MwYy6+4RLGDodwwIOk1mmO79kGO24LF5KuKhDnmc686mB8PyMqhshtSzC/
K/To3Gf+HoxyaYT5aIEyWYrKuZKQuG+cIrCNry5ngbW/++WEJ6KlSUF29UZGWnpT
rmjQFi+39Ai29UDkYepATpy9uYzXZ5NmpQKsbJnpRoKTU47ApoHx4mcwK1ULB/5n
DiiXJnJnYodZzpX4GQdwcfRarechZGjlDMo0nd7XGNLqiPojc8I8iIYjdqs2BjQm
IOuJNtWWhlPOgxFPYXoL6FGOYYaHs+CJtYCB/HEI/hZa9VZ9NUJckt6ED2p2Gm3C
Jw20IAOGs18ExGW52Vn+F5Z1VHXSuMQBMg1imoLE2j7M9xbvgF4OGtUdPsxpHALS
yX7euYUStsEj7z7doAaOnAgjbhhy6ieG5HgUDAOpkhMPb1e5NbCDdHi/8I3I1FRc
cKiBpNjbUYL8FmNK6x0tWhjsGbYaeWBa0Bg9XNMPfnwdul+hW1SBwWfyrnFgYUst
TeOfx7NXQORnOxbWC4hHBrt/Lrum/diFw1qWyG+Sb28R/hrLdkgSG20l6gu17ozQ
qKRTt27gEZwtfIfKJzF8UDOlRJALyxpHTKGZIbEPVEbGQTTFA2RM1XVs083/3ZGI
5E4P/iiMm9xRpr+fodugolMzXY3DFzUxHbnw2UV3t9pBG6G4MgxyzbsgRS29hPRB
yACTevy6BCzeltwiY0CW9Mc+NSV3pveG7x1/Sis3UtopCletKdlfWKqfs2CSP9wo
UDaaMsvCBW06Dmh1a3Ps8xmDwB0ZUECphr/Lkvl6+LFGXfL/9N7815rNYcEOAFrF
juKaNRiPMNjOMfWnr/Uqkqq+vhpEkg3ldc5Agqu+CiNgnS2humy5Z8ebWcGARyKk
qM+mk44UEIdlEcddzcGq/W+o72wbqwdutYTEgRZ3xfHlt+DT2kqs+W92EBAbj8ln
nIzbxw4W2Vb0rRv1RH4wfWOjer+uQLNJ11vO+zcb/SRKWWpBeoJ+eCyHC631nOt3
/woxC08+qmuqhJahlr9zwLJxtpdxpA9WlA6AfufIILWSymZMIuFmd2D1aLn+5845
`protect END_PROTECTED
