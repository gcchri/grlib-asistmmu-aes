`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vEUISeszowt1KcX7qH890v9TBRRuij/hOGpUKoaez8ut0fMW1wyz/BQh6ue9MLbu
FkAmjnw3vrB8zG+PlXkdH+IDfMy5v8CTQnXUP984G8TnqnpJ4YGyeR7I/WF0hp7I
4Von3tBkCZJMR+CAcf/U+79FJH0wop6Kib0a1v6SPHHBmIrHBRlgmJTIvaiBx8cj
JIHS7rqbbXrYZ6I6ASQL/7KlBQkcl9c5+PozYScpWZ86lRWvHp/XPk/9Lw+TMNoq
6nK0Gl4zZxHcDx26CRTRkIlvIf++zUHBw/qOaVDu9S6cp63twpP0cFILu8HecbrK
IuCHUIaaEUGyNgzEgpy4DA==
`protect END_PROTECTED
