`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ihH75LZtXIuORH9l7WBcd2U9f0nPn5DROpKEjHW8IyFDRSZMkvmo7U9T5rU4X+Bf
QQYOiPLZtzydmq1MNwhTrvgBQ+o2eAJc735p1nVGBfIpKQOZsfU79nXVJhSI5u+K
+x81+gf5/i3DH08JrPPbWmFhjMi5VAe7FjYy5E+uyKOHQA7obYxiWPALIw3CjfXl
fQ9q/eodOuO64aNmsh+otSnUvcN16QXBy2KvEoPGUxYESA+ofq2CgSyfSw+NfeKu
jjrmiO7neyBMSgt2U9kPxVsxLfKDM/2DfW7PDueGBXV8GBGL6v+AD9q7OCNQS6po
Nl2DU6b/ex/btHKi/EWYAM+1vA5kFvGN3qFojI+HLqMb9vs8X1BSgy17dK3DupRG
fM8ENbbbqbNZB73Ldq7QIrJLyym92RbtxW9/9c5bnwiuHn0eUSF/F2Zb8npG3dX9
aUu6XaEXwdcxyrpuzJSqTktOqwuvWzh6gZPzeWEwRgamN6ibdCEAdMMNisf8S5Im
r2af9KZEtOqtTO1uMpAtaFfSDZe4AkUux9WBvJwjbN1ivk3FV5Wo8NHLRnU5P9Vc
7jW+4w+1TmG0hu0uYpNUxt9jhz7NY52aFZrwTgMTM0Y=
`protect END_PROTECTED
