`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2vfdREJPOTw6sAOF+6aPni10lzO1ljyHo0rF3ZUzIWoFZ7HvpjxtZSZ50EzlY3xQ
JZNN6gzwz2SQP++QvGa4qLc5DBO7AxyNLFuB0Vf2tkOsCRl6WoGko/7GqVGgUIlz
5upwJCzO+q+PMV2p2sfvmPfm0tuMfZnHrTA85LMQ8uYYQx51Tw8Jobf3p54Kqr3U
O1RpVUP/2j2sPXyXGtBFegMdlojPRqwxrlFZFB2c7IhQRQL56Jw5rMPGA8dH2JXg
O53HCH+/QKHNCOgn06aT7x6b+2G2BZH4RsykzEDKjJy9In/VaGSoIgn5QITfLzfG
f8qI3Hv3MVRX1W8M5DLnkidd14iuhrYwvMMRa0MfWYyAuwgfoTzEXLBLLqWBHFEe
b8EZgW+sCWkfc5Y9tqOsb+FQRtvGePO5YUGsoN6noLYWV0XDxPoILaZfj9ptKNXy
KHpZGXB6aIi1p+EClMdw2JX52ueyMoipxkDV2xGl8VTxVSkWRXYwSJj56b+Fbyw/
teNSIKGsbsmgfpS+jwvffjBCmhsikp3vbpNQ8Md8fHK4oBhDtZgEn91xDaoTZwg7
FhIcSlv5M88dZvQz1ihhzNm2O3wQue/ubxOv7FJ32h3YwMd1Xn42wnQrasNhBiIR
N5QZQS/+UHfOcX2vn7VqkQ==
`protect END_PROTECTED
