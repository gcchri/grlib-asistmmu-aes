`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LiFXtXmFBxEuIKL39IunKdL0OHgEZrawojgrpEFIY7H4yR9tszDe0I6mYY1euKi/
AtsWbysH6cH9M6dn4WFHNgjrQOu6ZZOpDCz+J+tm+atahpvG2zrLHW8vd8C4KUZF
oiHpETlGjzE5VCiE1/wkkuT+U5VL3t6+e2NQBVnpPPo0xUKSpYnrH1/9X//HbVCn
rFbkiLQMCDLgGoRYDxCNqDJ4oEzAZApKM0CPcmBclWq5vbiI/FE3ATEP+tY3Eyy2
BKJgBE/0t3D1jjj16oqjmz4kSgHqpTkbaH/LIXw0T1TfqA7Zvujy6qcD4DessWih
x250Ep5mkivpBrZ/qvDZM0FK+Gby2ujn9O9qb5D8B7zq9YOkBkPRCTtKPXbEIcub
mm+w8zCQPu6ZFL8jiiEVNg==
`protect END_PROTECTED
