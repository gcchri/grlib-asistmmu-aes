`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oaB0kxsCWjDbFcTXCt0Yufhgj9d4SXJbdw35XfjeZtrFk2Cr7BSTMJx6MU84dAGw
v/nfp3jljDsH3AiNrgmMVfNgfdCA0k5CJUN4zLLG5XcaYd/SQBQ97k/8dpReFFxA
Msbk4DApK5k5YU2034DAE4LHJQdChHAvhb4znY6lzh93eGFTMNhkAwMrb8yu6Hkf
Ob/Rkyl7GY1WYifo0EW26DilFK4Cw0m+T4yFYNHxLFZj4UhpW/IgC5blKkVNIZaU
B43DXCo2LK9oC576WF2TTXuk3VStybIoerEvAsOZ4icxL4bmAgLhKDnqbnzdKf+R
VBD74eyo8RMVtF4dee6nE4YamgyWK7+NzXpF7c8/4poksnhTN76XJTcDNQc9WXXG
ecipdN2ioZMR4OVFVM3Uo9Pyis5HrxIP4iKdWZNCyBpK8NwgY9wp/ebbF/ukf+hb
mAhyRLgNYrMypAeNA98T7JfQNpUBGh96ROkiomHg5/P5Ad8bzMjk4t5wm3tRPHG/
/F+49KMt24ZpaNhCKCrfqriqDe8IuWzk66loMwgkemSafnm0ZKy/Bc5DSOn8ZBdl
uR9CbaIwjLNVWLemD1lDI/8QH7juiPNeWPhx+/ek+HW3CP4rn/W08OJ4ha8izhNo
zhPUnmO7VtdcFf634BBk5obkeaw7tKgjEiYs5tZeA1JPHfan7dT8y4Jp/YfZZ1+E
LSMmO/Fy1cOWuo4DOytXMJNlB9xqE+SsJPO/OvCmGWYWmwaQg0Ql4wFQfmBa4A3J
ixxTL/gChf6d79u04M+Rtm7WYeYAmBDJcnXtHW/YEj9HvJgIoV0xNZb2j0UNemGB
qjzqy7eDQTV8lw9MGH39pikvmJWGvVqxr5Lg8xcxNhZBhRK/vAqRWIJRH885d2SQ
6ZzHjuK0B6tW/fUiDq/alvhe5bkuzEbPf6K1jQ+7SONXdLil3XSdwcpsd7sDbngv
cTEsTvZ3fkLTzeO3GCfj66hLADgOW29hGu0GGoJtZXcsH5PlojWhOaF6qJEJLxYi
smiNN3WXq+uJAwdyoHgkeCd18aAwqN4T1s3OTbLSuGxHtuFCx58cGG2yQirstS0T
s5iLqfz/IOGXw7sL1VljlvqN/pKWXT5RTGFPS7m/15IxcQqI83nQ345VM7k/KxEE
QHpzCYwbcbXgwkgXHZBn5FFvigUs5CjoqAEiWsU0FeOiSC9sZcP+sg6GAmtLnMAU
3Gl4aTl9k5ly+taEohansU/Jei3SPInzsOZaP+eIYhYcGvTTD+3asnM3ObnROfB+
+Kn6n7ecDUPYgDNOwXyX08OCrU35WsR3Tv+ckos3iL1/MA7zx1JqakcGb68ixvsl
0AQhTIzAolGGdWfFpuGRGj4y8HznLu4IBLWZTGYY6g8tCOnKK1yxIuT8LrwaMW/l
ui2uX8FM7U3ifE6xH/X4C0DpjfdhrQZEcFvxBS54QywzuKhA9bYqldKpOi9H1FgW
36qcG89GiXj641d56KnlFc0ndkyu92xwFSIUWDSjsJJmpx5m2e+urRjNpeet/hW7
QqyESzJ9HNp2WzVph0bXgIr1GYYXctTeOIbGrNLlCbeYAzcfJEQYxmS2EGuzCX0m
IFLCtbrGN6uPjN4ZThlNVVHk7ougmXbqHLaMnMEUp+xpOfnA+YgTDV+GovH7pUwK
wft7imkBF4U6Y3Wh+1YTGI/gWikOT0DTKXu+/LhW+KjhZhaKPRB9n+6W2KdaytKe
fMu/8I6HDjKiRFFCxZGuePDZ3NRSmpGE3tg+J8pQleYE2Bw0aYw+d2ZvLATW0zO7
jGzse8L5ft1sKWp8ozNKWmAe5T4JTrnG3JdjHf6RwWdcFyQohZ0F/vMOKLYhQwwm
cT0gGo6u0IWPuR4zvOT5Jf4DcjFICQBJKkNmFSqDewPT9FCeMxUoYeQyLVK0IXVe
XEersa6t65b2X3gFyO9cA0kEB07J+o/YdtbuJaBDSbijCAOLtKyQ2SV0WfWyVjJL
fLck+tWETHCHuTRWkuXkM08doOsVxRqBFKVdBAEbG+2UzG4ne+9T1d7EoItpPjOp
BjUbByYCKN6mtgIF6m2uBreIuuexlBhuW4NJ0YUQ/FXvt/1t/VDL3bNCNLqifZcb
tPeuggRgAec8KcX0NLh2FZm6c9msRK9kxIFfPuuU+bb90v7n0Fa9X1flVU0SjGEV
zSDAL5oxQEvV8b0okohc/Z9VppZiU97y1sO/ATSXhWRR85YBu4KyGlHSdYuIEfyW
SeVZcR3R2gb1rAWVXHBKHWz1I6jyovOUNLlEx9V/Xmf0jm464R5RERpuclM1ndbg
mEm1zhGwB+uszjjmKt/65e8+w5D0q/u1vi6taywf25y2GvrdFMt/w7YwzwX1yJKq
W6iSWvZfHw8Ln8mYwvQwoOdgMMaGsDxMjzeDWbgN3bGNbcbQ2KmZ73H2V08I3LPl
4ATcWgUVGBGiaId1Zl3qzvw7uxOfyES6byElUHMO83+vpu1xV4fyv6xVl0KguTRr
QJfUFxWL9bcQtPNVISFyrJXCmNtUnktTDs57e19e6fA5VYNTgIV4tL1xejtnMIN2
Gzu3RuGu+9aJwoHXe+rhx2KZcPllHHQ/sTwxTBA6TT0i/id+walno8wSQQGaCDRl
FhBLz7kRFSc5QB6jVn7G2jYiVJ5c8yqNpOCv0pQEjuq6+yGHoev4PCgtKLIu66DI
1rsyp7LPl3aK89QWCorkzWSbExxnKjI/QdbxMEt7+l/um0uidCUhADY4ghai/QwJ
0mMT61XGInLRJW9lLOpLzhwEtTle0uiPUNi/dq8JdTyNt1CBpFAY44Hmyq2F3YZE
KW24uNoZEUJmZ1kAv+XVBDKNVeowCaC5Ay/Sj3WbLcmDV2VQmQm92k9yfbKnyydi
5vPkpFR1PBQMJ/ApRHVY7JPxYKTVtIJunFr4sEN0DMsBxAPsscCjuMYhda8GkzG0
rkaW68QeP9rga90kBShTxbxGr2n3nRxeBZup4k1TWtrO7OONbSGbun9cbM4wAspf
YtazDTUtj70Uvken5y0hZGLrxgZZI3deAhKKTV+z1MDnxSfoEe5YBUW/5uLHTvSu
gUOlrds/99csBQ+Wy75CSyL7YGuGfRScSRX1TWk7E/z2uSlVE69hw1H4n4ErSRj/
laxs9AaEq5Rxq9iuvpCKbiJxuaT8v8xQ5Tm5Pj5n7/goL+21auPkL6xbypBF261D
mJGo7DgsGmAaptwfMJOWSzBzuElOyeHb2XtryF6TbkkY8EVcNYm2UlOp1jFZgO4n
Kx+MztrRTMQqbqRTCPzXmc8XQUo0lG9mxAePL3fPzWPeWI3PsT37Huwp5aWH2d1Q
FyheXZjXmiD3nChhV2znt+Wp21BHYqR9ljWyLR66WyqxHUzLKMAAxZr84EKf0KYx
lb2KwYl+BTD570PRsDcLgqMzlxfa+zy3nFp3uQcQxlBugdC2wcmUnJoDizrngPuk
/h87iBIL1vOpYFNy6q1PK8qUWOEtC8MwE2Cv3q6obZRGoN3BYB/8ALYjCw5z7mgb
VflCjvy12OKt16G4yAP9tMrDZLRoN2TzT+698T/6JYOZYrfvdNlkQaxgO1MoamFG
kD0fbtXry/BUGOmwSNv8IcXH2RGw3yWor8L2WuLGlmLyuPvj37i7+Dc8j28rN0c8
3H1A5wfUloDro1JjeyWqiEjCLtBv22GGXg1N6nrY0XidMGawZbgs5b/0Gpu4fZ7Z
9oX2K6pMSep1m9Sfl77Y4H402DXkJukH9nrx/l5ixJQ/LNeO/wJD3v4syDMuZBKE
W1PqiNsLfI+0gjJYHf4rKs63pcFs4z+flpaUmJrziXT4WD5Zqz5HETIqB9BsIsCM
BU5UZ2l25EfT+SJP+q2GE8MOOIMCsSyDCmIC5IqQXt046nvlCE8Xi9u0VHcwPJWm
/7VV1sXySuGdnqACb0Ioi2NNIW5KvouWU+eG1oZWYyutg6D9VhfxHPCX6BCrodFN
9xI+rVeG/gZDK2w/DYGoTsfCLJY6F1swl6xJN/bolW4FdfKnXpJeI9mo/Qf4DICj
h0ee3JChjrL8/PnWsYe+m1ia3Zaj6uQvlr3hLRAJeoEJWsn4t4FbtdT1hOb7C0Il
5B5TA3smMGju9IbuntkAc7EmOlZOlMCXbYdUAhgLUhIuAOul2/tGhvYzMYjd3OwU
Y54nH0nLxl5AjcL7CAmU6c0u8lYJZXYf7DoXWOm1tWND0Kq0dUUBGuyFz8+//yj6
gFQIhyMVKeTXScmeD3SOEjL/Sn2pWP9OQnvqb/jr07McSFKBc1uJSP3I6Gdw5mpU
bMVTjpUohrPFdfQBnyOFuIS/KNY7CBkNW3q2BhhnWNO+Bj4DctHj2GWEyhkgCVkx
rybP/oN1o+uYaKEiBCmhbKYooiI3gjX2Wsx35kVMvOCmNR+aFsbkh0DOZ3gATjJp
JGuHGMn2HxkqbIE5XSmBoPP7CeYYAPiPhxILsdgGltcyMwdNcHH8kExJzgZmoNRu
R+175IpqnIiDU/LL75OmkjRiiuRdGrU4roesqD+S6cGvAxnSiuHOjA3q8IvAdg48
Bsa0q4xcdxO6AjvgAwNjHYChk2ij/fwpa2RttxTnSa0kIedco+2yVTtZqoQYxd5c
CFUgFUrw4YFcdO07qAIMYDf7MQSU5gE+v6OIq/sfgTVV2dYK3lfE8GdNysfeIAAj
Bsz3OmScTzcLeWjZfa2HiqzPnV/Oa1zDN5XnJOxYFNS/c/ZLPYVjTNRY30ya4231
gkERGB3VMBHwqXVzRpgnRIyC0SSE//fPFWB0jbA3FY4WhJZly2jcoRs+Vxa8QJPt
bbXAz34dLTa70bELUs1orXS/Niv73ylOkGkTgob40zuWStcrMNv2CQOzlWowU8cD
adhhVzi+zNQvTX0OR2wcOBtyV9SvRG1GWrgKYqACnWwKDvmxgTWzYPa+j3EIXSHZ
Oiv7TBdpPwAApKdm5y2CmoRdNmFZ0Z/Aw/VFpMZ42g1AkJ4L00huvA9w/jtvgyPv
3NOBN/0IeUnufUfPfGaPLx2ABOJTNXhLAfYMRSkR5KMjMWMdbTmjn9Jhn7OarOhU
CUxDO1q5pJhcb0CrjJAl5xx3yScmxOWIg4FMrmZuiUmwXDsDK67x+/sBpdsnXhzK
85T7PyCKzodqKsA7uxVzd6Yneev03WeNUg1FdDSYa+VdbvGw3nKkr27E5t+wj4So
FltvA/xBVGDLn5veKYhfP8VUUKQ93OIuZ52r9HGfUp3VhM/mtmdUNCoVnja974ib
xpLtNgxGFTrbXdC1RquEkuLtQQiF8inB+re70GIFcOsxToSDY54MEQX6GTFiTYK7
lM+1PHcEdhNXMuab/iaQGAVc9zFBCnjEQDjSU++VeRQgSt4UmeJC9Pr7xvR3CC1O
/YUQUSorRT/T0oxUjssk4pIap4JxJ+o6GkfWsHEAd9KgE2rEwetnZd5ptdChtEoX
RRiFAC4gk1s4goi74zRUfDytWpoEgJAOuf+70JJDpe+aAlThmaTxhNChcTzjWb+B
y0dZzb+3ihaQkRKyjq6aUX56j7eY5kD2xA48bHxvNt0cTcKiS2PQvjMUUFVFA2u1
iQ0Yz4tcwH2KVBjakLN2eAC/2mLYEdoD8RbP9J2Xzjs+X3zCnO92+qwT4qgjZk1T
OmwCsc5+XIRvxI/SDREWZdCsx3BTMwZpXRTRADMTdgAnqzjkHOKcSviElWQR0+uG
k+qWpAQqaR/0wlkhEWUH1BUp5hwG2GtE+v9j2tHgNhUAHcUfbT6gd1rAd2JL0RJo
Rr1WI9UqVsH5pOAFIRxzQ/v2kpLp0a+2IoFavsz3l3kYdbP4ZYFWc3nBLb62pvvF
Qj71SMDwxoRoG1l/KeI5Lh84jrpTaa67cjGWeIythfsTm0szI1ipw520+aPm35Vf
tzKtFULmvjxvPSQc690M2qtXn2NDL/HSJ8D86l/mzYZhFF+mVuzUmQ9ZZuF9PVdX
NMSQyypLO32HiaLxIjOIVzqmADdLdS7Jh+0GKjLOsyKL8wDgfLF/AIxOJdoS9RIb
yLL231cHUcn9tl/DXwD2MEwdtdot7LDPELKGHD84ORRZ7z0/dcjz/cWSn3PtLoX5
xeZjzTxNdJ+ge2Wwdy+QxYpkAx8Lyu+/oGMKywuICwVo952Q+Y4FhQH8fPC7Rfs9
FzvUzolAi0600MxmxzFbG55lW2762r7aAHKHqMjIrzfT4U81i7uJcELtGPttjFsC
8Rt7OacmykZgEx5jSjaYqLDEfyk6e6XINgg1tJ/X+fkFG/EE7NNtByd6bYIfT71M
cQT963LbqXI8GjhP9k7+9JaJyX9bTWpcXfxnynFmfSl3k/5o0dyRlJkxbeGRqk8p
map3VYs7NF6gMZEZg5bv9IKpfGvh1Pa3ly3C4F4A5RDZe5lug4hKKlwJVrxHWDTQ
VvMhzW5pVB7gHMBF7eu2/x8ihgHIMW6NoP29yCqzvySbYgDPCjYRM9ZP/EPHJRLQ
X/XO/yxauMFR71g877QACXD3Gdpsa9Apj1CombDRdeDEMqPBe/CQsRKWsD2NDvN7
Wb7K4zfO0tkOzrvYuD58azjkvUkBVbkmVkM+YVXeZTgq7957Wj/uwIBhfgRJ9g31
SosyPts4p9vzshJ4byDs3z+4G7afzfWZl1Zxbr6MNbE7+W0wfuMtnoKI8C0MW9Q7
Vg1yeeoVI+emG6WIqOfClKhFU2M3ik46uzUMH1Orqjpa/HZCkvyKxvs5CVKKFmyB
B6RgH2qZSQfOjoSAMj6P3QZqDWKDqzAlCSWpByjcYaCj+aAik/e6VvZKuNyi+lqd
q6s2PJVD/cPr40fvRRoF1W1pqJtdfUK0DDJlnC/DiWigT57iOSiBpCaB166WrO2v
BeaO9080y3WeSQt1QZ/NGAJlbZ6VB79l+n9H2JaVjTVivoQLGIl48gy1s2WCmMIA
MR/8ren5nwfGxeLhcvJBlddPT0RSHtJhXn7+tmgdFqOcL3bW9TlWqO6S6t+vsrv4
0w/LCeWYecjcNNrXHvPBzuLuNJzwUp/cakgig0V+O2qgZ6WeuIwmRPVOXkpyaajb
+3dvGJ2qHeMLX3fN7jq+lF9Xgzh2LrNUYl3xlfVM61JkCVaY5WIkHrqO09t0pdP7
77qfTB5sv4kRK0TbQtS+xd2mQcxC6kWw/neTKFMF6yGiv/PhweXGTdU0tIBIE7X7
L6iUUOlMysTKbUnwdmT2khwx89fuAGPtzv8hAJeyr2pScOqSvBBLAMubHNGSabss
TcxFvsf4gCAo19jLxliAniFJ/iIVGZf+3xI0i6SgAupRy6xhKhLA7z8fNibTYFIS
8Y4OROj+hiHJ+ZntMxffXbYO03jzWDRaJyi5r+xLi78yanM3d8+lcGD4Dlk6IsFG
gJgtFi5gKDRcaWko1uobig/CemcmXB2JimK0gHE67U3FqiG5it+ooUUl84azozAK
fma/fzgjaGZDKjRuT6UOmwQGIvnfqJTlN8dNcJqza1HuwZ4Ubm0j/+TzLlskCcHA
5bUydtB8mzyioXhbNf6fivHzf3x8tOC3sbVLbJu7MttLld2cVhqIr4+uF30gtjt6
5DUhZRnXuBV6u0vdYYgPYyzGio9/DrJGHTu9gHxenI7/kYJJPVpK/qVUn3TsQuzA
/scWAY+aK8fs6iMnmI0ftjTNQR26YOwMxB2gj5wyZ3PQuk1ZfAMggVJ7bh1ldywz
mUJfmhikzxMNBHkLtbYWpvIfVpqFS607kKDY0SvRFOO7e33MOaHcns/dYcOKzgiZ
EjCC7eX9cjD4nARS4RIlcWnIwOkOHSLs6kecYabkTFmQRDN652AZaXayK8uMng57
nLQJyAYX0zvpSdz/TgsBsuGvLW3x7Ytx+ZBb7w/24/x9nnCK1OWMLlod75dfxB4M
Q5WpC5p2qPqrHraPESYqbY9dLK1bUHGbDYvahPZArtTrL/S1lmQBdF4mALFXpc4k
Wxr+PiLsacvFnx6Pxvu2ABJg32PmzYX/iFJ+YGLCNn62rmEkQU675b7N6HH3qJFb
YToW0vsbn4Di/A8PZMgdD7cQdeieTxLDjxQiwCjgKGokrDUzZSXZ5jfVhW+QYH8m
kpRQerzqkgVFtM/zcaBiNqE76iWv6+vLDRF6igMK7f9nlhr1RAZDRkKbrUC3em2U
UQNcR3SPRD61WTG29pSeZV6L45U++T0WcLSXddo/WdR0qcMfXbMSs1LX10JD5LUy
RE/rNkF1zh20vAlylYUdtJVu8NnRAL9zFwWemc9LyBZz6G09NFMBmv59bK87bM4f
bzQmBdY3vrpaaceZxmtGEtX/eJ+zVZGkHEz9ZJyLcf96VLU5/+H3SIcK/UNqJCtJ
Jx5pg3DRiB6ZGvavgeWeZbaBN0rw5PLJmppWurPkJqQIl1Y06KChAYqrZn1ZyzsX
ym41E2vYzd7sj9i+0b1yfO38QCy5U25VXrPyFxEB5k6cfK7wvAaMD3YbJNdM0d8h
hKeisxfxokb2Ov0CjxPZXwzT9OjOfjHqlUHQTepjixg6KYJ7FOwWOgoo+Y34aTjb
WduYnOV8lLFEj2ItS0OuupEy/EL4183cMyXIE+30K89yfPXzy5J06Took6lQ2vZS
RQSftcH9So9wYeTpY+jdfl6U4XSHaGZr75uCpkWZWpLwtYeQozgxP6GYl/X9N5JM
OBxRACKHp0th83AGBHJwt5Fvwipkbsj8lYPX06n1Pa5iQeCUt5LVS/YonkUuomjT
KENg/Q2HDUNI+3VS2KCqt+oHLykCj111GMlxiq+d9TUOIwKEyvzOKuM7I+ue1zKV
ayrZo/IU8xuzyxAzG7bBhRjzVh0coANSQFNKYM8hpY2GMzhDwX2glr2wAMo0N+d5
s4zKM5fRR0VILbH0igpdJshgTUosivt1sOWNmm5kwJT5wMLPvap907b5XRvTxHtf
P+u1nWfxqMD8C84TquM7o5Pm0pTaqbyF6dYSqR8tukb6cunMhh0362IPryWtUkVZ
I9Hh0OgDIBYXDicNjVcKQYGsmxdCx7GGZmA26oE6q8iWEUdOvJjA4ghQKW6sJCBq
pa/k5F4ltYK4J0/IYOWOBC5KrJKLpjlf6zDUXzDU8Tk4rEYsksPYHF3vnIRiY89W
WKMrLnx+1jftX29NHEkWGaPJ8P1weE9S1HARy6ivFfS+KKFEJcLKq94eeT/9mbko
4cOctf69CyiVoef8QsrA5k28wT67d8uYrn36cwQB+kL4ZhxHojBLekncUJ+GntqF
ul9tTBB9as4L4pGkrGT63A/lD+dUe58FZ1ghf0lxODGnizxmf7C9RTbikgXNAus1
AGECkZ9XTCPoxAXGpVgwJCHFfFvsJT77eOYPMJlrQi7n6OOe7IZUdnK0QJVUsChz
6NHoLLuXTNWujU+i50OzTKtR1PBuN39Zd7NX+rhRYyuoF+HEedH95Vjifo9zod1h
qqdrgkryMdL+BZ7sqVorCLszJE5OrKYmrO0zh+5cD4qcFVfEXQup+KE9ELct1CT1
KbVzBNL+LdSnOovy5fzvw4wBi3xhYJLt/GsonvYAmCBggrJkhokOoviOxG1fT7oR
yiQwUoXd5fiRgEGHFRlj+u456/BhJfI07McJVErQvzK5mQgFQle0td37N2aefY3n
rLZ969PCqlS5ciJCt7KK6re3sU32yxeUrANBX5cXbI7AiBqpZ4CFiTx9BLFpWzr3
ExCRmS5XJncSXuOVyrHDglW05sYqnGlCjEWHHllzWiWnAYMGCm1SzipJ18LTHlN5
CKU5I8fZueJGhGZB230iU8AIseZHWiR4ZnVPp+mBXdNBf6y3UAJzSArBDzqDfRAX
kPTU7czJJXQQVZYJiL0ilNkjXwS78uH/gOQJXtF7Tg6yVjVJOO4nkkMPEo3FT09n
mNdwKYarIl4kJlA3Wl0v1Id1/xGtthzEysvSMin6HrThvSIeIkZ1u7i0vpoGy72H
pw0FX5P08u/b/JfYyPY9767Dw0sfxP8frs9WAjgzQKLoAD8ORo0Pl/EpHvzrt+Nk
k+hP7+jK3bgTMaye5B1gTEluEgmQqhrEppfKNHsOVS0IK1yxaXqPaS+1w9WFBjDv
LVCPYG1O3kSrSpwpvJUH9fFnyNIEmmgAHxwU/3SqWEsDKUXwpZHsFz7DvqTFTc+r
xHcpXhNZOV0CCzQzG2YAYXUIPoTdY5UUILajGhJbm6DWICcpYbmmWVI+0YPApDz2
qFM/ipaumOBH1kV1nhs5n7BmhkqkMR4UqTugefGuQC6hnDrrp4rcQF5K2D4zXtNv
fqz++BDNPxOt1QXOCMCyX9ZxF/slstP6p+80HlAu1wxdvRjccfq7PxuCxdc6uxFR
/TFwSWjgWTK0DCY31HNZShK7ihgsXXaHszjLXMxnHcgK7Ua7yEaFbeDivRtH//9f
bjCr4u4YCwLBlS1XBeqc45IDyfjZRL9Mz13xwZSmVEpMxVWeLPrk1aw9pmTbf5fs
j0NjFp57oIVvl+20pmJ42z+PR1ZXLNQc+xKa5c0vDF6/AL8teA7Q1uZ+H2cM7CZC
qcDl00P7tZRpVD79XkriNbiU9UE4gSgkC6jn0ULP2QHOo5U3XDHZSL1InsvUtKWP
D58EUhRu+NMgmRYbEjcRGI+x8rpXl67SKM/q2ONZMhb35ll3/jxjOAHbFLZqJg0W
5c5I+UI5u+GUqhwOc8NGipyyzEMXyTyaOrirOYsOry1yHZql7xtvgQ8exNpW0/N+
`protect END_PROTECTED
