`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UrYLqMJ7spMqbqN4897B9pFGlX2R5+8VPZabV/BBpYpqMMShrjLF9CqsS2EwAmBe
JYnCPrQxvmLz7tsIo/EpEMHK9+YmNpSrcE1mmXCkmSxTsj+GZ9geMjAR7rVyN2lx
gI1Kw+4bBvlIpCPv4nWOODRE7EDD6V/1cAzAxt+MobY+/G8ty8K9z5oSmKSf2rRJ
FSpEtSlwTp/OrXATrWc6uO+Mw5pgERSvdAcHbIMJkOxKhO6dzxNtYBHeFlZoBQ0n
jbJMzJecbyDmM1JIPbFDefUnS9WmXI32hVwCj0nszIotig5oa/43H5N7FfxmwHXm
J/QAmhQKcWre7lg4fbI7ikVjVXPdRt3CQa/V4zFISfcdD2yxQu608LZy5sxwMlOY
9v2aAsPt/hGL0aCzdlGSdxO1RRwVHC6VbNOfPXwqiLXU+CCXRbC5vBqzwHbn15tF
FuRfgX3D2Iy2DIGhSCbACmZ2eQFSnvmHELokUXAARoUuGsSLbuCRy2MZJFSDNOyb
GYXMv7XzfXPpsioyPmuJ2AItRqgqxHfIolG5uRBvwDsBfg1D+yuT1s7nDMKHSBgM
3bznraYGWQ+0I9DonOekIEla+xx5OVNVUEsp3eZEmuE/MciCJbLzeK4xYJO/rUQx
lBGE6oRbddDM7vVJJoVx9QvR5ABZ8izRaSloohvGxDVfo7ehr+vzPxUziYa3lPxL
cuMwtC6TV4PH+GwhMsqP1Nx5LuMnv0BYjLIx/0dd3659OzDh9f1e5qGwlDDChTfG
masdbC8lJli1k5/Lwvp/ij6vWuVkRygASkgo1FHvk1FaBi2MHAdYYb1b59CL5cDj
kfS1+cOniBN191AyQw9LLGjn4sYwE7yrEowvowYf8OjTeFktCyyFpJO7tW7Yztnp
VLp5XHA1ir4f5x+8RYtjXdzpsogM/zORzOnNkjFk4O3s7sQgGs+d2JfJXIIltCm1
`protect END_PROTECTED
