`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BZpETLjJtq5+gaBHYYeIxg0mcXvDZgQlO6BbMU7ce6X5Yip7tqAuyhQd/YjuWNWU
+XINczthnlnHTr2+XMXZr7yQM9T4Emin+mMHowbtzL9SoHALOk0XN+vcXWBSOa8H
Wrp/QQPtqtynk7035HMbdehbV3vKTuKjmOWwby9I6Fb+0BeTBati9PQyGd9pD5PU
5fhYobhBpI/wo7Y5nvuE0tSYoYAAEx9sdfi/zdK9usQdTw0ezkRfJTVCxl8vcI8t
5FG1yxmkzuko5K6EDSv+kM3Wbuh8JOTvXl/FCTH6awqdcQxh2eyd/bUcnWpw6yLE
Hyp20xjy+pdsj9YeAFd4EeKJRxPyagpQ3YZSnmLmzzSHaFgMmSqsi1jIyYdFU58g
7MrSiRcyemj6gKdPHT86p2brs/OqWczSz6htv38hJHG4UIAE/CBkSazDX/xfApZw
1QaBGxrk/zsvXoyUk52pz8qXRux0lYEx1vZ5ks/2oIwNL1SB5oVLdFW48qkO2zd7
D5gUE5ZukC4UIWBAn5+CzC5WCz/9ai7x26Bgi66N6EJCrwnRfbjzGS16s0EFZK+O
UaY0cL0X/8jxbSFiUHwq2L1Eh37zInEUwPhd0ww410/IDTQdxT6zRSAeoJOWP0iF
hQ2vtn+SJf/cHnMjz6V8GfFqW56Ce44lZlduuJ7LkaolhHoS9SSsEb9radyiaIaN
JjFjry/PUF9lU/SiO6Qpi8qR5kzkDx75DBJAjEM11xvpMyz7yfUTYwmkvfdre2Sp
W4GT6m8OMkeb6FaS99NmonVt1uYYpf1DpTo/WcFvQZAfpj5I2DmSh46gT+P8mqNj
0BqAJZQEeyAckHpj60Jn1ulyE4daF+Df+IOGXVefQrEDq2uWgDJVK0HX8ySRo6Qv
FFRVd2d0NfG6Ogil9Ki6OlAenCJMBtkQDgUQb33Ig9Uequlm9v9WU2vL4m+JIGxS
`protect END_PROTECTED
