`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zdsvsm76JvQulh0v7A1tm/t2qHa+2a1vpcz5SPbiPeiO3yHfuJd6hSQH4n3Oz8uJ
f1a/5dZILCQqQklUQix3PcnjBRX76QM3/Fg4k80q/8xEssc1PZZ8bVqqUpQZu31O
DQckGnlXcsp/mzj1iRoVU6L9Hra/E392VHDy8Fpt1Ct7nzbMBQsi0iMJoSQkXAd8
t9/TYhNId3jt65mPOew3wQj97ZC+tqp8IWoW2hTXNyP0tuB4XuG8l832FcNr3QSL
f0U3RT2BlhFEND6Ur0nB7QrascqFwyK/cdA9xKaOHRTPyVjOOqnbFU0LTaeWQQA7
lN/hsopTTanWtGRyZhWeLA56sYKyzHjo385P1Ud/L/sNRo0T62xr5CewJ9qujp9V
1OczjGzr8cusxHT/1VQ9GbgaVDafbCPnN228Ko/66ITiQwYeZ2dMh/4vDm3vz9vp
5bI7Al4+ctlzASJVS0k8xexV02CnESnbIRFoxwyMio9XvkVBSnHfePpzP2o0aMis
`protect END_PROTECTED
