`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5j1M4VMW/PPnWvHrTDfE1AzOimi7g8+Cri0hsPIRqvLS6NFul1KLRYJ90MvYLGwn
DXk1wdDCdaFNFuN/2nc0Gb0P4Yd4/ddQexR82JLWVvoH69BFI2lgM5BVZTfJg2KR
PARteORIzKS5vsL0VWyPOvfRKap+QEyPpq6yfva6JoJ5ZWvfkGiFsSkdQtNtD8+/
ZUGI0PVEpOAUP29hl/YafMwyFbqry8qv9Vnsb5OaMWgku47vEjBhyzrHfD6zb1kD
8RPIW15HpcocBOzKc713We5Yqm2wsfxhRwgTTJhF0turRDi3CVUhbzLXKM1WTtmP
C6w3ljA4DnE4iCumQ+yECbxVypwr0miBLYLD0VqqILhLT486rbSUADAchARplOEv
AjzQLoA/UGsaybjnc9ynTXdgdnlQ8kiBz3bu8BgebX0=
`protect END_PROTECTED
