`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OVIIDapc5fRVxL+Qoa0xh6djBFyN17J14fQH4/XvD4DPmQ1x0D4cWbgbzrb9IQtT
CE6STJiQTLS2SZ11MjTmD3E3zi/RPQ2kfmOIlSmq9Bh4izgkwh6Py0Phvrcxh7uP
/OscVBWGyALV+HjM4N2vVU+aIsP/Fr1kCyIAkLYl9oiqC8lbKkGEQvxX8Gyr2lhx
L7gBpisVa9DNS+b1ZEAUw0WhrYTlX8HxmRX7NfudNHnMuW/XOilZkwqCsQsNC00K
WUJb51pnnd/JJEHOQ0RQfBcABKs+odSx6zjN6ZuKXa1pJp6QQ+kc6+Jqif8p7nTO
CIw77sFQPC5fwKiz9UkOxDHzMDDyDDJXmPcMzt9iOnecuei9mzBR7rOGdZX6ib4H
CzQUJNgG/FwIcXzTSnTi0+PNsVvsXLC9fuRF/zq1Y1MAqGMUJR52geWfeK4cKolf
J6iQWDoGe3+Twia+rsJ9wr96lJkhi9fDtcs+XX9+08XOBPvnambzwABHBB7jpnmx
Cfb0r71fBoTWctznFhhq2FeboHflLns2BorhM7Co3W2x+Ry9IdpgYOUMCkudf8ZH
Ld415wHdO41cmuRb5O4tFNXjvfq1mBc8H3AYfV1a4HsczMpbVNiAdUunbFqoU/Ry
`protect END_PROTECTED
