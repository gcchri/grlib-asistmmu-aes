`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RySzfL4eIirZ4IlUg7nIfw+VSQbeYLksYX0Lq3JZQiYn0X3mVadAiw0UgUCvExcd
xgL1gV8w1QYu65ZmTYnlCoUu9/5t+lDnHqcnD0W9vQggPmNjos6VxE73awV9gnlE
EC25tauElaZPazYrMEo76RPE2KnnyPLObWCxQQiW0ftATNrGGyxEjXvPy2jXMsBd
xJuCHauYKT5BY3oYki99MLkKoK5dk6KjZegm1GLNoLfu93RGKB281IV2RFNrVTnO
jfkQCwlfe0wMN5oqaK/Uvu6Ud7QOXUwXjfTggir7Hc39ZmKGrcE8qnjGcqwCJOZq
lA2H/xKmmooginobbnU9nqUCNcvwjAaPe1xKBjgXFXxDphefQskJqEOwVLHTi8sS
ZnQi4y3xq1Th4qmmKDcoBpccbGQqU7Rn9daMCZto/0stGlbD/LSk0o8KNINsTbHj
`protect END_PROTECTED
