`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8eaRvEy72UVTAc33GYmRsYtCp3erY9eTdcEPcMAuST64uUBWy9PGZp8JSEln222n
NzIiHCB2ocyet4xN0cPAHqyfzFKa+J1EZciifZD81ivoTpuPZfBdbl1Bv79Uv/Y5
D4nKcca16uljJv5z3aZqBAEdgpIWGFh2JprhH++o7U0tTh0NJXWutHmXy/B77oL5
6P3AbOuvqjrLzbL7b3bLGAZXqDqC2/oFfphgVgdteE0DJN3vVGz7h1cXbGSQQtvr
emY0OstBv5xPouacD21rQM9Wg9X3x5xP+RjCvPEugH25ROCUeFyDmIvrHpUlhFRk
3CuL3M4OJbCScwL8E2eJEbL+jE1Lt9WCL9sU+2xCuHYIOQRWvEzlpQQ405pJcWGG
2EED4Mzgr02dSIQr6Hyz2u4sJ7fTvCjKnvN7kempw4tnKFMh76ne1TONvqdw9RVe
5xSWg7CSyNKhJByYp31Nfbod8pmeZcvZy2gEbqpSSCxSauOZMzTQBt90xL02+d+c
A0pP/Z27YsqCNXCRGgGSiOF7RBgp7qoE3/x17u/YI/9vGkIMnv4rm/NQYRU0HwYo
Ztb3wOgEvPIVRLoHHUpUK9AGvw2D3tHn/oktqvQKRpc=
`protect END_PROTECTED
