`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VDHfW1/tqj4zuFZoGSYzK3JnEmQ/cTGDsaTpkUgpDfXE/vuRO228aR+YNMdRgC7f
VM8Dp34l1eFQIsZ4NwCFnzcCUWDiVkyO/zM6jgy+HX0pSMetzXglBj8qJIQFPS1H
2AA6iEDHFcuVmIeqE+1/8gHbXaOazimbSo51g5N5+tVdoCBmx6rldGC+4DpbGSLW
RlyGA5qcll3HWDI711NliJWJRorzAKMW6JSNNZwk0S4F6fGG6s4z9Mq2cvAG0iVe
EwcfcgPL6PHke/O3gS82lJ6yrE+bfYCduDt+XsfVZhaJPin3uUyC84wOJZkWWFAn
tTkbPpTAVRyupWPvSqpvc1SAfxDdCyCqz5/Crq5UUANCMQ9EO3g5d6WU0TV1bI7C
VceRp69F2fhWVdAOFGAIByu7ghW1JV2weC39wRC/Z6o=
`protect END_PROTECTED
