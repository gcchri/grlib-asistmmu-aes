`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xokhKcBDxnUe0PnC8z2ng8SwhYMlIPperEsbYVHQxnu1ZEGW5jtqFVYp2J8lYaha
bnd5tw+xeXZZo0czBvRyZBTpsYbECMGgOKVbEfH8S97qds6QKJkisfmQV+04NC5R
iLx26XEQaFsjkNjCOb026bHkFZyEXzQCVE+IzNlyvwa7LGy01ytX9krp2X9suqkb
WTwXiB/szMcO2BCVpQ9tJVPFj3K2qWwSgh0tVSjISWLCuhAhf1inhQPTLiGW6rEH
t+9+OhGr4jzqblECRtiKLBEdrwsT8NdNakON/aenGrDASi6GBdMw2a6FgCT2dfqB
tAkIY2pfSIESIlKI5GlGAYvg9eA1XeQ/fyT5nFrvKm85oA+rCb9Qa2+qzggdQ+Ip
xE7ELfeQ5si8Vyr03UPfCz41X7uSR0Kc0CKwvsPbVs9/QV0NMERN/Jzt7R/pYr+L
DyEs8lgcNBZ8SZhB7dywhuf0o/yl58eA3xo6Cwbd0lagonjsuqtCAyZxzkHu+FXN
`protect END_PROTECTED
