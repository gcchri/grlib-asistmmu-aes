`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t9M2i8ccymNF/USTqJMwz8MqdISC40wwM70yQdsgX9yg732ocr758K6JCjURkqJb
YwR2vtsCQevaGp7uXNTTXR9XlbmmDMC2TDoG/rhQHaxYIYTijjvHb/k9kbJ0/cqs
fXEk3u2e/kxgx2lqr4qfgw0jmrxNL0IuapCJt7Sih6JSIxfrYGeZB/VZbxgYXeHx
oXq7ywcSfz2l6VgL2WgnWy3v6OmHBwTm8QNj73lZBi7uNGWYje0GPgD3H0SgHZn7
1nsmx0CHmlbZCJKtAmbfsWftcXRcnAibo4tn26aOcoeD590zAjUxhmHT2d6YSQhM
4HJXN9bebf3YXPlWEyEkzQ==
`protect END_PROTECTED
