`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b7Unk4JBZXZbN9HIDGUf2DAsb4NT/hDRNuo3JMZ2aY6fBEGlKpq7yfKFj+bmMcuv
UHcIysNljCkrh26bf0gEnvHNGBJuVxoCAjYw85+q4B1ho5kXWTTp/Pz6NZnxhMWS
D1SZsbJMVJoi2ljEDnd5LmPTP7oQF5YaonplXQsOzZ+NAB6wJ5VT/2B1H/obdISU
cuepNNJJkEjouRsXSp4r3vLTeidIruHrM73y6QIAHxQkoam8VLudOHbCV96P9/Z2
/oE6SVJa97FONVXeVusqkgoliaB1NUu99g8UULM3who/Oo7LpMax6n/NOlITT437
EP5/rHByGb6ok50b1JTIDezEf5dYicEgMBKFid4fgE7eDAzrZbPpir4ApTjDQTcQ
UqjA44sMrUPNszEvu8jGXEp/C46220ks9wbAnkr+pGlSNDerz6M3dQUlPQKo2Zz/
f8FMajzaCPWwrLF1QjAoLEoRNCQkw+lRBOUxlImew+JOtC1UGg5wdR0gm3Lg9e/8
QXw0pc8Taa1py1QPCfO+UWnxntLSVauwCHPHLPqpCMP13T4vgWqUWjS3EO5Z/ZfQ
vEfF4ek2fX402y3wC9fayQtn/ueSwCYN4LTMivn1811bevNozpILfy05+p+VLeis
nemaizE5P4I4jE0QDQ9loO/9mtQ51eRDq8NQkrnmuMk1+xAbynqmo7JXs+pPAFRC
KSEgxZGP8Uj/TRvdE5JcZeyszu6+wpas9O5/Le37lo6htLux0V7OTx18SrRYhGbH
5AUCgpQMM9K96r2SVhhUrmsHLk6epoini/wITpAvdtKI7m0YfzelkgOkSDXCe0/Z
Cr6J5ZrdJ+3ClwRiwBGyR7ytzWK/E91jGS+1MqtPnXl/+5tEIxKQBC2fClqry2ea
iyBAVJK4JklzjQRh6ULLorEIfMNhz22cjYv8SlaexwAEG9QS2bBkKUCJ8d76Hsx3
`protect END_PROTECTED
