`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RWLys36iWYXdSYdg/VR6rdlsbR9CvrKd8BnuHa+jZtQZ/TBEQ9SHLDQtVjv4/Q5r
fRM2YTsb3Svi/EsyFT3r5G+rVSWgccm/RhoVB0sITdATn8/410mbKPRPq/RYm7X1
JBMbYFLi+hVQ/R7OXehk5JDqKHIG26gLXbL4Nx9Wc1h54L4Tfy/yw8+ubmJ5f50t
Axr/ll8j1Jgv2oAiJl/ROyAF5uvYsqyqI2HvKTCvcibswX/7BS5OeWxXz9CIIRoe
Fv/Mm4bnQHvCvqdvHt0esVgJ46+wY84PZOM9EcfiUf0mbrkoQS3LjFnjqpzZyTdP
btqHdMoikcmw16cQB+JSAkUWlMBmK6Il65+Zq8jWqTi7QpRjrVCBgPp0bduVcNNj
nluGrxkW2zeKOJNF5uKi3KDl7YjHLxAPeNqcuF+nNsDm9UorH4PqJmFXR7tA1t91
u6B+tdkgy6fc6NR4W/zrQEKuu0dCTEUcrjAGHAaZPDfKyv7iQbF9pVTq5DE5NTkC
9XkK1Vfm50vTb/EGJvcYi/+h3AAvBWEzZq8sBJ/YKvOJ31fhEd6cJRUMb66gTz6h
QutnyTBcd8SjNTSvv+ILIuJPtmlvFM4gp1eqGSQVkll+oQ+tRmdsYE17w2oTrZa4
eEPdt+4ueKsRgKblpx0El2VIU09JkceYAsyHBIwZ7oJf7TpZ8JIEt/mQjm6Hi90z
XG6YZ6pK36Bo1+rCnS9RBxTbKDS833Mv+TbeLc6Kryz+uXjroyLI7vjPy7BGyrKi
4I0mRPiVFc7PXgKs6s5rFHVCZMMbK1WPfnt4KzJzJTcqhHI08WhW0PtPm4LhEoKZ
dmWuBJJkkZO3r3nhwOk7q40ftYyxmGm1A4Y52yL6nc0/wMgwRucNDNQmdvWXiDl/
gPd63HrmqpwsnhP9nw8jfCB2sA75tENt3iKWk7ny8FXzetzp/EkfQM2vEh75X8H8
TPq2Gxel0t0skPxmNvGDKA==
`protect END_PROTECTED
