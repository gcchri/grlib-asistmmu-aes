`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sFQyoX4ApHb9P94BHs+tNbVQOCmwCrUZzbg1B7R+ap8PKDTnLA96jFV96Xapbf9w
mSAwymYEPiNYXMdn66YlSVfVV19gNGzwPpG9+7/rPAOHRMpOozK/SFDSaqioWPSY
FLjsklorouZJR9F1SHQ6vs8RvKpxWLkj/k6bEu5C8jPQTG74wY02ba9qRd7+IyTu
jSjZ2939XAcobv/FreWMHE/nj8Z7sg959hf8IxGSIoluZyK/sn52N/rbf5KvdJDb
m6xzc/SPayiG3fUO0sGPsonSXFrSpQMOW0G06esC06pUwfUT1i97IErwXlnE7whf
isqv3hRSsGG9eKoQFcb1gA+4FoZazkccwvmWq1/SRRwbQVLIsOpttmahvnUlN7mc
/Oyng/B4IM78XVU8nL7wp+NLjvL2kApqx2UFRO7KgtS0q1eXfYX8x/+U52ijIb5r
NUNOZGrh2coTkZUTFbM8RyaMzxci5oFFuB3hHoBfixarbJfVt2KAeOMhpIHyN2wO
Lg1BV7sswU9kdCwy5nY4cDl9Q9HF8ZBB29vHDRDeZCMNDQzKzIj36gFnIACleFm+
9ILYSvgO68gmgsP+tUzwqs7ggxS0gOoMy371Pc/6TRKjhVy1FDsfpRf9TjJZ1zja
VjUOV4XdwiIpJ77ge+d7Pj6odQWBAKaKogoM9aYHBVgyYufftwkOBhVaMCt07YGB
ldHAFbxkdWvqv3tuaPAvKhyEANOE09sWd+SNCgAQttP6WKrrUTgfgbMdzeGewkZZ
M20+ZP7Os147TrRGHyWQJNZc2xRP0GwajDSG9dR4nkayndlBU5WK7xyb0dHZJxZ7
H+cG1pKgqKLVYurm7do79Y8LjqoYDOODIx8LEjyyVCk4o8MQb5xTPo4l8jW/sq+X
1eJTWL884UQ2P1ro0irO0ELpqhwWRpTq0Dx2PaUwSGPzNxzJwpVSOJeFhOulIseU
qOXVRbV7ZdEHdCBlSvWSA+6oms+Drrukzf4eOcTnM63TNtAOyOu+MRJoWK+lDPaa
O74wCVdqYg1EPso6gUEgo1ERohR/eGDq66eQriA6caI3zPQ6bzppfCwCPiKeyRUy
kThJ6OSUlfd6XmGnQ7rp6osQ4aKjAQ933U8GdFjwsWHC08hDRvcB3qT/1kKOmPyq
EXbJwnO7ugosQ+CIO304J6PX9V0TiTiLOgI2TbhLu7eizNdpb0tSZPlKZvMR99ob
nlLabD3FXsuxjvhuZ6vdIAEBrTSpbqvy66LR1iniJosUZHWVbw8KgIfwdH+u5mo+
Ne1ZWoq2wr2pfmZ6fFvR9x3AK5zunFNioGiG2/+YkntajM2koL7M+qEx0iubIXtq
fKUDu6gI2j0diGhmSWj1wtbvowApORw3jOXs7Bxv/L7fQRFxJ7fxLSSwA2efNshp
e3bm41E0FS7NLD2w4wvpuEey1RLqic30NRqHbVoF7eRwRiu93v2cGd17jwU5kajm
x1nJRdCArTm4ttDTEvYoY9aovKSRalLHjKxqIeC++XYUjmxqGvfvkCn+wLC7cXdq
hfnrNPmXiMgcnlz44XwbGp73/ejM9Q246WBprbILVkKL0ifTJrE25rcKuoplk2Fl
+mQIwxmOA3hcSLihF/IPbqCxIJ9d1QrqcUiY9AFnrkFlqmuyfEl/NyKR2q+kwR+8
nUwKmOef1c58MHXnZCaKTPx8jwN47G50XNxZP9sLE79GmmeTzwaaOZPvOU28Xe2f
Mhf3deZCRHviBWsWLWo3L5DxbuHDzFjdg2Ett2pjPyWejq7okVByEaKBDs4GUP7y
8KnA6pudUmVkMugtaamxCy1wUFV2Il9gjxNaqmjmZMsxJ5XmUlmLfnnAegYyjuAY
XEfckEdf+qzkj4DBZ1hF6v01IgU6KwYdtIaWFbO3guVPgf5D3Ve02TpxeO/lFNNu
Oy56cRzbUK3C2HYwNapLHXEEUkZPSncwZplYjCkmvbMFqrDqh83yaNuySnJhIcN9
`protect END_PROTECTED
