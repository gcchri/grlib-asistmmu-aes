`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Waldag6D3RgnSl0IfFtZNgIFNPyd1MlrgMm1olQOPPKw5QExBumzyCTF+78RP+15
6Idb9IGVYPKz9D3YUw6BTmBsLKP6Nag4/SOdkZbEWCdR0/bZLQr3MmoCfOYZUXV9
JQTUmG4AamGxxk72I2RJAki3+XFFHH93JtMrBLdfG8dyObc1O1gnOFR2Rn+/Oa1L
l+gIHo2E5UcZdMvvPN1qK9zqJlaHdDAneuvtAhhX4plQ136v126EgejSyHCRpz9g
QLitpuUc0qlG0xfPZjfJ4/H47zyYA+uxHzQ5Z2nEF/Iwcgly6vetB80RJoe6cDKc
smNqtdEtQg/2Pbc/QOvUfS1RjlRMbLWBTw3gNL6WDNoJfmUxASgbyn2aa1wpxWOp
j5Pc3CcllY2DXj/e5UGQwi989D4yNEYmqjiYr1lopOm+Y8GjN3YOSefvZAtb6R5Q
PeYGl5Rjpq5TPjhu+qGRxS+h4J4zSfYqjud1iZSVpRVGSXZg3Pj2qlvQIk2pWSjs
NxWDEp7W+gxi/PD+M5SFFKuRCwKgXZ9x1Vc6aYDL9L4UU89ThlecAfbO9rIxCn08
Xm4QFpL4BPwPYb8W+MrWU/XLQn8NrWzaZnc6lrEFxB2iCTdCi9rTRr5A7uLSAPle
tt1kQpp9OBY07150KtFZOcYrRSUFm2+lF+8zfb29hbUaYpI5X+5aq8EVXfLjgPCZ
4iOFj3k6eKdxnYkJgJpHbSMXAOXjSVDKByHpi15Re58pDAgkyjOKCN3ONxvShkHn
r8mufY5Ll6Qc998CnJnohFGANtieCSjEpxjlH+W2CSgX99+21CyFDK3OSuFRiFYP
u0aE2e4a5/rrClFl5P6tG9qAXoCmSfHyktaIKMnd1fakEOK3NrYwU6Ch4NCCeE/+
MdSFv6rSss8yyQF/CMFxttVGxxZu/QzLe8CZztXWNm98FlfRuBWKtWFHWo9C/xdW
IrTLPlqbmyBtkjRoDaIFeHH+1XBg3CPZRGoFexaznR1xk/9oBjgUOMlp6EpWq3d1
NI79gUWQDkFQxknfS2C7u3hBm3Q9pD4ofetUacSRapA=
`protect END_PROTECTED
