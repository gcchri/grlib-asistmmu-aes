`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ubMe7T4klMHLAjkXtPr9J9xo+A934HLRBdpz1/FWhGp72+Iza2kJn/UkDuR6P9SN
AQOXIxSR0ssDuDBYmrQrNW7JtppRLCB5enj7P7/quFYtD1inP4EZ5ltzCIliW1t9
bDRyXz+0kbP/cIIS/kbuKlRe/rMY1zRQ127zEeskSmu+iKHP9H++E0xbkEnRNzQy
ZkpFgqqwYPBE/ky/k6ad0fkIauDWqi+c+4qTUO0RJJ/rf812uJlBRTLPNLBNmHRz
KBc/QzffnarAvkXpS9jpQmEunRRM7Q6s0oyALdLdgTa4I1c9qe98YlSa/KF5vr/H
c9KCVt/yXN+lEZJ9BduvmgEpxLDZH7fhQtNcObqFAv9crl040EfVHzigxuIe/M2O
QrEnd8KtofH9vnnCB97NmvLU2JxlzXiW2t9jMhUC+4tuOpdzVPmT2IENExi84xLp
sM8kMq5HYc3mtg33Ktn4ET5TJb3oYpx9PahIGROg/OQ6RzI3bpg/HbthdT4atDIk
tS3+aP9u56XL3CsZUTwSzM78fVc0oTfZDxknD0yUGSyCVrXjoM+LheLpeO62CG0R
psOF4gq9RBzkZU8yZgNf5SDL9UNQGip/8iUu/OPUJ88mRtE5cXIrZtkf7nVKc70x
jPJbfvc46SvLWdlH4stgHxzKj2AEvBbSGtfFS40huDBNhFpaJDe3geuSLhaI4sBJ
8bb9FKZX/jqN0mKfis/ayLs6/c53VXOD/FgRFHw0n9gI73V+CNZPIUc+0NHoNAaz
4e7EOnVe/ObeBluiBh8Muvg4QyKuqvOZPDhVrhX+ISIyBzU8e8zuLDWWHPAuLhrO
FWOHBpYxVdXXxVdi4kz6ho4ann4b6FXP/2AHWCufIajlWrmwxglyQnyMwqm/8KeO
FWmb2bfAnDE/kS+OHW7e8xhZN6w7PDMtodz1dJ3tNeuWgRyiWzrjQ28bA55tmSCs
YEuXwp5H2OM9aPmi5uUPJGw6FpCsrrmtTLEx2KueNedTBg/F4iLJ2XUfc1s0Bysi
/8qLO0QdbiDeq+n70bc8/ntNBH9nHdAPdgEhLHB2iVOM13Gl5Mvao77Zcc/6A1Xp
hPYb4N8QLSqNnVjpQCEgCiDO0cMYBjbc3jBcbd9jbOpsBcpkglilRTUcH73INfwj
BgZtCZEyFzEdWFgLrmsngQ==
`protect END_PROTECTED
