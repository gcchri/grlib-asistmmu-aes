`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ULckUQRCHfdWnlczro7qYcs2tGvaY0lNUSETuOfR1qaCC2+PqW3jI+5od0k7vcr
Znmo4/ITNo/VpxBi1sO+mFVwg2ZZ3MQKNaaWwiNHd0g4KvPMk1zYdyIlfg9+Txj5
r+6rCEE7aOnP7NR7clLtlSurP7jbzFTRaz3sdbtcbBBXd6CFZySx2LiAfh0XgeHu
9VdKG60pVHpN+dsbqzybYYybsOMXxgOz/t+NbhC25cgPIwLYz9c0g1N0iL3UWB5m
pPEsCeOdWVQEINYjN+rgGgS2pn8WCXee5/ut/Trwg6Pf5G3391bcRzmSgcTHqmVE
p8CapenSPYdCa8Yll3XaHJaZ7QjP0n+nPeTijgOfXRy7XFLwvbnardg2D5alSLN2
scHqGeJRhMChpBGZN+FniaNHQ01Fj/VNiH5FEbRIkKe5CrzjzOXG6WVrbetISPWT
iPRGRvsMNegvOhUej72aNfbGv6lpX6sshUrbNYf024U/jpEBAEBVMi/w6FBS3pgT
Tb12ksN5cjTMS7VqsWrEaSkVegTJ9joQ2TgpV4nBcKZpIBrcWNp7QhcqKpe97ENM
`protect END_PROTECTED
