`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bOkZIl4Q72hzZXeiwJk+e2074nYdgp5IBQ8uzywORoAhGyIp1cWwMdzo+FYhyWW2
WAH5Qcyk47uG97Pr/ZOTYGftWvXoZngd7PihQkbUiggx4nuHx7PaomYcwucKE6N7
rJs+XFe551Z84PtTbNlloeQWtLH+2ErQLDGj/eD6MRwRd4hGf2HoSV73MWCj9+yP
ih1mfOE5nqbmKUzPv9L+mNnZN5L37iTdAIdI76RFY81vbGG47MYK/5QcX8Ij0KR5
QES07ikF9lmqfNhZpC8+oi1P6DNFoezBXhUFs+bD7Mq4a/3sHdsKsqsSFA+dM/U+
X/7uBhDh2TyOranlP3Xe3YGsruMbP8+QST3sCBLhpfRNHdoTxCGYTezAL/O5JVkX
aSXkiSFn4qqNMkUcnn8zj16oPqoIPSSqCAQZYSHLzBPuCLm3EhPnOdWSvT5yaRi9
gxrk1H4JIVfQFkq82gO9CcSsQpDn+kZr39R9HJnBfNTsEQNC0slvfkOjawtKfojW
ia0/BLbtRHWoyChvUnBwPyEajUxCfPD4eyJoRhN+eMdVKL18kXFLRzKwThmv8Gxp
8gqWrfR1ySmj7Wq0T81pe5htznfzMpG6TG5ODcgkYVouvkNW7KVe8gTGCj6iuDp7
A1HNblVvB+m94/Hgt7YlrA==
`protect END_PROTECTED
