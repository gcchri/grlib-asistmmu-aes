`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jhzO+Cxu5qq0TGQpIJsRHQJV95g9aVg+LytSdVA/pEmlyD95rSzST20LpSBOtQg/
OPxA5mdvdtcXCMVQVVitCZb4wbjNBTEA5OA93wK8+j6FZu4nEq34Vw8vkt/8aa7i
on1WygkECFSg2NlPrJpXnfIzXYm8Lld5CYBlzwSScWdKeCLFDPj4Hdg8d47tI7sp
39s51XAFXhgUi7iP3ZYro4YgrtWGIDeR4oLzes121isn6lPMA//xNJuKVOdTkYwz
j/ImFzexXnQvACwK0B1diGpKAQVUeAb/ENkVEWjIRj9kojZOF2+TwK5hqTixDowQ
YgitgGwemr1QohliRNlLjZCotO4Y/3Gcti7Oc93+cvSeyscPH+7XQ8hkROTzN24H
gCxmZvJqJLsCHQuG0AGqnmjn4yvQ3NmfQrNElaaExAwBCD0sEH/jgpMmLDAZXHsc
/eCcz8WPzyu+YMKhxnxpYJhNWluihauuvpcbjOZivnRbarEDAL3ul1Kf3yfvA4j5
mbCQaqwzEqJI1Z13fM65miFGqj0biq0wppXgMbZsQEB45292c5luRAX6KnAsiUF0
iPuZYeonEdOzs8OFA6D/x25E51Zx7UxLfqOat26UjJM=
`protect END_PROTECTED
