`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XUOtJmYCj0GZu46qsic/XRFYu/5WrzPegBEenSe+WvCIpksg/4f5GObsLxW/wu0k
7aAnc0gAYx7fqpQPETAF9Qiw1kOAZ31/51N7kb3QG9Aczx1sxXgS/mOLK819TGmB
YmC7PuscErpoUBtgrglqy95YN7/ZHs0V5sdveODwAmNPgjG4EeGYvJNx4XnxTXDm
EkZoaYVS4M+qMKOww3n6xryqMOdcz/L6op/VmTByRvNYx37UQTLtI8TXNy/CjCVw
3xxiQdaBsOmY5REFpbrI3CHYykKCh9CUAaHUIvm1aCFh/HcUCEiwF6+vVLJ83S5v
hLrr9J4Se9h3TiTV0/w1oeTQg/x2uviGBsZVYfgCvhQKCdk632a528BYadruDgef
mVgD1l3/3o1mUusedeHtcY/K2tw8mXkNZFY1BknUYq29VyDHZE7pwNlZE3q/33Xw
flKScR9scXqUAQ+tL6YKMirYllhLLBARimp1no4h7ynrxHQOUBzdCkMKBnQzq3nZ
6mPXkTwl0LYWQ2sf0fDaoZpIfIazgRrF8ibkz3ses8+eSZBfAgBTlZkj/KkzDzjk
sJCAHTRxUalKSN0/hRj581E3w3b7ps75B2jjHvBKMlNYW1cKrlVTshEu5jpSgfUD
+i3XYCQ9WK7id78MEAwUjw==
`protect END_PROTECTED
