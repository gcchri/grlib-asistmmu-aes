`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/R0bwt6cLZgR3TxwN200angoALH5K0DsXhmpcZRkqXFtWjB5qn5S8eyIh2fNfgp+
ZGfi9o7KzjdFYzNx90ZYiKJz7Zzy401MDFS882QuuKgrUhmCSzHPxH0JzDWIl+xy
q2OdG5J6UihKuzQEIGMt7VOqpUyUZO0lfngT9LRtOKIYFo1fIudChe2ruN7GV1UT
BO/vYERdEaWWqY2je30nsvdkl6AB6/YDQzIYrp7eE8ggX544BmCAM7oXXT7dNKj3
F8zxUT/MN8tHuMPpXPdx+Z7N8K4elLofdSMakzYfzQ+cnYGmgAL3CTNB0NzmNZCm
t0YZcA0axQ+OSxdn/q1hny1t7CImFY5iEl8CMD9XkoGZkURAGUsavWDLcCpVtSVj
0BtbL4QqG7e9l4JY6fJIwUQm7Ism3G341MVblM3jBzzMd1Eiab1hRSTNEtliovN6
vmb1qDuaq4YWMIedG3FLHQbBP0NHuUKaj/bIe1WPAJo15KcgIKj3B53WRJ6PB5an
+p2bsFa/djBiVzRYWXf+zDAKM9It+8F40w8yMZwnr+T4rRh4y/n3PWhnNCrz6m6E
xRf+8+PRVEMuiIaZKTnUY2w9K/HNRAUDSVhwY64zkpI=
`protect END_PROTECTED
