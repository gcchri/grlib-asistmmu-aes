`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ws1MJ32gYc9Ns85jIjjuZKYfwyNU/U3nNvhQ/SxmCu/JTiAVK2rahVOyQdKiCSQ8
wmYVtny4Na54VTw60UM09TOg6Qx1LJNFKESO5i6vF3xQnDTHF3gNc8k6a8u1uH+I
Pt17akQB+UPLWRj9Qcz6Z+mIxuLbGqVVsqXp48NJkQMoR/P8IwpsaZBtnqKVxaLL
HN8rrXorrs8Zob5ettDU2TLwffEM4bn1AcdritbTy9DnMlIT2v9JWaCdO9OPv3oJ
Xg1h/v9TzcvoDx/pW6b1K1qIcu8J9Y2CLl2MAKrM4pwjkZa2Mz/PcY7JqXPdxtC1
QZXYvOo1r8WtkBIDs3qQjS/aFK+KKkSp/vAOj/hyY0FBzdrBB1ykWs9DnSyiVgor
h7mO5AMcKR8YBysSGByJKcGwseBfR2soI44YUjTb7zc=
`protect END_PROTECTED
