`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+meiquC3wyMy229DqOpCr8r2B2LkA6XssasiVh9+5ImDstqKcutkT4xT6dBRIxxE
e3PCa0JKxSKpEA0/nCzUdgVMgBogdnZQfAsN/0KuM+aqc295dLg11hZ6nhKwNPjC
wAZNmCN53IVxVSbbeoQq/C4Ol8GqQNSdzpF4dPT1yYUasc0c0vA6DsVmvovXaW2Q
ejQGbjm0t7+idZxQlA1d6HcEPXRGZmaGrLkrYw+OYzNpXRZfGu84El0MwDAOOJER
Oof8da3Lbvyq+L+vsU+YSN/y+OmkWeAPfYgH/lCLXEkLlJa3eEV0q1dw2SbJTAOM
fRDT0+7MoUzNjeOLCOiuCyGUYQS+3NDOulltf8CbjwNJDFM1/i2dov/uz9nf/7d6
vyczw/XWNJzrJEMduGOrThnct/VazK2Jj0TZBpt4DOFikleC3uppxDYyoPGlbTE0
msO6M1rvxVvwFDa4gVuEJJzMm3sc3r/0aFxAxSnHlymouKjalcPow0m6RD3fwuhQ
Fe+86wqARA+kgOE9y6UAJU+H9aQIKW+vzH2QgXm0CT89l32Rjz9PCgAZEoPbhVZF
`protect END_PROTECTED
