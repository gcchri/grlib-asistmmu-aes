`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TY3atpQlGGbGwGyTnHlQXZseH+Z5vYOMJpn/P0Ao4bBfUyLJ8DvlyaK6eFPXHgfr
UqzO9teBqvCY3tgkqU2S6oSrrb8uKfQI9uVoU2UAVf7a1k34NwUlmQYu2i/tYy6W
tUslJ9DiuDlmoY6cHAKXBjmC8oyV678l/hz59tcKUAjSYlUYCZGW6goJ3Y+QgbtN
QZRs3WVpSdiEUp81Dk4C66jPCZyZbHIfXrLYalLgUkImjl/+Oq1XY0HOtP4CzhJF
VQOPSGr7ko098l2i1yTEG6kKsMBHfvx+rXNKRe7tkJzpA+0kPEiDmOtUynGyFocY
x3IoSJJoQ2u9EIWzP+xcxA0Gild8XKpHn+MNHiPv1QKGUMU/mQnq1pAMVYh9RkW5
KgY/rZYtWjF8lWxUfruCjw==
`protect END_PROTECTED
