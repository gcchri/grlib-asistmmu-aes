`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qFIeJfVLKZVOomjmK1zsdD5MH+kBpyUy8GyaO5Q7wH0BP02UUUAi2UryIiB9dWCU
oQZvtuJo6TZyE10bfjbYNEuPCgClIVsnaCT7ftaMFa9SdE8RPrumwy2lkZhwUSb1
vjHdxKmyrhzsZ6ciswebGSTkKTuaNGBajC9CMT6ZiKhbvABOXGGvmqhxSedi4+dy
hWNqOfWTV+nn2xaR1XmcVM0L5s9NL9Wx6kFrvdarefeeCW0ulpBBFebLEE0TZ0bI
yeGHSH5l5SMx8V/8AhCYB4UmRVQjtoMVhciOoVGktS0PD0tahRWo9B2BdLI95QMH
7bWFWyZ37FdQmOkTE0UPejs3Y4ruwDhGpt2Dpio6deg1lGnlclZyrWVbcXNJpsOS
jus1o/kSYGQlPJu1XABzrb2fCywfDfDFqhLWeRWZNmAP4Znyk3tnrfDk6+3sR23t
4t0i2klNa/4qNMRgPajr3jXeThOUA+LyLvXWbld5p1I=
`protect END_PROTECTED
