`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Xt0ErzGV7WUEW62+Kj++1DOdkOnC2NorOhPwb8i3xU7B9g0Y/LeJErvJ/h5u77v
XCP1ee8GE4X2UcPNte9RNj0BVXNvjP/GHiHIUxb2nVyXgiIz2qiu6usRQKnfCT28
BvZLKF7isC5AKZczFfjMFGyF0u67u/dILqS9gMpkuT+8RN9fCuMoHL3tgqiqTS/5
d9twLrXAAYpb4twro5rLZa9fiS1kxUZ6qKTfS6pGkUlJiVTdeQ7b00r9bv5/mhi7
q3eJ3hH4bOe2MP6chxGS6q7xyVi6/rFyoldA8WcRp3K1uNf57UNzKOGXoOo9Pvwa
XPjsSjtZwuYfRP/hIaUIxnf0s775EDPYw4bsZBvngnEPPM2gRDAAOj/9cYYZBnQU
/HL7BjvrcE5OF64bwdrRf6TeLR3VPqxdEhuu1ccSWkc=
`protect END_PROTECTED
