`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FZMzblrybUfbm6mbOXNhPFh0u3bHWSBcdj/bnRTjI3C4q4P6/dSrdITW7WHUg8Zs
X4RNoHjoY/LMK++sQJC48i4GQBqJK2VTSSe5oik82YH0iUG5w9qzwEmi6lUhOCNZ
udmurt7dGTav2TBvTKZB36mHWckHYc9u8WloID9MzQ6eYNbOgZMr4M6lpfl58ZiI
XyiPV8OY5RTEy2yWoZY4B7Rye1JT8Yd0AJ21bKuM9mjbBgIoJZSlIFy2wx/MLTk7
QbjhSYSRmEmZE+J4VaG7GgIDqs5ZbPQ5V9Ynfs77UAPx9LgV4qOBO/SEheL67N2u
29ReEAnm453fYQWGUsD/mw==
`protect END_PROTECTED
