`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Az92rPP0KGpISwTQMSC7QleFDotT4Mhsw+8zRxBF/QbalnoeIwpQ0Ztg1SCdqCcz
pNgXHvPzi2hzuiGdc9QghkZiAQbZQ6a36Fdr/Ai/7BtJmsjAKFh8oqAtpRhBjgPl
DRuw3cuY73/Yg/LpYw0iapfC5TiX30gXbQMjPmSC5pVe2a3Z7SCTQA4z4QXfRdzv
uC+rNyiB6fNYmIT8GeOS4LQt/K+pTs5dpUWC9ScyZRfSjt8M0HffUTVjhiGpk5yq
a1u2aYK5C1UJiKFBLMXMyWw5uYz65U+vgj/n01A3u3ML66FPscYoaVyudhyucqzz
En4Bp4DKmAuwS/VGbBQxoywekjtnW82fynQ4L1BlIIWARzoTjp4tR+gDracEQoiH
Q2DjMuO74XkpYxZprSA50mAIS8xq2e8pi9Eu6BNPRTg0ygwyCRucbhNxHE+DQFcr
E32FrmqILZa3vY91J0QVRaGI8XXdkwhsr/KVK0nH9TaUOKs5hitP29eA2F8iDWly
7JTO0MYnaJcbT/Fm1M/FSYZ570Ho8BZVxmn7QbGtNXQ9zxYw72+4f2FDDrWhcEtP
7769Z7aBHswksWBktfSS80IR0sp/SGE/KOMql60S5jiwanPvg8/Mxku6fdnUrAGl
vJjSOfgfNrF3XggYET4N/LIwBJOsJqEZrcbbVDvH6AOE/Pqes/bj8n6ZftnLBwM5
SaZgUSwmoseWy9QhQ4dwOTOaiCfRd/iRrQrPSGyLbMq1go5GzV6twdIExRpapNEa
bVD94Jpis4Eg8Jmo6NnWwLjQhjXDjkZVmg7T2NJ/1qqOWOkMzIYyIPxikfI7HE2i
2SnyYZsbDUruHhqCoYYNOVaUZMfxp+dCug9LtFD3RQo=
`protect END_PROTECTED
