`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BqUHjSfHPq5R8bVERQ6A1yh5POZhEifUZDg65Cwq7hWHOhjSZt60SeZK1zUoCuO3
nmPM7q0kJBpH01fpvE/a95iYbkCZDcG/THDhGwW0+263QRkQF6Ejyf02gwSQ0cDz
UyNlOLBbbxrL4GkWbJCFIPT3RM34t47/VcqwQ4yQpmBAuuXn0oscPgrFS/8jJKTX
E0F9fRdK99XOLxgT7Dml0cmjZ7WP+I0odeabOe4qpMCY8WJAE2lHV+Lria5zZWj3
xURLoH4AUOG7HMlQULFi4w+lDDHKiG+jQpw+6CpxV7vivab2aEvURjM+/GnNZCaU
boWMTRiIHbaG+k/SUcDM3LT/KcQdWdERMGkVLsLnWLvUiztoSSJ+bFxOCJTh+PZV
tR96dFktqAiXHHJC2QYG+O/r2y8hV6Zma1pUb2Kay3V7lTI9fOaPHaGQHhoMMlJQ
Yh4Epjc/N3LMrzJJrbnOP4pwQWs9MyhHjY/qglnvd2/SEdiW12rGaBtnyKH0Id8Q
qm7aYkuzePlcVY6KsBinUg0e/hRud7TPRPEJM6tH14oyr1IMRkI+tnleNJBEEoxv
qgyHCfI+amWTaMjoOVCRv01i+cnIz+7IlUXt+9HNy8clEYrpXK3OX5Qt49P5CW/N
VFfatpqOjkNWBCj/4V36ifA5LgdBS0Aoy4WDMTRqOrp1gR21XqzukIZgESgc5aTr
PAYXF9UFwc+y0LR1siH87no9yPG2cqTW1WcuWt/ZX2RUQjPjA0N7BvGHv6BqxFhe
YiKlpKVtsiJ6nsahTTHJo3aFyB9EtjO6PRYiu1yDAgQ+9X9Ki1ey3O+8gEaXBEbH
vOkxIT/NgMx5gq51GfMd3hbxww/lrFum/0iLvPdckyA=
`protect END_PROTECTED
