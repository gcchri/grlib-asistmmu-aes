`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fOnwRcqMefPd4AAGr+RdQfGxYiwbRsVsWr1N/5hhnb0o4DYyX4QC57QqnQrNvnUR
M/BH6X5gUZ0ENP3233ULHjUzHO/3wFaR4UVn+uQCB2Rumo0GMGzfwwigf3h2E+KX
0DJFddyzAqsfAYyKKIZF9x0jJf6+f3ov683vbaOCJCuITKRUx13lAesMaM5x2mEv
ly9pD/ecc3iqMTFI+2cI7HGZopseDPHHHLZoS+NOT5/Q8u6nZREi+ORfJvGF+hGZ
TqpFW5ZPuCw8IMxB0kw8eG1D+jrWM/fMPMkad7nm5syP5tSp4cSlOLix90o66mdG
WTGM0Px9efWhP+4CuqetibMnP5AiiLJbdEDPkOLW06mn5QRXK+XAZdNdXK6yGpgT
pREw/GXzXHtS6Hmt/AoBRnZ//yDh9md60SPnjPr0K9xGtVt9bzoNYaSIXG37JaM7
ockwUZt/4OuxBbma1xqEqQSmlBAenYWwPhOmoyCCY/6rCVV+xWuBa9D9L94IyNWe
udFePmSFCZnRXIMHgFD21skGYdXMGJGIG4N3Mq83IsOen5mb/EXetDvL5NRlN+Pl
K8xcJRQykGxnt4J6QQrVjklYvZaAUXZoOYogU87bj2/cp53Gb3w6bAbcg5c9zoM/
a59ByXyRgqcGkUG+ybXtqpplJmtjr+WyCN2al5of1WfDwhfX/FtFmISC9UyHsvXr
1864XQW0ukjDzqCk8n/MhIuJwVuNa07Cr3R/UofnAqYbqjeVCCnK2awhIifEt0r2
sfVqFWOHpixtnY3HjzeaXoC9vrYXBEdRZxAR1wjszefXngpXVm8/G4S9avRzVz+U
Yt0k1vjwrGGYQe/C+u0lo2fxI02nY5wyc74OWIqrt70OJG6AKWYojbPyW0P30+RK
s2gg/Tln3Fd7m1EUKJEiMP6giXw9uqaPQ28IkwAGQQY=
`protect END_PROTECTED
