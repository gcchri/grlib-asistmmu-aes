`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ctO61zaML1D3jtAQ3Brz2jkYEMd7qmrHSUYTCRQOqWrDsqhHd1MFkiM3soZG3J8o
OFld61lDn8xbA+ZkZFaOcxKfUfriI7KnOb0lLozxSEiUYtS+ezC3oaV/MHX1Ph+r
c4cc6g1nq+ozENA/2qi9jTfJt7f1WI6BqFdtfoen5zUvtTP16ApljUJDSprtFs8Y
Zj1Mm7cTS93/XPBiPD2UySho84+YUVUtHa2YKgrAp+9aTMFrNniYDLU4c+6/0f0t
1ZjHr6fhoqLW/hAPLf8DTuoBGtnIesFz7b1n+wUEmKoMD/I0Oq69jH/LEnvDlPx0
uu1gmYEJOc8s14X0rsJVqLT072JbHFoTyU5SAdE9UxTkcDFIDVEH2mCYMOaqV6N3
wDohwIyvYqAPEIsWqfD5leK/qr6v/Kr7WsiTW6qCVoov4M2i5ri8Z6cUIuaXaY1/
`protect END_PROTECTED
