`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g7OCY9KewGSSKk2hZCMJhGD8OEtlK5WAfpJsGtYLSp8VLpxp7KKDY6lP15Jm8ylH
qmu9pq2R0yaFeqqG6KRn9h3gc0ytpy9IifTOinx6InoareTyNWZZwVYXrGwdQe1i
+zRQXXoJF/ZrixTAr1FB+KvAJY6EXg8Do9fB+/UfA5zp7H9bP11iaFyuqoPj/+7H
dQz0g9sXTfhqDP0T9HXCwqhdtmdnbiX2a2ZKEbbNKeP32+RTUEtOZouuIVckpuOd
xbJmMkDHiz6ZRlrCTWqUlmyX3nmkbaHtrJG3bJWSZDEg9F65y5ZzHHyGkjRZs8vV
lolNB+MivbV33d2W5ec1JX0NPgNeCtJlDt+Ui53G4pZyXgdDKnvTnjg7vvhf5v/r
8IUm0tubXMvtmMQp4EnNRXmkj2srBRLiNLlA5KgDtFJTM7fe08JZNNgAxTwkRMG/
FhNlTH83q+yioAPutkKHrEbWd3V2tFFhXcFMTy0KsY9/vcDO+bzyZt5kL64UfYCB
djKqOeDiPoavOCXUO+aA/Jp4P6c5spKjXOijRZdvhxVFmgXR0RuHC+7WRx6xZK8G
dyisHcELk/MgTO103sD2h+YSq0UYfpuu6UFXYe5aOga/3i4nAcD/LzVOlxPqj/dw
MtAMDuXVgjhyCbqgOUiVJVCTzLnp1jIwkt3BS5LswmAqQatOOEg4aYEdIwx/bHLY
KL+IiFAprrqXVT30cZpf2MBSTFZOzEw8UqlHzwhqP1aOmEY57TsXQcVONnutj6pJ
sTqemboIIgIDhHL0MhQ1fg==
`protect END_PROTECTED
