`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t7PVjG2ZGOXbcn8Eem9IAcqyE5/IfkaegKSVYl8onUKlQiAVTJdls4FMTt01Kc2d
P/QBfOun9+J9nd5/HcP+3I0jpduqhcgg3WE7am8ukEcwH3E0f0R7eBhxl2ivFj9v
NeReGbbj1EZMsnPNPEQcmDuC/LeMarYfh+0UHkNw7aArbHJ8BMjhCfmxoEIZp2ae
xXxZT4RFfM8UOUTVzuL5+PY5azNXiNuoIFvmCBIsWXTZGIuelvQddYozj9tHwC7N
vMtRXfSXVdx1DIQ1PRkq8t+c2jrRjN2e1SVSCLjGs/zA3IPjsqfIIbLOSXXehDX+
PMfzgvC5qqy9IDPUuRBNwBNN2Top95BmlQN10vLxy62wRKb/Lfv1jWegdCZXYLm/
`protect END_PROTECTED
