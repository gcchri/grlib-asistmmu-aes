`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R2oA/O64TdxEKclS0Rt3Bd7O/VrJZsHTW6QV9/AzyuL+9vHvbT0HExjmzPovt5zz
OVUiX/wqY/cgJnZj8mupXp97H1+bWUPN7aLPPtd+ELm+JUEP9QlUYVxWFba50mcR
TNMiS8WJFkfpzkPSn4RPl8lqJe7Zr8txbn1GuyfTVn7Hm/UhoWR63vU3PQye7EG2
vR4zq5eAgYMG5maBUJij3waCED8//IdRNAL+TGQymAB1AdOX7+Bc1mLeKeL/c0S0
ixt0vZTSWF4UG6bX4kgE5gldPTQA5785WHGPi8E2a1UyoJRw9Wt55Ti5izHv+kJ7
q2JQezeRT4PNc1fiWKhpNXiR/y0gNu+5DPrKczTaBD8jpu0X3aDd+s0EdxIqlDZN
5FrbeR1/eksVMijxY+DxU0Y9UdA9ik9l+88yrY4rirXatnTgGaslsBojC5kNPt30
MN5BSORD0z1omUD9dT/PmcEiYnR167jMnT1hPG87Jcx3nZQ4BUKF5KoXJ8J5jsV0
JyzLg8lq+yJZzXcibWGqtGm4W61d0Ub1UnBitMKOCcSdOdJujNN8sxdBjE4Q+Q4W
kocIEUSXo4SWgJyOOvz4J3J6rxIFKZDKrT8fVTc+S6AR7X7cpYce7xmlAiEuXEQq
dIVD4ZSFwBtvKNLUPelyDaklXE3zDpTOJSPHGt+coThoFPgBCVW+eRxAtFjTbLgP
SP+EkpNK1PlAqiiCE+Dzy9hE2vwq/OCvwUDPFm6vVGUYnZjCOBwAOuBq8IOGzFfn
AaW4QfM/hF3+AvW4WkwGtMTMEVxRIWqriPAYCIHqBe9r/fVSYCBSbC+7v8ruUX/s
xkhAtm1Bfi6ZHiYiCyUthKUGzg2OaBDzRTh1UJ3wqaNa9aEJvR7D9PL8sXYSgvvk
Gb8q9cm/UEXyoRkRzZ6G7SQQBXVSHDV48IfPmMrsR69ucwe2NyCroEuWDMY0LT7D
0fOoLAhcy4orDJJudZ1AQHoW8xuHlqxoqpdJwdVH9KSBFd0KNX3Z7QxHYg/F5YRH
e1LtdAA9bbKOJ5yNu3Ecx0upfEbjFc17/M6Qhuvxo8H826NrEXd6KF1/MHjc7l1f
L2sMFxhRrlxwRoRrs8K1yzcn1n7M2cSkbihSHgxBamdL33U3ICsDN2AoIOOclCaM
e6lsJ0GwCk+taT2u6k82l3b8VldGjIY2BqU1y4By9ZpXU4ZKjSkCvgfWqcFY0I7o
EIHMkgzIb9aRYeeAilMidbsq8HDdieag2JovyNp7Wc6MweqUyAaa0QRK0uGlYyxi
qGUJ1nJ8RxBg7Fin4qEZ9POB1qz3CmTPjOE79miS0wR5OaFfOZpBidgZHFL0n0jS
HDdqfTBk6QzKHEhUvfVN8mF6E7rQpcHKl27h0VlL2TtfzKbjPoAGetBVv06a44Ag
sNZ6XYq8aMhYKdOzWn2m3o3JF9uR+jPlQH1pdmtkSnRASjBkL0UaTGwWXy+4ZYrW
Bnqcf7ZQ5iuxKMRoSYggQ1RNT59eEsq5Voh4a8ykL76iWZDrNBX1sA3Wg+jRf3aS
5WGv6Xhv9QHTpblY7er0goLUxWgxCylvLYdHDiVOBejREGSCU27BHXHmAzWdU4Bc
tVQ9Wtb2hQa4v6o209Vjc4dDEDal+hwG2u+CiuMvdnDuANkPiAEbhoup8Frg/e8R
iC1RBY2bgOK1dSqS76ddQjZb9SIKWXWbxVaCcMntHYPUSHdebape9V9fUqY8D5ZG
42pk07hb5z9Ir9d8Ta2wjftvKH/58VZ+RNl2sJPtYHQKr1WbzJ3PHYKBcIVJlngQ
nrFx5PU+KP+8Gqw2/ucGYNQzllktf1CRo5osjTa1OwAMiJXpIAt3dOh8noIZZNwH
Jn4uhdcKR9ZVrt7r7id5Ely7LCjibLBU+DXwqGicu3BqXe6HPHbBy86WpBaoZ6pp
/eejjvC8czRxN1e1XblEmx7gG/O0dFGNg3v3sfCwg9xdeHo43YFtyV3jNpTRlE1z
x8XqMb2rDNbO8VFMzlsfhHuJw3GvJXtup5zscJnKp2Z45dk1jhcmGwMOBWO1kJbh
fUVbtX2dizI/ZZEupA2RSUnV85FQCElzJil0WDZTbOTpWsKKUywdbw6d1aOSu1Us
LpTUBnMtGxQVqGr+JqwvBJrmbrGUUU/G1Q2mG7zsNCK2taCju+imkzC2bCkbapfA
20kRcT9DvRAFGMuJOsKHLUKjmev+32xP+P2693gZGdsiSWWgHCuR9AIXNt94JRxl
cIuijagd6tcn18yY0+bScZD85d81YGFZQ3RgjWhDpomo01J8TUMlAOeyUyvyV+RY
P+NDVrSQS6WOD9Mx8DqcWvaXI9TQTL/uQX7xwivEnZR2kSXkJgeitFjmy1Zmp1JG
kvPc5gnaP7040dnNsv48rnW69VffDnUb8FVjCNGQFl1mOJDxnj25+HaUb16DMoZO
hjjW1L74em2PIJGWA9HC0XTk5fNjnl77Um5+s5Z2xMqhmzXPQdw34YeF6OP0e77x
6ll/zuXjuezew9oWQ++1ElE64DcTyHYk5rhAgE9lR0bOPC9iXlzVkgOeJP6o1tih
NZltEWCnTZPeF0lt1rR023ridz387SYBN01inUBpFxvUbxXSKTs982qbLj/TnUwz
8glfNjpBwOVyvvpJz/neluOz+BTAr0SlvPDlhHXm1DtCOc10T/0kbCjTJZdYewbC
auAHvG2xDo69vaXK6kChlEwsyNuJFME5cGvlmhzHVQsEvWdgkhXVtF451xsy4YEf
PbDMyZKgV3qrEIw9bRcFFDTG1ryz0X/devZ1amHV1dfKrdJ8RN9iFA9rSzlUzmxT
Tx6XTlphrAQqD9yMnM/aLAdx+M7FW1zHQDfKrtxkhWU4flzBFfQ4YHlkgo4H9uWZ
cWzHC4rrVjx219kymmWWS543UP0ZKzc1FSLE2YDfVVfAGnTUZbgg7cwsbn/GxnOM
+7RP/eIHyNvnzHHM7EPgNwDMGxsdixWrjf1e7ifCShTpaYsaPnKDj1o8BqFxwTzO
N9Kj29ACwkjVF8XfLk60j2cX7vbsH9XQU86Dl38Pbj+jhP7uZxJIRb9yGCY0dAWL
Skfz/xsYtZcXYY4EqRkj03R4h9stThXxrwu+S0VPpkDwzbs7WwWj0uzQSPLqzxjp
Hit+47doHdva9kOM6YHBXkMSZbWuyEc7MeY/kMJqygdQQb2TLATHlQ1NdMaXn066
0My+b/uyzvf5L/czoP+8EXQ+iNycdyzEEQjZTZy4LDs7DeA0YIgQJGoRDei69s3Z
ZxJAOiUghlfbpAF4DqCSUFXeIEjqfVV69sT9M/0VqqduFlkAJUoEB5+lMNETw53O
Trpq0KkqG5GWRxHDJX837Zup1SOvN7hzbhz/C8fh/mofsWuBWotuJ/nzpqNgr67B
St7cudqBsswVV/Btu/MVGrgvvO6s+naCR56uh8AGHXeD/2a062sk+UpbyyCg02qH
BJpyJDUbC0XWpLT/ljG+bBx2OF2S99tC3IRBC+crkzhILoiWAElrHKJtkWyl3UuD
Cc0h2BtWzmbuyCBZjobACNrh7r09sOQwtH6B4nvsM5WLK9RhSDeG6xta+atyibCN
kWI9J2BXg/Zm+trNeh2L1xZT9KuR6BE9cXzDlpfK+tWUfYgSDX+DQMAsLnWm6aP7
g5VIOHlEsKqbbPRNCezo/rLtTqj/ht2xQPRj2D+s46fuza+awerfVrX51P4lTfcZ
GaQ/ALHFy0T8xn9CakiQtXDQvMSdOgk00rRBaE31rrz9ofpn4nTgdjXFZlPIxkYW
mniPR3X1PaM/TxNDAkWBO5MvoGR/o7MQXAvfR2W3lm2i4bg9Zh6ZFQwevC6bTw/S
0ICcbn1xP4J5cmbhustDfcTHmR8ErRP4A8z5y5AgHk//YKptB6HTdygNpYimcZxK
75Pu3HFG1tZsb00e2rKw3ZJ2zYKa88ffClFiwy04r/su/E3JDwnQn/xMEnW54VsH
byxWfhwKYgs87OflThICV3UDVUCb1InAyJEccKzeLcIZlJ5wJpjKIQAWBKEQkEy9
vJQV8bOjupeu/CSgt1p0XWOsxLIEW9Zrm+Ei7feOR72+1ujvXs3M1dFNu1rqoDAP
kJQsaSs5OOUb8EakQwfckZ3ffoDL0SJtKwZukLxc6x7WASAZ425+WgXEL15lEQaV
UAVHfNqZzg3cAnFoEsd75ff4nJMRHuH613sDCHlUbH5VZy6HMc/mAYrXosApFT+n
A4oPnXJ17TEtzQ89fCiXicjpGgjEypBiRMaiAoRXeGZm3MWtzo9UfpLBCJiVOSOF
9bnWAjMwMDWzr9rWRvK6zoZSwShVtEI57vW34KZnZcBxrVrXVB/EWlOHmwZeElRK
8EQ9kYZ7adVKDhokfHKxLRot7vuCiZEtAAImppcn4L4Dd55Ap0+a0TfZCcxP+upD
pGWfVfwbNqTVl9lZIQts2WEdeumy3N8UMRXoLFpyD6BCiKY5gjyKEvI8Bj85fb4l
1PBfJMby5vWTlKsNkolSKeyA3RpoVxQkG/WzKAjgq0exEEB+EPdVQcx1UFWk7lPz
G5dnlkH/FixghWYkheS8+B07ovhNXQ44rEhywfxGksHJqfneheDffqYulTDM7+IH
e7EZuQMRvXjEhILx3qi5FLCPb8CfOSfkTs+H3YCLOzKtjB32Tav4DWvd5BVQbmDB
m+KV6RnOx0UJ3G14kw9JgsVOdc5xVYJbdaIjvk5cxjB3HJ85u7F2zN6sMZuj5OcS
R12Secbfmmyeh91WEY4aZHGpfYoDIbyhitTLrX+06RfjrCfQb+RmakksmEzdYFTy
ciMi1rez8XRC4vj1CIfgR9S94T1IHOZ3ODvxIT6xvLU3zlZOFZDkErGsGANrNjwQ
eql9hjsxs3ix7P/LiZ1RPUBC4rn1xNAi2F64Hxi7Uqe+kuxeJHsjjaLNRr6vxF/b
ZtpX4+FWl6l/Cnm7CkNoOrcpiPfXLApaMrDq7poDDSDYWKbJ9Zx+TKTejHVPgE8W
3xy6zKnx1zuDITE7DoeODiK/eLaFV4Ubh19wrMmVkebUghJSxeSiAPKRDO+/K7v4
ELkmprNvj3CbfN/9gGuFcRkwUkyn+9Amg8SO5Ci1T6VNJEFIRnPPhiNXNeyj8gTZ
LDXF0nrXBD5pUZTZLzaE6BJz3apgQPY8i6Xbrm9a+1obtC9RsvZxWLMiRbLy6J2F
m5f9rYJLGmoMnj1B2RgOXX28imjyhNC0qMBXr9X6sRjNIn9AYUhsgcP8DVpH1qX8
0gy1ZJDUKVWJY5SoBMOttXcHAQEfsyVIcxcUyGRlIfEquhdsXy/xcpCxfthW6Xqh
u+SAwIRf2VOS9l8OjB345b6orkghbD0leLT2bDgtDN84mDPyo9Hc42qSXA2sApzp
7E9bCnyi6euBDFx3GV8FLN+dBct5uGMCwqN5XGWOA9F8OVPUGep/WQj6uaEEK1Rx
Maq/TONR2IY5r+sKNTaIl1WgJtijvHb1Z4XzuSR3cE1jueGJMMiQffct7UvMzSi8
kj1G4YV1fzsKl54ZoSRlD7L7wDyBXZTBWIJlKfKGDZ9rGO/es/5Bj/qtwME7Pva4
2dtZ6Sm3wwzIZ363kzaL7tT1CBFf+Vt3PWr3eGfDVtz/Z6zLNtdqqd5KrCZb836B
OAF8ks3EdlYrw58hjQCYXk160IgOWNiAKDxiw/9KwG54ED/VtBIXAjFJkmP6kRZR
yFZnv3qVdgB/h+xGMIuB6YsG9uhb9r3MTC+5Y44H53W0Ipr2C/+W+vdVwFRU4a1f
lSMiBrgFgHXBC7mKS1v3peUbdCCfszUA1ACSsspu04QS5sCFTSWhNKUwq6djTbAU
b7IHaGAWuEvpOVhth2qrFxzCZY1xUquT8iRLwl3DeAEC9MJOP11xyAPdcnRQ25od
MmqG4aPxK6sK77GAnPDViRiK8zwJfbVle46FFoJ8z4hqovzPsOO1iVO0Ec8SxyF/
i6vuJ/v4MfNkATAGwRhrk1MZSwzvhv0CtErKduhkyXDcIhh/BWqeQ9QJgoZTrerJ
W3H7UN3MUFPd5Z1EEC1ibyEk5iJUAFAzNdK88MaVP3pIEzCfTIkc23vCvjL5Tpbp
0yYmNhUgbxpMpYbi7fpqeiqRkW5uwF0xJcGNL2kIQ6ZNsHYz40tkwMawBYTC5BN9
aFiW4Zqy2qxBfvfKHQ7xwPc4lo7VwJogT5IFcVzh5yqqYQ1EjGAsN7EuDMvrOPTM
XkIuOZCNVrqv5bH30MtBHCbY/sy6M1bn5eFEffsloj9jKMkmUzipePSnVbeN2cI7
LFgyfO5wqco37C1vpvXfXGiTEPzIHDDQdoB/Qv8lLffj2Jt3aoHAxpVOJ+2IRE5z
haN0wAGVFQEUeqrk/oA8VpSd4BDluEzBnJV4KGd5xejnGbF21OtkTWVKomBCHPu6
OJTOb2awUWxshzUJ4g61DAt61B6fP70KrVoAhZ+0Ab0Gcoe/btN3/JiKUpgqHVDx
mWcvjkbpV6gEJ+4QEUR67hkjhcsaHglRgnIHF9TUEPpWf5ZOxstnQwitrM4Zja0x
2titu8JMWcDCOadIySXxUjYhru+JwBpTzjpEBd8XdPd00UUPZyJO/eSa0/i1CZk1
pf7osV37zLLRI1IcsbftUwwx1mRbrZ/I5A+Tn0nPXRFKz37F+TlByRw2cKRFZs0J
ki8vWqtyNH60VB1LFrRZ3+/YpQEs2LU6sR0PAS9hZMPxuVEbXzeE4opWoe3MqPuK
y20bZHZ+1kSmHM1h68zvP+7L8tmLMIz/fpqQsjjiSlUubv2rryJF4JaXC2u4CACQ
66L6R0SueD/wKaqUAH/ScnaGh+GOUNilwqa4kA+9WcYd/L0TS6sPRjvyoMiuTwTT
Ejq0zy1j6O879sfoO9SBqkVtF3AnC2oaGeu6RkIsY2OxybIepyY12hwgZL/1LO9K
eo6l+V1EhUWpG34jH0XR8c64ywzbTt+wA5u021Ny/jb2fW9Ux/wHwJRTpXPxH5QU
tE4NsaZpDPYy+lcZOjmRtZKDYsROt8GgsO8Qn1+yYatimaW0Ww3ac7sq3BSOL4et
isxAs/taC63+A2S1e6Sd2/DaYruTa9/0h/O9jd7t/w53DcEo8EGmvnkERvVVstbI
3MsdKitKsAKC7RzuDIkn0Ar9Ne1br6R14uCyOJDG52mlyKePhs70IFZbidz360En
9d4tZFq2p9jN+085h1s5aJGAV4iuuJqRjrpVuoYrJa2GfYqOFP2AgGfCaC19ke64
6imFCDfwnC1R8je6JdyLN7PJScUxAfbVO+qYWF4axiOsOkCM3K9LD/gz3xEf52BI
blrbwb7cgr1Lmn/63DBowJ4+hvpSfQ0K89LYZgK53ei+lMUsXt2uRhsU1kjUafo/
Zyxj4F2f4TUwhFxdpS1av/L4jNu86sY6KII7kN93EXKGlp95d6wBvD2ht7T+yXnK
Mh6aIeeQYQlbdA3VnRxfC2rCRoeT1Pv0IhzaxoJfpbmLXXImt4C9RqDrYYyqhA3r
hVxu8g1VzFTHVjt01V5OnX/S7suLwsFbVkgRuHCnMF9766L/aTtfqBNHfoZmYYuc
atIqIb7k7/Q0XS8CqnWZ/BgB56F3RDri3jKkLlDBe8yakhyMzUGMpB+lceSr1kNI
xVHKyr4uUmJHY2fuZ+ENEJ6mb8bYXolEF7wnFYi0ca2k80taJZSYFf8a/Z2NlT+q
mPGEHdsV43PO9f3Bxrjh/CdhkiAikL/p/QxQrTlfbwySnbIAVp1Lq1eUfwrwuLbR
qrbzJoTlC1axaG6LcYtELCDzvneUzenYhmgj1VQ0nMqZJtFATto/IqFVtfkTAtx6
bYsCHqjYio7cl8SpY2TxOPIAGv4HZOhjEmLLTOmidMzppIz7pmvNA4IXByCF0Gyn
hmBHE0wJZfsQTUIznm52AvwXHFJTFYSShBWyqfoJW2A+fIQzLbh6gdn7GMb6TvMJ
D4scGx3CHIwkr09VOwG57ctabluRqNfDl/nwcLg6xvqM8yksdpApJQ/LoD3OCHeU
jFYArfxMwYcxr5c3B9tD4eFsJrCPOaOIG+98m4YsFwD4/YR1UVL3NZKsIbLgj6h9
CvpFoz/hxWAyFVIxelRnOgAH2b+jitkknWL8gt/jo5zii41R6PofVMCq4V7FKd/+
OeiMBkTR2jC/vsx70T/U9Pw0Ha66gbCKJrcqrdje86058Aes0a5dYP84/4ji7Q4U
lw7OAvtznmV7IgdGWiTuwK5TxBy+B1W8nEdJcvsL16+YZKhAmRHXHY2Yf6DiB0qU
wPyC19qws86qke2R41ZkjzUvD+SE9I2JAbIElR7/WXT5zigLiMbR17og5lJtVXeX
NurVS1Ar/ylvGXiJj1tb+BXpBjhJ2ZxKAyhZrlP/wLQqjfFMS112sdG91oIlaNxj
NT7a49DCG2czY+Lff2Gb4hdCgW/5Btf3BG/GUruj8AngheiTHgYWIdYPdrqlX1kI
+PcoaQEB76wN2D+ZEb9dgx1eZMKa76G5dnuRsvEPTiwYssYYAHP9EpE//G022sW2
mPRqcuIXInjiQvVyeqFKUqaaNU3ADejrchuXthD4wR6cBnFIfQS7WWokKMW2jaY3
ANT4h0iYBCRXErhSxjMfyGB6jC/o32C0M5vb3/kX88CgPPuArxe3OQsblBi8LaRZ
sSee8oiCYTIH2OHn6398VxYzMuvJM85CeeawHIdTt469ZTDsNmTJsFKLijgMX13e
5lr4lU/+zdtELdFRgnsVFi4HzbIKCct8N/HJuVW0rNJgXIiJZ6wFAm/+R3V6tQsq
8Jw+0Uu6II0u5a00CqwmK1o4U6UuOiL1NuYy+x3N3dzaVxzlSCdmKNqX374fxG57
PHNpsfhlnL5WX4lAbcOgfqGOSaZy5H6n7DHG2VmsgzBjXCzkILu9R4iHwBtb9ke8
2geYxV09JMaGUKmTv9yicgO3Kq9hDrIX+Px0B/AMN9yHxLWbPZH/YgcoYQBMeAhl
N+7M2LYmPIniqZ6ZjemtyFFgoZL5OIPEU2WlKkbuVnjazd2LEIkfaAGlC6HXJBdt
Q6PY9h/78gwauBJtsjZshftvaOnwazLV8cZ8Y2KRUCTyvU4AxqsMPUQFjjnbL9Qh
GbAn+Y1UvRNt288uKHNXkhAyKpQOY3S+20N/hD/88HLS4OGjDtVnRkkiRIvBHrB5
jDegRTkd4FqoSOQ2tK81j21of8Y8RlfBx0JVkO85NqdysKXNp6nBwxm/HJbfWt5a
O/LxH0fIqUDkXXwiyFXAoD7ZhP8MCaWytLQTPc6ExFe1682KYz7xGNr3mLZ9Fc1G
Pi/ovViopbqRsVEvIVw4pb7fHWJLWABwpxD/QVkXHPnUuNrrCdcgQu8vxu6E0nbj
woqeIwd7aNoHgkA69pF23+vyfJDlq8GBG46pYSQlkXeRBZPyW9sHMp3WIJ7eqyTm
k8trldPsc2Tg9/J/zJNNgCF/gXigTciQiUwwefDt8h1p8y62AYA7xjF7701azSCQ
QdmKe+J23NA6Phg5nqYPqTBQ9ybYK9j0QllSCUAtxfa739WZt/goxeI8mjUKJTF3
OfpWmklSjFLCbXtHNFbEdAYDXNqGfGc+nU4wToYKu3IKaLichJFw3W9PjIU3oCYi
7V1hWx7DcN8cw+LS/ubTjTistdxLgdXA59UtBJJuk6AxBfPZkAqHpSg5rzb7pnY5
wCRCJDO1Q8BjcThXFWzU37K5PQtIfYgMJykf6x9CvJnFsjZtpiwVJKahGy6gdfeP
Ytn1Z/+3zJqLBfZNEy8u2sQlJs/OHAKKif+XxjXCf8/qyhCTcJsx6PxszArB5RqL
eugPK3FT7yAYcKE/niz7T/hlL27YkfM6aghVs3PCIBbntemmqYGceTKGsTjnE6nJ
gCyP9vDZlELbx5//ghC1LKZpew745Kf/Mb0XhbmRh6lC5f81TY+GBdD2IpxCg9oG
iVfMRxzbMWc53oDw1WUZmOdJdSEAwLDlz2pGMjoAosZ1JnleA9sG3un1RWv9QGzO
OhN/NxOpLbH8kDjKH1vDlK1pga65pZwEQUkvtLe2kyEohCN1ZYf5JwUnFL251giT
R1IA5hnGmLOLEc/6LumnjJVDmIuaAEX+1xRsOboSTXWPJZ5fFpqgZ2rHX5kq9euj
9TAnGSEL7Wi+bUMFqxlMGPUgfD8OPZ57jWu3UPm2Jpfa87SOhpDIsX/UT7Kt2x45
FM0ZhGcHHOPtFQY8GJXYeL19fU1iQxk40AgagUWrmQeLWspqaUrTbanuv9BU8eU3
/4+DksHUGrXljLMZL0drkQ==
`protect END_PROTECTED
