`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q/gX3hUYt2/JKuzlrDSfHY2mCAR66uB3zNrwiw5jVwzFrG184yco+k5SAAh8DbWy
vtsBYl10F1cZpjBAupE1WAKRDLLDKFntT8Jnipn1n30eBH2Gc98HQ4o7xuObIAbT
JXIyNsTYjcF2y5zxjPRuQZTCUvW+7vhl1T8zE7RUyfY+kj7kDvi/xpuffws+cJid
h1csTOFAl1GZAZEKN0exsT4dC7fr/cVqBsVsHHFacuXJEcWSiLjZLhxjdwllt056
pU8nAO6IFu3iNvk5G9ubhMHmyL91BBKo3y+jGWIRx30MkwVlm8a9WiNbCKUb8gXF
NXcg9yC3iu65+PHSg4MLxLTUHRm6kXYn+Iw9J9y+/7ldIPPTOOdwLfTltuIDzA0p
YA6w8fiBd+fa9gg7Wz5iIOcFbTRaS9ZTKBOckWsCqO5uPTYncrhCgS9uHOC4WAF2
qf0so/4fUhvgbN3okZWD5ZaLxdUY1NsS7KmRDebeH/+/OnL9dgKijZhkcye+qdXp
KvkYqMsnPIrLx0J4/g+ki9veo6mC4X5T/q1leqx/FLqWPSvj6IbUtj2VgacfQGlB
aZJsUZInft/u08hViHKdvQCDR+YUmnI9KWa0KovXkvpIAEcCvHcu+idpwLpUI0oO
P1Jcott6bV0j/DGx4aeMvRZ7RS/Rrl5hZEromm35XQlp8nvQpCvE9zrstWCitPv9
K74MvMJYsROXkXRaiJAeRn9teG3T6U4eKVQaS0l14to0eGSXT9A736ukQw/v1g1v
DSEV18XNpXM925PpAcCwTtU+OnvoSoA6uDpJmxTz01KbnoRX6wH98aHMXojaRF7v
lE2SHe9vcKiKv+8fVZdPwNDNWFoNVX6hCQDHb3TiUzvcV3/vQg2oteLST49op/vH
6BnOhy+6vfJab6mKHuEYe/B395MvjJwIl+fhlccUe9DPSekgwEynlY8LdyI4Cwdv
Cn+E9QDPO3rHhbyz56Ad/Rdu+ei7kbrTsr6C0CChPIcmYJ/pKA8dlBj2kD+AeF6F
pDIs4BuOVays6NNxAwfCCtBcB+BRi79rB5DGEESR/b8hNtZXc/5oSz9tJT0MFveQ
q/0apeFy1QwD1bqVv1JZQogOmL5avJ+W3kcnGwrcqP6PfNiSLr3ANzGlGVAY6Kdx
sYlYy48lIlDz90/wqz7sdfqXmASNbDvs6rJaau1G0Iw5jKcpLIvRS0Li0hT3AIpk
oa651boOQel08wrYjqKTWjM5a+6OtrrSIuqUIa5i4lpsLAihdSp2SfF1AzEsPHw5
gGlv8yaI2+MGGv29P/JBGuzsKHLefsBCwS1AZZvs+mjicKQNKL+ap0FdUWyGY0NJ
fjnkKeh4scbRWcFUr9bWDEZdMQgWq37LiTsse0z5ko46yEQMinQp6pcGBTmItHNB
KG40gWAswHq9gv7+ZNXQRsy+hlORmzwyDX+OSlnQya4KHYlN0kZseUpAEwRQ8SDT
/2RC/axOYpdU5+k8IjV7Ps1ZNjidKB0vTLIsq5VuM5fFRflCx1VXuiAUrwqPLV4C
pnygT2P4hRjxY4WhmJ/07CJYZAccl80fqOrWoHJDTFiCwW+Nu3LSyLkU2XOttQt6
9D+4AHKO8K9/KgS8ocsp6wfw31cPRewXMkhBL1ybdPFu0H9/GAE5S/7gJDiJYb2s
yDr8ePDdW7k4wrvxsW14usZn2LBFvQaw0HBjaivqxmk=
`protect END_PROTECTED
