`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QvgnJ7Fi18Y2PRBLvHVccBPu3WlBENWaOFSm73/IzZ22SptS2f/vbau/eLSsJj8L
1olLcowvEfFI7875V0PJxx6veh6B8uxO1IzImngESh/1CxGVM9TsN6iwVenbR9Cf
TUR11zhDC3gJHpTGS4uMzJlzW40ESclS2tALMvv7s9nevxZZzFFaEbZGczVvn4o1
ECP83ob103N3wLk0lrGrcS4jDewH5Bzx47snOsD0EslFYGtQOq64j7U3CNGuwFJ5
qCrc4gS8lxOgcDLJ90IJxsBV7iKj2tr/f186ICxiND59I6o3EvCb9xFVlVlI0LmL
gF8ADA4J6mOt+Sjhtty22GVEtno4ijsEU7VQU+kGotz0nrS/Hee0TiAX95qtLABe
82/0tv0Vj6jMvdJCGCTu/PaiOsnenQ92C+5/HlXP/tA=
`protect END_PROTECTED
