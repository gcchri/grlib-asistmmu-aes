`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SkQbIXO2tcs+m/V1vgh1HjLeU4Dys6Ayx57gEo1vM0UWfgrjEtUxMoig871ij65k
l6KgwjsCja6NZvHb7lUzQY/CSVTRjJeEUO8rQkLSjld1Rnpgs90x05RTNw1xtnes
Q2y74J/5OnU9m534wvxxMvyXtC+uR+FAd96ZAxc6qCV2AhkToWv0TvwRT8qm/VQc
oMzC99Jn2p5x6ma4vHt+bD23Hp+uyopdhio45/jaWt9zcy+fve5mTVkbM4ZlAChJ
mvwIHmDLimFqDFoU498QO0+qhH1IsLhOhS5TNmmHniv22sl2gMcUHO9chUq65UUF
S/ClByR5tloTbRWN8ao0kBu4mgOnl0LMnHkPJAgATGTAqx6+T3At6d4lb0L6gVKn
7QydnrEMtQtqwVKiTTN7FEmr0/K4UdMAN+AYwZCcOV3Ghr+9XzO5Z3dnUzcrpjRx
1E/8LJfBTpvADrXSvESgpkjk6qYFSv9DxZxLCxRL9h2PGXPnSzm9J/Lcpxw14UyJ
DEH01x3kZk+C075lqY9I6DncM25AsO23AOQtUiYCKtC0reyodFjj+Yh8ykND9FVK
CfKi5hhHgYXb7kGONC/9TrjRulKz83hYtDOPQ5vCp13aM9BLtya6pVHhsQJ7Ep8O
KlUO1mn+trpE632mHYyogM7xaSUBG7xqz1eizsjrDCrNfg8V4+gDQQ1NQc2oBTjP
yz4s7ZPNjOD0v1P/ySDSrDlaqRkvky3lkKR+WgUzRSL+kFSpuCjNcbAKxkHTy18i
1vi2RAezFijaOwmDW5tfpeTJRYGrVDAre10fLQg9WNcKt5SSE9Qt/boJEBQ2/zI8
YrRdra/wuMJ9cLcKUOL94T+1t7xvQ2c38tu+vn2OST9q9xmw/1KQodKs1gfapi89
GZG5VZZvjrTeiZgYh9qgig==
`protect END_PROTECTED
