`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tun3z5LhtMvCjcJkWijubucHcuogj6MLTjdtrE/BEeNYdaTJqbwarosLd72MSkiU
F/v5suAhdzK8tE9vIc9sHE3c3jUFcM9rPc77mKYyil9rDDekKcnze81bpfTol43t
w0jetD7VGa+13gaAPJzO1tcR8sCAbu/LJASS5Qhn7SX+aPkeeH7mds3A9Xo0321B
r4y8D+yMEDPQOYyWn4TPOmCA2KLpGG61XWyAajwylLG0nwLCBxh+SdGypxDGgrER
wIFgqKfqGcojmjaLrjQcUVERdVkwfJw4+CxbKA+pKNw=
`protect END_PROTECTED
