`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ARQMPLkkqO0L6ldrgV1Kg1kpDmMhSYDlaiY0WCUhhhTkzQiiNHdCLGaicrZwqww9
pP5NAK7Xp+zl/jmvnsPgSvfsfQDUK1Ht6pBsNfpDanb9YW2sNQqo4uzng8jft6dF
McTbkSH9/6hqoIEYIbTxddQjfnMzhZ+r64TQoWsQR6u9EO7f3ewwgmXIOVTL9u7K
AKc0sQtLDJoLUv5NUkec7P2ZOabmIcSe+bwRV6zBC/A73eFWvszARhPplTD3UzTe
xLm+vzKjHnR/B9NPlUffI+viPytFchMCgxj8L4vCxHxZBc6UT99WMXyfJ3HQs7xG
AzZDbJbJqLkk8taRZDzGw28iWodTrI0/QxuCxPeTAp3+g+md8fF9KrD3CqMcaYVn
S3hcEIXQSYvrcIsf72uGHEFGg9cDdu6ULeeZMcLWhgLCLR1cUh2vx6bvJQU5t/Xg
W3h7Rq5gV9zKEU3yjfiG97fI0ZcjnElQJvGQentcJ5bUn6tRGvxyoRMjHLXBxJl6
lWt0SkeT/yosYFhcR1PQYn0o/xFQA//Qp3yfSL1lg0/tXvx60rL70m9FyKpwyIcS
6p2IAobOgIN2yox9Pyh+KPpuEKzQRcTeBuMY3xwuyyBP7GZDd2kBLJoYJoU+bzUe
zpy64vwZYVTLCZhHuxISDZ216uwPS1aOkSPu+Che4D1len6GAQlo79ebJcvofVrp
lnjRZp0XrFqcwgoYsbGpt7ou6EIc1MhEzbOf/q3WMdcvoNCnRXiJnhwmo9U5B3JD
ULI1CmuSXcyGDvCj3a/d+GT1dDCQT1/BAVUfEO9lSAcAOvakn0RzIIJQNUefPLfx
QbS3YORpPmc/RTLQ/m9Ed4uziuXeEd0+T3nhJZO/yaOSWtm1FOJ668uAKnu/ugNn
PMQrT3os+PwEilk5CuqzSHbmVdBb1edcLUeZcjmc/pm+XGM90g1iGqIUWX5R2ouD
Pxr14+TrVv/xgBF2QjFrofPReKY0TvbIddgNg+xfjvljENkBNIr5XV3dZ0Q1Er+7
iDnHKDM5pzoz8g/6PesvDYNX8FWInagQoJJE9CkZFJinCi07UAHzDrtnfhTlULDR
Jd48pDyvrsJ5oR94nC2AfZ4pa6BNJHvGANIaQENCBGDS4azHjHCeMwxwC9K+Itwe
ZtQTVjTgrUVeu4smgU7LyPTyoaCDwe1/EbwmtfX27YzWHYQ0N2TQLQCHFl3/ZtXz
JZzGKfrhwpxYmzSYLKI7vnSz7fz5Tt2q3Q6gk849RpAYzYqfOU2SPF91+sqz0QHW
IObKKsRVipjtVSJN1Lwy7eXJEhe4/KTrybwyvAV8yHc4XbHSgz8+JyUODJ1SbvG4
kU2wyXArE6K3dtlm4EBAXVW7UtiYzxdjtpQDoJUT/V2VjfMmTYmvgDlTdtui8JU3
L/V26KPxBUN+ocr1F4alDY+id3oe1wQMvgtrh39PP7L4+UCBIgibS/usq2jdMKhe
jBR3YnxeucVJqxW9VstOmEYopG004X5+HBSAJirB5DWMQlekIE92SlvqkYQzpzUZ
SrC1Y8yK6q2Db0/0qSJIX8Zu8QVXmifjK+7E8YjAdrlaxJVPyyfLLn1L29z9ExL+
qyirue3VJr7z0mJERR6eliLpq47keR4g/kkRKyGFws1UzYKDIwt9GuxpkKT2v/PT
99jPz9pu9BAfChwVZMuxtOsffn24CTisyYLBT/GvUFJstc/YDhsXzNg4n7SFoDHD
Lfhau+Elh3jyIzyMV1HSHnKW/CK5WhWntZuIXPtyARvyQSdPMpCYBBFCbT66us45
uYenaNAAEr2A/iNwE69l3NfpJwAPafPUPIHLDpXg7ux8Snstr9uFjlP9fI0q8UqN
uLoBeF/jNcUkeu1gKmllmXN63CQlYSQHxZNvpwtcXlawg324t6bHBajVF+ikqCiT
8rqpVb+ZjHTuH4qh8TJiJ+K/FYozW5sf6Wtp9yG1bCVRf7fzu/VWe9mpbEiUGjR7
Z3/f6t6ayNJh8CVjzgr1cABbFkcIl2pz6Z79OToTa7VpJMOPwoKxSsbY12/GUrcS
V+z6eZOeWyyQNdTvKaWdThMN6uGNFfS0v45V0uMl6aZHQ+HjkYNC7imv3rXBD1i5
uVV7fi4kEGRyhV2hpeMsL+TOkBEe5bf9KsIqGR3v1nzwwuJ18yhfFwel9cpiM7ak
Xec9fg2NO/TltFgEegSJL+bBl6OHxO98s+bw9brlAJextXSJFpBVCeT0XptAtEJ1
L+CHAl+8MiI00DLhp7OP3w4X0l4i+8oVa4UQrakEl4ftf5Nk9fFNvHwjbPrOcO2h
t+2o7q/UeackmTEa5XUELYBtessRPrXNDPQ+rFmG38Ivn99n0XIUY6bx4zomicRy
elTn8dDtZ2z8xSj7wKAOYrMnQBwdIaWNGe0s349FYVugxu9w6TZZ8JWsF/L4nsDt
LCpDR+sVkWApNKWJ+XbY1pjpRffNklb6bNljqvBRWkpB3ER+0iNglofnqT86pgzw
cwy1M1YRcNBgwNC/+0qcljMGoAqfVgYWavBnb7zAuGtWcnwlUZJ39fqDExGp8X/z
pwEIZVANGg5VNSRwYpTpf4Ewn9fthhjvvs07GBZEHQJaz//7LpLRK4I1+nO44x7v
qqLubyGbDsL7QALqaZNXODSUhhzZvNaNyKlNIFMGN+v++G188c/xJDlqjf7uPv8T
giq4mf4tORNB5XTewr/MHps/RqbtiTjp8osEGb+BNDL5Wfh+ClmlxCiDHGKj5Hts
rxeExTw/GFKKyYc/8oSg3TmwqtDbXyRQxScDzWyFERXzejRL4qmBROQmmBLm4VFI
8x+Iz+CYM4nJtCJ1sv3xC8g6/F7xwmaSwJUWlIY21DHusN6kXTK/Sk9cMcm8A/nt
bGNbBwfoKCTRGknKScGa3G46ii3ZjTkhxzx7/oVPU1kh3b1uOxQ2v8rcARXPyXb7
jcXASRp8VFN1ECuzCAyW8kbMq/klZIbT6QmlLwVK3oSkTnmMYRZnnwJegm0XMXKa
KYq3ZvfsutG8x6zaMSil/1iedC3ZtFEdk+CEvDhsH63vpgoYynLawI+lkXLSqEpO
dF9e7zzFaWa2JJgsElM+6lrIjL1KO3qSC2R45tWHO80by5sF9xKaGO3067fLGl9W
PnP6RS0Tosp0JpCoSWt63K+Wyj24la2P7uB/myWEsAINZt4bnH3FlG0kDU9b7E4n
PCVPhoZsUdVna0BFQEhEygZiDETRpr29JBpbngOa7Qz4GLFKqA8JDdtzRMqL/SJt
RlcVrYuUb+PzL0ti0MwQ+pkX/a4kX/RSjWSGPWI3n7NnDqrCQS4kvNzPkbu5Dh2F
9UvnBckiTXvoVzLkKWPe6g5t++HoOfajwH+MEdYMnt6snbhRzvqU20F29aBOeSO4
YgHl7AT4LiCjqVJakW937D9PiNI8L3rHB7nX44fXTBpcrRazPcMQ3vlMN2tON/ik
q9y8uHDhfGjzkaQCqX1Ia90cnZSuvEm1wCkgkEhtw/nvX6AGaGAKCcToDuMGKzn2
AXBFige/TOHenioQAmbOLY/VRaUWj1jT364SurCaniAJk1v3uOC7rO/6Knp/z0iZ
e1TgKOgaAQASXQZjcEJ9b7Y0EHFsXlxfly+k4jCww17MfgELdXHn6N1z3FDKdLEF
VqMeOTj5z/rXSfIKPG3zDHHeBVIMfLZSk4mIWoWsxvyUpnkV+oMQY0baAML8dQ6C
h307eqk6dpoPu0eSbMbnkN04YKTnwJxU88/PaK+AxJYie9udl4FEgK/Xxuj/tkK8
dDvXv4b9U839QRVjHUrj04gOZ0JhNkJBhNfu5ySygCbDNOOgEcocWH75y7sA2U4u
1vMQoM2+oreDqvaXgLZw5ctx0ET/vwyUfcIiUSil3X+9JiqlYdT5HLdIv9cB0hzN
omb9lnkPW4fbD1eolkKCl22rM0788/Gwg18k0JC06y2d1M87EvaBuGj+Pqy3gYl9
UEJaAD2v98LetN76a4a9Qwobo6xwI8+dGixCcNvYGJ1FcHo/UeSvGCVinMYZ+MMx
C3aW2ONyCqltiTZBhSlykHUmiH567muuqimgL8mLOx0JBl8PEmnRX82IePjzyDsn
dqAZp2IehqzqPc7aEeQNNznjjnREC0mvqIyYBSuZ9GKb31krc2tDetw2mTGIqZPX
8YGOPYqJTgjUk6owEpMNbZ54tX2tIczOVjhAL4iGENtfSaqfqwjwCzmwBz0sG8kv
6ru1tk7pdAJ6pa5ehz7yD5GozAxmH+mNoTtdQXhaBecxiqyrLSDzTqnh0WbO99dn
KbDVD2cr+xxn3Xb7cJOaHnMQ5UnfGEKNkRF8ML91LbGxrEpJHLXvAhTN5Jf9RVeP
yZMrOSgr2MkbS9y/07fsumMnFBF+/rwQRPzbsiN4inJDLtdFdg3B6y3OtfH3zQkS
2GTtOfnpXm/tXTvIsisNmaOhc/GQwOsmfcz4IErsUsXBpJ3sDuAIAimnmLlw0srB
Qvh6n5PfOo/4qjApBAKw5EzODTiiVcsmgFNFM3jjgSHzhybWkYH5JB/iSMPiWcHY
8fiBh+1cHZkt8cw1a1iHiXWnW7Z7XYAd0h8nC0xP4MZtEYqLJqF7BC39MHksyv4a
RBuyTMAVoSa+jnrte2gp6b1Z+8CHrbPO9F/sViFAAeLfoYwzdMx9/Q6MtGOa2iZz
Tg5zh7qhyD4Plfd0IpPdEaaXTpmkC1GF2ryagTTQMdyDyIoTm0lAdlqcoJeapN5S
+GwlhCKq0V7LVEvhpjliWIq3nDfEj4jUIDFyaIsxnjkB1xmjwz2X+XISaMXRmw5h
nYlHMnFk2XkkAAaXtnX2F3O0hBL8Lq2CL35u2AQ+tCbPSCCRB5x26hHSaIt4x7na
J+vRYay4AzXlqlNoS+knlzqcWj27EP59LziM7zpkI6FBWiE6LHPub2PQJPGYAz0O
QvJzIwM5ILm5bNnobT24nwZqehcJZGipxi+PRLnFhN2pUhJ6lpOgiBx5UjwGjtur
Sqmcqk5hELGHmCyJMFtiyfk1sI+m0PHQrgTaM6tMMKP2bC2eOzeE0dka/XkvMula
VWU9BPUFLIFgG4Zd66ASXl+JwfCjh4pey6xdiQx+HeO0GETt76ps91+Y1XQEAbXx
LYqf1c0HTLO5S7nGavG4u/LE6V/T6UdexpES3mmIbnLHly6WKcfLKsDujkCnUwoY
6d4eLeegb94xmDuFhfT2vJmmYpyq7yTIaGXha7xz/eTDiHFjFnvDFoHICsMnVgwk
B49S60vn29GmTjHD4D9mE2w/C2b3wVHJ/SD1r/GufCPK0EAiyf5mIVCbVe8e0Id/
Pn5QoUyvgbQW1rDRGTKzSJXtbb9ix6vx+45nOwdKDrgrAxurrh8FqkODtoXhjFDg
uyIHWKrjx0RnnFWKec4mwA7fl5GhYddhxOcsifIpQXFjPqnJm4SkqrxaZw0V+VjZ
xkwfFdEqhChdi93CYQSYPYJq2FC9r7fsGNxmskC0GCXF85Lzc/TREsoIjX/7p1ai
XEEYBjcnLD/T/lvvTJe9unfkzygFVPKH6GfOFRFlTQR5rkvy7o/fFds9cwgfdvZg
mL90s/9pppPitDtV3NYglK3RtUcsNwQycWofJUV/CgbryDi0+Zpk9OMs1sVpCHun
XtqsbHgpolqmUXd0NbKuc2ig2tPSJm49wbukQ+1I4uq5GGscJvwhyEBOSMl8849A
La9/gmD4nxgYGC0D4Op8wUTgnjq06fHKrBV3BaARl03sajRHQ56wUbAMByJOR8Fs
pqkfiZCjluQojIs0Rv6wNpWsVSOps4WhWUpajWCdE5w7k59AFiRtxpWN9O+PFNQl
XJKh5mHJZhLXFJTMT4WGpmzIzvZn39JcqVfzBvRu0alCcSqOCiNCrk7XSo9y+o8R
xH+m1jyxPOnadOndM5oOj2B7wCmnZ9uIskGFsSkI+e+svfZ0fi1DzhdSaKwkx79x
yjsA+FXq0eLn26sMK2wg6jCsjICb6pGSgobgNaZsRueD/oNlm6YeYPYUwUJPlHyA
Ved7ihBYxcfEvubNaBaoGi6pYgrg11ndG47JSsty8L0wJaFusGlH2qGwDmKzgNP9
EbXMbiIsdD2Hi0AopQesUpb2+2xQtiA3gD8bnrdCia7CQnMOGqsvxWgGlWc94zXS
DEoPzpfHXNz11DSlGxDz/XVkJTTaG++wzYdfa6adaH8giWChE+oPBW3OUzyWQHSk
jgopvBHbAExCVZZ9c81It8s2XNPn6JwgtHsbKeZx6Da0zUIwWMB2eunIjn1+DvUP
rgKdbtFaeZUqWpl4vbJnBaC5lT/AGf9VTSeFTLUe/vRPB+RhjEia+bX8KeQD2fwY
jjA1dg+f7a5ZmwjmlGFFYJC4vm8+uVksHeweE2VJclaswcsx55HEsnb6vZPAXeIp
TwRbXPkAsvLTHKnvTEIFu1qbDjEgVZ6OqMiXj51qp7VFm/kHlXD0YxK+WSRF/3TF
nSYPbR1TMxBBrixYf7a1tqFvTO2OH8oZ3Nzn1bsg1x/LaUViveLqKMRaavqwbp1E
5Kxbk8mkQgnTP2v6b+T4lK6pF2Ck9qaus3pwvQXiTfktHx5l5JEW/0AENt7QqnOO
KQp3G0ynsU4QQz/n0tf6470fi09dmPmtHaS28j/0llyQ8cd6Rh03Na/zI3D3PCpv
nP0Rq2DSyXxAlPTMH3q+qnYBNTXlJBzYuBNgPo90ClkjO4ULOfPfB+k0CCod0p2k
4jEfmjr8vY1AYul7yrLd4wfoWgZL5qS4QpWTaY22RoO6z7z3jM/rzXHeO0EHmYMf
lV2FCiss2fS3iWwU+Hn+azrlDGlujzS1ZpV7Kzc6RUm4QRapr9Ir+Y/OwRQkoxEM
mniJ4ofsmF8Emyi/254NrNqfPF8kf8XC0YfVlKLRlFJzxoms2s0t9LqF+MFXBYrU
f0jIPmtzeG961VXPqkZTUrTeqo1DcjGCN/ra4LHgdpxfkpnf3lNqgayJr4r1XV9K
b18yYmCU9YQ+CfvtZv/ONUfD3DgGo59zROKNa14dYW3+HhmXtFSDW51jhBaM+NHj
wUbr1NT3VgWiHMSjjPpyJHrxipzll3sBRvNnM9yLCK93pzT29cVgRyrDHA1oveYx
reZYqjoBy4+leXKZ830yM29Ofu4rPh1iwO1X8dw1zWqFx/zG5l7Fx4DCdU4qqAMp
9Xdl9LDEgz8FJZOTYm8DjheUW+82CZUscl3g8YTYmN9E17rgG6DDzplAZwl6IrjW
JFTnQB8pxOj81gYybqFW7oMgh6jfc1YE6dmsr2HxxW/00pxjcBie0NtJzzoEoj0L
KSfrsaHh90hERHEGJVdCPoF59VbPPgj0roxeEOLC8Jrwcs/gvMvvjliA5P1lnRj7
9HU66lEW5pk+Q3upDnwU+YTB0409pT8eMt1/i4jvxMuHKw15DI3qh//rOIvgD3/+
UDNhluPF2lTjdUZJNnWHrxRRQ/FPIIfh7iGhU7KJEfspo6umkYpo2sINtFv+ZQqg
8MkKCGa/9JhFefHin81JkSB8ORHSWgesF1sB9qaH2IB9QwVBov50YZHSniI0l9s9
1zc5V479ejpDqR94wPY2CbHED7GdNg//64decKFsUZXTjoMUJq8+Va/HbshoHZ0x
u2rgr1dV56aPyl15f5hZZobs2A3s4xSZ5nDkvAHd/RelMhsBdx48r+Pq91DljZyF
A16ycDHVWvM/hrFMDnASZDvC62DAkIqgBaf1mcZi912gd0kZG+/qb1xxRDP29fHb
tq7lid9D9TvDTcpbFwSKPWQ5+9Z4CfjXkARQUKErFzdMYdTgmhqXXxb77oq6w8/e
wEVBQ6fahjdUIitcOa+TFaMY+I4VwEKJxtoQGBSnj6hZ9lzuHtr3lasKkKapYvI+
I5IWAj6Q4rV/ZTQfaNmLn5h5pvzNUWJVKWBOGBRQXc0twKWb8oPnty9aveCjh0Ou
QwXXFgCHUt2vprmd8DX3i2ZYukmWyzzu3ZV3e7CaOuyre0utRKi0C5+uYMnxPVoD
LGcTjyKtE4sH4OpDCpknBF5qgkJgGIhzLW8BhbAyywFatu+sqwQNkHNFXQYXa4t6
eHt9fByzPWxSNXsF/m1PGXvI/Y3sMxLGzGuWIguWeXbrrLPNSp3Qr+4Y4LHML1ti
Rte6ozgwGw2aZyr514DdqO23B5me8qTfBjP4izE9x5DDd1Jhd7ZpgvDPcq+V5mX8
0DG04uwm+v6iPLhb9/i0zL/v4SRKfbfXyAoYwF8l1/txIvEYzvejpyAGNdWFSxDL
iJDnCDjEyR9GH3qECDOJOBWMjftpAXFPBI65GIBfbkb3aPk3/n1n6diUcUBniod8
JuYP5jtgdlZdCs8zRCpDvn2TJbme4sLAZbfAia7P+eARUXS1xHH5g6Qtz8QZ+cAG
hFaFG/e3lBtuY8vfFNkh38kNHEOIZpXY4mkJKm8vLyo2nXbTcgBcpB/vfv4YFWrf
pzbpBQfnLpWZ/7t+NkLbyadR3Bq2C6LliM/tpK8f9BbXCLO84qXcb6vXNBRn6bmi
fz9ygxRMXoaN5lekuFXWo0ABlrAhjJ069uwJ23PB0zJoNbK+I7mY09iwswPKQHgS
Cirvfzk2kK1iUxR86C/b0mxOQ/+j08gZrksO2sfw1w/NZW4qbNJQicoVY+k2Od7L
lTwhNWZAu+iDbJTnyKksIMyyr8FCxG1cZxoDhf73E+xVrDbfQTEGCDOvxl+oOnhE
Ib+vxaVEtKFYhlpmr4V+qQdjvNot4i6t5qlKgJ+TiRgf15BjAQNNsbNK1ykOQnzM
IMB1SH4jLonNzXw7MKM4kVYd9pJQCIbD94uWbIVdbao+La4/kdOWvBuHW7Ws9szU
ZlE9PfmiL/i6+ZgPcIgGR1CR0WOlRKnTCwK/xrE6qyKNIk95W6+by+9Mhzm6uB6c
O1/XAo4rJ0Rtu7jkt0dPH6hhpQHijiCiEJ6ns5JyObXcGGXXpiyqqpBYanX8YP/h
9rgASB1RTA3PPKuvOKgtDkzRESUTdx6nCw3qjkOqi9fzNJmPPcFNpp8Yp2kTesV+
qwVjUmXo0dKzwLo9s14wFSVxZ9WMESoxkn6uUqee3AHBOW3Gfyir74yADTIj5AHc
57xBG5wSpHhsxvZGs5O1BoY+MPVR/OSiu1OVj3JCfANGaEpbKmWQOvbeYHr7gQ2Q
cjQ5yPCLwyc7sYZzsev/2rzD1cA6ayrMmb5ZohX1CssqoQ6TKWFPxTt7wBQ1SOUO
7xBkkZF7b1aAc+r6G3q+ScXo8gFffMcecyqsR7E6CUk23y2q+Ya3weLwTdn5sxM1
juWqf3NLLgdTp2zfn84VBtmFpNEtjMEMgzcxxPyyXX72OCPj5EM3YqvXyT9V9RvB
ZcLKYXfFv9eDBCQBzvb7eer8v44ZdA68/6wZFM1DT+GibIPoKjZ5Tj3/TEbhkZxl
1bwnf13gbgP7nYGNDSFYgqvmXf10W7K0k10X6Zx5Dpan/2bVKUUIMc9l1Te5SC+g
RQU0J96GLudk0jaiCJA10Gs67+/CE9XWWN6A9vHue0PrdsmlbDp3AeQd2Btnunfj
ydBZqKNg9Cn/odnv3KLhRtMtD5N3vIs/3YUovvRy5i9CKjKnD+o3FkqaaiB8qv/a
AgF+wViVTjbZHGvasz0BfMKWlNhI5ExYeuWe54JNL3pTZ8ZQ2fu3BfT5EjXbpKzH
EBcKSGnkIdCyEDETSwwrNLXUfXcwe4iZC7E+RgiCZMXa6jPBWD+RO9PjpgsWsPp5
xa3rqxjTVgW4xl6kPWo8LSuzcKTsrQYUeGDftvedD9XAo9/mp/Djv2RuelZmHLuo
hq9BQSS5FyMQyrbZI0aDhqtbWl+/Ey1Orr6RXrhcD8nceas3SufqTaAPRFuD2HAh
5VtVYyh6rjjP9N59WfMorcXDsR+9t0ic1yIaArltper/FZuR4biIvRKCsRu15blg
QhJUyTxN+FvznDQ79tOXJNmszVQFz+6erP2m2V59OY+OJJGz3zhkJIW1PPNBJIuG
9wLwrFLvy1/KU5Pd7yvm15WD+Jyjt1kmGXLIBfRvGXzeW0S8LIpFX+OazIQ7/RfE
gmC48nPyL9oTmiimMQ2rGQ/VNxL46N+8lFQ7ofPB9IJnvgFZMzoxOsaKBodHpxlx
iTtvJ9j+vC/m5CsE2j728thjpW2glffZ3zI8oHB0k0ZNdFQDuN2+nXLEGXsObxQN
08LA/sOBrUUViQR2vnccMOZeoZy1ze10EEWxLBz5uHAxwQ6rdzbZuZYmD4LNgZ3m
jB2P2BQtZx5Mo/bHsEwSMrDJMt4ryMh/2bESq9qrWSF2RURIwR03TlndsJvXZZtp
61dTiTRNqNNvtvAbPijM84PcE/fv6AjnCfz6Gt4v0i/E+KFHRKETuZ4hggVkaCG3
3fuCk0eNI8agM3vzNtutyMGMVN6OuCrmgeFCt9P79ky3sdCAfwKyI+055QoklGhC
qTZeXNUjvn+ggNn9FD+FkxQv8W0RDueEoHLCaBlZyidwXRtkZVysPs2s5TuN8xvW
tLtNJ+Cxh+XyQu+NiZi/23waSTeRzUsJnDcYFe/N6/VSNsmZfxYE9spyGC70/HZR
tUnl7R/5wEivSiYgKNUAN1AffxsU/E1WFtPYats4LVDlLZPSoqOt21kTo20EZ6am
se32TJFBo1tLZnBKGAdOL5kRR3h48Ga4fMy8dNMt59nG9aDaaxUJFIXU2jHj6n92
1OkAJaNUE6WBjPsHvjR543ZtSrWS14F9pRNSU9mP0KONzQMc0asGw5i9rVbA7AIy
MTUWCf+Z/IDUO8bA2hqSS8KejdwBMN4t5AYbLhxNPGlWlrImkUHC5O/UX1RNCxRW
NbDo0gcYgH5s3Y6oseUOjKMfiSkW1D60J1w+b2LnIGldbzyrWyG//r3xVH1rWnDe
Fu95DBJVQSUliI7eEhYShM0nAgp8JrCuV98GOpNK6qaal6n7yoOHoEEMwWwHIcRr
9C8Tu3Xa8cyHSCTJp2Yj7k887eg+W46CRTFbx7zWFv+7Fludyl55nVPnAilc22Tm
QZ/Z3I3vDySqSbjUjG38JA7GZSWq/GLobx0rlXxcc26txrff236/rbnCZNj7PX04
bwB95xbRMBZyzEVZDrdsNZN5fKDPjLUbe3n3ohbVAUWFW0UPSjFAcW+goSihGTL8
xWkhKxYTF/yX7g59IeF52qbLXtJWMBVRhorxbB6+0G+v3C9afQmQXzM3ApF3YciG
7KwmVzwIse6miqWuqr72zAeqAgawrUBJsWztXVA6/dVhRNbwocc1HbkdvauW0URG
k993rDA11OvW4XQq9YaXBdk2zmDO2UHwd3GHUJMGZ77hhHrZwBO5QDvzZAr/bHxC
/g9phIxd+lT9pLERCSy78gn8h3LtyJZmXaxT4svLRn1oGXhshSlC6a75/tJ57a8D
nV8+vT2JX2SQjt+LSrCBuN1MdbUK4BgfeTLHmVhbpDcWI/abNZ65jp2i5OTr6OYU
WzGvL7Syj5+79eHiRLhekRrT3OZ0HbaIGmLbFnI6cL1nCEWPw3DCmsgoDseuxQ51
2ANYdzJk6yzDLOC4JoM/5owMRhq7ODHK3GC9ftrJOuiQIYlZijE3/nI8rWKVxEm8
x3lEUnMQoZ/q4PQ2lVfYKwcCRxOYe4p0ibrfHwXYJQnifJuALcUm0UPXlOHtzla3
4fFuESJ+iwl659MKqK6zynUZL8Y3nDbiRI5KdOrn4n07Gir8B565z9PeqDPxyqGw
ryzZG5nsV4Kt3556wWhrpJXJv7113v8RL+dNghTeZRb3RhRniNC7BCzUes7lkKPE
s2RiAj5t6SIzn6y6W1k6I8fNujkZ4ML0lFidsEFMcHLKxbJ2EOUqEvCR1vMB9wfW
/vU1vt27Rm9Owd1uaZshEV5D8O/9VxABGv22/s+Vmv5LEQH2cwcz6JghL9Tiug+A
m+TQfJZa1pv/HuaKuxG4tPhrV2le4/7QdWZ+FNhN8TxxxE6naYDaokLmjT30XhSA
TpXXAmlhMECbE64LXru0icgPjwHH+Lm/8UeaUDFqwsC2EB7VM9gJpvuTtoHdKVK1
o+xG1+UB1ULFoDjpaNEVcLK5KolxRqMIUNS+kLaVifttn7+skrlLuHOJArO3NA6Q
BMEOtrEHSCIhb/rEz65rvdhyAiL68h8A7SWu28lEPpB9wa+iwJZx6MhT2nj/48OU
UKzr4y/LgXjqrKSn9LuSvn3Kr6/5EN6cGSas0Umr8/UnKbmJgD+VXsJWW7vAdbLJ
lgB78aRsiRMnGp6LKYlp/GS8wzP0VsXj5OEZInaJPkV/N4yZnjkcQs9HZs7yrXZn
K8WEXaj4rvpcOSxpfz2xE8w6M9HjWNdyFGXklym0YsV/p3UbHSF+CPBAjZuMYasp
julfuGZDtDazt8PLAJQMcjmq6sdLYGrLjp+w0ce+w+9+5/YLSjEIKaiDkQ1EI8cQ
Sr5DNXyaHZTywvhPFOGGr9m5N0bmhg0w0Yv07rQHhqkV8s3T1ldRhntKeUI5Ay4Z
WqTHZhv2oO1PcXd7ZyyiP902Ak61pUMIyPZC884NFUPWFh2BRs6c/21qz349tsuM
PDfx/Q14Lg4hNktZvcSapEE/1VGfRpjMzVH9/+tCgkcumai6uXCym2ksncy79sqw
U3xGCxhg0uyimb0q4R7oCIl+QZo72dBttY3N55lFz4Sn60biAwRE0gjMYWmVHM05
0jEPDm+koAXEX8ibIUdI8mxjdmI6b7doe3rIZIMpJXcoXabBirXoyvBhPC6kqUcM
rjJH80w7Xhzs79/92NjZVmqwxkgaiTyzaRU/q9jYGtExRJ8LNUXg2uP2jF+k/1/o
tOCYGZarlOZWgQdiwPlDO3CCxXDcDBsvz+plIfUeZ4kkqn394FxdRpC1rcZHr6ON
c0b8TrFL7o1gnvXeHoPF5z5nkHhxuj7CNbRdXS2E//6MOdwGW4P2G4/JM9n1tBze
kbzJPacrrv7EsSftIZ5INItjkZbdTPq/yn7DiSsdQ8cyuXbg5J+IKMOGhee9PWJ7
ISOgRmKXviHb8WUch0TMOa79YwAP+SM6Ss84KIDZSM2cQmgiXrcnnRqob0ACBLTI
+HaXkXwBpG2WT6IMPuZymav0OD7sPX/u9p2tK0+vxp+dXoi2RYiHvfI7LMCy3drV
rDEwdiqE4WdszkGUe4RViYS/MDqWles+jXPkjC4tXPk=
`protect END_PROTECTED
