`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R9Ei32xwGNsvHKOzYXLYCax5tIIi/d+XCeXVv2PdUx3VirXMOmd69On4wsfRyW1A
m+VcRpMKU/SJ5laIiJacPNBA7HLrDNkEC+ZsiAoSRuF0O4c7muu9390fVzPP6OJw
JnfRSKACZbbdc/Wb9erNX0iN1+aK5jX5K169AVlfax2QCrMLgDm1TSNiT7MdFW3F
ndN9dQklTy+/nwiZ/7qnJfdU6OteBpb8wmcvMy5T8nw2Mlj7f+Td3tSxecouWW2o
`protect END_PROTECTED
