`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NYnZd3+gd9OzuhF3wcY7vWVeIujZFHhcJz7KlR1A31tJyXeoIuyS8dfMpYS5ce8O
Aq8JS6EY0OhPeK/Y4T6hOChC9xcTymQOBKtVZ34efP7eLelpRNAwwPZtHM824r7f
nN6L6kH4LJ38df7n9SbhckW8OzCrn2iGU41gfAgZJaVFAb6x2KVRIehj5+kYtlL3
ONx8OHjgrXB74WsPc48MOcj0oomGC0/F6xkxw9zlyf+Ko0mqZpV/HiOgDkLMTJSr
NSeb7WW6chG1MHT7+4Bk7Os+YI+7Hq8f4hz1KCNB/F9yMz2L5COhwCKH2T9yjCc4
7VsXQzMX5NIygxqTy8p3odMorYDA8sTOW7/Mibpq46+/R91Z4d3oyZN3zAEd2sm3
`protect END_PROTECTED
