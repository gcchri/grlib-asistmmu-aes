`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TaqnXR/vbnZr3K60LuPuim2iHXbddzj9QhuYix4DGiXFyXQjosMzJdKJqz6lkoaJ
GbgudiUcBeGw1mCxbUWhN4i6ZXRiy6j+9cjLxDB8R9JM7SBuFe/YhJYo40acZWH9
eithNazfPfwoJpEK1xb0LpySJlWNW5LZs/NgfPl9S4lKEmfPeKyMqUitLc0QDIw3
EkAeBYwAZiFWi8r+hfo25LEikxUHRGwteSqefdFPMOvaAbS9uaxgZyPTGjDFshtL
tmZ792pHzGdHeYlZgDdxewjUByJhEi71CVK7k1LQS7FL/fI9rR2gxg+SK3UuvGqm
pqyTAx2XMoUSGXcZyIkXSNNC+8hf0xOdpBp53FSvyuvxIebYhMz1WqACd9QaWjXZ
7wbag+D+QNWmWghrs8yWJzoHxiJIhFXt4XRHLL5Ipdi6Qw5R3F0TBfCXgVLxSOUu
j1iHYKIMgREyaoXXPxcKk+g416iyj8ZUskwoQq0KBHJtWciK7V4FKUGDHmRoU+2F
gh8hbuwIbgc9EBYeA7XJ9yx/LbWX9RVshM9Mwk+gfhVZpslj1OR1j9gQCEWsM29R
nv/W0Zd7IrB11WwAuKkH7Cwleh2JuMH31vHvPUHxtheDVH74bGEW3OcmuGkJ2xfP
WdPHRNm3JYfLe8J/+1VTjh4GPSzSQHYR5K9i3GEapBCL6BYfMMh9O+LwTodhZHN/
z1O5n4cJBUjtwt+qXXXbzvgEBicUWYy/czpN46SziGnw1f7OpmOxlJfQuSLO56JI
IpeEKhFDdBMxIFV0VVw+neMG76YFimf1XtxvTTDx4Fl6XKIPoW/1BnOMP2RB+++h
lo9u/z6ixxNLIIaB6P6Ug5atstQvTn5bu9kZo0vGjLoRiwc6P+19lN8J92igVc8N
B/E9pbtJjldMxJ2nFZOn1EPIS2EzaSmjdXCWASZI8JG/toGMkUrpYo/mSuTryYu0
mZ/4Wbgk4vvsRHMZ2NBRsAZf+F/8SYZdRPUym1kor1m3apZ7rH4THpJfuL4GG9sj
PZp7FimzQxHIrbsW5R6nD1Z5cQt7leid1xZ1rqwcPUfe0fp0KHF/HUeXodfXnAio
ckNuLLUMIQrNUrwFo+QKxbcxuaNIqivOdo/Fdn5Nej+fXz66DIjFtN9+L0q/4V+s
VE5T/GOg6R7vJYrvDtNEyIwRBF5acE8gWRfLSXqSdpC02tZqDlTrnASj1+ljfond
p5lQJ8Wyeuq+pRIYw/9ci3YU/h9xOaZ1P3YFP+lqW/qPcBlI57iDvD0XjTk5U8aH
8n6qAza4ga0MKkiIYL8Ig2QMYrMSClWl1QrPAzfftKppkvXjOjQOIHoTy80GqOiT
7KLNgLAtaRRGzmbn9ymfjMCtJ0n6d8Rgi3P+RbmNDnsQRct04gGjqlSeUWQQ44vy
KkRs9//MhwZN8gq/ReSV2qoMQOcx3CgfG5PtN2FpIj2lbgSUInymK9EUbFbKvcjD
yRBNu6HjdxRkBm5oS5sotuxJL+o75JzqsygZaT/uCv9WajEZ61n9grC6i8fbPwj2
JtfyfNuwLhMVM5rFadKVrKO+niTj2sFQg0rHf8XwLv8+uCJ5ki1E4DKX6EDbMgyr
ESCvLyT1wcgm6U/Gbzy9xwG/Iza0MXU8+1LwoJWLgZvPWfqF6rWovssPBq+0PeF1
wMPWaZzxfUWJ20vGrUmlOSk2SW73JoIPAZ2Jdv/kXnb5+ps7wzpbnHFIUTbiPmsd
a+GK+S07v+zNruIHzQd5vpnEG7ayHvcZwCJh6j+9gHKosDiWVlzPvrSbW4AOl5x/
HaxWBIkuYTg9ynjDkJgtueJJJTSlS2NZsvTjfkI3QvcbrF7Kq0gJXqxOHLX2XG3S
imUzvRFWwdXlAftudcZPUtaTQottUD8LLkMQfJLVNS05ccwftfSaUeWSPSK8IMFc
kflHruMTqH7pHG+yANg5AXWHblYwGllJh1R/wzR4GEraRIzGgperOAw5RDSBbtY8
erRxZcRmQ6p6DFhmVvD2eZqfoBgkp1bgMBw3rJdXACjl5MlJotXB+PM+3x2TYmOm
9YJmB5zHhrP3Q3FTW9RLm5UjePsFCbbeSxgfuo+uwO+Ng8oUy3LZ1or9+lHkqG/i
LDOuKq7mNS2PH1Ha1w1NUw9LU4iYRYX4ladrqOAoJwHEhO9iQQuQpyXa0Ldd77ZU
dy2A6kKgo8XIZFZ2vVOYGcgQSW8Py3pZfwlMnSdxBQoKdWOazIu53F7bu964TejI
rj4pGLDNOw0BOmT1zBnNAG1aHQNoh0SuwQs2OWUq31nhMf9ey+Hjso1lrwshGIyC
6F78PyCXI+heunHcGpb1mw/D6ROgDXieG+SRIK3z5CHS55Tocabm69KRKp7Pwhn1
vQgjHv/h/+cZt42WKefa/Wnr6hEgf0F+r9AJaTxLTuXsqPYkC2sKv/WL91J22gdt
5i91Dt8qJOU7Jk/AOnYZWcl47XK6N7YYS6L14o/SHAqlTGMDfVvQJuwdH9BbzYt/
9wkSJa6GLnhcvz79a60Smec6ww+7SzV2imrPsqx1nb2zZp/IeXyO7G7UOUMjXspW
uWsfnvF9DJwz9qHYid3zhw5Y1TNVXjzNAGOV6gv2BXi+XqZLqj7tPiN1sOfxTiGR
yIlLyjiDCexEXnmThLYUlD+y8s6oGfTbYrXh6rRratvKD4pnD1D1UYoGP042h6ju
A7MhDX0Np3o7BZDwahBM1E8I2YN1uJ06jONAAWvoARoVR+NNgJmNbik6UicJZ4o3
a85a6mJVPcLu9TU917jsCV4sBpkQOA6fnJ+tXewhLZtYLVioalY6BYAwr5ZJonDA
gj7LHvDm6pAK/CEvTVlv6dHBc2zDAj1XIG1byWJ6bELEzGZQ1uONHP0UZI8p6t+k
sv+DlZiUyfM1m3zQbdtp1a1as/tCyorJBDzqENbrRTWNZD5FZT878SrhPq7/ppwk
79exgVyWeQMIAlTXsBAO345uUp8yB4oYmlTF3auzxV5d0plH6LKAoTKFO31upmS8
ZcncEgW3FJkXAqAhUS+iefCx8j7xHsxc3FhuE6EXGpxbzMhvYxuH/G25ZE6bxlal
2dNEbSnBwwtxeVm1CeUulYjTgHg2Lckg8qgDD9ieTqSDmVEZbz1BBs6GRuX7HiB7
Tu3+rfpe5A3GG9/0BZi0Z1uWDLU7HFqe/h1NSPlDcT47iDIkv2XGJQv/V0vCKVqX
cULXrunsWJdnbKT05oWMKftOfbMinUjPctzYoMqrYMQphIXJe2EgUMtOGqNutFH+
wmx0gplsCZqbxj3m+XNDqAgEON7+d7puRjec6vAEjR/t8htFMpfOT3CaqHmbnK2/
xI0UqcTaO7A6bTDJSEZhzw/eblRvzAnXMPE/+tbSP58ulnhftB/S0TINt/CPb8j8
W1b0PjVwjKv3Aak4hE5xtfypU/pbpPU4W7D1uZgf7XMI+Ac8XsLR5E3BwRb22XGt
hz+vGAC/+biMUi7p1DcbLVCjPLJcv6wB2LYGU9qALCe2RKazp263kedje/x7+QZH
+/gKTTUR1ETQ8EVvF75HWfVe73QYpIS0MqcGapDAppuWNnNifNfH0/zzPSeo2dSi
K2Vd2FZVPIKFPbl3L9h5aHfBMGvEojGyMwatR4w3QPhYLNhNu9yO2aBFeutvfd2X
afalJ3uUE6CX/vGlQTEwrSb/ZhN5iFpOPkde3P5u1febXwYjo0k9FFV/2eQW98LE
4ulnm7yogk2cbXBepNBfJZimmTBJLH2qyHDDmUUDqD3XTiT04viK+ncWnsgQJ7ko
eangpdBSrnntNLRWlEXvj+vqC4Im/ckNAFxGTWYAV9n9IKEqlNWj81yDfK3pWWJA
gL/ZDnEvecu7O+Fp28RF32N61+B9StBsNiS0XtbF6TS/EWn5VOJ6EyD3CVlaH1IW
qFa6pmI2aUhC2m/3ItfP6zl6TXpKn/TutJLDZh6B2khy9y9VnjMcvI/I4V7ytCwc
M8vsAYOg5qO8V9b7ilICxAL8LyovvjT9pqLsxxRS/EupCOk1XwbPbZdTOIvfelCZ
vewUarGKxfrnR36zY/pi2gZLHLrjr9CmD6w45RDb5FU=
`protect END_PROTECTED
