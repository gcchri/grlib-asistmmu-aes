`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gwxXx8KLpyx8rm+VblVOskr671qMYUORjok58mMSE9PKIh/1MN15nlUbskkV2/t3
pCZZNSjEqQCOjCay0rLLYYiY89V/oMV6p2s4t50LIBkdAX5jQR7I2jpH/UbHaIn9
VzDXD3kFNN5zpMsHavSN4+kpv9L6tUcqoVdfXSuiJSm+73I1Oeqha1qM+qGpafDS
4E3NiCgSyqzoVomS8JWtahbOYpArcAFY0fr27np9n9UzCoU4JZ9RtPBqzRHYnBSE
IwJkJGBsuEstS2rlJqq90RsM4yxroHWkMumwkyrPthWLTfixe6PXOS7wO5kfwGoM
NqwRGD/WCMc5j3x5L0z2nO5H9EfaRjE4oiQrL5l/8n2gk2iYv04wMtrXOGWAioPy
bVKvpKrNQ1s5FtJDeqarUmH9699qQfXSqXF5xspBQ2Tk7fowmxt5XbfQbw/Chmhw
Vv77MHPYCBLOYeVXgd9o1+Ed643+O8DRgdQmDeAL7Zdulmy/jAkalbX18Y53X3o+
84pw2/tqzQ0kfLPNgSxvoowGkBWHBXUvrQE2tUVm6WknmTbl30VIKKRzOHlgBor4
/vMCjIzk0ME/FcS0njm9xXNSqIP0zLJQqDMYUy8jfriMhw8SK8MWtKZMbkrVpO5z
iBmBnph2Q/4oNkZVoUacK67+iLmomjHVSzLwFJyg6Y166qoaTacCgfCWmL385+aM
RIJmyAVdj2OqkyvH4lnlN+9GX4S87RHr0Xa6lxbWff1dd5mlpIPsNF3fpN8puUEg
SGgjZUeyQeT8IBcYX/LViUJxfSQKKy94+VvtXA4/Mlv+qX31N29MXhq6YQG/4RhQ
F4o9ddLkVi8sNmybwyNUqln07zCVVI8yGvBS73EqdNzA/OEjSnf6p8btRDH4dPyN
O/rln+7ukhHmKzI7TEEWvqJcAPWIwQiyog7MoJVvRL+nAW5N6j8rrXDYklklLLvU
mWZ1PJcyEGQqZCaapZ7tBRk6A4HqqRhKWGnRNtmwy37+GYGLB/xaOmeIqDlybO5p
8H+WJCmHP/9ymZtiItCInDPu/4C52GZKyurYLgX+tY4SqDj2St0PbGk+TGCw64aa
eAoqqjCQ8Wd7RmPEsDLmuSNJk+oNXZMKw+nPlaVaqmmfxMHZVi1cnvS6jrEmHSDD
XVDWESuLEli29fx9cyrySJ9RVIejdkt+jQ6sH0HOzGNCivLW9enMbRRySzQYmUF7
vsMmWdki/gREoBcJeGH/nR74ygq2XQXNuYcvezeiVmsAN5MTYLHpqea1KMvQKlVY
8x7NCm3nGNPhTNXgiqIPeWDRbJpB3fbkhDp7ImDDs76pBSZaZMi70FATaSAmL1hM
L3csyZQodwa9ulJ7xvDCM3RrbMrTuShXLBeUSHSfubKpEy7G7rjBc358fMk/gTQu
Om9naHrNwFvDSJZQ8WEzcx7qw/KQYYNCiWqRfH2uNLQU7IQqP3Nk3iB9ccIOijD4
HdStB5C4kVq3Q+hv8kSOLOv8BfsCN0ubQBItfkjWkT44pl8GoN+sSBSgGcMHVhkN
K4Isuh3GEDB73t2yVew3UyfnlA66CH7/oALbiaY3g53/bO9eEK0w3zWt3ilLBbEh
LDiNx2KrUtJQhnxzUguxI6DCuNfmwBGFVMASjJyZZR4j6V9alvZfyUunPKRMvA4L
loFu17SSCPxGIpyeemVbH37QwOPCTz3cN5ttZLnnFSIAe2zAfQFndloVh4fSd7wk
rxrkSEvEcrlc/siVngrdmkPfvvs1FBGdsfEOE/NcP74TefGj2rK5gUptjtt/COr/
Z4kBC1hAvZWw5CzhwydxZP3W5GmeABxg6nVyuqQzFAAtvEQQWpY//EOm4OpjpW15
ccK2CUeBlyJmoIaY9NxD35Txu5PCQNd6VRl2gC5hykoWeQ08tbCj+deHEtuZ5mF7
+nbyR1VGDpY/MiaZ+6OeH6mXa68qtPkRgACOd0/QrChvpGoRgllUg+w7vSAi+E1w
LWaV0gYdri2J016rLkSJZgPQjvWFgLotAu10t8F45vwgXgLmjsgrlPkRDuxRIbMR
sJ5h6xSp9fmUY5mxfWPieNBNdKb+2kEe4VkuUDnj3XHDWHPyfuFGFd3FzLMnnYI+
GukrZjbmy+IpIATOtyXVguguqHevZdRrVUErV/HDcukOibYC3EP5Q32KCyHU7bpy
eMSRejKbHMeygqjkKR3fpRaqELAwPFh+EjJ5wy07wRnG0xrvVhtzobC0+KvtgRUy
S97oWVehD/gjGAfksZ2dvN13Xxppo9JzrmfZtuBIUklupni00rJCKDxgU60m/Ixs
rDgHU+qw1SquYHv4HAgCRpUaWbOL2RKsoCE4gRj+KhB5d2HSBXBHWuFAZAcVQRzX
geH8uRpQlV/205JYhgMujTHOfrCHxB112/mv8tSmCW4kBD0HNMxobSEb/fa6umxO
VwfzzHB5cbMIsf9DYPszTFO7VS/CdgjCPt99lG/e9WcKUAfCXWYi1E56PuL4fYvZ
ZgLfed/A9STZjLz29dT+dIJdLTzongFhMZAEeu3XTIpeOZeviyRvdtGHjvjlekR8
wlUBYCGgDim69krjGJUps0qC91tt7jb/e1z2LL2/KBfFTiNJ7pTCQi84dMz2VrPC
Iv4TqH8oaHCPJFR0cKzinvNVjHVu6Pmfyjuqy37Dd1yF9debEhOZ4c2H3izALqqz
GCUhqxOzmB4mP55dmCUMrODh68Em6ioCU8NAMXPxIz0=
`protect END_PROTECTED
