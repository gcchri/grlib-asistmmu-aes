`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x4s/V8FeF7sTUWfb3jY4GhGv0YB+CUyW4fkI6qmmhewZQZZvaw01SFOGgbyDFbri
A0fCFGfxwM+8U+zUIf5cNPx4Mc8I7iTJHAKsiPqukW2JgC929lQwWnWt1uWEvciM
xOh23HVOLWBiYI9OuQHDuvy3HOHgdyYadC1YpD6urZR3Cq3oYjJiUoUFwSn831Ll
yAek5TN5gqQye7Y0gL+O+MEYeD/OiWxVySAcKnwr/Ueay2gx1kvd8LSPYOnODmGR
pddGjBMeaW2CgsN/ApyqTFIe/xzf2Y9aaGNx8iz8bM+10erD9hLo11ne5YGrKMRo
Wt8ps30AAJZA0ukkku/SfqqvFrZr2edrbDDg+iM4ZuyjRA2sScQAbTkjvh8SlqC1
16OuA0yra1/Y/TaeNqp20A==
`protect END_PROTECTED
