`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TeVCuJX646uIhhWT9y2n9n/KnF5d00SKP2Qg/Qm3qLfr2xGI2AComAMDPAqqTFLd
3kMexpx4FfWY3SRqM0VqfADi0uZ7a48AbHdGdvVs0E9Wx436g9bIqZ5mkFte1Dqh
uFKtjmkBwwzttmVvAchKCoUDXZOovO/dk7kS4ISAf/vMJgmTuuIgZwTAScFb6VRh
W1cxnhlO/ziLa4fmf8GCLrcF9VDwQmxpOXbfF0vOTT/HFPLNd1aR0zAux6oj5Axe
2wRAMPqCIRPBwO5MrUVh787pZImgv3EGpNTwe+T+8RjRwWXVmOz5yQXsdLGv2fWf
f1QteVvqwripHUTCnqyyIxM3nbZw62zqdE90b2AEYkPmr3vhmNe1pK9gnclDovM2
YJPUzXZIq80hf4QVYqNL01r0/chG+I45xp4J1vg/PwnoxfNibE9ypb4nTJH8X9bX
+5VNVUQuhrzkj6jui0WGTZZJHaZdzUzzbXy4mh9os59ongkPxheUHH0aSn2OPp9a
1K//oa1B/YMrXzXyu1nlWr+xgqCHaZRb//tzkuwJuGONC2/dOY6hUDH++pQf8jAy
2A0oxG3PeakHc8V8lGBHJX3Qpnww7TccKcWmZiZHgiFO/xUGOXILShVQKqpS+PG/
h75LQk4qtnpeShy7ekJo/MGPBOaj0UtV31WRc35nGqRagvcj06ZBFNAFjrWH/+Pz
OBo87vcU/lFCrUPU8y0abdHXRKgylUmHv2e/ePG+8AHJWrMgYKH8i6hCdA12m8c4
HQVUgXXpX6ROBkzhqZ/MFZDdSgBZxn1exBNoCLhNq4PlifSBls/rsJYMgxo+W8s5
aSYTxXNyn6wWeDHBZWDrgfiv/S+ZGvyARFs7S9XxbPdjMiolKVR75xtaKdRXLV9V
u7UoFnRfkT5PQoJFmK4Ik+zwiVbkZccrDMQXtpxh7FgOAhNERID7f711lsr11URr
hii6yRn6xzmfUzhu93JH5tbFxXfP5jOBmfHym2ZYbLuFQLQGSNoUv1p0u/xDUsAO
2LIQgLAeGBZhfzcnA6Hw9xYKxuYCSFZtgY71sRiTmjjGHrwabQQQxX4pjxUgII+M
sWSlCvH+qbW6EnRrKjGckQUzfsijawT21klIu8Aexv+AuPUfhlJZW32viGOeZ4fp
sjW58RqZeIilc5WJt9/tMG2FLfRQfpHMfpXNX8PV1q7S/E5XN6y4zkZ2Ugslf5/q
UXuzJBq1umGMHUmk1/i3fhTeI29qGQDdEvQOpID1TBJgmP9iuEGwLfw9GHW+4xFv
vSJXwrkCnVwmlzTKWBlRXhVnPMuFh8roDD/QgfMZUFsp9ITvKvh0ZScsgZC9r/EO
HaPxUNP4qT66DUB+P0el50HETiSv3P5ad1Kxu5PWd4K1+3Be43s3ns94exxF3oUG
2id6AfyVS4Eo8wXPOLO/WKMX2sOtlwX8soDltfbZGMWWjELUARLeERCVdRgNaRBp
3W3sg4GvjBbZ8Q5thr2Bp/UV/XqcXNfsSisKR0nIAn4X28GBj5JSU0c6IedAirjg
d5+xC/eEZ37Olmu3ih7JpZ/uGSqskpkOBrzLkKmEoZK1+enW87v3gRZAb5gJOlxo
y1y/Vnl4v/YbquICNi1Vdqkht4tnphO2kNd2I8fHBDMjXjwc7PUwpJSaEmwaLObl
BcKd43jXsiok71JpLE5gfVH4dTczG40RWHqKUVtHK85FbBL43pkOv8yJ7QrFVXHi
dSJFTJjpqOGXMIzVtlZfeqmv1aeP4WMRl3pr1cdfDTGaZQyqzur80etI/jQXRG5T
ahEgKJwEcTXPIgxnJ5p3+tPZt4TZ2n5MdX/eTuimOXcijuWpNRNqJsjcCTJNAyFm
9aNYfVj4aSIff/FZn15TLQNFjqcEaIa7Y2EEdJLW+CsbFcyu6FA0xT0qFQqunA4S
jxqip65MSA+/0VhTFCpPGX3y4+8Fx0zVllQT46QkWVSNoLiH8g4nJCCGcLX9pmGq
Yykd09G7wT9XCdZmTBqHZrYeF4SYdWzy2I1v/6YTD0vxXc7O7w7C/a0d3M3dgKhY
BhsksAfdJVRG0mJXV+7L2DWTl6GPifKo1kuzSovcX5SKnpigDDyrELxVGoFGEHw/
cuM7H+r1azULWxywDlJNiCBaiL2/dAoDndz4JsT4PY3aUdGakz+w/L3Y7+z/Afq1
+/VwBwfTToHKE5E3ZpA4d5WpWwrzAuihF3icQVqnjburJDboLFdZ3B5w7LWB1uWc
RrNBfZdyy1xNwbV9IbQtvRzIC92La3Sd61gXEQBBJ+u8sSTyw+BHPlkIOe/yOALt
pa5cz1POUKVF/qFu0NvbOBnaG8kfKaqYUzGZmfHayGJyYVY3ql/TwUb5nvTyR66X
ha0DvQ9NETKIs3UI5OnqHpxCU6nCkuWW6toLMZ84EiTEuVVevnKLz+ir0klAbIQM
UlqNHQuAXhofag4XwRHWWqzP4OL4jhkQ+FiENinmzOcTWeiE5U39bbYic3IGLHqd
9/F2Y9i5e8t+4FH1r+0QB8LdibEobYLoLHINQXYqE09w+CrfXNGc6q7mh9g5Kwd+
Ycc7hkhXvSjQWmO5trHEMY6koGqdok0NyVy7o1bcLcOkdt4xWpDDBrxAGFPw63Yt
i3WuDiR5xVQ/FzgqlF4KDGYqCqsiZw+zfqjsnkO5I6QASUcahtYBDURN6VFWkncy
jQaCGqFpW1/B+crKwKwHUKXSiwmVxJvR64lhf0Ld0mfFUCVahOiSY/jWdL7DwJoQ
0P2bLVhMr8WCjoLTR/cZUZaqUVoiODywmGLZjExwt6thvZX82iOGem4dD0t19rf5
iKTVgdelz7RJQNu7yacca8U9ixitQjxEVrsiPEYRaC3pqsytfq1jSNG/m3V67NJL
UbOa80CSAlrtz4BQQiYW2KPqxM/AhTqOzXEildgdfhcPTx5Cp6LQXi7/j5XUEc+S
HEYKB+DZhAez2SdJSPMoPk0/tfTf5VS93tuf48nEzuwpCvGJfDvlMudjqt0wwnpi
JUUrnVknQb6vVcrQNuBdTQsGGz3ZJiKAkfRQdVKwsHod465C+Kv9wJKQPFfdJMmC
X8s+1rew2lZHwawjvorQypvTVBAFhy4EY4bCtOrkMBhOf4QqZVyGwAxRNoVhRV+a
+AwYhm4C4gLvS9/Qz7cD8K4Afb+kEluAeXtg35tY08FGXyX9uf50khnoE2Sdt5XU
pcJqARD9xhaLSWCUMzY2KWiq6QpQi+jCClKeRW2O2hS99MWTHJIj24XPgYnJ5bFs
plTFpiPBsZE9/yddV1tIAp7TnaMo4gdhc307Tm7yPLLGbaXIeRPF/2edxYAAxoh7
6LXPv2krzNv4YNxChR2MFpa9ZMTpQMVAwAQ72ajE+5izjmC3apj+SIZpJ1s6PBX8
CjckpgY2EGGZ4F/LLUELTcqSOLOioBHKvwKJlxjFSyXR7tC4tmsukBirGyie0sr4
HesSMCKWl1NvkRcuw5J9yIj+yqio/Bb0+tz4FsXxsZ84UGeeyKctyzvH9jiH/H/X
xEmlaPU0rmwDYNgGE65wGdC9SMll7Vw1rpL2cWIJihPNeNsE3Qt1ZM3taGJWLEUu
x3/dBM5PPcYPKT88KyTLalaxj44BnPk5cjPBJ7wgLzyN0Ao/ykrqGFV4OlddQb4B
Q17nHjbN5EjAMqwn8A3UMrGD+59Pg9LZBNTo9PkGGJ1nrlREYKnbt6OWlMIo+W7i
9Ai3Bav8op484gbN6aAYZrxIlVGRKCX1sQepvyLYtTwTdljRn5jMzoBrPOVCW+5i
iqRgJx9o9yqs3qkqPtrqoScJcYZfYMp/sPGdp2NppYD3K6WihLL2x8QkrdSAyPq0
MN98xAXfrocGYQX4KRzuQnv8zk7U7nGXku6tcUsXsejEEueZtj/SKG0LnH7XY/HT
2599r32pXO6TcT2WBzkOOhcZxFmXRZY3J+tQ2P2dXtVWfqy16s4hI75dcSiRMKWx
vSKf8OcT6jdPp2qYhrFS4YBIB0My7c8Yqqc+uhsu5jyJZaR/nT16E6LfHB9hbviy
7J9YwbylVCSfmIMPyNnh7pZo7DLVgzUZ0KmJbXNrLDcgRIvoUdxtFXRWPOnlVKSW
ZHkhbRbR9savKzsSpMh2n4NRPAovuwiTOyMMn2/rZDendkBlcGMjCcsDn5HDfYmr
5GiJ3qf4fkbFg0A3iI0ABiJwqdXLNCcGDsnARSgCC4azoY4D2UyHYMUIcgjLRcNP
VknRAY5Xr81alczelvEDdBA1iMT1FNRLHcwPDAQPkxbvSzE8rUbF5y9nF6vezjhz
zLfZCpUMGncqBKkMmO3wBiPxODPa7i9N3MLRGV75Nc1qm8e82JSTMNQA5xndUvho
vy3Q81la78Z8lbNvvZi96SkKTgOiCZAFnrBxqvJk64B0cceAtBcjFzlR1e0De48I
mVpNNYCLxOfC5BvJiOvmtKzptLWJRssMTazpzFdmkvSNFz2K3gop0KcobkC/mdLa
WRjbpl91vPdu8S2FrvoCN5KCvQYe7QXnN6rCVAkWPOL0/rjmVuKp/yZL2DWxluNx
c7o8JiJO3T1CkBYo26iyy1tJLGvGgjcTnKxnBfqhOBJIFLsb6GhF1fa22KAn21WM
FDuTCkRnKkhKxk4pYVlOX6a8KJTsBU/z694jR//9gySSUoxdzAVYWEcoIZgWqmng
C2AWgHgo27BuPFovxoZCFfj7bIevLvBOgZJWFXzQZEiaESbJGja7em9c5HbL8y6w
wlxyH9GP+ZS7GZAk1b/ymCDJeK503T5XFI6YZx/A4xWCuOsm7Gs4oPD9juFH0wpu
/dsX8a1JU9xHBrh+lfjQSfNRur9PWl6FSK7ucmX7rcuiwbqOftc9xw15FylvLfjI
2+isDx6tI2uusCa1IPbZRzp89RPCXPy5QwvqXBhEvkxfnVcOzDBKhSriJGLMM9Cy
lqFqEn/0A/EsIpr57vZBJpl54RenWMGTvWhNpadTRuVvuskODrkHopnEn410g75m
NAFJB75jmIieWAA6eRd91c1L17oqGgkkJpKx0dPUQTzJ0101uIt6qijBBGij1GCd
2NBXCH3SmgERqAo1awqGwGBhKGV9pZnI2yM5X/gpLZcs1guhmtmickFE8kBGrhIj
4PyYzxlSKbTDCtzTlVB1cqYk14jwJyP4ZNx+tAi2y3XPFOGqT7knT1P8uxBc8j9r
D1Gd8FtbI54JgkMhGZb8k0jSTJmWDzL84sSRQeXXqH+XUhdsz9FnzWwVLfxwjfh/
vplln3iF63eZ+oGM99Wju4JeP9MKsZhLGEdZGEuLC7XejFEYYi0R6xR+E0GdQjzY
4hagNoANK7YSuY7YWPqgH8iheOmez1vtjev9/t8QpwkYoYh/m1bTotkdgGNs3EES
u0WOeJCa9ycDN6LX76F1rM7Thx49D3oH2P0Rn3gw1fV0CM2R1RURl9tpmolBhrXv
AdQJuvnlvtOMxqgBnvN5Pr6r28G7jaWR56aX2lh2iBlUsy8J3iNLa2cST8DykvRW
QthNCSPI2lO9xyibOudxrZ5iSK5PtsimaCtsXJwG6NrFH4zMf1qLZKU/dPPgnlqe
tRKtqmdHeiz5aphlclsaU2gx5sXvjk1lMhPEdZZ7aODQXqwa+M05hCWCzew9j+SR
jPqJU0Fkx9kzqsEDU8agL4ZdaRoZxfxmIN8T/NqaZICcLQLHJhTnHVXlfZPkrOjM
nAYdF9TvssFNXF61nFmBw0MIuuFjUmmQaigbuTnLEms39ffBs1ZdQBB7/iZRshgz
6G/jFoXafD+sGSSCHGNPgGjfZ92i/gqB33A6w+a91ccE5rTq9LSSx8UZfAEdWOEO
R0qXeu0LINwr0TSHWCP5OHz31NcT6otiAqq8HWq6fpdUrRdKtlUASN/V+qy7gUdA
gEA5n5Z8Seyqo9kUytUgSfJ4B/N+B/blyxGAqK9lYjY1Y9yoLTwRF8mg28Qe5ICz
ZthlUyr/a0rsFmQRBuyxktOEpIH57BkHWX59pkexq+OuHAl3TrKhl2WcIspwAKfo
AXs1CUmrO7LIPNB801viWsvGN8n6MRh4E6CA23QfR1fqjUD8P5HKi2TCxrCPx0SX
A5ngHi8Y1mm3uQtsL1s/UIYgJkOz9dZzuhmUzIxENVlSld/Y0ErdESYFD3fKZuus
Ky4FxbCWvIIjxp4TkcTkxw0SHd1+Fal84OuAVIipSFzL8pLTiVuWB6FCyaWL/oHg
Oy2X56F7AZoy+u5jqMwF4vlvmBghQ2oSj90Hw9QO5fzouatstn1qUnoLSIsiktIb
NxU4cIyY1fGW0//Osyj0QuZU9LAR3EaA4qOArvf4wa+V2/rcv33nDXGL/oSn8ugb
8aVrxqEZakYWI1lUo7MzIuLVbWhwFch9f1b5443Y2W7/I9tLNWI0WKx3pPybcAiW
Tpn/6MsTA2JUJFtPDyhRV2NEm7YX1acNAUTKVq1WBuGMc60mbb6LsBGbfjb0bRI7
g+tcEJFiIlbWjEC1Uo8L+idASVRHj2B1Ucm6kZX8FxgrseqRKW8m4/xoiNRzo3Cw
OpCx7uPjP90fNoeQQm1Od733kTc854n1uA/FsRcd+7xmGOIxgeJUonfH8zxaoWu5
bYtTw54sUTd0V8Hm0Z0a84ij23oOWyCJs4AaWH55vttng1WqoKpmxs/c906UJefe
o31Kn6AHOgXqim6YvWQTepBq+4x+wi2Un7ysgEmE0ouQGHHk5Fo20BZqdelqjifD
Ue2V3qVVHFCDdvjJnANowC4o5AvOIjSZ4bdk2UD2HspE+mzbKeBXKBq27sc24fMo
V0YCsEQh19wNoLKT5h/27mncqO8l5zSNWzYurCJsftWkNMiuValAriPfNKCI6LgZ
H7vfxe4kEaHHwInKvvQg5zMYbKjI9bJ32zK9F0OALDSf7qPg15n0DhToTS/TZtkK
EpefJD1EnxXdIOcstjzvNo1NkEIw2B/1+ZJTB8/f+i3tRrDhYqAiNnkizVD8Ie4u
cmqcb9Nv/XghyrI98hQtjHHft377+KyuwsdesTELtdZIjJ0vm8cZDZgI5Nb4UYvd
EMqSgN5oxu1caQbK7HWXBxA4QX2zi1HW82uuijlah5cKZR3G/3PX6lNLxCFfC5xV
iA2qTymTm3qgRydxwtfaNTVpjtkoyo0wft+x8U6Q2NrbZ/Xe7o2ygB6fkVepxkTK
M9PFqzt9pvPHDortA80pLKFhTTNa51vuxxk3BFupajz+mlX2Rq4LBfyDWq1a/swj
zojK1KNru38GjZjhY7MFJBzs5kJxMjxik3WrhLCKLXSFUEXpxeQtk7Zv9fntby3L
yWCjx9KrSU8bCQXYPvGp0pnmjCzYshHoSriqZlC0D4Oki/U+ZLfn8v7HD01NuXm+
/teTxi0Pyf/KzQQRhQlsUI0ky+kprZFZhk1GGAXo+zsy7kIb9Rawr1yk06uFvCCt
OV4QOxQqS7ak8e6RGJqvvU6m8ss3wZuhqCYxLhpUgZs=
`protect END_PROTECTED
