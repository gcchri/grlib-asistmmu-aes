`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T9TQkKDShUKzbRBXS/L/TRkIYa6I7FtFyAzm0ANByvHTOW4y/oRV1sOYRlt0BDn6
t+DBPKiNagtJQPyceiA+JHIc7y2M73TtYgOyqXPDebgBWyw18XvV3j8W63eBaxfq
3IbRQLSvU2zF+/3RiBkvQms0Az1KbgdBa+OyEqjDJcScgHtVU5b52hJL67o2LEYg
L5bZ15AVZXVOd/BErJ9Q4tYZSE/RYWLea0bOkyEUTU+0nqkeI/scYTP0yWdTyIFR
TyeMY7voGA5mcqH1A1NwdL9LIeDXbdZoqBrHw6jQNcPJ5LmeeZlqrQQbLwlxMoXu
eCx/A+SDLJ5PolFs478rmXL1ZWAZzm1aBr62kzECi74bPYbtzAidNiBBiVrLusU8
i7Th76KVz8JznvYL6zzk7t7SBJccFLg/wpkefA1sSlW38Ns/MBbqievUGMGUxMd5
EK6YGI4ZLug4LFLOOZ5xy+HUW2A1UeaGtp+o3RneBdZvxnyKoG+0OLoYP70HUwa8
SjJUFLXvFvjdlB6D3Eh6dqWO9TF2958ddIuAZhDt+JTAx5cyme3cSATPRfCJ6yVR
UFoufM04BAeafu6L+XxhScNQmiDszp6qDglmr4I/9csTGTR67Kb0Sc81j//Q3mM1
nr0jMgroiURHknKzJ+Vt6BnUbBdbBi9FDpSC83fo5CRA7Xdqf6Ic87uCoNxHONN6
XXES0RO1f+rvsDPHCGGcFxlVsj2GQ7S2wlqwA2kEAA5HJ0FVRPhM5zlKgTNtkIXo
NQHKYfB4wSe/jVeijcJhwROgIxsSC/r5sgg5VYYS9TtjKUBkRr4xV5aP454LfovB
+58BkbDNvYuOg7Vs31+cxUiD+Pv87CO0uvPx0qq60Gp0p6KAcgJ4kkyYl2UAoGEl
hIndexYkVvy4/zaomkF/+i84X/5hhPAMohdAx9r55VRSK+T6zMyIKCJMoVM6U4V+
C1ltapwg1VZUN9yRhWLuDT3Pr12bUdTNvZjIeYDL9b/sLpPKd11iKATSllMfSpQN
nCv96szfoKmEP5ue0QNeqJSKFy3+nwLDrH4B8OmIpJsxQjZU/X+GokrZSrD8mqjV
Mn+Yntv+jVsKijrtR3e8CDKhzmCAECuCY4u9pENTJNkDkslDesxfFlHKVmkvXmMN
eqf1QSf/DLOpnm5PnPSoLQ5+WExGrGOHvigfuvQWzb37vSK5weOvq94/GKvHepCw
CsjPaRnI8mE/9eE1xWW3BL5wH/kKcLec+bZ3vNN1zaSfYuRcs8oySbOVIsBuQVou
8RVnVYtaVKtdjfgv7US42PT6wnWsnzlWX+8is+uc/wXbMGyd+YUp+7G5gdR9yf0J
VFo+ll7TnzKKWD/EOTBobVlN7oiz/BMJ74PTXtG1p5aMmGhx5VVbRu2cp3k04vBZ
XfUgTwA5pWaU6btu1u/FdstWVOBILwi8af760MAD0ne43BhGsiAWcpXrjyl63pn/
CmV1oY/J9l2DzQ5p7Q1jJ7NUofiJznL2m/QFXPCDRDmJ+WbJBEFj6nwlXpgXUqx7
kyDbrNc7v94caX61ynPYxBRSsjMEUXBLzuFs6Hg6M9eSxMttPFK37cHJbSLOicDQ
6Mb31gx4xzpe82VMgRq+elQOsm7hpZOxjiCvDkQJxZHSomq7sB1QHas/OYgtAAHG
8raQ2Ak2z/oxA0ECvDG6Rr8VLl7IKh8pgFZzUGNKlc2HHPE44O+BLYNLRze+6akt
Z/6JrJzuG+4tQ2HTJxy9ws9IKKfmgTtvR/TXuAZR5uqgHU/6UAjfCe3zSFMD1nai
uxO59dAAIRLVjfcCqh/k9gLLnbPKLlINTn4hPeAeNJ5TMERFSiGSTH8rgCZcsbta
9gqhF3HOOrz1NYoXfFmpxv98JlmtD6a/snvYaYoRBw5UZTziN2xtSWzYQHNom79o
aDRvfu+wXvavB6K/amfjV9/9uGJUe956Y1Z1vNPGJt896tvoBgQhsg2wW0f7tZVn
9ZWRuD/NQ7oJE/9tSW50UPv1EAc7z0sjoDk8oMB9F9aPUgzpyU3epop/qXFJuO0D
hMtd7YYFOCIg0DjK6NmVS5pqTpgz1aSIPPwvB2ARqrvLkHxD46uz5XcHyMl84FEy
3Z/pCjqbj1g6Jkf4lrO1R0Is2GvXF8ulBb6rDliQVH3ENRwraus61iOCWveeVCn4
uCnCZL2qzcGp2unQDa58gt/ldVJqyBG/G20zvGWJ2gSuip44wAZ1Z+EE2XFa57/N
dT0lDmluatPP70Fk+O0UtlOY7lI1RYhTDeaCB1i3A5uYAYsNIE2x+9KM6N8ii4y+
81EqCkcslzHlHd4G/lRg2X0cjAfaJbWdlagV+q8SHP33wXDdKShMnZzHmXb4yLRs
A6Oyol2pHS+/Qp9c02ZC7dqZFu7JyJaP4vKqTdyolJBJ0cRMSCu8jYvIuIpBJm3C
uok7FiTk12mzbaa5+MpRKBg1US8sYaDlxDTwC2mvKFfOw9A+UpzoiQ5fm/j5g/zA
PudOELi6VxM/MpJTyvrqNHnVQtjOnYpVLKdjv3CVQ+B7q/2hWVdCoipQ1zzVUQWv
AyxGLFC/k1qu854wIIdmrLp58ddRFJRp4ZS1KZyH/YW/5reGHSzHjG+0nfQHAHNq
hX8RSzK1/foUMVHg92OJUSx2J+rCFaqCtCx+WT0RZ3Rwuea5tnP1ym7BAsG9iQ05
MqZpkveBbsxKwRJOFl1xww2V3pN4il9uo49n6lEp/xDwDhGYI7yI3eHgoYn1Apw9
FxjkMWxzjbpH6kATBpCra0Bs6znlbw02S/39It8zLofIGwWwdzz9Iknm+hyDtTpL
wJRBK+f33CThxdzyUPppBk6eMndp+7beO36Yc5l6YZbLZ8VZsqiE1pEnVI/pG3qo
IbkssJYzmTJcgqLFJVHukSuTkS/srwX+iZQqqhElkVGD8PT36FQyfcSjWtv3yQp3
Z/6olt4ETV6HbLBhyZTAaDB8vpgVRrdSA/TQVqgdLA84iJvzK+7WMSw3+lIHoXxl
5c5nwXemIbDWZ03qxhztrp+lE/7zG4bu/rH0TQ81p/oA19NXyiVidf9NJegK86vH
p5oeCrBY1aOISHtFxDGSoFZ1Vff3Z4uxtkIpq1StUeeJoPka3fXtNbvI7VYmZyco
l+CM4mJiLRM2uK7dXY0bFeigd7NEnkMEk7InBpHzXhnZ8Y/LjvyDthRO2MT+FVnf
+ZVTst9YxCXG0IQLPUieessXF7x09ROC3JXSEcKurRopHD1of8QBB8RmeVX5cTZd
wXIYFD1VAeT5+A7z+kmSgmpiqOLwTRe/ycfUu+6C9hewYGPNwGfomDNpR8W3kfP3
CLS6bzGcHomC5WVY1XeJj3yNILK9y+j18+ifslx2ByRQAbT2loImzA7qDqbTIXXA
8oFxa9I/cb4OqqMuJhH2DQm6Ms9Pz1fXnT+yTiDOz39Lfjjzi4S6jEZ7HsXnC2on
T1y4oS16eCDrtYPGx/WW3EoekS9FdU7QmNn5sGVejBm0VxdKG8bw7xuKfTmKqvmH
V2a0fX6RTGQqxGH2hyoihEQZPpPSod+YDxXLu3r3SXtCMbcNaDa9H1vb5Tp5PKiD
rgrod2/yudFn/NfDuFtPwQ==
`protect END_PROTECTED
