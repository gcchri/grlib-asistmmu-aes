`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1J4WnWwyhE2A6javkPptsl/qImmx6CRvxoAjNIJFMdC7xJXZXZZCbxNU4ZCSLEvr
zzu8nfRBL/Cin0vpSxJ5hLhevLGgJ6hx7mHyQ99hJ7JvS7a6WDoKnntbS+5DaLj1
/QZMDbAxPd87cC6RRCw2jA7C22vi+gnj924MSCsKeCc7jnNLPFkQdJvGpQqGCREg
WOtQEjsCzkLUt9savBgnP52HWzGHVm9YDSYNeIKXTlpF2LWIXXhjvN6w9optpNFv
68x4mUh3EtI2HjDcFxgj++xo+WQ1VTaH3aJRnaNZ8oHCF6xXXK6fEzz+YOaQxaYt
QSYFGHHUa8CM9DgPUCQ9rZsRLRkBrrzzSXn8FvYbke50Q/tUn+fXpmNJx6mtXU9O
VCRydq7Qj/vbofiqwcLUs4Sgc8YqtBDqumDl13ntQZyA+9mS+5HRQshDYOcM5Lc6
BB1vyGYgH2hLSm8y/zrCcSIAo1CKq6c/nVK+aCyktrDKMfu+6W4XSOuudmr+PD1r
`protect END_PROTECTED
