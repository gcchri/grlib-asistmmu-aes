`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J9H9mKSo2iFwi4TSCNXds7n2FeWms6cQY3osIDsZvyqS4vUrF/kAihWBJgtmO8Lz
vX3mKRslZZ+0jtEocRk8UvmNTXnEr3fiXMel65eZQD/je29f++tRAzJ3jImTBQvZ
T++5lO0Z9JrchXJEnC/RLvIZXjmH690dLs6uN5oDPFiuFDGFpe6X+GblPzvgZiZx
E+ad/uk5dunq7bL68BerOlAzebyHHb99MJicA1/1BFsg9g40fNIDprATfTPXfThg
aZ3wceCRgG7SitB0yox+l3ejDcf2+wJcMBYs5SfpT5EAbcKPrLkz60g7B/p89+RL
qxDtI+pgENiZ2aXMI4YE5GuoGTZdg1Ra4skxe5VQoNntp++hUQ3PKoeWePHPwC9s
Wjr54BE6BgvqpZpDLMCKGZzXyiDn3a6KBP0fiiE4Ip+Aga8rnir3KYsSmEIFkZA3
HvbnJWuPfm/9oxVrDI2SQI684e0Y8j8qVmGAd23OAt3PVVxAh+kCTyOK9aFSPDYN
t1wuahJyMVzFG3SoaNgOM8RIxsW/fymb+PnvyOIdnbd+K6Vs7SyAhC3s7Oznv17I
jahSnvYc6DxcyFJ1dMibwvLdodtWfJqhdNwioffVIZiUaAePi2POYYYDJ1e+cQMz
lolyi5mpGNvzMpWsqCRczNPj0gp1GpvTYx+YRXwV7sVRhY8E0oxn/eT9lfo7P9yr
6Ypsj12h385W85o4vCPfcOWAV6iJeY4jp5gv2H6jGb6e2mBVmZH8s9YSGkyjmcYn
YuTWTSuoO1b+J2U0rlrvavcbsqwDEHou8OhtlD8rsdOt5DV+8WuLjmwL5qrLsLt4
J3DatPlzXw+42zxWIaLZCIMbbQ7U48HP3hWnHR+TX9LTBMpAbSTKzEpvVX/eLbIo
swsAIt1e6yHLoCrHhQqEL/v1tfNTO0TP3ShIQxSNFUclY/z/hjzgQqU6WxjYJuhI
sOdla2BnsSHkwMsJqxIlcUSRj3e6rS163qgNLxxpo3P6lw6ffthjmEsiO68I2/rx
Ru79Wb9lZEHgvMPVzKlI3u6ci+9x/VALqAju0s/IbYQNVqpX69cUNE4iEjzW8EH0
XEwt22h6YNs/YWg6RMmF/p1GXgxCNjv9Cp5dO3bbVnp8Oj+8QNw0IiakvQmA19f/
Vevu10ao9IwCDSmXoLmLTtL23E0Nh2/5Kcf/QzndLMlA6G4tR/YjPE61rpXHrK6x
ktuXZDmaoYG0JEKnc0LNedVBmEcRdlkPBUbiF6kBKjVyQbj6GMySjOn5zK76x9vK
8xCoaCwf9WC20mCLn7uKLkXGLHqJ+sUrL8ibNFH9ixvvVuK8RDE1dGj3DNdcLb6H
ds8WuhrEt/Lf8rAJkR1qr5sbzhxGkdMwi9KAkz7poT7sHeOPe/ujCQalcye/3VE9
XVz+EUO+jUcGVnF6oDVLOu7N9wgDJUTCN/EGpTwJA4x3nizm/pAKxknX5GDgjhfj
bJK9aVpfxUE81hNuVkzM48TGUk7dl8wI72QssgCc9FNFHqA4Gc7H6OzGIbQPDA6w
zi3EC1thQ9LA7ndrR8vG7ejRnNgEehcGL5uwlquBRI+p0lvfX5Ui43aOuDfXwdt1
f4jj+wAaPar4zjzgNeCLo8iDibrsryx1xW/pNGn9i41YsfhrF5uUaNlZ3HyuAsE4
ecD8LeO+qUVEdvY++GELN6IfLYD/jLdgtCtn6e4M7efXuLAfIrls6BuDSf6Mbw6L
6vbhlQD5eFPNe13dNyRSD98vMWgzz5jiask1EhuUcpWykRZ4Pth1eqBPCRkQ2HIZ
rQwZdMJ1Al1ztXeT7bv5H2ZmQuIRzaDMB+mNXBUWFjq2jyMN9dOj/215h1VCRcn5
0wEYmhvFDaa+FQZ/oHcRVmVSefiYLYpeB9n/sTZxr5LeohwYUfKAHjYgvZI5TN1/
+2HZmJGmDvQIgEtzVJ8eq6rCfmfdkuTAKvsUkcqsv5MOcZCUuei96ltfc7sWCXGo
sV6XXPlLnfOv8yAlsSKWqTUkTbWAarrjQSJEjGuwkTjs80dTgRrzzLOVIgd+/5A9
rIvkX5fGr2xeP83l+dhLn8emd6T/OaTr9UwemJRQrhgcd7T3XkArHj0girOF1vVm
XbIkmDzCK9r0AEggT+0aMJ9G+PeKbhw9YIbA0syDV4M9e1dsMZof7vHoZttgtcUz
MFCy4TyjQ4rGD80qIfvn39tyPHuIOlfrsxmYMUTe5kPb7al+srv/KmyWJb3X25rn
9zsZgXigVnozbd0IrOJmbuH40EifHLf6ZhY7XDuP17fAgSyQQ9jPjQtHuYFa8viY
9a27HvMjeKBuufM5z1tOff1byI0xkX4PX5ywr1Di+Irr28IuGnGVyNTNdMfEOvkN
nGkg9VHhCLaaga7hY70GGHKIYoNlvfNOOFQ1OIjE8yEw1s7xFewXguvHK5Nt3Zus
M69PV9nwtmVDcue5WH9PIVY9qxTD5zeDUz3l0/Wida57RYef8R78G+vHZMqSviX/
5N0bRkwJKxE01cxjUu3sl/LiCP6OF5HI6AAGAYR1spPabbLYAWcGLpqUMmz2WnLB
qmsQmXqU5i0MawkyBGtlUD92lRK3gldYPjrqiVszXaA9SGwOjVJWq63wbaxC5Emo
uAsxc45h8N4f5jae/xckcOHBR8YZG1o6AMkw0es5QR5t9A0qJ1B+1RrtwUDfRKFX
nDQud0qbUbcdReMcOjGM8vQsBGtwOLjliCg+rAYjddULOs9+PWNnhVZ2lkl9dlse
AUV838U0rMvISXTRgE/aL/nfw6Ae1VLvxRy6WlzmTLsPF/mElR8iXsDRkdmj3iQy
IS2xFLLzcVR8JhCzBHWMzXGyzmx2Hsev+LLWJoztPBuDJ+Yl05H3zctHLfWSUrvE
bqLw/ZoY47SZ7M2tDnSDarVnxbCBkM4eVqB3QKA6e87Mt2vhDFH9/OsZUYlKWunP
9ZHZAKKm3KVwGwV1I6nbKB05syCcsR0UBDiWlwWgoFbhicZd2VV1i5tv1XEmQkIn
vUObHAR/9A37eZEuAGeJ/T6AxBQ+K7usMcZfCo9M9yjhOUeC833xSzUXl4dvKUE0
F3RMe9F1A/YyXAM3gz+jluwT0amu4X1Y/NKnebFgflMh6Yno+P1KchNzj3hEoKF3
vnuCmdGpiE+nhvoKCtvDRYQv4tXQWg4HNkkFCZNotZ6qyqJNfRtX+76x3zw7ws0I
1JGoGCeHPXfzLFRp2PJ20BTbXzzjIHtgj7gq+t52S1L2KajjOTk1x5OH7CSgM5Pe
95UHUleRqDnk6mttQYC8boaBgFWEAeWYGBmy3nI70ND9XPdWoI09DoQP758EFJlm
FpgisX9NYGNNtfGB1otMmKi/iq35UcYCpK4Xi5dBAmPUPB9ylX3YpuLHpaFYw96E
AsRgGHSGChM293pFWcz9roG8qp6VrYhGrRIhGTsmAI5eL04tccMGj17vNTbZ1El6
SIDC5OL7J3t343jlrBFhMPLR1+5Na9x/mWkyTr1FU8HOWYaHCZLcnDuoTpoWgHZV
h5K8bKC+u2xn8GL5zUpjo/iMy1vBVuMMiD6hpEnQyJ1Gx/83cbplzVrzMCL7D7K0
/1HkwWcbwb2YnQ173Z6afaqO4ex9lLRFa/n0yV+W/zw=
`protect END_PROTECTED
