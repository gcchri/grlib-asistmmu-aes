`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/EyKFdVLSjTcvYxH7m4AfOnp9uV64zZaUroZemnVAsb8CV79IsdmbS/4pVgEHMUk
DZ3l1HZAQjzFbCFxHaGVUv0NYGDJm5P/sbazrhEPvs5PffRYnuRScg8X18rpaJP8
ojAT37BeVQFNLjG3ji1uNQyrqgSH4BmTzhj1jV4UGOjRdv+ySJsphAL0PDlYwW38
mMYgkxVs/eEgHcrZBzJX7C5AZVREg76GaFGR/TB+z+oGn2A5Mug8BMaKBCUrUna9
yb4QZyNiHm8xoFTvyIUHLaUU6HiWEU6Hvxr9y42veU6k7MVdfYdMCBkz1WobAgu1
iXlsYpz1vdO/5NzS43XI3pNI1aGiGqphldbO83exsn0RtvutmoHPF5PDXrkqRC2M
QHQoaxoAIXqGY/qOrtdBo9M1OpI+guzFGt0EgLrIHpYDOrTxXoUVBKEF90dH0Rlt
lv2ZBLqrEad5bxjqVqVEVb8JMYHlpGmBUnxE+eWX/1+EtuX1O9JBS75pGVRi0CYo
Xe0eislwZ9wQAp7et+5Emx6kcPgnWcFF38UpSvpyK8aAn3uk/SbLpjIR61tB9dWQ
rgjT2Ovpr3xhNs/n2kRlyfB+4yg9E8Q/higiqGnb/4XJC11Q2vjYJbxdeoc3gBQo
Z3hat17FrBvpUxiXo7bj30zpL0eEFeYtjkOtWlajaEiYRLqhzd6iJsh0SrGEOOVs
rqnvg5txm0ZrrUjhsDeJpdoqIe5AmPB/TvsD5dfUGmE=
`protect END_PROTECTED
