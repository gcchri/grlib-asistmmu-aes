`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NZsTGE/KqYk6+KUOk/oijmFVhfI1a6hhu7fcrFi3a0Pfyee9vGqbcHDipiyI0Bm4
kN+khAt6/F43c1Z3w+GWThk08/d/UK4Dxilwat9gH79Q5XZgrxhgsMDICTtiu4wy
hEqzhrooNQ5Ql2Xlu3VM2Y+gePfog64HgA3MDvnh8lQrV5wa02bUU4ZMoK3naO4t
fRmuexxVixUcIiVH/5VspHkEN4SXndxBZtmqqVVjeRODQm7TT0TwyhJpmdCrj9aI
Q5gsv3Ge1bNBAth95YvGLMXcm51FcDxRPi2SYtzk4UzgiVEMAT71wz/tmIOABQsg
OVfgrKURzJUJ8mtivl4Iy6Qw3cXDQJK+HREY36FOG8pxTnVGHG/cWdx86ayOvnr+
FyDY0DKT14NM9h6/1FbaYUmm7v7YwQJcW3Boe95WMoN3aDsc++pTi9e3EPQbgj7a
ghPaVoGB3zc9RZ5qoiZH9s+rrZKWNhqLwJNQJLGoJsTYOPFXiRsfIsgnX+AzO4Rf
AGZBhqnj12enM5lGPZFUvQ==
`protect END_PROTECTED
