`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CG658Lk5bIXI5duT6LFILq8PDm5Fp61Wp71Gsx7UhOTWuHxduTzNiYoeL0P/CDtD
IuRNiQmADKip6pzeSSNIVM+Yf31vQyp9z1iNbUUqKkTMBrot+pX7MM3+eRqT4JBc
LAx7ZpIJNsjvf9jlJl+mH9vHBnRvro57MUGPbZu3A3KhSuB+HldpPVXpGXYVHRhJ
YE2KWa+3Fs2gaJKaIXhrhgNbRlyHAeMolqt8ZPUjqpqJPYJQFN65N1wuE1lvIrU1
c2IgtHrlXo10yVfEgdqoJMJXoYIg8o1bRUvkTlej/0hT3mGtxG3FPUuPLHmmI8+F
PjubxKRvizUxJZXkpJFzx/9aKh8rW6PN5cs1SGItUEw=
`protect END_PROTECTED
