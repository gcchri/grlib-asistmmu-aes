`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KlW4y0wGfZ9Bjt4NjIeN5NkhQNrAg5jCJHxS49yM9HEOxMk42LWbHLjMKbLx1vJd
swGgK2Q0U6Hp1UW6DCccb6rOf/4+S9usJAZK345J/JWgNKHqVrjGqYUQVjt3yotU
mipy2WTQtyAkzXxVO6yzz9MAHUgSVgYDgY01RbGNPoV6tJFxO8UYTAUCABB0nGmZ
MSFlkmXw9CUBhUm5xeCFeejzXrm8xCas98hSFZzCGx83f19SsFK8tLac0YMZmozn
s2aNXdc8Y4+m9hP173QMWrt07W6NDr49ko44ZFstBMUZ6WYokNCrd2MwrcYobAkV
RMWdAq1NUcpTgGXzjfBKsYqFA1KOwcFlQwOPaUkOd2h/hoNO8aMmnPDlvGAUTDWs
qAKYNkj81ASL4e+qrqIizr2Ku7VZieDYT5xX6qKfQWFFHOVU26J0CziA+rro+IvG
mwyPBqDZ6IQ83U3XkDG5uhVu1GQ76ePOeLuIQlHuun4MOUhl1Ka9JAWF9V0cs76U
oXvvMZqUBGiEt/CldDRLi0Z+rEfY0wgKF8N2TyHsRqlgR+ScwxHpHc9gaWOXL8yi
kgxZvzONYwaP14p5xvEj8Kh1xkkEa945KYGoTBJmTprCBha8cI4LAjh1fsbicq06
90r1qQTnhWuFaRKMgp36iaAbEibspyUZmNcjQKr5C/x0FmJhIjnxd9tmkARzLjFF
aqckP8niN1vpq4JEz4OH3JEVJwljLyH/PKd5NBJU2XmXKwspn6sX47udWeURtiiJ
6YrSuY4ao2ciuNtgGOiEYFLddiHxlQGBoNi4dBg6BlU2/YxLj1m3NFuTGYwOo5a3
8jSjDljHN1kWjmYH78YwnJcw2DTDiZKy2xvWbqCXbJ8aXse1NAuUgUXSIIQ9Elc/
aOaeiEG6EZ2N5Jy+iD/KOty/uHlIg4c1ghu6CQgrYXOhw0PiZq2dsFL4aPCW6WFe
hbjEtoZqoNaRxnVo63JNk3HAgRy8lF9zUlm3vj/eVobXDYXDJsyWgelVgkEPNpxZ
4+jBRMc2/zALWzgbLGlNNQLlOyBKq/kGEX1EDrousLp2TG5pMwxudaQxsW5mEUS1
tRpibqHlFzNqc3Zji+FH6xs9q8WvqGEHFDu7k5kJ6Z+P15EwgozeC7KvpiCbOCOC
B0Gi5G//sFedjp4mUIkyR3Qs76tOl7hsMRYPL1zvrPReQfqFRfLNbQcd1ShAlPQw
8/97jprHFBdVSv6kUPMWPLU9bP7D+GVRF+xdfbFVwYM6AnM1eGtZjOqRayK9rVMw
UF1GIXNdXfeAUD71tgB6C1jEp6oIHsTsAL31fBvx5jIIO/caf8uJvHOCgBBd4rdy
qbJHVss/DHH3l3hP7dUp+D7Z5bhGFsmz3D1uKM4LGJ4oAIzMq0lwJuEdq7q37q/G
GkBwSd1eb+M6ZxNNRIYWNiFrMaU+V0ZBO8sKE4epH5GzLu274DtL5Y2zgbSrhv6r
16CI/TR4W3zAYbrq01GQyRMcEVDOH2Wvs7ZsEKVVYt7ax4xLLo0DorXb13Osramv
rPzzObXkeYdOD59yFYHeq0z3HSrl3KNCIxNEpRvZ83EkPPBX3ojPpAUNgynriJEZ
St6raiTgFioP4bHh3uZ3zPQpDwm2keRmoCbEmJVeED/Z+L4KvKKieST2SzOMIDLU
dJZgJbFFaWCPJIvOaEWUHKrC9uolXXDv1DA9KXMWsOYULJg4ViSfVl2w+m3V2e3B
72oJylG8SYEa57+JnlPDZ+6OvTSfv7h/VETHts2TDBukC2T66eyDjz4i8fTRAZZK
kSlSaNhnrBIzKBDrcxasBGLipsiMZ/C3pmdNsdvGW7Piy/nQUCDYWh6gCjNJk74z
MeWyrxWEiXZkJxf4b7sPAY0VqHg+Gqj1gWOes7LdGbviusyNK5KRWEn5PwFPfdXk
XN37ZDHhmDzfd6N188OIdjuQIasL0wJ/ewut0SNAsHuDMx2jJee0uT9Md3GpYP/M
SXmUh1ZtbYL4q22EFp1RwLEH28M9GVY8bwqqDup5YbVafev0+bGoq+EeV+MXtNzI
Ghbq5iugDOes6O6ZVF4e1dz6Le/eA85qDoH4iqrtkjiWZzWhT9da2kZViflDHzGB
xMBLZbuYMSOUnMEh7DMEB6d+MNjcqFn/baTTj6cVyj+gd2akDVmOsnyXxdej17TA
IJw7yn3zHcuhUoh7zp7eCdxtfjgSJ0w1uOGFFbtOQC47iL0vUe+Z9T19fhplbYL9
IwEtY+m50JiWe17yxueGVqzSu/hVymwwI5uHpFeWwKfqYC5oqWgzJ96N0QAteZgg
88VZnB+WcLdPHfhRFh6nafYZLzhH3S79NUCHKPjmjvpSUbOSvRj/8SfUwEJuEJ9e
df9rF9uy9QSJ+1/3F2vvhpGBd19+GweW+pv3V/n/udyoKPQOvWSTAYhlG3M0uEG9
XBlm1Y1cvbOf8sFO7PVTuWJog/qa5nSgKangtGbpNX1lFvawWFiBg3hd+dYwN6XP
SOSAMhLYZEHeR8xpThc3eQ==
`protect END_PROTECTED
