`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vOt0DJuBTlujkOkqKPiOJQD1y5iS2TqJfvSJSFxBKEa5b/ohT2ULikVRMZYKELBh
ZxaUMzKlND8pIaahs6WRQ/S/n8nQX2VgHNFtXWdt3lPkUkHP/GKtX0rlhoGrZzzn
dEPHPVK34yOpLuS8v1rVxMhPtsWn6VIs09AfYCbnjZou4LalBPXu7tcYM1JUqpDH
sJiAv3GFtSI7JldzMIrWRBc8g0JA12kTC9jfhdWhz7ppIlNrahe0Vza7ry/bWq7d
u2QZHMNG46RzF0C7UF+mpQS7vmnOIvis4vrN0CaxR9RmHswA7xd7aBE+DUH+3LqM
k/DVsQmmh8PW/Fiv/a6Fgr9S1TTbtv9sYGpbkfB/4P/k1L8zeKMYnPPQhOzFmMvS
Gqt99p7XqPsJuPc84yv3EX9UI7N3f7qh+dnkN5sZPATdzdbyNK/TXu40EiPfqRy2
8fbJJBxxE1bd+aR9OqmtxCHoKw45GnJ6cVd9HTSkkygwsS5GW/1oV57AV3JfMDCx
hPgUBnTrcB1z7AvVcJL+CJfPrtMPxyLw5+qCLCzkw+x92hc8W8EakN91mHuxRINp
cFK6ovGtsDr82wEnlcIfy2UDhHabMM1Dil+4WBhGd3iiga4fx04AycOYXq/xdKlJ
MeYjHaM8wLlRpU8kfBZeTubBVSWQ7wSY6Y6GCo+FrPNX9ye9KJi0loh8OAWb6iFN
P0iEKhyDR/GP4JvDWy6QOExi8WpX7rQkpev9KspBGp9Ee9O66u5J5RyNm+E9W3vV
sxXZCrKROddqGwP92R5qTPCdqYeizBWUD54aioYuwLRk+ov1A/swHImxMV81FWJb
wj/qmT2WornebIVyac0ksqRrJjhLr2Q1e90Pw8UpQIlzpYJf0vMDQvpQh2Vk1Ob5
mct2JCKgnjsFoH8os3B8nP8qwTMtGzy8M2SOFRNh7sHj/2BCE0a6RidUjFFB3esZ
HsHcGcqxrRwME9sAVDLXlddFXibslMpedSbU6XSJH+dqQ3jKfv92G7/bSTM3okko
M4n8huvfY73re/+JPC+WDQ==
`protect END_PROTECTED
