`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lDkrcOv9Am7rfkZjYDnVaqa2A9EnaYc0YOrnPI9h2MQDAWB4/OHA4r7ING8raF3u
eWL11TGdiKx7wJH+0VINE6luixC7oifTs3NBiWpEefTw+VLCziED6luzlRvHHVVU
oDhcUzpoi0EfQfMnZFTR01krBhLRKhMJDBrulrWf6+YgClnzMRkj627EhguhJz6T
iwYVzUD0DAvOQ7wQ/PKwZi4fwwNheDwBO5spRGJHe+QowQq+LUlh1v9yKsHnKJCN
GX/A7VV8gMd5rm/h5Lmij2MJ3O8ZjU6jK8FUOVLzSlXIUXzLIP1KpvBtBzZxcHte
oerOGrKbiMlX39br4cqhjeE4FRwnhH1SqpKpigk+ZdynAsMH6jz/QJubpNFvYpOT
+lTvnoWIZI+rXPQS/5D6cm55u4+lAqtQLPO7+5T5ES4myd0GJGt89aWwD9xp4Zht
f0f/ott8xz9hIxk352tYC+0F56wuAbnPfngP04IxCA7TPnMCoZDG5TadIMrumMyU
E3MrKNvnzFbEzcQK9d7EaEYWVWivaAwpCfvUU3gk3TneW7HmOcK8wHCulq1XtffF
ltOC0xZ0/jo+e/fapOyV5DyrdWVVac2HJqWPlaSV3rGzFm7IFJe3Ttx4DWfPi5g3
RdkpUAHA2a/5KJAyNnQg5+DvChM8fYdtGMz2orzrfMpuI7LU5TlHaHQU/oXQulfj
oIQooBqgJIO2nYU1DaDdr1EQKQvaegYJkv7AXlasQyqiq2WkOTGfITJWDaS+TKSD
ij1COO9pkGU0O2hrXvNZiZ3h6jQuXu40V6lT3mwN8qddGp1NtRiNYIh+q+zzB4Up
PBN21YJW61+piigAujlKFsmp3HntYU3kBYQ2pJ7xk/FuwdMcnc1tVryAeuCSBYoq
rF4zTZ3TH5+ox3bVtxVQJaLHbdfxDUkzRkKJjGkdmwRA/fNsp1F/Kp1y60admV8t
uDIV2TUzPFsihoLHMc38zW01umcgCisWQFrZh147b4i1bvwE9RR1IvdDpvF5hsb9
eCxD7dNHrZ4tFBGaK8099xOnJoO6noBGdS7i/c/jE+zpzrAzxYpd3dEsxnZCjKrc
uPnrH4PsFiRjfuQMV1vYOaxezLd7feO7u8X0DhxFqdnS3Aj7U6gWaQiBLxYXTAqm
sbrHYvCXcfi2xHrdAgyEjY3IS4O5PfTyVPv6fJBasER/kAP9/krf5AaEzdBWILl1
F3v7eNfu5kU2RN7OWgcqn7puv1ISPNFrhKHeM7L9SMkJQ6dWbLqvFVNTt5Jk9HZ4
Gq3aIdy+g0J927CC2KPQFrqfu8u+xF40QDhQ6BueTHTSympdkWxMibr0i9TthzM8
fzl/VHsNisjRn+y2oPRAh5utm6WsHh+jmye59mgqBwI5VwcY7SpOYdt9j+4INGGL
jTfS1qOqGKg+pZddQ5MNufiztueOXN5bnw2qOax+6hy5OF/hXHmaN/wWHU3xLxNO
3VcZQ7u2I40FVkMH5APLfJrlMgYqxRLfqG413LLH/CvbcdTAZCJVdLcHxbS73RkT
bbh7wsqA1bJiCQ/bLMtvD4N4McDRTZqslrLbN3y5MudjADev/aHLWfHiB4whJWKj
B1MiQl5NzELVZ2rOb+SwPJj2q1zH/JMnW2+Li3vfMj1y4auECtAQ2L9gqh6D70sQ
Ve7oxScxVuODnInG7YOOdgIFmRTHUAaZSTyFe4HkwE0C+mG2wKDxOmNvc3Dr5CYv
eO0zFMz5I0aEmVX+xX0OQ8MnU3+NBUgo7eWI2Fx/jP34pFmtPO5Hpr30VGOuvzg3
ZysLkvVc/1aSGQ+7U2k+FtjLskj3WDThXcGl7kuM3QCJoRx/E6Pt4qqhbJS+s9wc
54a7RRKFx42tZGSL4z/H4o5fSsOaBrPIddyDf9lYbwwlPZS7rD+7JWy5pvpwA86/
UvPbK+okZZv5t4JQBYo+dk9QFH5aDldr25Ez1LacRBrUpfGKzKfVT6semdqrAfub
ZlhTkoRMSr/w1CrpJ/1miO1HM3B1NfScOor3vlfkSvC8jne6KchvLRP5dABKAXFz
ew2Di4V8W465+9w5fXeLHl+HioiMzkzvF+wXEldnCYlO9uGtby5nCJV0ZR/3O29B
zzPpciW82gI7Cqb/i5GKxpleNepFLLKhZxGsEH8/dAiRj32BDxdi55/bD0bbGmdp
x7bL6BVFRZMqZUFELFkq64jqsHCa0Q/dw1Bu2D4S1KhCO/lt1jxwtW4ig4weFwK+
yoAb74CVVl8N/VHCEESBNoR3wW8Vy4kukgmO0Eey8TkXSSNkTK+K9IePoSG5liEJ
0tu8/AqZ0eNnB46oR3+lSAQZyPM0F1xft/WH5Jyir/DJ01V0+1RHRxKIVyF0bdaM
o9z2JGDpdI0qE6VBZryz9wbqDhIfSZrGQK5P15/ItSpcpToFVujUaOEXQuEsPkCH
w7FBzZqI8b0UDNx83+i3S/ursU6TKuDsK0hcevXME8zIhhH7YLD9+T7XFtkBV43D
CLurw4GVFis7E3+zm4dNTkfBGbEj4WfnnRwWglph1WuyMqFYn5SmhhmjW2sza53e
HFhESbVgJiGkRZ3aXOJNZfkfXZbjNOpnD6WFryTgLnYT5fZBvCwoOOsiqL3/Jcof
f1ddcFa/7NvJ9uxcg+eE14NRV3Xj0v37A8e8W47zU3eWRaK7JKHyg8dykgzPLrTB
o0n+HlVEI0mfSL2lCQHjQIAHPQdCcEbcTQc1r7FUHuMclISAp1W5oXd+Lqcgo3Sz
R0nlPy0DfGYaV81m918CAryCROUJo3d0O4oQAdoVgmdO9fCLGSB5bfQQCw3PAW/F
62opsHmPxGigYwM+VV733IrGBek/acTvhkomhrCxi6tAPNqvzxVQAtbbBHW4Rn9w
yAWDqh5trvttB2esPqOSF30bNU5d16SAhlU0tsrzoim1IRcQ61eJ6a/G0d0hRfyB
AZ/sdA3QfEZRQY4ziVK1CpkpZ5K71R48f+UdXv/n5IyFvE8f2Yo/N/qZjSQ/NUee
hRCTNCahMb+mBcuZoHRLY3v3msbOomZ3pha3V02wDxjCH71b2OSEcErzfRk/qcuG
lHRcEZYTbK+aMnTAXdGBbdfV8GdBp3oOkVvsOqWPGfL5lquAzr86Dmru1jMcxFbK
EzWnUb01LaRVWwE33YJwNbsKwoA377MVw9AG26TAaxq6Nihz8yvRAvjh3yQhSDAb
9DcK1fjNP2lz2llFMi7jZfG4K418xOQMHikooKWfY2nxO1FbP+v38ieWGjoxCNCL
VHOrSk+taue9LdAAb+Zy6+pxW/G9sCM4s5Q/PT4QxYAkPhWXxIbp6ouFcWKiNQsI
guKfr5692rY2ZzAepZO+FMrIO25TgB5E4285YTUTw5r8IyZ/BpO2LRdnADS18PP9
k55UZWSuRcKcr7UwIBMJSnWjWQa84iInieG9KAqjBMZrGe+zZDUspThYuMRsbt3L
ASMe43Q3a6I5Ezdy5jWkrj+OZ2ik5ys3z1nAr/g615oUEST06jGW3okHgvz6gSBS
d0unvdz4gfaHeRF/7KV8NqAX/IMrsoyfuQQ1BlVC0bcOBSPydcT6AqW9Dqrpt2h5
oHhyRUjCVgOlf1LoRRTZsywD4ySlyY7BArdg5G0a+xLE5sq3rrvyfcbnr9UOJ1GZ
ONtDm+ltyBPQsqA/sQ+gv3rxzJ4VWQw1qR/9RRdqBI2waPCY5htduKAiPjRcuYTv
0MWSjXH/p5vQbJmGXMwcKVpt8bWujnrLjILqdw/Hs2g0pFfgQxAAvz6v8de1xki9
uGCDQFUkB9Y/S124V9EIem6QUY5gwb97+dSsoo4p8aoPWo9Owa1ODZ+SByL6+DMv
ELR4FKMDRSa78fimrLFhYC3wh82J+OAH+LYSPbaqVglb2sRnocl9W8u1g4TaEET4
K1JcHrjwQlGTI1KboqC5P5HmsgjCmkHkhFBkGoOzBK/qCe0GuJIEV1AqwPrFT2gU
lQn/iHN09jti0L5qrHiElUoaozglS1ANr9kwyfdx4vE6sbgKDik5ruslHWTHrvJJ
7ucbybZIH062c7S+Q4eUqBvj9WLatLSBADwk+edcJMIKN/QrwkFv1EPPIv5rhWSe
ShdtXoQCofVWTwesah3P4rMtVDFHdkpPg8XDx/gYn4zMugZo2GeZnOurT1ErLChV
SIo3NlYtw+eEHCByh7Pxf4JmHs6aa8qIzriPFwl6MF7HMnplntixYoi6wt3OGb7D
Zo5l0YEUEZ36b8o7RDQqYKw+/nO3JdZZvicYJlhGsz9EIINATCLlJ0ABsuakH6Xj
bSmIPKF+XXmmN9YIV5eVeBcA/iCQuPdaGtpgM3khj/556QoVfUFq6pt4WKg/SWfX
NkHcCmKrbr/b6YK5k++bnvoG6As2in1XZ9HkEzEkp7/NgE29BgAbpk0ABpdhbi+T
q+lsgze2MEidQsVOd3SAam+LmwxtLCzNnMWPwqJ3PF8oaN903BQVxf+HtjQe3eXs
cfs5JoDiXhoiaEwJx1hCrgC6Toi0UpDmdiZTZlYTXew0iZbsdvRgtKMHrV/a6cG8
zEB0iWX2n2v8OB1PPk5ATdX3TFtb++uKmPayIJUggYjVRpOW6250T57TOL7rpDT9
Eb1cE932xDyiOG6rsn/WZzQhFZ9f3Z8opmSD6x0YWTbDrP1LN497NVPEOs+rJFiY
rVqVqlhBEZkB+o1FdbCkKxIeAGvNpj1TiBhEHwTsmAEp7MwPJxL3T4vg1V8E6MY3
S+FQfb0T5wk1RNg6Saz8G63z7axRuPQAGCIydoRGbdBLf+VGcwnCDxvXC1X+PkOp
z7uts21iUicAlRuE1FdkHYql2XxJUh8pB+nE+eFRF5zepC0eutViJKy7JN2us7LS
nUF0KBnyUPlHVfd8FEycBEki4w7uCOaQCAzedtndbKRu9nASiAO2ys/r1owG4fPD
FBnXUc4TX20niI5SUzyx6li/SYLUOoBqrpjb52eLA5BLmM4f78kmzqg0SwUVVxl9
47PKwVSYZlXNguWh4rG9x0N5EOPaDKZbplY7Zyf7ce0qHYwCf2hA7fDOG0fcRxKl
BmWDJr12odm9s3A9nnNPJrQPVMqYBr8Hi/+NYpNlQvUOgvRahdTMF6iJ2awBUnlk
7+W1VKGzodqdQYuOxdhO4eRSclqyrNCQYo1WzTHjmFXRu4LoRBxHjSw4WPDHx0yQ
tY9oIrLFc5bY9C/NgIPT5ShnInzIclKEhl0uVaxpGg/lYQh/K66qqYBtEeDViLh8
JJs8tnTsEfXqKHWGcD66SNfopDTD+iTJuF1wC97i6t7QpgnDilo5inxyRgVa9JTK
mXAC5LIfZHPNlWfIpt7UW1nd8fJP8WnGS6j8rBOsxOHugJ3DSVPJfWI3wbDJVpR/
zwuAwCy6+JvKJ3Y54QLK16BPCKgMmIGv/tvNSpwKScDsNkvvzsvoeLbjadAJ+SCP
z4T/zy3u9ZPveaD0GpOaGSdp3140RgnVSBJHfBblPQq2x4L1wma656x01URU2+vp
txte+W8F3B5/vdJlwKzcF2spL6uXGVCCdQr77WdkQAcSUdfstJoIyFeIlXXatgVe
EwS3Ody5Tm7a93vtvFLhY7KF0BaHJoOI/WrNRKvT+N7OQKMWkCO7DNoLMddrMdYC
/F0BNZ12HtHplOx0SCYjc4aw9Sge/eUnPdySjLIBqIvraBMereP7c/OIYPXHPVEH
RhoIzQL9Bw8YVXe4y78h+ehEUya5t37isacQZSDNHv1xF9ELwJjFxUcvmY4FOx+W
9BZe6hPrsM+PSwBLsboMP5L6RLIbWxRc5aVectEm3osmUAldm/nZui8/7zmBS4OZ
cTv8waS5AnyXDIgi2RhQB48mnopcUvIKXxYR1Wvx2e2lXvXqsAUA7d+AJfVySHr6
HIPMqBg3qyq8L1/waSi+ukp2nrvqje0/Rn6tnnHY9i3pQqBOZkQ4hbmqzw6nsKxb
5gh6t+ilAvDDwIJj9YAmiLKY8R1nkwTzzK1OaidjKQrZR6ObBtPE2aGu+7z7DcNi
BpUhdAw4Ijn3upE0WQRPhzqXTGsVvEzmZfUPzHqiLOlGj/4zvj1tDOfGr+v7Fim3
TB8ikQA68nE2DFvi3O5U3JwEq1YKqOewIZOeXTS0aoglkAoeAhLxqlNQ87PaeoIM
/xch5eQuMy58ZeOSsvq4qoTsYNsI8Ced497JHZdirbXrm65+auSVAVqOdGQi5lbd
+CW7XNN173g2aZGoP6Fol6wQIWgjBsXACG83rcA2BwG+qjUFu9046vDvWvqOT71i
MNFjJoLX3bS+j7q/SHbwO+xP+gerMbIoxLHyemtS9NF0cCDuWQosSAxlkLPz/W+e
D/w09eGs4LIw+CPTqrLsUN90FfmBFdCCliYdH9slZdaYzS/HNjVd53CM6qpLirt7
lby1WVqm7UuMvyQz4M6tJz8UrPLFJ528YgT6eDdo/NsDCDJ52F1Q86vSqCAC67vO
ByR1MWAC0rEhXRPEV2h7huoaYdayITs6e5sPnAJIlixzQ6BUzlcdHzdpdSLn6/Pa
XYBfJhDXtsr4H+pA/VRoC+eI7i00Djr/1F/iJBI+PSbjpjEeGqtHAADDnOFuv4h0
G3rGWz5sUhBEIMS/z9ZNB2pm9oZMVLsNRvHPOxtz3FVZ4rHm8sLcW9XvcTV5/ZnL
wLnO8XrLvf0oqZIkB1azQcT1rsssSZPo1H8PMxyq3w3rsfgo+peXHDKooj9QdQIL
3sDHHuoAhVVwWw3wxjvD+a70Gd81y+g/k/nyh1jQoUBs80nwYzFUPa3wcvnXgAkv
j17WYkS3ryRl+6c8rWJZBGgA8WF9mMRqB51G/G7IXaymxw2Dxs2YBa1K+3jd7Ual
08g9NCGaXjX3Sx+5ojxNqWZtz9Kg7Z3s+neDECFZf8z23AYjP7KILztjBxhTifSQ
RKv6xg0aTfHwhPIzXkQL8HUCJwypqI3EUNCJL/N7zg6NxR2nlRqeYOLRjuTzujhj
86XcnY4jHjO7JU4ulmmj8Jq2qd4WSn7Ht3saNYhBtPPO6PivmA+kybAevWIhxi7f
wvZpf64W2JqtZaCLpbeRi60QvXHo9xKOzU5AqwZRx45VC8hT+tgA5Sj1YzpGF3+G
BSbKaJjm+Pze4Z83CeaS/bk/uasfaZv/WqEQ2CWGkSvFi0axM+sAD2KJsqnPix2z
EFFtEFYLpkB8WBQL/lVPc5gzKUdd99wGt16T4R2C+Eu7R7dp9kPtdsJn8jJ7ZS/A
9guA7CKxI/3YTlvhqmSwM9hlHvu4k+PJp3v5Si69XOd2HHLGtDTH1xGpMM3/vbZv
3M31pRczlDpPaVn5T9tzNiFX8dd4tKLtpbmsgJGx6sR87FV4vxAPEpvHA/e5sI64
0doPopcXmRixUZRftqgmH0+jTYGW4bkZsXqJw0K1iLtwTss7nJ5Cgutz7RUEAnhn
DMwJiWOzKUgavmz0f6vRViJBINfx08L0TtAPO+VN+TjT8J/D3sj278r2kCdAfkj/
C9ZC7TittA3KeNbGZEzqOgxHqK/c2mtlOxOnU3Qcnsv+x8+YTaN1Rgjpx6l7/J7K
MGc8jZQ4XsV5/867IaMLV3VqoltLArT0qlDT3K7QaFe5GF8Kom+ofX8AIxTOOUsC
XIVt/ES6o1+vNwbxAHxRFmEJJvPvRQt92bSXwXVT4m/wz6rkiug58ZqkaXIVnE8i
oZ3m8qkQIH8pWaAt9sUBJpK30xyoZ5dNUO6OH17RXH2gp0pw7UGAlcyLkv0xhHuZ
HrmvGgb3QhiitrL2tRooUChBUTEB8V37FjaF93/ox05ibOytJXDf/D/Nm099Z0WV
Gx3bLjGnFBQ1J1ZGTd+6CJ/JGqnbHfM0IZdU2SLrrou/1n7m1ycrZq5qvt4QJ7WZ
NedlXJPl83Gs/Gyvi1Bt+IYsvd6qjJS36DgCXgJhb1ksdBTQFQZv8jGRh+F2RTH0
UqKgznniNzRc9IwHX4HloLqsohLoOiRS0imZVA3olyR8KYcC3emYAcYK9aZ1Tl43
yScRBv0VyuF1UwltsH6jfhLoXQdSuTQAr/hkTSaNNfGeW8Rrmmu6sYDTQGAAjEmo
V2PLoOwJdTK7GL1qpWnm/5WIodicqgQxXmOG+Y0roXdOGFDrArlMez7i7igHPLZw
R6i1EPL6lqCzNR4x+LVhNC5GpgszGq7o2Y9ZJfkqINU=
`protect END_PROTECTED
