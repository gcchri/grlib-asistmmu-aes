`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I/Bai3CrqHp0gjC69QYZx+yfp4T8AC+PLaUDVzuWlOFPc/cJWVBR7vXX239JX7De
4oQQi0EC+F2r1MnZik1PWDq66C9vRmJyYLa2CNaj2DtAGFSDtvlVDDbqz/zMCurx
AWbgKHzINX7D9SN5sBCYlG07OWGHfpLwiGtax2lO1jKbU5Hr7qeYllVMAhWp1WO+
o95gIy8Ao0W+HfCgC4wMy52gLwnNOyuyKmYVxEbtk6laI99AASivbr8/KM9fl+Zt
Xx4W7jZKx2mAXy9Mq9be6B04UmIFc1fTTx2T+OHU9Y+WxlYkHhnRVSMKvftm7r4l
cTJi0PyCksOerii/O6h+XCbinRiTsVvSql3xI9N8heMv2KPNi1GIq55q54EX56ZM
eV72Ozz3m27egEFSqWs0PlPX7jFhBpdWHRtL99axWphstLpQgtwJleiykwpNXaGg
wXuipP5lV41V7snU9y2THFgbVYYSK/kzZSKo2m6E92+FqpwqbcVaDyWkb211l3Rl
i6B1Obs4rdg5JSJaVns5gOauah/yFMAdzpYklvKjeztAksi+Ys6q3ruzGdcWydTv
ENOU76fxOnfV/84KWmBE7l0lhNWW/Nh+Xp6M0su40mawT+rTRZfqkNIypjUeAfc7
chcslydHmTKqiPc4XHOh3QlvndQ/mEWUgzbu68KExnwrOZ3TsWnGNREVtkWR/AQ2
ydtUNr1lC6yTb9WXHg7agJ+wtcxhhhbuXMGmoevjkHam75GV3sT6wVAFbAHnYG2U
EgVFdMn8cbFZtW3hQABaFq4215PoXb7Sk/CybE2nCOfz7iVP4nJC2VlN4qzTBVtJ
`protect END_PROTECTED
