`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0t3rVP/cz0Dpa+7mxUuVZtq+ex3O2FCPoPrESKDh5lz/yyInHyrSz6mNkI2O/Gs1
XH0nNhch9iAUhZoeCQvST4zqM9Kwr1+wjha3HL9yCMkkGReQgokYKB/FW6eO8qoY
7/E78q71IW+S8wmEG7Fa/SIWsMuCG+Eck+Z6G5TSBIe+Ttg/FaLtcheYH9/VE8cG
VWFbxcwicC6z/2p4X6EanmDXEzU9Qtui0oLhFSp12TiAFe8LQ7GjGykUwngc5Ar1
zaMRU2ZFs3qG8bwgtDqimC4oLASGoF3bN+HOXX+mC+3WypcXmvQXoPFngxnlY/HY
yxrnpDESxeK2kFq9usJ5xDUuKiLneGLOiO1ko6T8ri4=
`protect END_PROTECTED
