`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i0kF3/CloPCKa8vSOhtHi5GCb8XRXAGaGiI1zJ0RwgLU/JKXuqeS6D1L9I35fgBj
rPAlCkq2xWc8RULFUSXQ8C6OqXx+x9Zf1zUswU+f9aUHHm01vvm+iCWsAF3fX9Ia
ElH2BQSft1uShETRU0jGlViDN98DB4v7e3LzAZ8nAj66zNtuTE+ojgHk6CRS2qRU
uAqZSLp9xj7E56HkVQTDwvVeQIWsOeEfNIgCbpDC0iYeSXwiYNey1KY8uXMyIl9f
HiaAW2We+0oxxTtWWEMcDJkanOmg06wzqX39zDHZEi8NDbPghGNkVniKxvQcnexe
ekubzBBs3aiiyCYnOkn8lEFc1mjuxFuOsi5Nn2Uk560XofkO+m5KHhQg/CbjFmT5
/LLYpNXcld5zieHAMqEV3OumhfAbN362qN3ViH1xwKttGoCAHp8HOC+q5jeGZCLp
rA9grpoVcG8Ss6/wvhv9U6LLkNG7OxOIrT1GL0qC+VjVq9PMjKj+Vs9BE8eLt9co
ZyHOE1LukPrB1VYbAx0pT8XosYEAEXIeVPGD8Hix2Q7+gDVQBzqMRXM8//zEUjfo
mRwyxdtYmh7zXDohv0nXmmB966vZ9X7asV0kiYbWD94yhWZxzDs1V3lDLm+LMvR7
vrCs2W+Pp5GiKHBATnmQAA==
`protect END_PROTECTED
