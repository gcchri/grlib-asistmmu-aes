`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1V92EEB2Y/Zhqe0DTKplnax1VPjgjWyKfiCjGeZevdNhtF2fKsdAe4BV2lNU4EbC
URSRmXxE7Bj1m83dY3Kkai2qa38tiu+p2nknIlrfok1sowgQAP2ciTV7i4veArPy
uS5iC39wPiUXHKgoAuvqcjB5V/vzilM0bkhCsT0Ioju8S0X87vcPx0SEHeYNBa0U
8YDkULE79AgFmAdWTXskMUEgbXEktt/U5OgMPnzNnr59XaXCr0ctirYMWbuhM1MH
6MVF735wcvHYiobhUUzSxhGAcuIIGM9pIIioQ3gip1jGr703eN7bUr24v8FdJoqo
ZYye7CsMkEkxc+UelwpKzoaxNMgVsK/7GeMmcil24za7lLLq64zd6EGtTMDVCb59
HFEpFiJ5n7PaNW0L4+yaOf9taDFf6SKTnx1SwjYZTqgLN1dlMa/nL1RxiJIJ9DyE
fkifP3khZ54pCpAs9vUx1YY7seJT2DOYX9YspeahvIo=
`protect END_PROTECTED
