`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UuwtJE9pie+NN27RLc8pQz/G2bqgshSaAHsy2IHobl0hTOvyaLtWciirDYhyn7XW
nI/Wyj4aWM6pfQqXKSz471XYKXJWJziQsPperIhlwrYDK5vre+zzKIh1/jtj8yf5
6uJmqOsdePdpT1lqAUojh30kjuFAggHMVHYkXWp13wR7QfhDg1oSOCRnyKz3wOdV
9HPzIT63lShcUXxiodqmUmz118JMQcVCtO0nboHnjr8yX4F4vAEmc/8oyLgLjvOi
HgNqLr8UZzdITOT0dmofjA==
`protect END_PROTECTED
