`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TaDvUyRZJn6LXdhXVPmqOE5F9tk6jUreikYp/PQlbP8BBsldp0qXd0JQy8grIOQz
8tEwb11az6JtQA8a9uSiJ03RH2cvHAETRDxedhLhC4h4csUHf/xU3Is8VY6e91Yc
klPLHf6kz0d7PhQ1gtmCltQAA/9kGBaztNNic77F6s42UxnQTr+W1m7iA5tFYDrQ
ooummPmDKPkkTQvdc5z/07a7+qLv/Cl3xc9LxDNZ6dMk/EmondF7KoImgnPKPPmw
g/8T4uT1KSaHyAJv+ckuoBfrS9iY5y3G4ibD73hDzQ2QVxNpQpCevYY5YOnu4YFE
0LKNISDkDWUM455JEa3znM+zZ4ukVq5EeyGaez0D/w4Wr80TPNGVKpm34jxHtq6a
uBSch4Fb8loD2n/lAEJhnLzqPYr59+TnN9Pk3MTDEyDOlFA2Q6nZvL4T+kvXRRuP
JyVhoJY2S/oebNTBTtWTALleEZRien4dK2Fh3C4Rw7cCAtYnI/jdvorHEDCESVGG
lanPxY+VN6Fgs13DPQ5LHuLY7RX+srx2sJ647LpiEm0=
`protect END_PROTECTED
