`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z6SFncvyz9N306yMf40hG7BZfA0KAg6vMx23wgJ4l6B9tH4gIJgVw/acj4psZ8eX
Qg8YwRzg3f2IN41K3OJpWcAErs96ZGagY4vu88mBMXbeM9bBCxX4KKDu2aZqlFIP
VDVmQCAMQHF2wW8e2Viw/gLiviSmDKpEEmWI6FReUioMJzjUYQ6SL3Gatb61a0C2
sMik2sj38/M/sDkG8EslnIqHTJZLbgNbBhSSqE7ntjmNUzSrxST2lHBTI7rSE7CB
ERraKIkatED4lkZbpG85pKJ8qwjFwhpedPrxwT8/qULM41Jo0y/SXDaSOMDa7kk3
PtJTeI9VUEa7L5qa2oLOokYUVuGcQBPgmLlBhiq71x9NCLsm6he0VxjFKAL7IWah
x1hRtk/MdLud0qY3sCa3iw==
`protect END_PROTECTED
