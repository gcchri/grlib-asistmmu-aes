`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9KYbPPGgaah4GPwKlsKI0Q8KuqFvI4pnh9dfEUfoVc7XTwTBFBH8A75SwH1ziENX
uAq3IT+4rRbjEn9BJqqGKWSDE9Ryj9+Fo2huY4EbvEbClSFEA5atVt4MwKpXoi1R
G21kOM2JNHLl61nlgrRWElCO6/YSwyn5ZLmSAr+u8ERec1utLJIsl1qTNuEGFczf
S4+Z+47bkK64HV3mbzUt5ltxsC7TqbEIlxdHxE4Khn5V7BBcbmORjHGq6T7PcmYE
joraPIIOgFfk6bg1PRweyOKG+SjWN4XDenoz6BdHOhapjazH5Pvl7RUt/K71GWav
fqwyL4j0xHGh+5jHywzq1EMoKrnoXt/284SF9CYx2S79thYa08FaYgWqcYJ9JBG4
Q6kxxwG97BseEpmSIrhuctzxEMM8v5QFmRibd8gI8w8xKD7s/zpWZhCXwCEmIfeV
`protect END_PROTECTED
