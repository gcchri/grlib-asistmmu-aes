`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cvbpPV/JyDYHv53ilUlLkvB5LFA+4wfI01Qx9vlDQ/aO6UY1c+eZ+j8JsA+lNUDk
qDPYYp1u+n36XFlJBvl7HnuctxaPyj0AdwR98UvQyxboJ3izLWmpoX5nI56gra90
s6QuiXH9XZiY4k1u545eY0iiNFKnt+RnxEoqGLKskZgYBDUt1CglGOUN4GaaqewR
OK+D0u6DCoUCbYUv46Dt7wQnso6o3vxlq7KXlSeIVeEFcYt1d9X3mWFcOJxEG+VE
nxSERfzmNM95/inqS9ifwgL6IguImASHw14PUKYr4ePoIcGa9HoyYK5pQ4LEc0uy
/xJTWgP6JOuJNEFKoSbsieIRy7oypCA3K0MXBrJWnwZnyUV2GMcGKCfIrgQprnsi
pVWGyhQ/IjqLIn/oEc6D3dXoE14BSC4CcOS9rbvIOIrf8eLG8/B/ntOPxSG0ZXwc
BF9z2gqUwsgihVejUXkJEKcRp5aZ0UBOpHAGEhPgF4Josi8ml51T3DLLNFZ7K3gt
QMEtmCiYS4yQGNUVsf2IIQzlbonZb2aZDLImvBo6cpEzIbog8RS590GYugO5MeFc
Po5h85sgdueOA31Xts/HqwDFoEdzYUJHJn1Rkqs7B78+wW3XPWTb5BPaPwQBTRgH
6wXLiOLkSlRAZ9KFS4rjETLHGf3D/nGv0TMVP85Boj1jeFL5gsqnRCZkNn6wd3IH
`protect END_PROTECTED
