`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GbHklUpmL1Gb5XdDP5TueU2kqRbZLkYKf7U2hv+B06qkNqRaPsHK3AxVWjimzJMf
CC3ZtcXG6OtwG4yv7qRno6ujPKhDZa8leneXj+2i/nfvEyX3eU32kEBMWAhxEcRu
SCYW7edwGaoqp5CP62OGgHJ0nEcGQcGOwv+cu1SOlCvzt99K8hb7gtTlQLPqy5gl
HZHRUMs2J07L/FfpFWE6WpF9baoHt1dqaOF6chnnQIq/rqC71CILgxPUuXl3xPlq
mDJzMP6gCJCmPpfmv7iLtwmvoemNcKk5ZqU/9k8qeti8OzEyYhp5gLBs9f/+3dAJ
qLsEvv1k8viyUyMwklLhb81yBoFd5PPQIKBeWhvwOuXDcvaOiZm6b/Tu/+ErrxHA
sfFsRitUVOzhG6eOFHqfzv9nkIzWzf6nfGr63N+rJAW3VPd4jCFws582/Us2T40f
QZ39dbRim71a1oxnjGIDwDiG6GwZuSquK4UdFPhpcpGnW0WGL6gnLQ2GQJOqUKzI
f+gumr96QKoeZt4lsnDOPO+A2PYsdW/r7/YOSekISmRNnZAvavSlgRI7o0qiF7jb
p2NEolMvAeuQ9qLlgc7i2TOiUEz8ZlGPgNmPLFePI2Q23m4pS9vVPT9KdY0CbkQ7
dvcIvfKT2CDWYtfR+F1ng3IuGeEBBzFMvvWzckK0whrLesLN5mPM2p8GgmDTLQwG
F5q6g12czrmbGtZ/oHiHi9ZlQfiyVXuqh9z2K3qb8iQ687QkSscJhzjERJ0+O2mh
uauJwapAscjyyZm4kRKzSVO2ooqB+TMQg3KMF+SLvx/q6a7ZCvh+SP6hSVlHnn9N
Pab1H56c/32JZ7U5NOrkhHRqZY9+pN9zMu2tarriQtYNQ2KBi9hfl6hGiX+mTh+r
SWfImZfUiswYl3wRvSxErj4PdNQR79l5c6UbRHn1jNUZGJn8PGFiv6Dml9crqZz9
xOKYUNtSuCsmdW3q29x/kwbGyjltExMu3vwauV8/vRR+nWQ7Ql/iWP0SA3kNC//K
VVkbOQDuK9X0kLIBk1Ubt+y4On6Nb9GOMUtSfNXMERJVg+ZFH4j9CoAMtPqyXgtA
47Q0jRx2pbTFRMQNV2YfNwa1RVbRUo3AEVtH+dxAobWz4bM+lG1vT5YSWE05rL30
yypKDU3bPNVDhZ+QWi4e0COnKUyW/TxzxUKERNGT9S8uI/EufJpPPdSwBIr0kQJB
3uQbY8xDPTbxEs5E7NhMpt/VFSVo5XcsObWFAjjzFOhHGjwQeuF8DIKAGpRLnm+Z
0oDuNRSrXVqzSu9nxoj78sPobfMjRNGX6mzTOmbsUJsU6y4uSbnYyKFCp6YvgID3
fnfA6sqx7bzZWRieHTRYiWxZURaNAPSl4wBRLRVOoOSiv7e4aVBtjEvfhvpWL96M
fZY14kmY/jwVPP5C2gAMU8HDqASOeRf7XGR3YXmvk1Nlq3Rbo9Czrj1dlx8dHGbl
ePiomIVwcwjdniLLyTLQCBcrCumXkWdAE57R9MhIRHjWVtngmMylEuBksGF1Ccsr
BB9d1AzQmutp0aPQ4AAD9T08tAV0Ypb1IusUn+iXh+1yIkvk9pNddVX7TMxVXD71
5LCIAqCDNN+jdw7JV+CfjHdSOSdgt99bIppGh5piQS98S3RX/20qkl778Vzq42jg
c81TV1Bwt0BeyJ5iEr3Y3aU6DJBCEiiOfBgT7L4RlIbFK9H96zt28CY9n+tvSY+Q
eHeIYqt4qG3zpvjEjb7CnL1+vGLdqBc3V49UQln8/c7HWYxR3+7k2tkDrywdPYhi
D1ArkkeVpcSctDBU76Lbyw==
`protect END_PROTECTED
