`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5WQPA4W89e0ztRAnSHUOZGbLulk6AXITwdEQqnPYOaoLK2H6igTovvGMNd163C5d
JcKFkLlE7wrMahDlaz9Ub9LLLSUitF6sNG/VQauvLfdq1RjFhUcrjuEMl7VUer5u
8rfrv27uCyXBP1lYcUypCRW9wWvz55mib1xgbQWVEYUtj5B7sy1qLCraEbe8rjtB
nxx7l7qsq0/tQ7W7TC1xCbTaJtsSEVva6KOo4mo25aakDDuEJCOgbWsmvmqHVTu+
Son/P1xkM9eFHkzHqChldSHzbzQf3NgH4RLcPRKTlSer2ePrlFkCVUOfhiOKZZE2
W0rmbsjP2hJSmsiSayrjZrvecPBvA8Klm2xT1oIxoZjI5c18IISM6Xrp6bwdXLz5
ko0rPoc3U+p4rjE5mnUutLrsGEton/w2mgpZDIcRgkusJTUKZwVhO3go1OAyAP6R
xLW6W/HaseUAnu08Y6QtOkMmW8XM6pSW6i2VQsA2FsTM0e3yYpnrP/SHiKQBBQuL
vefM1tZlrTa2O3NA3auqmvHsuAUHrRMXh1HjJ7hOd3S2dfWo//hyNuND7QPICpvY
trN6++8EIHF8NRdnK1JDp5Gs05/PluPnBOO46qTkQ4ubdjk8wGQYMAp6PSjWjTGH
h3UXooPpMHMYs7sh/IBt7XrFQbSIQHVLUMRUU1oWglnCWf0UzZfUSFq/ZjviNWGD
QpGRiZphOcM1R11dmHiZ31WMpEO+18YLYmxIZfUV/Y6zhj36qSBqknbft64HraJ8
gjHmC9Nm6HwtqY5K4dX4w6mU+Au0yN6bWC4hfwWHoBHyO7YzDkRpINtRe9E8QLMU
qka+2CAtt1VSdOhj5jfj2Uf9VNW5JNIPFIg9F0t4PIVbW7aMiGdxn5RLCciXSj5l
QgqsYkWkiVouil5jbVvRGvHt/czqgT0vITaGp0oLJEjGfc0idnfouWg6+aK8tm5S
E5wZ/pJrFXOFmvNp2LdpVE8jPMnxazm+lJZio7acGUncK6sRrO7EwBKYNP7dVtBM
`protect END_PROTECTED
