`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nl5ChwXSfKKr4JTM8yuLLsx2RRWGNSkfI3wUmTUx6HuH6iG4xb6aahqyNhRwKY42
pGjyNOB1yXblZKuIc/Cx51sNVPheE+njtSL8mmgLhcFxUFcoQRRL/YyWfbnfeyvu
CdIOIKJydjFwMcsXpjjZyaPfo/Ik0fVLRm0iZkLgmDp4IuceC+OT5tvlvaEJ6OqV
tVIrauZDDj2aN+iBZ4Hoq/SlZuR0YXUGkJH5wC44MfoA76URl1RdmcRThWtibvkA
6bNc6EMripDe0c3qJ/WN7wtfdMvvEmND30qDMTTMYloeTt6Px0S2/Ou0yBinWMtV
ds9pw63mzxj3DF5HjypyOTNWVmq/lmmzPjLRd0xC53zV4Yrny3xzPPXj6K9RaLEP
vmiXAiM4TP0awAD5Hq9MtEBafFYVNtPpbcG3ffU81hnkST5SUwbf84tAU4eQJavR
aJFzp+8LGHA66hLytHrxE2L/unRG/L/z4Pjo+u2s/A55iBThLSXjeHR8MH7X9VN5
H2zEfM/6erVD0+ow7jELK7r7a9S+8M/Z0YRxO4Bt3VNvuL1bsTBlIPAZYaTRXo5u
iMfz2wQgyE+pbDt3qoEn/gMCTybVhpsSiaXaBkmL+n/6C4SI3GsxmFs8ip9GXJgC
UB1+qtM61gnGu3eOcga/N5Be6CGmd+qfP4aFRGvPdYozNDUImp/m2CpbO9h1WWSt
6Wwyqa/aR9aLtR5zL8y+oWGHdWhCeJL26+fIWj2RUV/0J1VeTydVPqneFgb/JSDc
lXFJ2gdFs1EG23KRG9r/VM4bNPnQwkCwxrOin5J+QsC4RTdU+rToBrHhZ7lel4mw
rrKjCfjGSwumZt9cQVy5/61clSPaXdQ5+FNbVg11COwpQ59rH6XGMTo+EloPUr88
PLJZnpiPxrVPb9g6feh567de/5HnTjltyo/JO3dti7XQyoDCOBBLo3R6TyAgZsU1
t27dgIOGz3e4Az/cyXRTms7xxgpv8Qe6U+9jLO05LDU5AncokVQygumIqk5aAMxo
brm68pqet5jh5klyOZy7XTD7PoRyh0jqT2OKKzCcuyX5LkSr+1RgnMV+8iH6x0GI
oRuzF3eP2JPJ+qWERYMSzA==
`protect END_PROTECTED
