`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CJMQw/OzIdFuHtdLDT/aXZQgt4FcKacA9LvegOnLIgtmE1wpb0ifdayJCdsbOy61
vsDw6+ugDxUL/TupPemp7OIZ6dns5u7ltLehPm91kqt3p5/46GL7qlQURRgAbO4r
eh9Zohq1GcqciuCBtRZngW0vOE8IOsMiOZ/KAppdm+9A0tUjXhM70nOIYAbBPAyG
8bWbUJg5/gWO4HF+UpELaZh7Gzgfz4+cwPxiHfLxVAChBy5CrxGxywxIkFOLgzlb
xxqv5PZQaLc4N2UT4rXce1AyB2G3VCNjRMTcKM0hMvOiSyh+Bg7KaM8bBoXZ7RRx
Ov29/fI9GbteRpXqeZOP6f6nF6LpP8Rll2QRy1sfy+GS1z9oyA+SQ2nmJ6OcuZq4
pviP2mzPgDtX0sCDtaFyzdByZy7HK/i/kS/FCn5wFtxk1Js2v52IbRGgJw57DJDg
tq+J51Sb4bYKWHk6YjiR4904vQodYZ05A3wgc24zLCM=
`protect END_PROTECTED
