`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OUAxtMZK72padieL49puhsoVw2jMl00jswGTf4Fpj1XhkivcBGxR/PKZ+cpEV0+p
aOVZTFXUcbZ6jmOocuH2txFXumtiRA1OMN+C1SAcNmOFPmx1xjrdQ42ne+IgEP9o
+d7ftvzug4LS0/OLthQSfqBO6WD3YmwLqk1bZTktYFLE5q4nkFIWQ5pa+G5683eM
ABGEhXNVYNtX4ZYeJoKzF/6P1QbOmUDBhLC8T9bIKXZBXSZIvj7ODB5odExaE6fj
jLtDagTLmm3Anm+U2MPCLpqNOneYu6kN1y5bNzUHXzSFDn6tSV0oVb+wOZuPkpYt
xv4KKt72o5bAlb169UiiNFAGWI4UPk8OvudSZ0T+XEnYcZCQeNmYMHlGnjl+FrAn
Urp+z5Q+Q2iCx7g4SLWg4Q==
`protect END_PROTECTED
