`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mbwQAIret/PFrcwjpX0W4Rty9/NOBsGc6Ld0yqTJYp4Vs3m/QJYRpoUtDJM+d/Qz
ekDFukpwUVCiNLBqdec/8cG9WlqUR54Vcfu2SqXnBrR/mFiay7uz9RyTE+RS19Ns
joZ5VTmnOxi77pUimRuWpMXHQ0eViJjGhu5hNQec5azUYzK0zqpRFlSHTQwep7om
w+8WytKACrWV2KmxEJ1TcH791k/h6FcP+/Nd7eGBJQyR+qHe0IGBZc2tAeuDUxLV
SIJAhxeFmQ2YSdiPjjop2+ozJTyYr1ZP+yJ9IHBq5V8=
`protect END_PROTECTED
