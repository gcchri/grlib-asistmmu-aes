`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FoG+QYZItAHqSIeYS4quHLDl6D0Wlys35oTHkmKIUMc8j9UDKtvvFZ7m5NXnfQy2
rR6JgyYTZh29rhTkpXxgpUk43S5kp1CGSkm5ra147YeqITqD8NyD4q0u8Wtms9IR
b7IGQryC2f02F9+9NEId5sAAG2hQmw/Kbai6Vn9WsRJvBY+b8TmLPHCgqkzEcPvZ
eAx5AB/yLaS5tiDVfHjWQ3c8b4Ggzvb4RT0euFQ25tSEJjJt7QOpkenoCoLSAzMy
q84BUlvkbyW+8pS6bH7m+0G/ZVQ00qNFgxggigdDkbnqcuUOv7z9ZLWemzC47lFX
Bs3bk32/8Crrs1bB+3TJivRUX03OWxiDTZfitJc2GUrJt+1IAlawUGrxwE4MGFKg
tmdoONbGPOJ8Cy9MjOYGk+NaFshrU+da5ADsWkjeMGYzne5WLpGV2Qx2etILqLut
Lpz5PU//ks2dKbexFXx1DJaou2vsCEukFfhWVQheFNgQ9K4pI26zqPqFOM5hio+K
uRTs+jYXkBkjEOVvW6/gxH5OVFivg6JPq2pxhynFe8y9OTLoHKulBggeaSxMtsh6
K0fvleHSr1eFAmpfKJsl4YfMe4lz8Y1KwF2wGgImGibZYy8pf0vgJol9V1axdmzW
/ijv7VzqUUyZi3pzl8o4Vw==
`protect END_PROTECTED
