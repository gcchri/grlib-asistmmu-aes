`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2rzuwh8KC8VjGjrwk9ZCb5PRRWdY+g2zjmAhjbcPJ3k8vomEHfajWotIzqN+M53P
kDW4pZv6MeFOKmp9y0y8VTpOcsUKJXORrSCFB4CKBe+gMVFSoOv34lA31audspBV
SmE8wGiexAPeoCdal99c4pc/IgNL6io07G65iu7rHwpQpz2YNTVj9QdC/N/tgBiw
7hHPtPTU7SYONeVk3+vhP344FAwbfE7pyiq6i1kiPdYJGLi2y6cGRnT0fZPnVK4Q
XQB9C34taYtqRrix7+idOMaZ1gka0WmvsxZD3n/9PgmvR7xbhc5OalJI66TBpZue
8tnKsoT83Oace2Y4Hh5vqjZTb5R+V5OuSh0k55UgWDoeqtvu+oIqZrliFpE2+YY0
SXXK+4/5KDPoKLqig2qh2YUTyU0CmgSBSYZMbKyyzVILUvC8NoqB+wp8Byh1emZG
bLBkyjKPy9FZ0vIFBv3xUg==
`protect END_PROTECTED
