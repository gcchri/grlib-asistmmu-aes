`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JuiA9dBSF2Zw3e3n8VsETgTT2i+wM+3x5XXUdd9TKkrxJu3Shw/4e2UGR4+tvoHj
weCBooDMQm74vyci4pn8Tj98YlFYnE3agY67GFZm/UBKIku0aCf+SVYRKooUTDPH
AXbJ30xfza5GWbih4k9u/T/mawAZ4wRgqO/cuUQYhQFoI8THOrX8B3Yl4grjK/G0
DcRwXPKFp0uoLo8xW0lJRZTpx8rUngYZTP0Hn2tYH7yN6kcexvX3b9gttAsn6xhV
gj/MHT2uc+7wQfA71+ULCs+pPi55zrervjOGp3tbB8A4DHnWNmTn3MhPT+0Q7Z5x
9cRfR3H7hH2UsEfPlZQ6+7DIxHoqOtaF/vslkcJcjHgJNr0XFy5FNqSt2e/5nw1Y
j3lgX3rt3W3MpfW2c7XfbTo4T6/1D3E4TQPRnAoXPPYdUaHpRuGhFWQfh7PuS2SG
T1U4WWjDqEqW8+pZUMI13mTlAPrkf4fj5oq11tu9L/zbqk0b6bo01GqUtxJJKyvD
QewnNNGFAT5uC2ose/tq+H83WaTj7yKXKBkw+ZCeXC19EBI+5IqDWkM/cac83tn9
`protect END_PROTECTED
