`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWOb40RSW/cGRKqwQwyxP15hhP7zNjbSnJlP0++otSxIOaK3tazlan0a9DBM/S8W
36+yh4MpoLwz6VbANLqwxIMTaRh7N9pZZFuEk8smBRObL0U6uBIRfWCcNVWiL81e
00AfxwV05dPlYCJIWALFDT42Yd5EgoaQ48peZE1EY1ctj+J/lDnYOISrdAwLgFAF
ZroZlI7TCTrAM21uF+r1AgftMm9CazJgD93Es+2xmprFAUoOuSwK4k6bGl8C5gvQ
sLicptDX1qvwRrBaGKA+Oj1UVeVgwj8Nuzcb/ozkTky7DYTyCL4+i2cUaLordHMf
nS9BL4P84/XNOpv1+6SsTGI6MojjNmmRfKN7IsIED2AH3ZEYlPhD4fVxP/4UlfEe
OC80j0gDgyoaVSUn2+KhmxeUNvLrwPFyxbBZjb3e3fo=
`protect END_PROTECTED
