`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vIP39Jb7Qghu39SM5cutVVEH0OFc8BpR8VqdukxeTCSxDZxWRlQrDgQU3/Q30AJi
l473Oyte9LmFjEjHglmPzJIflXQm28eNi9Rful2x0rgXwR2+A1bFyMMC6RJidW5n
cvdDvnpGONiEXzus473KSMitJH6sKjAAANFH2j0nyXyLyNeOqGQwbtpqPboqoONt
dyCOjAMo7eAWovnRF+yO39Yoj6bSYFNWBi+nUheP53JgoKTFHEe86OJ/bTDBHypf
dNXLIXaJJ5dXsF2cImt3EYSDUo7Hw7mR14Cbt+0xx//w66Ze646IdBKJMuPq1oTP
0SAbIw+GzOHz7whkLnj1Ni3pe9hicTl/Lm07VMQWwcrW/JnZB/9+RXknyXnnN/vh
tRVMaV6PtpxeZVab25E+iAY68FNiKXKcPZohX3QJHA+0x4IObe1rDHYAwZuJKrux
J9hZCMVe8pOQYAkZg9FRJwY8JX27As8zX0IgHL1M1pZg5qklqRaQLAZxvCtbYjIY
2LMJCvdtfBqRfnEZRWCRKhWKFuR8ifk6kRx7N+ppqYXPynj6qk8KlQc5LNIdrlh1
CuOpM8ZGu2EGAxPEwGhYCg==
`protect END_PROTECTED
