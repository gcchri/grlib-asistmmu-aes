`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3+IbjUPg7pG54SsoiuJ5Orh4cxA18LRbrVyezvCyaZqRU3j13vTjbXj0dmgt1Lsv
MolXqXJS/tAKtnb2FIgdlvEmS3EcHaXYDlnvAW41a2aXIpUoDjL62f7M8V7PUQJ5
z4UZyvrwh6fdTe4UsF1sEhnw7jXpMfoI6lVU6wIp5AO/9cDJl30KmTmLyNwjC5HF
YtyoAj+MI/T7Gb3KCM4jqPo9twJBISC1TRICSr4kKZjkpIXkUarvsdck0HnIBfSj
YiVVfCFTomuqkKgN8RKbOOaQTIebz0BMDxTkNOdvtk2MzEHbZbIQtcNOJBUMEqHy
7U3v6zHQv7ORsDbEaQwBAa8zw5qVNXfIRVj6vRzuo9frBarQj01kuIXTrrtMQ835
4SrKIVm0pYzWm6WZlRuJgg==
`protect END_PROTECTED
