`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZzSKz6TTbIrx+P9xPgl0Qv7G8/mS35Vm8eP3PApKxhTppIx4O7NqlgUqb3IWK8Zt
u68utHmrg8bdU3WBMmWFcMVjnuRizlcBSKF+9BmnIHmGzPyw/7s20snVDEtepaV0
QMr+HgPtDpxjG8YuVu+9Z9jbL2srWRcfDitwoxaW15+qDAOJq/SQu9+RtUXtqUXw
wd6HCbr9IkVT/qwK6g0wgXSwxS3nNEgV5A+AnjqGexG8pD7gmj+pD5AZuKE2AR0T
4XrvbXAhH8pY49w+cn9GTUGFhLAaI27ZWXqcnPmvR4bQTC73EFVy7EVNWJQlpsUD
kY83zXJFfmfhpgR2oGAtgcre3gi486CiQs0HREyyMcIAsr91uSNaiIDQxxa5Vmh3
D5dbW06GkqmqC3QFRhWJPoIcEzv7ajJimtS/L+SeU8y4VX/+3R8P1IAAF0BU/Jp3
GGXtX2S4I2+fEflP3EwwRwGYuj6CO8Es3WXzWbaRA5RVm/8zet23qRLkrZxo0p5G
aIspme298YuCq39yZdFnPamhvaEfXpS5xvyuPVhP7DZ3hAmocZvVAkQIcgWzbdQv
cUFSIZ0GccfZYzvT6PprDFnj3xp5d+iTS+Fq8DRMUs0Mzbt9ckWwW94v9U8WJk62
`protect END_PROTECTED
