`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XHUs8A6dOB8VSscfvrTlLYaIydmFdHdbHe1440zJZFRILvm79YQcHoBQBSudVsYu
+ph4vkMYB4J8VTl/U42HPA6GYPxFq+NUkc5FGSeWgP+Q+pGt2PFjmAZoZAFakWHV
q4S0TK8wxTENVvcahLceyKiV6mkBXohOIZ0AHHFcqkzRUDLSTHlqE1RnwrID6qq4
31YCHU3HWHe6yhvvANRCM799XJ+zXesFhoXqoJJHKEh/l4/7ZhvpUtNHqsqkVNiK
b6VbF0jceskkblSiYErt7eNep9MHAVVuvjvzu48HlsRpy0IU+RM9SYw1HSgeWol2
ic9gdeToqgbxHYMKPer2ZWTtlvjtSbCw5PF45B8/4m8=
`protect END_PROTECTED
