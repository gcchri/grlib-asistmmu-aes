`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xEzCa7dOMMFAQ0UJa/YQbJn+pPTKwhvlMayNtIdW/qUE85Npdv1eKuaAuKeko9Pr
9pwHndWKYl6vBuIBXAv/a0YKlcLeCFd8mCNlucuKGNcZNsaVHKm8cA/2HzR5neyU
Qx9wbungCBxvhH1/KvxGeGXPdRJ5tn/p7Wxd1HPrq7IgbeyPz40S7AtauxkM9QR/
4rTDj/ppNWZ6k1y6aLGw+eaL5dijzltGzc/XZ4IptTumuD3FAKj0niGGyV/JwtjS
VoAjjCI8lfAcMiIrjA2z2bKcg1cXJ6kqtQJ8gK9DXLh6eSi4G1HKzUlffjjDilmU
T3sEg6G7ZwKk649hSQwHpMxgg0a7WG9ejSxCGolxIUVfup5/KsOba8EVr0U4Ovqb
v5YIB+6IHWy1v8sXGY3dKos//8hAYQVojY/NqpI1/pxXRQrZ8NdVlIqNOoNPdo3r
At6QfLRuoa2FRb3TaMT85PTPF8ThTSdyhdgJEU4ZXVHpsAtSc63oLWn7gPbuOaNn
3EtGaBU9saHxt0H+eWLghRv/krGJRAtXLgGnl16iiKdFiCRGAvKZwhRfpF1XPMov
`protect END_PROTECTED
