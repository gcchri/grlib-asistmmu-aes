`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pBaNMZo1K+M1RFQqHscEtmK7GxKlNkl/DINpR8/A5mTmgsg5OonlxWnzRiigSxqp
mbhiChZU1OAp9ORYS3ooZm4vZwU9PEYLr4JZBUnHBjcFcFX5EWi0QCmo+j1wEXgf
OesTweNjYeFOUGa5+quH9tvJpkC3/TqUD0eqPXCxI7YIeLXy6JxIQIXcAxSntWRw
VVCV2dG5HnLrnXhC7/LDlDjdEOhogcaNUSMqHF1ska5QLFqOzk9PnJd39tedUsOP
VOkY/kwNpnRh87JALqHRNqUPwtGD29aqaDcRsNy2er6h6coNHQ8ZMxXlVEZeNIDi
w/OdfeXTxCz5kB6DGiJ//7NCkFRk2LXFR5cTGs1sE4aTMGRCo9BAJpTUQmAHSMnw
D7yP3atACOsq8qSkGaSkgJg8mU1RhLJbNUU6HWcxx6Gn92mjWmQEeEkNRwH3J35G
f/6VPyWA9DzeGIEUIXMHNwErL9Si9zB7A/2X0/FWHqf5/l/BZa0zZvC+1QYjXoH2
5j6NQ99WRqKc9OabWXkkHS3BaYCnixPxS6q6yNlgwHK0x7sSeIvFFdgQeIAxZibj
h/vdQvLfQ5j8DtzJxPrqHv7Sj1Y4wyCwqLdgTVmWCM9muy3RPRxfOu1odgCqb9Do
HBftK+YNIX/ZuFXxdwarNUU+hjGOmYR+s8JPjblabNpf7SIUby4iocKdGhoJkeYO
Y8t5NpX3CVn6b7i8meY6hYsfD7VHDoAZCCkZOh6nD/9xb2ojlUiGayev08GKJcos
nY21Kqha28dGMuX18cPN7NZ0vPrMVDGG1kmRczbSouI/VH9oisC+FpzU6KdMJNmx
ejDEqIig/Psd5UjRlgxYzhrCW9i62O9AWMaGRfwbk2vqUi+bVvcTnaWfqf+afxGp
SBQgasfAudiY0Lz1d0WudQ==
`protect END_PROTECTED
