`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
34yyplcWv6dLssJw1x5ZVjtWog/e7RzYvyUltIgNQUskRPBZOlHsMPgtBhvLQRfE
7r+DG3X8Wh0iRnAX97s8ub3tcYZHHS2Ktxw0Hd7n+sC1BV72wtDoQanOTLp/ZK7/
bDsT5TRrRedI0D3Rv81n2BGU5v/Fl9lnILXcRwCFGQuBfVidCD2m9AUkaOMQsAgC
IxaikRioCuYZh7AI+LRh2+8rYPpL6QxLqolZUw6OpzXm1PPVtHUfR427w6MD8xtr
lbC3TS7kL6+UJMN3KAScWVj9MkuToe1cX96DlDOXGtqfXClFzQP8xB2CBSLQGOlA
YR7J8x+c6yYIoGQ9ILu/2n4xnlT9KIoczeGJExQrcOJon1v3Jmrc+Yid1Cwa8Q7X
LMWL/V+WPhtBlYIftdn+7zao2/zEOH3KMFVusspZYPc=
`protect END_PROTECTED
