`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3Dg+jyslnE39SWHB6RJeOwyWeH5L5q1BkAWwzYU1ZcCI2oL3s4oPY8q3z45reaA
MMnuSUpivFToyaOnEy/agGF411B45x22guu8+FBxWcEW7GQEB5gw/lTkAZOPS5PJ
fpX4F2yz/Sl9iKu/e9wrcxn5W13j0Z/yq4tzNyb7Qf6kkuYaZJkhKMz59ZtAFMBg
FLodP5Ui2WriCeMZkbEltnujrDJe+zZYO74A/rSNUrK71v9N+T4KD8JsiWQn6Paj
ke/3x2rqNx6cCHd2zFDvWiujA4pECF9iSou+l7P0J56GcWTFNt+enL1vCxXcdgVH
fiV3AYkh84jCNF4k7em7McGnCl7CDBL0jsJBnNE50eOe7Z1yBRDlL1jhaO/GmErc
kx2SPCTGNch7iyCefB4G95of8PmAyTr+WDS6Sy/5uRA=
`protect END_PROTECTED
