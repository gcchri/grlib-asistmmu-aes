`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yckpeTjifBWjmqsQrWiwC7T+27fylZrIU0Fp7PHMopWeVCJ1y0DpBij8R0BFxiXm
Cj1gO0eTGSr8/yRavYGWC5XG0hW57YakKiglgpFXFz8qTfWvWK5ih5ARpuH5kGPz
TeVo2vpv1hcz2vm2UFpbep7bBPnHnxj/qHMKb/8tf8YNxEOrvoKyXOLSg7AsVPGM
E0f8OPZb1ArL2jAD4cTrFVuY9Yyb5TIMXV+sNf4TuPhkYGwtMhr/EkjBResdSL32
yIb3Vhj0TiV2jK56xdqDAqo98+NdYCHnkalDyxN+yVh7D5ssISKjzEub8bPIOmVR
3TfkZYqMTlnEGJXF1lJdRjrNwt+UJE3HBRtVTM1esV+iH3TDnSSxzIH8qw5M3vQP
bKBXFzseRKJweAyyKpINaWpWWN/zCZTqFPSDV+jnGtwgBFgkcYxBKkyS+3EUIr34
J5NkPqD1G8GRqDAJMhPzROv4huX+QuLHH9Q9VrXo7Htux25eMa7IyDE02l57Gh0g
N5/2OkXZhxp3yQ6HhWrCgPePmFVyJ+zaWM0FLBX36mx8pfOnM35zrgVFhqEZjrbR
PJ0QojCGqDLqu+d9EFYLU8QB+rjWw36ynXUxnQ6s6JnPXIiTYA8Cjr+15T63vvBr
DIm9sme2LrgVtxKxhxrP74AMAe3+e372quG0t5N05y9SjUWxB+OK8CHLRJyNESYK
tJqzewf7PABeeRcXeea0xK5Uv1iPU4uXhD1eStiEZotVgw+KG8KEC4XbJJOYxDZO
PmbB0/wKRTaI6RBh+tBlCA==
`protect END_PROTECTED
