`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
odDX0MGJgf9booUVoOcyjPtIdPIChAppflN7UD7xv1NrKyHcUJTDWEvgpEMzgBbI
fP+JUNkzRPRmr25ooIH/dBZGE7ukb9sNdqFwqno+BQ3Fwy7z1Cfdu7yLOz4UYkyX
J1fvykjmS7pPyI3qEOMcUxo729euMpSBguYlzTOH6gpvRbawAxGmwYCdKfnPvqxc
ZH6YiF3y1INc1G0IoIFnggYFxrNBjCMoAvaBSlGd1tcqD3+C/L0ExwksOKj6VaBz
rGC07GeBMkVujXNnLkKKSK+Oj7iq+2mDd3UEc2bL/9RfeQVUbfaTYNWP1PxaFXHK
`protect END_PROTECTED
