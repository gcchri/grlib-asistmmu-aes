`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CHWxEPYb0jmf6xeANxIPpTotCwpNOxtCY1IY/ARaP9svGtElDwAcUaUQF0Q71R7V
lgn8Ne5eZDtcwtDJVyVPkvK+0CktvWtcyXQT016aFl3Hg1BT4u279pDhVlg3Zf08
bljdKO4aqZy72tDrJ4k/yjYyKtIjlMDUIGp0wNBsrkOfohpAVKFd1Y3jko8M92Vz
UWRCp/6DEAxjhIXgspFuTzqV7xQu1tDClWnQ0Chi3IjIFIdfHPqqxedQw9nahGKb
cFIFb4BBWbgysMr0D/4N/hjKAKVQpxnFjEylwB3QMlEWQsry+1+H3flBTldrt/J1
tYZiumQFXvgd8oVJImQX9g==
`protect END_PROTECTED
