`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p7wnyDxjEndnobls09rrFcsZEzEM/DekfBEDxzJGVORD/jYTEr5mvehsY6X1CfEL
s5P5EiujbN2VXT6E9/972rLxow0n9eD3ueXMndaLQKGkmAbiOVcyoM4KgHNYhRGh
R9l/8LITrXnstAKTNt/wq+RU4MOjAQEzRAo2gVEvHoEHbnym3KiG4UDFHkNzye0z
ti4lS1FPZ91CNdm73Uh6si1QM1by1qUE/S+PtnCSihrr0754+tZbJbEiab2miY2T
s8vN020OQnWPrbNtzOIs+BbpSPLwzcs24pEg2n3QXYu0LVCUOTFRX8LykMk/rPFm
DDrWnmraIphz1tKxwyKnWOCyk9bTdCAQEYthXBoRZRUE8fVGXCu+5uaBYcmnukOi
l4Y0gkYESJAxwVI9oqWRZKQbGI1ZXRmbAsWpv6RU2g8dJawAOqQyzQ6DLe2n4PI2
PdEhqpWikczVzRxp5p0fXTQld25G0CDZjBAk+MpTcyPTtDBSDyPfd3ANx5GB+aLO
LcpmV9gcO8A8Taz6wXIuetdogXoVo9RSOlguPLibOfoY491oi7DwKkrLdccR2iBH
lpixrf16jiNDPCrd+QEhgXErBJvKxKtvzO4FLZBLrJ/hHyy2n406jFq64PxxGxnf
G9VBXGaLnnPEHOspwnyD9oYnrCaOkFWGzdCmb7jNWcKx5m/xpDlsVAZfKUmgA4Yo
p1DRyZhfe1fRRWcUbtFBORjtFu0K3MnSMM7ReeOJIvpwDvbRG0ZoL4TQPlNv7FJg
8uYGppYoRhTuGnkdewNmwWMGYahVq+oRdVpKluT1X+1lhISLfWQGYS7Dg8NA7mWj
egkeaQyrkXNMhr7YL2C+PlOAr7lq41fGs0k9bZLN+GqBBTSZykdtxlgUD4cQoweK
pBBk1Qvt2kd6bboj640jKaGigLNZ+rTNitL+mwpKws+PDcFz6TtIidpTGurMg+ul
2q+M11I4evIC2fbp+kWJIJZ773o0BgM/DpcGiHf1H+/brx28RvFOWF952qtxeUTw
1JodVWMk4dazURmYGHKD3Hu+gq1tt5s+HgnEbTyNGodPpCx/C2xQT8QFf3DgiRRh
brmGhf1MPZ4LTgH3kcgnAZnXb+IsXpOVAzYoJCP32j9csVyukJnPGx6RuYWLJfFo
Zglx6NRNJDwQFg6sIXOiBZO/ZPZhD+Rbj3iwekexkKjQThHwkG1uy7MR8Ad41HS9
`protect END_PROTECTED
