`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C1ANKCQZnBWUz/wFHueZBxSJg4BkHNd1WeSGwYxY5yw9wMCA9tX9YYRM0I/j/IBo
wVYXivpP05y0xzZsmMW4tu6sE+a8DVGVsE62wnU66PyXNc7njDLwV8txZ0UGggnT
RRUt4oBk5cxkFGboOc+N6PFn+adhWKhDiOZmYiU7VAKBCOLnBmHviDfBBjbg9AEX
UPR5rg3ULJQkWGtI665RD9QM39edY4fInIKRZukG17zCeyTI17zExPhTlIoFGHOO
+hYdRZLT262hb+xSBsZd0AuYYYgDWaO8ea8pSSqcNwJJccqlnJfRlbpjI2oEldmm
2VsSGcAEL6+hNqE/hDv5t2KEBgJTh9roqM+00vMzLxMLZxSs7ODUVlz4gQC3Vdzx
3XTpMq4RPESKtx8ZV4NcLo7zuOdh1x7LJVisUTgjIu2tIWcyEuiCnhucWlscy5zq
`protect END_PROTECTED
