`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ZQ6Q7waMqmSpNrX2fEQTbzwvANN1baTtnO4yFGIDqynv3NCCMZNJczNApJWAiM3
M5xzM3BcFUFeMbEFSur49HwFeFHLXBSDRgO1TOCpPnh5iM3Tstgqd8FfUcloD+ek
hqiOYNs5M/fCuSqXbIukAJQO5I+7W1VSl3H505tbyRZv3AkYdH193Au8AlAUF2+j
aYJBufqAGtUJ75yzd8XEUxAQbBQfAaY8/4HsL9CxDtnSgFsmk6MAvPcpbLBIPoxy
eqL2ivtEKe6uKIpSOXO8rKBRYMYIC5eckOUQryfiuqjutmqERVHK4/nmytE9Uyyv
abtLgDMaUpbFp2Tqdh2s1qGb/vCxHkv9xuSYyhpbtDz0WIg0r9iSWj1oxByuuLpq
nxsdWgrSTqjrPgGBC1lDMO9HLtiCyuIJGQwdDsLoWAYDRc3SlDKhQa2Qg7RDCJRX
VtaayIa1qUn/rkw6polZ3vio2i+TSih+kwJ++1XF9jcvR1N28qHU7HN2Wom3uQx2
T3vP563WJ9XmmYOfTtrPI5C3MFePWSvyuGUSteP5KryBr6quXJ8hPQ2RZy8arQBB
L2SqKAIpRKM0yktWDG0XUezgpa7f6QKdPh8j6gYLCbwN94seOXMbniWztFe7mZxW
OQ8RdAXV4yhxCEVIhn7W/g==
`protect END_PROTECTED
