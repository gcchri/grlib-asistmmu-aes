`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hPQ49AjnCl/pxvOULwPls2wSHTJLHaLS5O/AcydmP7VknMq9x3fs426ctyUK6U8a
2x3X0JDGtEEYRyx45GFwV2UCtpbuVcs3sK4GHsIx6DnKcjy5NRxE1odKjjMtRWIf
30sm+UhCjZfcwPwG58ZFKxM5L5MYq91i6Rwud5LXJoRHWDODNLRJuKtGmJuZlUPv
9qjQeAwTOqEpO7/AM8THBAdGMlZyNIjitxnXNKCQmd8oWx7n4X70gSCTshd4dQyQ
gDZRgW3/OqVtZbr0SF6xA8QY5K3fMCuImpH3emerm4U4HypXebUN3JAh+bt1b2ty
hO59pIwU8fwkbYmGIQkO9blm4tiKTVxHQPa3AmFw8zAzHszyIIWlNMun4WL02aUs
uzo/UpycVawK7+aynnxuM1VqdGCJnPLZXemA6NJYqMEZN42xORUqCqzr9IlGX6tG
1K+eXUIGa3S9mM2NGSdFD+xtie3svVWOrdjhnDjsYtOp9qhjIq6TgC80ZfkMER3e
o9OrlkZG9x1FyYEDiORI27zm0iQ1JzWoGRbSz0yY9UDV1fFAO84rbtbLI3m/bmyB
tgWbYlX6hkbSCm7NbB398Itz1xuDpH6+e4WlpoTiZoUEPjeoz44kzii5cgQVX4wp
F0tL6J9/J7iNnNMbK6STPQ==
`protect END_PROTECTED
