`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K14k0A0FmHYg/bAt8v3Nk3Xk3OOajP8SH+DdcOQPrsfeEiFBbM8AksxzRKJIxefW
Os77jZrrqm3qFDncn0DtnFteWJ9aOzH2zaRghBGMNmAPToTgQx92nvEPobcY9FFP
6Rmk1TQyeZKU+fV2FRZ9LffYxsKrG+J0eKN6rENJKNV0dsAqW5LV22DxWa5JV0mH
HNiuHHiGxisjBH8OV5GZxQuQDHFwX2ZfG0dfQ/9231IJ/T2Gp9OwfuWHBUqVQYrK
Sma86GWw4EoeKdgYyiRDOZ2udct98MJCpifrwkQqKUaAxZOsPrNy2tIoFdWMuDyT
eeD6c9gvWzFFJNX3ndbDYQrBtIIrX8U6fX4jBPVcmdF15wGKmJmY0JNr371wGJ2k
PTIzIbX512r4LDT5DnZFbN52CkB9ASPEHnMrEZ20xCfpWBqjjJeTrJA0zIenQbtB
qAO0aXE9G2WuoxO4yK+AhtRYw/qkclrc7tn+6NxP6CLwkwlbvm2+fy3y/KAxn6fg
NVF6YnAjvjCW6W3u0Ft+lWpF150F10HBmTaYyY43yMSsCFH8I2PSWD0Fo3zSnsCP
+5VO7RBoG6Kk2TIzlftnbsGZem3kQ02avgvRxk5DXEdt43N/IX3Lo9L0MrXsxh5D
9q1xR2o6BxN3xrKLog+Nl59gUl573HTsJmfmaSZLtNBGJGFoch6K6dhdXc4NZqWI
XDYT6oVZ+65MRCqDcA4nzKfk5EISuurf9JRddKJXM9hRNxUbyV8w/zYd4x1oJyBT
AEIzwzeMfQWuwnUo5INpRijkuG52mnQFDvRtImGk8f6mC86SlFqo8/WTDAKHZALY
T33Wd6BXrkadGZpoC4OAqvNhH+32Xisd9gGAhIAVGih7BvhqXfSQ09J4+Rc81d7b
KDpgdVX1/GO8I1Y8AktGl0eKve6ynRoBGYT5XdUi+b2xRbOwGtWgRyNELIThhnpj
mhwPJD7wvcB4aVtgUAvw0BU4gjBTfdH5qJARxmEFZgSNed6Zjx4ZnFbc4YlPbPSR
94P9kgD3rZzqmDwLe2IW3Q98xYe/yFCte+6Kz/tYiSaoK5yLqdkKxtBBvsiU5Lnv
tc5MjHnZpLttR8HruevukZgcKKhNlqZNzq4KTLhVgbOE+C7dPpY8dUyCJgFMZTOJ
DGPGkmHMey14+SbfMVrSZFVz4A4wQD8Ozp5XfENyL3jwZzmi60LAHu+hv+GEbdv6
00raI8DeOPnxi6ECGIYUSuy+6/YZSly2FWnKYCYH3eh82uxsv7T5sZmAd4Bb+rFf
Xp9p9NAj47mzSxA0ZIY3oKpA33AvQrCiLJXjlo1nuv4qQS6CciWu5AwQzp2y9uiN
uo10A4/ZG5b7RNRlpcziKZoOOsMCKYlLOjhTWJ5QaAgmB4h0+iAsy8PKOLliVQsb
gHeWVeZJvHKiTr9rfOIprq1HYH9zsSsoAoRlqJ7SziNcnWDO63hIJhiWbcdJjHZF
hy3x8CFt2sPTKsG8+sFHA9ewF/gzB6qs9QsEVDOTIKUBlsaaFcXRWj/P5JGdssmP
3UEU34ZgY7lsM5pIfpG6u57TI6ZwYt67tEzECd/dXps+kA+Rgkh1f6OEcmm3C+0L
8P86rDVZvp8AKVeiCJrf/ob1QKLRigl63cKddPYJHtOgCm/Iyvf2G9+HkudzIznd
3j93xELWh5zXC/ti4ffSGIt/zf9AMzPZpJb5KROmceo8ZGzPRm/C83KPOgr95o7U
+p3GOsA3qaZ4lxoscCGwRbGZfHkvbLc0zUCpZjX5O+q64U8GBoz1Qg2LoOGP4Rnj
cbkYi82sTrlLOLJ01wmGwoIP2JuiJT51LznEA0LdRZOReXA8VVQ6Pz5pBcP4zuIu
FULSURyt6X5PMmXaT44Ftr2kc5fs1j3tLnTh/hvFYCeg4IFvXyUqOy7V0lxEQCVU
/D2h3tarHGTvvhLo7r3DeQbs1E2FnKxv2XKi8odE7ds4xYXuzqtfAClOdSPBCjjc
nztJbpSCVrdAV8X28eU4mQ0zF+IABpKgHrn1HPZ/iluxnGl9Livvspcqj5WI+WRu
3epZoovzgg7fAGT/sm4rHQj/PPjN2Q6iObV2KKynhVCA4YE84FvPBLSSDEvLvoT/
xunqEL6ULPakIBROmloA6aZ0QcJb7tVz15FkWhSoUlpV+jej4Vdes8rW6Bo4f8b+
7O9hS018QfSiC/aE7FpziTP22q6Q0aQhR9PunTANUQ4=
`protect END_PROTECTED
