`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5DVWr9HzWgHma1QuhuhKSabyqYc1BvC3YDT/NyCl+YsqfZtpqQYWuKq5zKh1qExU
tv1UFBLa2oDjxABSE4PYbQYH6vYM3Gwv2r3xLsf5Z4I+RUh+yoKE4cyYUPLXLFG1
HIS65wDqZmqK+wMOSOZKb37OOQ8VUDrCDvxG0VhPkR6qP8UCod1Jv1IbFR7xlsTG
tE0IkXZ5XFNPD5ogZVXD+wXdyLO6xalhQ/IxlUtzmYrirQjcZ5QUF15U7BoUulFq
Un+OHfsOcRtnOrv+bwU5MXoFSVtqgg/yV7rNuuAepbuoVSZwmZkrkOGh+UOlpcQi
AbEyo5SHvrEU+/vZuRyKjPwmjvQo9/swt/3d3/jCNRQ=
`protect END_PROTECTED
