`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OzwaXVfO9iCWib+QfuGFj+eB8KdRT6i9NlXPojMRMPoJ1hsMulbxxrqoh5SLv5ck
hGIanv7IrT49YPyXZ3KH2tGCoHY5Ip3YTEbthT1ucSEAi3PWcobt72A+Dojab2bB
lOdA3itl1H2t/qLnHbhh8a8rcZ+COKYuiZ0nvDynmgN+tG8+DDO5LJgRsAsEWQ6l
IbpIf5zh86/qcg9Yrp1HLaJ1MEIfr4z649Q42XYKrm900zRH8fVt1/4boRz9ztMs
dM+p6FodSxaT867Bc935phfVRQspV7K5miyYjghbDs0CAJHyKCu5XUNBsywj4eU+
XkRjwOxfhfu8VeV3yhT+OconRE2Fm0LTtHrplmTHcKC0ecjxyQ3ddnnJVxQ3tSJW
DW3nMEE3mlo20cl0NzuaPr8hiUXHZ3MHp9a9JWTOAzR1G9O4QEX2CccSi3UDGHIX
7PoSAvBKjFgGAgq5mnX4U5crCZ++EVntp81CiEv847lJqvnAXeRrwSPHjLtytRnk
gr4RP2TaezpJQRGbRCju6qv8chhuz4O6hShADEfeSJX13/FLg8SQZ2YLLW872+lU
6M+Hb5uxeFci4InlwVaTM3erGxg9DlzbsbyCmzYeay88DGZCYXrRjl8qH65I54i/
5gnttIAGSnl+rnCne3gT5mxd1arnDPuikBNCfeaT6vA7sy0WM1U5RTpatbwTTTZi
Dr+it0iMLu3Qy9aoNQ40rcWma3FBA+BBic/UEjgLMBzn0pnVr6h68WUWo9+3C/y4
gplmpme8lzPzg5zMbVYhhrOs19vsmy8Zm3het5u6xEiZ2gLagCFpdH+9ODghRmoL
ryV93ung//DPy+BA9GPn37zDR0t1LUyZfI28PcplUs+dS8HOkN3C+LbxakLqUcLN
ZOXb86tlCEGFqXUhdiecHX72TH58cjsqeJaBHuurY8HLIyG02HzvO/u5YRK6IFmj
ya2+8lYW1DYWuGfAgl9SFv43Ux7zEVv92Z3zhtA6kQ2b3JCePutzO5i9JtdUOxuy
Js2+Wc0sKK9C7d42Dr8FJMswViirAdLPbpUxM0UrVCVUeGkqOgxq4G665k6gKFRc
DL6DIQkI807iJXVJNw/na4ocNnhe2ks76zxMgUS7YyDzhZFv88KWPW7tqOomdNQn
TcWzTBf9KPLPa8NByxXueRfdMNKUGn28/pzKCAjUgaA04jd/gCNIS0VZ/pejcAPt
L8tBXDwtMNT678h6M+u2v52SQm9WrC2Ziu8OyFS+kOo=
`protect END_PROTECTED
