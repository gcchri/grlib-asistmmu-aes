`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GC3EOXyyvfFHWewcxcQ6uFhtCd1e8UlnbHv8nJ1HivPpRbowJXwltmohmDt8UW18
0V5kLyi9ma5d9NFrM9XZJo1x+K9o7U82CKUP70h+pFPnS4WkV4Go9ZkGAdcYSZqq
Eme7DAmclr7s5S+qNfcbrw48RqcvZwHD5+YSuaXiky4lbhEX+cAuj3X8sm/uzv94
nvG80Ih4LtlP4fB+7ZFB07CD+dGxv2VD5ACUINgs1rBww+5pM2+0759IgSGkH5JN
Y7fNleEAx6QNHgHmpJi5baL8GayqLhIgPj0BW+pOWCgg97kvoeSn31bhwtQ/dcRq
itYhxTqL+6spifFxwTyoVLitufaLWh8ZkNJSNqlBd3WmCofAs5BtpMs8J3y8cQrS
PQS9NdIge9/VdyUo/3cMKdMSN/6b2qjj+vLPxGvXZLwaJvxEDw3ChLTNjYPOBjil
XDW8i+QQjtdPX5pjyYhqIUKSt9FvAndiXpKzY+Oit00=
`protect END_PROTECTED
