`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N2fI5FnauhHVhDt+IZAEITzO8d+t6XNnEUsnlPMrhNoUZCuCw3Gq9GWlZnapCBST
hTFJXZYW6RNaVfHKFb1JRWO6yRKYN3x6SbWOZ9RbINTsHTtsC3ww984SgOLdfMjz
aUJwBhyW3GXQpCw32gAJieWk5dfnBltIr2lZtRZ//zbX+0scYFVfJwE9UTKWUgaH
dG3K1HzxxS09wo9TauFoVlbk6+ihpSAfjjAj8Zq5DFkdX1zwmiyFDmpLK9ItA2I4
g5LVll9+di+k7OY/wipCwwU0hfOz6DcNne0hW9nJYNsuh0MiiuQTExTToKCgLfK7
xRvkwo8u4mfBLqMZ0c1+jw6TUG9tpkFmw2lQ7QrqiV0BaSRYNZpxAS4R9/i2KctR
lmbnIxFRBjqGp7b7hBEPZW6p2j+LE0H8t70tb6rDIXyjszPActJTC51sJZqnGw+3
GEkF+t3zF3z8+dgnG3Wp5qD9Lbmv086BJHPdv45cv5rZ4Oufm5s1GbCDfEBfl7BF
`protect END_PROTECTED
