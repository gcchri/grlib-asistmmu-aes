`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fueIiv5qEkb9pKaTZc0mwKN0DfwXWfVnLFVSAB/RXuI5ypGiTU08xbotP+QKjgWw
HWDeOZ78Pz6QISeeVG4Ap0tUKvlLyUH41MQhTvnWtlnHCu/QPCdLgDGGQYO3L7fD
jrvzAa8PUHCBfHu5mqn8LTQLSYeEdPjMEQwZiWVN0qbS+LnDlGdT9VeEish0Ydie
LnBNfqMHnK8eqJ05VA8NyYY1EscAaMgopHJp4gAN/sc83N9pGkfzZN0c9waTeM7D
hQHvPM0ccSmo9BnYSq2x4Sq6hepYaWTfl4dNioF+22CYNlwsjONSql08JO3F6ZIx
RT2CYfCuVJGKBG0Xf1K8bBL1yWhfsm9S8canqvRarWYZbp+fB4pxy0/8SUSa0Wld
j50q+vq9Ah7PXZkS11/TiQvXyv/Ax67HsJsjvxQ+uj+5EuBtzpIlHn7nZDbPbMGN
Qw43svNGQXVhD9cFFwQsuVmMLCxUT5JEFQRfmDv+5m51KMTyXp1+UwhDO59egF7N
OPmZIBTCLEFs8M2fNOaCsrkV00HIJY755K93EDf5Rf65/+yRCJ/f1UOxIQNsxfou
2LosowTCDf/nrlN1zhfisjWDMb7I8v9IjwZrxKx8dm5sA+4g1y9ojWH6uaLYmb0a
AdBX0+WvxfRabfmtGJsJD/eSMotgGOcBQo0IiPVd17n273nEKwVZ0xUZf/UlAqW6
nPUoMwnS80FIUHlU9q6nxddqAIpq0PkrzTUSFisJEvBHqXxPj8/gRVsiEp0LqjbD
YQ8gPA5Ij9wIgzrglv+GzzZDY4hNVMNCda5TDRgmzpQKRgRpxQiez2XZVqACRHRl
YP56xotV3ccrglA8J08BLY2e8kE/tLUZPMFMddZcfKwS9nsfUq9mlijDGJ1rBq3t
hdX2Llo5V7nQhXgyw361QyAzABs4bdmW2eKQ1dunPWLga/xui4xKhjtxtPvvEBBa
`protect END_PROTECTED
