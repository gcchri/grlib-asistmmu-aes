`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SezRK7lsdVgGNVjF0To6nveXGRX7Plg/fNEMQtthyVjwapjNMRqhAnwFWecSGA24
1rFrv+gcYAyEWWZcrsD0i93F183cyVuGRa4AMO7UCwZDRIA2GQBQ4HBERVSQeD1t
YxIhLoKchv3sRIDnSKfr3Yd7oli/4nLiYM1763H+GnodhmLO2GQGDEB9TW7RpMGi
swzBDiHz9zPcsP928EZKcixnYdpm9/OSpolBtaviYp+RKIRUjcI0PthU6coR7pqb
hVM6/pcK4UUElSH+Bx0tioSXo0kAmdtGZZXQOVZ/dRzUWHiBPkq/uacn/3JhtwUy
/z2wkvk1o4StUA9OllyTBxoSjoUdmA+R4gF48LZlTlgfZk13JbWFFbBYLil/OvBd
WmRISdQk7N3sVWwhMrkM+u4TOFKtXCUnygX3X0DlULNk55IuuF9ok4asXGEAXSmY
68NlFsgvMRynBjYSocB6uFEhODh+75z6gyXyo+szwoi5b0MuTbCi2yGqWOUcaPVS
tNncvXSUcCNEg9uxBebuvHVD9oOSvcBWN3ApvTwku9gfcY3zI60qX5Ikhml7qKws
LWbvAV1mYmQuNfTkG2lIOgbc+20d/5JNaLP5Npf8vEuThuHH1H4AEJ0FG4qZknoj
mreVUINgghIVQYghcfQplCCzAzlcR6TrO1q0ZTfJ0Wt4l1cJ4cIPF1/3oEtttWvE
PoqZJOqp2BgT5P3KTQ12T6txb4g7R8I9y5SOACjMC/qybYf9hrXBWMw/xcbkL1Rg
ipwCaUyEmvT8gM6d13m1mXtLZxTdwFoAc5OQdZ9zcOP3jIOEZFwdsNop5mr3BBmW
08yWFkeMsLKIiMoUN19b2twJjnvGY5bhTT3V3gdeO3PxasGj2CWH7qZBEDDWb7Rk
NwEy/8tMCKgQIzUUOvG/pd8WPGtuMLaxLAxeyILnBxB/bbb2MPKEHhF7pFA4LyP5
K02grbynVqi/nHuUmK4D3pDcJe3vHY5fAQT67D1yw8HryzMsPCyTdSaH/g4WQOsy
cph4vQQzNPDlxughKIffRkZRMTEA6sHHlhsM6rjpf9vF9UexrHleBn3jhBbAz6Bf
RT56uAFVC/5Q2oMx8bThtft3nZQvA4e6WN6ZmdbfwhTIk4lVR6QhG3fByXn9wj1a
llPcQxK+UycmbNsQEVO2/4PFUzt97z0kbMR6ah8w7IEUx5hicuWM+GviLrKdpRmX
g3mdGehtjYatbq5hjHdrDpiST/W//BJsmvIexabFU881SyiQcIbQGu16V9AInDCj
C2RW60GKpp6SVWOhx/3n9h5nruRpg3SBtZq/1DF03VUAURd+3jvvfpjoYfYLe8AD
Hw+lGEWpt9xn8o0I+BIv5jPQG7VyArDMiyLF/1BhDavnEQrLFVX+c1U+Of7aiWYS
I5bLcrvIzkxJForyTw3GRg8jUwe3k5feLvA8gmXsBaGKjYm6psAoXw06JIWEki3h
d/ARw70o1eGC7IhoEUDgv8hJUfFDvufgC9nhS8WJg63pCWLyWIdW3ZxHKXleVlNS
UruqCJIc+Osrgiq8HbKa6vMwU65jkei14LN1kCdDnABGbUM3sMns7Qu3SGZ8Vare
zCqRLd8KjKRpEwAzL8aFbzlX6Af3O6C9bwzQqhdoV7Q=
`protect END_PROTECTED
