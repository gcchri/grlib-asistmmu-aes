`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2po7PMBC7VDRsHTq4wcEH85XX2uGMQWCNhc07lPZOcgAfH/PvS55d1uEbjNCUZWQ
ca5sae5lPf1/nn3s7HLXfhqzrLCPj78HqwnGf8LuhTNvt2sbkBOfcRys7zYSXnYp
0HDR4a5JNF89Qp3JY3spAi8siMGmxC9y79vJ/GUbPCOzvN8TgcWigoWHnul/XSVt
Acyws1lb6o4NdyoNMeXHzw3Rr9lRACt7vBvQnQcZNvmcXU88Ou7GdPFeAqfMvbxO
pkYk8DDmMJTB14nzuCHnZyJ5jNgfiQO3Rt1sXGT/yHVuKmPDNViYgfHi8EDlCc5X
v9gARjW75tHokD+MYOyrtxGbWn3oWq2Yc5TYnKxxi0rlsQJVQ/HYf7+Miq6/HMvM
`protect END_PROTECTED
