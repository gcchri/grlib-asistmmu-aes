`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XAl18SjqeGAjaCf/2nfdsqwRTjISgdBhQ/UjhUPE/zaW69JsCnpWzGpWdx+f1YG7
H1Vf6A0z5d1f0pjO2oSzFSe9CtgGmIOdfWytFFTmhm0O8MP3J14NIgx9D4nlkKAn
k2+5QuBapfV53T+g1V3qQWCbXRYg4NnS3cfdqvQNI3557EddA2r3D5uozXRVesvs
X3bq9agbcJTivHJSPekDcP8QPEn8jIzUnNFN5f+ATNdy32/dbYr28GEZ8o77GvgF
4G7rajrii4GUBcea7YO0pWmpI709AQ5GMjjTMjuvjJ+hqhS3aS1l9gL8WAdJ2Gqw
42dW17556itr0LootsV+OVgkdaX4Ob8eiKiAQaVoRSU=
`protect END_PROTECTED
