`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fArSD1hgVpQqSOEyDbK0S+V9RVwqo1akrwgskxYnYHJa9q005caZxqhJuZSBHLIz
sIQA5sD1PnHH8aGdJks3dBUrdlYzERxtbxD+ewIMyUU5y9HjhY8I/4U1jcmvmbNh
Ug2YKi07SIpzSoqGfCUrXeGdvBEc2RDf7TH45ewwBt57xxyX1KkdTk7hiFuCCHm0
SmGSr7IqIBHz40oBCf3gyryGEbyTCaEp3W2/BpoJLKLtqBjvH65tvBudn5vdY39Y
CbpjhhhbgeRCuJc9+Ba7fTZKTQfdV5HLQLA4DQhZu6eXFjQDYKShRKPz700rV1Al
NOJB6zOBuJyTtp4mqWxJpDXzhzNXG0shCOCQCK/ZrBqIViovqbn5SQva+Gf3Pa9Q
SozKcVK694wcC/tP5CL0JwswobOH5yCQT7e5v+ZwNLHYPpdfSTIo38iBLJKp5jZs
wb1o0rkSGEsq4QsxxR5DT3q+WdqeXGLYCJkM85GN0ww=
`protect END_PROTECTED
