`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U/b/LJlRVC89Sl7h2w2VqsHzqcPXUteD9ueUnBP++WZWLPpS+MSaalqK3ll4l3sZ
9qIvl5J78uhr7h17YzDH2EQksx/BEMAhNAa72jAn9q3TD9ksfuFJgTfw2c2U8KPa
rm1N4SDCyUvgvs6cnosUKyZ+61LDLaoqS/xsWBMvusOEaJKzMUeRvLOGLefPZQFb
pr8+fyXxKmd4ffym05mU+YKT2RTayZZRJJVY/cDQo9X5YhiAEQ8NgXa+DZU2naBG
7K7jkaAfOJiYX/hwOXA4d2PYOH3ZdEvhRTbLstPqcCDOnZiIV40XwL8MOKfvW09Z
SwxI8R5xtYVTwcnTN6/AEiGg/8qXS7OvNIlj31KTbI32+TvNg+5WRFaLRjxM+0OJ
cCzni60NnnuEgXfMcr3sGVMyiBDcGngyC+VK8JQ6NxARrqAeCCLo/M+gxs3vIp+p
EMBUbrc0KIsGIZEKwlGjgam63jZQSokS8J4s0N4n/gQbkxfkqoU6PLYWMVgd7bhI
aV1hnhMYSZRc66WAT/CQRjiwJtVkpLF9fUs90UX0ImeKhx8XyPbQ9zvCY+I7t10M
H7Vyegc9WMq/iY/BGGvF+Bn0nZB4R/IK2YJbqw7g4ZqSpiBcn7eaL2wJmL3IxmQ1
hTbysI/sNRlGok4tIgvSrpmeNE6xlVtCmfRem12HvOv9zds+AP+yS3yV3ADrkQzL
gmkjaInEW5NUbRqTIwwKfVErN92vJecF9Gri6rRDjzY8vc4LTlV7tNFROFQcU7Vc
0a0Wo3YxniAw5JAZlpUSfXUhFL7nPkagWpfek2+ntkdEI3x23yj3CH+RiIc6dRBS
XxIVvnRjWlojTkfp8gX/EVU3aWg5GtYtjHHLHGxfnBjNjyPPkKlm/PqnambFKvnD
u3b5Oeawk/JAsi3e4TmDvhaRiEQDRf48bx1aPvAW0xEQZqM8ahp1zx3p5T0I0CXZ
`protect END_PROTECTED
