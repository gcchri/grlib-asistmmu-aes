`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
swbBLDbossy9XPRMc6KoBMcv3ikKY3AMITs1dzy0E9hNP0z2NvizjZfv47CQPF7t
gbBjAgmsoPG2okW6s6q+wXCSEX0d7U6qouYzRUayLbu9XIR/I15XPuPzNRFuDL7K
KdZoypRIQtmbQoUjZ/bkboydOlJEyWh5ZTvbNFC0iIZgkk3A9XX2SSL0dy/i5ae1
+mhAu5CjB8DbOElRAtxO16F8kNxontxACJ65zKkv8rT3afFSMOQR4TTJMv+CcLzL
jG/56vKGS3CPJ48/7Bj5YWGI6VOJ1EFU/lq7o9K34+N6zkMUIEu3jDzANXQmicWe
ISAKU7i5BATiBAopl76ejFlJV8jXcfL+iyhyCkKc8Yo=
`protect END_PROTECTED
