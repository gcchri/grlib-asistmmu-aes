`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pqHwjkbafs9j5IJPxAcRsj3tfJ6qfvWbGDAMW58b/jwo5PjSYgeuYDvemqx5Z32q
IVK9anQmO7Dxu5xfsrj4/okQsI83M9qoxaq45Ufk01KpL2MwC7+piDIT6PnCoh3q
tgW8RdqfJwt/Uz9fCcg15qkm0OxCqEumAFyRt1VkxHSdlCxzcxjoa5evRh/olk1m
YLuirMOarPXMJxsAVYCrk39rXXn7DYAzMzn1gyzsPQ0KFNBaKaybY+L4uJwOusb0
OxI6eS/TLDzoEbnbBBtEIiGFw3JuSlW//Ti0q80QWCUT5VJUXS9fvy0nLDVCvyxv
lkA8LKl3eY/4jQjh6uBN6mBX6m3kv2DyFnmLGgoZuM6/A2G81wsCNsDSqMXLi/02
YkaCas12GsvOV6yGQUHSfkdY0jLjQ2cyFBCqAN654NjbVujFe8myAqlfka5WthD+
+C//66H4zjBXtevPxeiX1n3SvDNuzgX2T/H/qAivbFKQXirzjSea6wyeIpr/yATe
D+6gi9f2wrpoEB2zQMmUXoST6eK1s0ohayA82v0x1Xdbgf5dR342MXjjTryMmAkk
hiYrVdX/Oh3eWs1v9UT5rte8iWhBblM9rL0V6+lI9kINACvrN780RXp4dtdjzg8M
400Vq106+zv5xMIBSRQO4IQLkEbHXrQjO/ZYWhP6HCYtPpW683mDnehKvjsy2dHP
hg1FdokXbNP68O0ivilXS4ahp63nBnVSZbxpFPnTXhizx/UIqyU2WC/tzPfwXUZ/
Zu2IAiMtxlQXhapA/ndmCQ2s7i0BE3nz8cTnn7UTCwPac3VyTuQVh0ukFxFoKbUl
ftIsroLbZXWvbQABCzvaZvv3ov+OxF7EGVt4WdeI7Bst2+DQtvLPgAGhOhxWGg8/
Jju41LZEZmTnVMi1LOdvDg==
`protect END_PROTECTED
