`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lFXKA3oSBAXsxNQYub4nGHeU247Vv8ymR6MuVNxGGGk9BVmL7IP6Yw9/KeORL6lE
rBJX8iLUBLBY37xGeYxO+w0DYNybPuRoijsjxr1TZTpawMqpYxqmNBgj1pburGxg
E1p5KqX4X+M6dlrhx4iJcHN/o9JkmouM7iQ05lmvwSiS87JOnHxDJw3a5TiEMWyj
IzmRYy55vxid/Updqk3eg/mtt+rWVj4t/KQgFsC+nCE/OGntmrWs77C5V46iiATh
EI+M4Qs4OOzST96A6JeFe46YkKi6Ddk7OmF3hNZQ7+94K3MGoY1QDDDgT93q1LtX
AODpes9LPp6+qeW14DEnTr3vv6eodLyu3fqvGQUA3Gfwa5gqdWAvxblVbt9nevO0
BwAkDemy/KPphRn8V/dHB1Kv4N5OxX4YAxa3D6pagzZZzJI3CBacRvWynP8YgNty
73+xMOofyH2DDCpCyjE1SdSZ2VgeZvuxeRscbrQ6CbZuFzX49IBqI0VpImjY3uKR
QuYliP4r7dQ0hrSzlTXum23hnuddJSzWFeOdUngR1DDdMXZmDwsXoQISDAHG4VEO
oRq73B2RZnaEUq6zCRn3ZLnsQlM1RhFyjAPiQLjzsd5xeIhqe2XY2s9Wg8fzuyjk
c4pVD57iijnW6+27JXnPXHGj8pW2iuZGiq/S80WjPRQsltxeZdAgfPTf/34q+IBU
Fqgj+oaJ+p/6B6RTqUeC5jRU81hrAG1hzJCF+h2JcqMS70wua6NobNd+6X0xYhOK
wNYb3Mh4u6IChAyT/BPahq3VB4Ebl6cj4TMWY2mElU2szcQ3aaqL7FLzwWueCNKm
mRKQJ4Vf2ftd/0V6rulAANYWhIaanlhdKuA5ioFh0JJEjkjdf7nUPK2nbij/3lnz
W1tRsz1WPSpZGfP8BCas2KKRtaXofVqmE7j4Z0KY7Kggfu10g6XpeqW+pIXhhtCs
9iB6aORGuIJFWjqBBiJRDQ1HVJ2RDnI8KQNzx4cbYuqj2dBssOw34/PS3jak81aD
mXILwjcJNqnhN0997J6eomKbX8Zc26qxsypR/n9vv1T5KjntgH7FNH5eHCvmezSb
2C/CPQTjeHEm2SQ+5cs3wtWLzJdgq+lHANs95KNEha38NUp/LNMutQVxRMLxkJoT
duTj6vSFQ5zytKQA1tpZ/5A3pA/kqsi8oIs0HhhDTBYx3URc5pmKqX+xkd62i8Hs
jdRyHxc0J8ZGLCBUtOoUy/lGbof8Nf/3/lBdK2TgvvfqTFJSbVL6nLtP2EkLenYI
COEIk2Vk7iyL3fuQBwkY5Br0DonYr1sXLPrc5L3GyhHVnyL4EB3tdPMBjb6bA04P
/548b9QZYEw62vYXEdrj6tGBx8fyaYqodYG1257p7K6XO/BH1EHacz3jiHJ9RgmJ
+YJ/lUeLtSLSF7PiEAXp5NcqcBstHwzJLnUu40OrwvRIzK153Nm2fRkYOTGiSWSH
XJG7s9VVgKGn8eNdNAcFxcFR4+H/cvPyOYI0qAyzWwXnCby0qKcmCbyB/xTqYueE
+92j9Bbsg63ie+dCIBQGIJONoN4MqKcNlSfZoMdacKS0QBF+Iu36jKJT1omIpPKJ
XJXPiCHP9VrYGSAoTZ+5hrWs4iBx1iPBPr9HzwyVTBQtJylkhQ8hv413WwAS50Do
RUgxeIDZdVck5U7fxBa4FVnpQF7l7f+zBQJzlrQn2nWsApkWyvhE4F7bfNAP+WYr
rB2AUA5dZvHIlEJj9hOHa61H78hSY8rM+So7RyHuwpEtyrMUGvomSAd4Qae0g68A
B5IZVr8nSSgxuAZyNV2xmlLoZAMrAuttkTWK4WjMZ8e77Rg6MAfa6FwHujda5QXj
XHYdg9XUvisjR62z3FGz7KetW20LQmHyiU39AzCGWDklkMIoWZ4Wq1pQiPYNazGi
g8gWU4qEDQF6h7xb0xxoQ5gHRGouMQOYkpA4tXAs9m+TUKknk7BnkJQ9PMPtoWc9
b0THPQ9rDFg82bvJJvXZ9gMH3dOPD4rcc2sr8VxsWTr/imp7lnobm42FU6xTwuEI
05Hktw1fonuNXHcVebjbPoCSwNYdvg3YLs7u5x37b0TfdEbtLeQGtr+1dpV/blU1
FEycU73b2WlaTWo1+PGl/1jgkr0ZyGtEBfF64XGdtJ4y3lhLPwAUpCjxogTInz1F
0LFNK1ZWMh8DGCAbL88W8y+r0Cu398YwFb4Qy6dk9m6KwrrZWIkboD+lq1vyyBjb
2xNNuN/L/0tRJ9VJ8vErdCT097Iw/PsSpmWIDoSqB+Dzavo+zq1tdKJIYX6uxPac
it0fa19Tn7B/EWrNfQEkR4wbXHSEPFA36Bvxvx3SKc7dL2r77WFRmSvCF1/eSSvv
1foKH+9WyPE7QhrnJjZlTCJH5oER+/RDVhT5VCGAq68C5RcpQ2sXgLBqDq4THAqL
hJRleFPdxRW8+svwR19VuMV0h3x8OOrW+2B/y0wJfY7x/xCsEHpfSlpyL4LTXVzo
xZoGITo/wTIM6+CklPqQA9NO1SCEE+36vKUAsREencfgt39VFfQgDqJAztmcsrmG
l8iKxigW67UgRLEM/F2QQYw+UkzslJwPdmxT7ijgIeFFczvjxWd/VpDtKsOIPb3I
0Q68CB71P50Tq1x2ptryTwbf7H+rVG3ub5nGz6zhkIs47g6BAoq2xKkUFHw6uAQw
GW+imzKUBuzRcC6DVqWJxKecZmQeSCQdvhMRylhAXeLv4KOduDU51Q0QyHkpUWXX
X8Z/D6Y220VnvkEHWCIUgvaI0FOOJY6YmFa3la5g9/7x6yIe1AyGWgL9jfu1WN0v
DEeT+43gm3MnVhJDMXVngEyJc/1Pu3UQi2AFYwlaiNEA5Y3biMyxjC+7ky+AvRjN
yyoVY2N0OxsuZkucYPRwpSZNPEt4xbEO6/BO6f+n48H4KmDw5fj9VNSN7bnLQVyS
pSjkzEKa0xAqjhIE2C8eNUlt36zJR3QZg3SC/4CF+DYIYwAV+rohnaQh3va33UWG
GM4okHL7miYXn0iT+SoIHIOJteRp8zZf2G/go0IK8atmIpTVc4fBeRIDcQPDj+gU
YS+6ILfQ1bS85SLzvETcfZT5+au0Ju5DrLgPnkbcFnDR7qyS/c9ktKrznpYiowQs
DRoN59h6+LgttRu+4oVIy/RCiFkRZ/XBdnFyNOvhTPgc/gMlDwF8a0OdLkXL/kc/
Q+hJEYjBrdmKWOureK0dDWQ6QuoeHuXZtfG/nkEeWhTydVpenE0SDZi6kCas5UGR
lqcxXDdZyPXu2ceAOEQG5GCU4sF3L96djDFsO4xrV4fQSYkAd35k/chakxO1/1Gp
Gbqyz6tS8Ta7Dn5ESjeXWW8TjHJPGbSRY8TVLjhzwWjZ8bnVUBirz5skTJLRTdQb
oyz6CO5nXYSV4NhK88mRNyiHANZk7jB0Po/afAZ5oZjNqPabf7PBKvBUQ0BJ9F0z
R7/d6uozQip4izJ0nWl1KHkeN09dlOfQW4FGjDmCsxtVGFX6Alq8qtZBgYy5TKvO
E2pkLLrbTRcqoosEKXTcJ1JbDvQHpCIVTAwvRyZ8b17usFh3d8YQCKvlLExKAZEx
111LNN/TR3rFwyoLT8yAnKxo8xafx+y5IIvR1b3+YZsxZNi6jnZW6uVA8SzY7d9V
vS8j7t2NDD2CXFPGnA+O2fzQK5oCMsO4eFBNf35KVXapb71iB5ZmdI/X22sVJPSk
R/BShV9yIMs9l1PFd8ctkzQtrybD92J8btGQvad2mAvrfJX6l3upxKmI+VC9+Oa+
ZFANU+WKX3MKyXttVAM8YXWY01AhthvgPanQbx0+QhG+P3pnKrIe9ZDradQ5wLnS
T5jJTfsBIVA4sMJSGdMbP4MjBjh28Y4Gwn9dwUrr/u0VDDcdh0ul3lIUQQMx97Kl
zmyUJKKrqDfwSsQHevd7YCD+jA9vVI91hFE9feY3Hry1hdlzKucphZzyuap6mv0U
IZdKl/n9B9TrEfd3qAhqdMObpcHoloMgc2aT8cn7+tJPJELRMg59bYLwV6SdqHKZ
E/xI6+91YfFu8zq+CVdt3i533CNvqH9LQiW1PprtViwejO7RbCj+66092MXXoTP9
wMnKHXRYP9WSeryWpZoudKT1FggnWrPbfToRXylJJGJx+DolWA+ILmsXiHNNroH4
wp5BaTH5FKStEJbj2yLM1VdFaROtKWGeD18dpEl4iEilcPGORbL3TM2TNK92smgG
/+hWOpoZ5RUI9YcLuaE5XZXVY1tU+KAj7DKiefb/h/g5aeaqF6HXiZnUnsdlEGig
35efd+I2V3DidOq7Oxdw6NvEF78Jq7yfL4MfAsEvyd0frU//CDvMMhhUqGBPqZBE
q5bSqrFfreMQ75td1qB4gd9FWngdE5ND1/LudvCDq6ed6vnkZDfHX8DwEq/lNUmQ
RChuEQ7F/c1w/2zL9lXNoPa56E7xMNnJJ14XM+UGiTaszrkuxTOt0VG6657IEvBF
uTqmIjt17gOwipJXt4A20MFPYI7yeRaC6bNeddsBBLELnb+vPiwAcKvb35sIqw05
WO6G8OXZYsWIhxBti8pRIDD7yEROwco4rY/OCEd7gWdenRoWvA53kkxNsIjVQiLO
u0aXFZqSfPEN9IX2+zbNwDla4DR+YR0vJckafJHC+hgs2szP1D+LXy/18cF5E5O4
o/he9u5q3bVygxfR9Vx5G27ToAePcv9UjTR5XNKwPMZ54W6pqGEq+3KnN61c/rke
5XlAQ5mX/46A4QINlVVoup8BByluP+beQA5tUEyOmx4zhMigwRcr3+148s4xzrw7
jidIbgk/2oi+Yt/X0Q16x52oht2cSkPuD+IXHLyn91WozccgPElr1yO0rnsIFx4K
KHhXaCho3yf5oKML9nlmi2pdeQE2fkn/u9a64S4t8bP3LsyqWdVkQlUpXh4nx72u
LKe3BTEmLsGb0o//r1qr18DwPBqRhiKi4FkPbtkSSMYL2qX71e3FCkZrVZqot4H9
U+Dom+6ilLPBMR4J8S4GBye8tyOzjFB6X5XyMVaDpwVvk6+YOJmzpZr6wrIbI7Uh
hp72jKyHB37nkwuQi1mM26B9Z4NSpYiXgOWiSmtE2wBkms3KWf7/A2CaATGOaK6k
Bv/hIdkxidlPlQdb1khmhk+Y80wb8WEe1OTNqO+md7rWWvYCdUEpEPo/Ok1ahVhQ
0gUOQ0+6LC47OX5mSUHXrDXtNOjG6DF9mG68EkB8G9LKo8GVLpZEoLUYPbc+29kT
B+z3XyhbkpxLq/z5BP26o9QUpuJFVpD1scjd56akO8zUkhjMqKreTuJA7wbTTqKK
g5rX8v0vLwhCUSImicS+Frhee5ZUHuRRBY+1flxC/W2JExTSyMv4uFD3jOINy9uo
tsaEIPeutP0sWlZgigpkpsOwE1iBj45bAI18o5neFyG2YplwETXpnDAIRHHcMMOL
SVNR1JU42N8yc4NrkQbqhTD8l5vTfnL41Ph8HA+xsnroIE3R7D7yGQ4ErPPjQysY
j2n6UaXGsKGmzWmI8vvZQoOlqvGuAzpSmclt4jRcU/2Bvfo8J63mi+UN6ASxe+2K
23DJxc7pnGe202ka/yPpbHXG2RmW3H5IeG+KsPXzpNFTDhaRckNibN0K2/ea1WMg
lM7VxsUDSnL5AOA/2E+ZPTjwovsyX1xVVURWrkvtOT+sedQgPUhJqePgUXA5Gart
eGIx2ZfAsX+DncjGk9uvyAYH/0i/b7z8HtM9/rfkL3MdYhFMs+AQadtHvwwHph86
Q9oL61ggefBBKSzxzFjRNawCAh90423Ugv1+EfPiSgrJ6HGbYllqpH+DkMySsWdp
37kGD4xPHehQ6Nfj/JBZOOabY+zQW4ZBHHulQ0YpgRppKWHsnpqrL2NIsYic3B/V
JQDYx+sOwkGqelwFL2VUwoo5IZLM82RNvo/TL1DI0ZWc3xSbIh+haV2NA7iwQx2r
oeIYD/y382nGADYGAv6cK1rfA86TXgHvpm452rAyABFAou/OamvcdM+anr+2PRVm
//+8MNti8dH4fpDX68Su66jYaNZsiVuMKnefYU16xLDTom6gcQSErX7HML2fP6px
nBfqJcQIsz4CPHnKcFGE4D6MebU0nRqTclyLpCnzQDVT2tu6zenz7vLtNt12+L+J
wTWXYbrrHk56l4QwE7qp0y7BxgfqI7iNouKgJhndIluHVo3CamU681bwuiJ32+vG
l4n1jaHgzmupO6BrkF2ikgPqwa3XZpvJeCTe09xlQV6lTHKiP5lqqdgf4tPYuZZO
CxpuJ/LxE2nw/SI48MwgMcLokRFTEQ41tvkr1wuFQHZOeUjTGIaDvVSk6PF78YBx
av3sikpK2CjfLSPUY3DW1TQq6XQlfCWkPE04eGr63w2UafzA6tuTvt8Ho02r16k4
LUNuuB4PgwabS+1wo619On1zSPGm41ZTOef19aL/asL3D9mFVPQpTkMOHgpKiZd1
lVXMPADy8sZ0NOJcPujJA2cd1GBERAPzcao4lN2QqCt5EItp2kjkH+ccKv0juf1O
10n+LatXlqFK3OdHFEtHSlgmHzQPTIxTO/01vz7TaEicj7fWz9+QsByc8OERd5ia
QpbvGYfUnctVHP0Yuk+UNGx+YgBQsWAJlX5wIUecaPKxG/J1CgNV6NFI9tXvXmpg
qdRIZXc8bTbR5O/l+osTs44yrLN1JyGue+0Ok0LqBwtJqo8Fqj600PHrQygDFQ82
R9HpjrQYmvPFLXW+Yzef6z8jsXfkrkO+NOwHv6vS6TUMDUgOz+YDBgrTV98JtqG/
3Cx2Iu3HVp9oCgH3gqPxC/dg1J1IJjedopXj1If+uMmhtUK316nsjAJhcVkHkO3I
MOqSrYkYZMUCFCzeMlZDrWOH2LLd0yUuhXNnsWGr4QjhlssOy7noVA59qMyAo9fn
GRtIEqA7XBODbIqwLb0Xjt9Pnu5ZAHC7KBtNPg7bMOUFUKTJgQrByVgcsU5h4EeP
LeylpL1Z/6II0WGGYlbkl9o+UHLlQL4v4C6ww7b1kpXFJkJDJR3zos7CjZ0SxK4r
X5myWCmRDPQue2f51ZtN3kZaZsv5zYixm/s+KL1AS5egDzWKxg6SxsXb8IxIoCKx
uoOxHHPyuUQbRynSfiRPPzBGKASfD6avEIYugGUSn5GOOtauX35uoxDMiyIH3Y6h
3hrj//45xZENRFOGg0pO2w0odI5olba8drV3BG/trWSo+g7C1+Obrlaled04J5ky
LqKBUVI7u/yUeLjFWD3UTqlX9o2237MoHbF5LEL3OIoYu7ADBDW2iJwnSCzxWLRq
L7qH86Bh5d8BqArNlmOMxYFWkLvc1EDwIdVFHeaUv9hs4vcwbipDaofu+1N962+8
NInUrpS5HnxKS0UFItPCB5NnsAv/yrpHeZEf21QpqJSR3jnTqmdsm/a6yC79b2hU
na0FVZHvFxkkiBzt9krOevM48J4bkPfWX1Z+ndYeOhBRcTl8w4Yi8o/3erqmq+LR
3jC9OeTTXv+X0NJ6MNwS0GWA9VOtlg5zRvnFZLFfRLIZAP8pS13YZ0OexNEi9VWI
BDhUjnrH0Gung9hUijmSb87LiYOL4mx9//a5xwSxqoqlofvbAOUzpO/7atP3D5Co
q915NxXPZXecO68u8ZgwjWf1xjuTUI+LEdV9dx/12z4YfV5qmRBhwsiWKPyPTNXi
l0shrxDJRQkzeYdXad7O4G/APjFe2NP67mASIbYJqi2TRBOo8qp7aqTjtPfiZJMR
4SLhdxk8xML75FKChWS0GieOF90zXTSEKaqoJDppplEjMqM3WNKfPKSk4HSBHyp1
zYkgceMwsKqvHwwPi1ycLGzRP1+ZrRvHgU+PS6gzDhr7eZrscyS/6bfz8MXGzNBA
wxtKDbMt7PcQOwXEwelI4yMHgwbv0jBO5k2qhxO/lvw0TNy891GELU+BkHnueIvs
EUkux1KppOJrZvhC54MNXk5sLrx378AhWUqrtRB45upa7d1Cz997I6Oo4n+7qdOF
kjuiahnuffPBlEGv5P/DbEJPQBOIHHOyVMCfMZ04+zbIY9438xjYdGQ+bOxtwP7+
Z53OjS2KrlXcvB54KWzMoniqk90tmjvk+1/D4KmUPlqgb64zr/bXslU2I2C1twJx
+5iihO3HKlMXJwdG8amFhHe2s3tvakVlbuC5dCj81vZOFpD0FOmyJpxJuu1477I3
ZxtqTS+lZRYRu8ZbjkDeSX0y1ouilksDQjrMFG52Z7oKLsUIfgzaGSsgfSaro55D
n6N8HtJZNy2fj9x9iYDYVX85a4J5y1onH/YN2gyom3j0ZD0ulsE4EBjRGWEsbDbj
m2Oz0U5YZvdX455Ak6jNMrl2azK2LWQLGC1n7MYSsKqjpNXbVrvumNBIjPKHOxfw
BiIOMUWTCXtk5efV3ZYlxTGcIlrN3TMD+L73GI6bDRECl9I6NgzXMikZLcqASNEy
6X9cUJy17kAEwifMqjshsZrIUjvTFHCC/Ed8ywWkrbctL6eK/OG0L8nV09IZvX3T
mHbFgufku4cxwmDu1l3njHBUTz360cSSjb/MrefUG+p5pRaQH2rAQZldaYyN1rI6
4psh5LFSZvtXJRyYeDz1wjsFQyuY1TAJW3VEvV1P8Hf5PdoQKQ7qx+9fy3pvic3q
yx+XJIvNWqWEGU/SqSXZUokIbivh+rC8Ax1F5cxg4KA5Ixc2tJmdl+ndt7dNIwm9
O8hyJIDeYziBIiKffET+GUYZu1qUpPkoN5AQrMOnzcKlleH77mE/Mg9R3XiBweSk
5GoXkLQF+jucBuMI/LCfQt8OSZj8P+l7S/1f7RlzUXAapBpfOgBBkfBUHMBnGJiU
1L04fglaMm4U6IcBb1vSaA8B9bpob7ZDmwYb3hFXTYkGVQuO1uI4LuWZVT4GZREI
kTJ+LNTjlpHRwhwCDTj+Jammjcn1PLCopakbQfzAm0LH9n+SKe2KLeRZo6ZInOFE
Ep2j1IQ9V0H1IYQGPt6J+SkBxKZlG1hDumzBIVDTLBSBKm+InvkMwdkGwnv15uIP
sMjpw7KUfk8Pebw2EIWaaD+TrGAVmdF5ts9W8z1/FBlG8AytGipY2af+ZlXjn7bm
8b1a14z9KAtxMX3wZ+tk5YVEC0vmfegi0svHSOmZtT/tU6CBjJfFyrr6ZevHbJMs
TLRvdgq4sDyhU+V78sLJ9Px3p8O8B2QobJ9VXpC2GnY5osrcbb/3nRUZdW+wtFaW
51dvQHGajzKzfnAnA/XPOZC0zcwNTTHKBD3QKdcOTGDSbr7WESI01V/7ip24MdtW
OlpyiXKEGrRcmSatYeBn5DuhklHfQiec5jkbGHcqvY5bthMaKh6pXg8l3bu5Og9Y
POttllufFg3PRtg/uEq3v5Nz30g2uHLuPWSFeaSr2JNpvNqy87W1nWDfX1SbJLcK
BZiQgz0QSoTJUl45S0D2ZcimW9FgUb1MiZJlMdCebWCRHszvuQ+3a56qfZv1kioU
Zp+WqHmGh7tl7uXCIDmob1s2553ilODDRrMfucDQtQRzQYZFXdbEUK9LIy5oZSnI
R3zEu42Pd7NM0oQTHGitcED2M3aY1Fq1su/BVc/8FTbIs5cp/YwuNHr69AC2Fh3c
W1uCDSlQb5DzzQ+zPlPQSkKn6RycdfwtUn3m00FEjJ3x0mumwHjmtL/MlRwl62Qg
csfPNLIVjU34rmRHMdPbF0N8tEn9VzPI4Y64LjfAoMxMw5r4xUQka6/+nAFyqUPm
beKtPKWpz8XddhyuOgKMPdbHfBRvM1a/g4U0DoxxE3IyGZpzfmeAAccSVz2vJsvw
w3TcIAhpiT1cKPDTsK5JChqT+K4626lx+/dvLIUtiRA5+5SlbKiXNhD5mOE8KiEe
YV5WHAdlISwdMtuei9XF0iNvLsnC6yq/jorGBOoWe21qtpmCQkL+DmbBn2eIFGZk
R+oH3AhtWWH+T+j5qS9Bt0chPeiBP3ADC7HmoV0vM/UHvzQitT/SeVqEnkjl+KLW
pTqcLsWnvgn/2sqkvduUX1pl+f5GIpYyWe0Lq/KAf3+tauL6nvhhIyOCtQnnw/aT
jy8IZ8oa4ShUubDeHMV8bYKgD5SKgSCav2OrllmSeiwfCSNKnQDJnJCCW7dh5BRj
9v5VtjI71+Q74QgLx68qRDDp5DIHxdoac0jWq6u7vXv9vsQTBQpX0e/L88vfxNVJ
wdo2jMvkXtSM3DMKxbHl48nmXMzaLulu8rP24eFxhcQ6rlYyoondUh5jAbZZfGq6
vVH+ziTw52X+Wv+B+8h4JAJJGGCb9OWOw9TuT1pQ0vtUrCVlw3iCeEtb9d5Ns0u9
seUKAk6rXL4k7HjCGzRVUuUsWEqrKZIgFLVTQOduMY9uKQBjTfmImi7OlSNnigru
+jitUfdbLtmHzSIV+ZtVVJ/FMcjMndKxMWoos+ZkDoiBYxULG0o9kyDiF6m9fDhQ
bPeTLQsFx3T5p96aj3+g0eR7kSAV0IWXJbk3jQVi2lMqbVIvOnJtc3levkVBFP3v
dCKMggylYt4bSbQruD2pavdhwVW9cAaKvmb9aZ43AS1IzBuvp18ztr+pZOOhuXM+
x48JgSWtYThBBjjJ6/7C4C7+iRi0d/V9JdD5cImZMZMEOOoDGjlS/10Ms2SLR2XI
qO4m8hyxs2t9L5HaA9XmNrkL57wxMjKLi+rOD9lzZhEgBZ2khCbLokGRQ4CGnqwy
ZYIgpfo96SDQHmbqNSqrNkWrUMhsUY1WRS5FOqpQ6pKoUPhqYhBQjxRj3prgly+S
gTpoi1hlTujKvE73hsYh3hdLRkEnuGka/RbC4IZoV4B8gsnv2kxtmzygWgZpxPq0
fPBT02on89A6ziMVFisLbJvlcmAA8tVsaWUoKR2vaROnLu3VY0Ypt67S2GFL2pZR
Xh0b2p+l5B1bLh07KMrjOlDeXiwfvEJVKsfz2hMCaLr/hgDDaXfOFcPb7lvHR5lI
WiaEz2TtskKPqmm0y5bRZ5rKgGYeM5RK/QPJ9tsI0LQp24mtEGza63DUEIfizcnW
rgOXRbSwJu8QmtG+B2utPdog7defnTH64Z6+JUL5KykmNujFCe0tuN6VJ/vwdJC7
T9tivZxzijsscfAIXuyc6BQ1ltLMGsnAsabuQNTiXPNxpKy8BXoed85RN58TFdOh
b6d6hJ/k2zfYu70QDkJEiRVZ7/AnQC0fhUwvjbuc3vH36dTxnaav3KWUlwVChCzC
fXLVlbBcANhzqRcHn4xbupKrIbZHEcKJQjAS4Nw3FaU8H7xJLE3uZz4ScoOQ7pFO
slXFZLBq0Ncrsu8WOe35g/S8+zN/1bv3H9gXcYwy/p4oBoT4muQQeYDjz4wO0bDV
Lna8iBIhNpBVBXqj/IPDv7KKnf9aqLtSYEJAqlDMyYKMMjsVUNqQ3/wKBUgh3Ref
6XDRJD6kAG65W8uEl/rZ/pyJ5GkggiNjzF3lutr0SDCUD2mJG6YK3KTmllxcMrap
Z/OcP60uGcT944NQEDM5KkzzRJQE+neIMvHdttcDDJv9zzCAJv32swtsYVYrmz7Z
7ptDkDvKEau4rMPr8JS+axqZ/nIkc9gs1nzhZM7okeeTPr9TNV8d8I1651m1wcH2
csgewB1mQtpurjXp60kmxCaP+lsoRLGjNUepWkE26XLuargWWe29yBm9oJge0ZjU
NZ0c+/8gFRPSyVS+yFmZGLJuBk22qxGtr6/sdeWsv0YR/zd3QlaXfoY2p2Q221gU
w4poMwgHvVwYgLX8Y3Z1Aoa+/4PbcbIQCYUydqS8I4LXL+D9z/Oi0VwzrMwlBzHm
GUjebk7aTrICseeRSoH1F51dNueCCqMhYWylVm0ebGoevEOvRJTT26dVEbYwmLUj
ed81rVYmGq2P7x0kB3OY+XNm8es3OkCqvI36QJLc0gtDWVVYHRM5cI4wq/jq50If
sZBcrUyieAZcByn4k7XXbsYgzgvTDUBZd8DY8CxTfCmVPP97KoGhVvjm+LBkIjbG
MCs4/jcqfAGDiefbqCKDoIlqkPTvofyfRiw7KZC1RFX+RSUFIZNLtuctcbf7mq4l
lJBm23e/iM/Ggs0hDg11d4gNxxqdmHywTlYVZ9xeJMdLdbODNhIUdnPb00xqFFAR
AgmEf6VKxJPgyiRfe41XL5p+VEFIhJ11bnl8eY4e87P0cjnBBINXy0o5PpyC8kSD
pUOzNMuqxFV94XRFodG2HNDJZPIukKw+V19tg3+ydOXxTMOhh71SdXouxOH9yi+Q
H1UMaH8jba5qP6tglt90MV1/20+9tTLB1r1tRVZHVqRoZlj/QslYbIvzQw5itnhA
mPpfK29wQk1/KsnwecFndYdt0tCfWvze9c/kx15mNtNo2p1WAidCJyGRRER4gEfU
7z/jFcmV+W+EsDDtsl8FzqYXPCUfRbsVAyZF4UePPwCDc6TgEMKpkCT+AUQleWk3
Lelp5opRgoFC0TSIzIHWGfGA7GIBFD0ElU/T13nvKsJzdF36WSByb+pI477z5XWA
BS+G7CUIOV/hTkp5Tn7tp91pszVmiTVvruX+WvOcrGrwbk8BM+yVCOTX7UIHiZ2/
6cJS9gbTRps45/NBnSNW/GhT45U5f2J4OUAD66G8qyQMuH77/hWHOXj2oCqEBaVG
mQR6cB39aJgH7sqvKg7Wauxx8H90owAtUiujf65oAtnClW+2y/EcDJNkvAMnjvpk
bnbPatD4RP2VVXVFFf32wMfE6jM7mVU8Zr5zZU4+73Inq3F6YlAjW3IafMBmJS7V
+mQdXsEUvRWW7/QxhXLr46OEnQx3qLlGH9nzASpXkgPNYP1kmkVKSYak4F8E74mH
wrdWOOGgxYcHVZsPnJYU5YJUyNjfvHHRSHe7JztwF5fCWMAsB4ohT+pT5yzpmgQX
YMSE9RYaExe5Wsw2Kk5yTFT/lfrj7nXfj5SmcCVbGbHxAPrLZxfquo8qL5+taOeE
AqamK2vUWEuPQPPNs0yEqCHhZNn7DycGzdeLrd+g4gy8/UaPZCdVMCfaclGBlI01
W25D4fKeeO/dpbDCF8s/k1BgsGJjMwMCSe/bzsDUhXIXuMQ6vzirFHqmfzvhdyPm
hNtzCLiKFPy4vFdLJo3h4b8r7msGhHzxdcZjeKVR0OTZmw/YPm0rLmXTtvvLTUsb
KLFFTfAFzd/7Y3o0UwKSt+eos9YTgj+XjCfD0S5RNzoJ6to69BWF8Vij//SdQ0IQ
0Bk5BdUW5/S+05OCqHRT6d9IuZz+Hwaj4/iuNjuwKtudEva7b/Yg/btP2sguVWo/
6sDLLMEINqzZWCcwTU3h2JU57SJ7slg+Me4N4OC2lYYKAYYGFyUpLaSspsjLkcKA
C/My644CVMaNnc/3ELf1RqBU9TdbljQn07z9zgk3WeRQNc8J3BmEPI+FjPFAsnMB
Ifu8T4+bhF9/WOaKAm3YdYQLWLxIt1fUg8SqIdMyjak0dP2GrE6VW+oBjGShoswW
P8wESg1/ZKOpjqlha+avuJMwlEs2zqv1TwC2hsw7JiQhkbgLG1d6M+rnC9/Rrw1F
q0qCV8ujNwqvRHjd6L7CflqftYuxrn8Cm6kgo1b408+YKVonIuz2TsTq2hFkCS5b
IbyilpCDc4dhAca6+rn9VMiAyRqW3ER/ZXuvHYmNPn5k6Ghn3gKgKl0Io0fgweo6
V0fon4XPgxouRYEXweRKgTrpQ2OZH2/ceUawPzNvY9XrmyI4jMNttQ1AoeLI3tTn
nnqhvrlYrk3eZygrMryR0LyFMH8IRPl66Q8kzUGmsXRbe8yKKymnT6ickFRvC19p
cvJvjZrV7vYaRV82x3WMshYvx+hex/FN9v/nvyJUqICapdD4qRdI6YUJlr0w1Axb
GlChH7tBoYTCsdEHjp6Rd52tFdVFcScktw4pWn5nAatQ6os8TbwDxDhjAFrHrClH
RPww0wlxJps3woTOhD2116H5PnjmJMYM1AHHctX3kyvmzUmb/yaGeWSzBKKTpRc2
9wz19x3av1kjAGu1+BZngKSJ3A/Pj5Of2vNWR47Rigt88qcMuMNJUVhYUV1DPVJw
DpGeIWVVyq+Fx7ZTl5LIf37aIXL4wBOof8K3Z7TdnlpNM+kOMRe0I3vOw/vC/4oa
+ngpClfnrSCs93fHkO+afeq+N8BYhG/wF+q53k3t6IYW5WrJRuEakM+2F5xFwGKq
uctIX5NtBJDd22JJmweDPnrSLjlcx8JzfSvl//TAfeR5ZiisdITpe9JrkC+mMHnT
/6xwkO8R4gIj3OXqQVoSWDM8UhPqbYqrEfdC+AchzNm6BgldU5DE72mvQpJZ2ZzQ
yJAPmC8FjCwGmibdCsc7kmos5rLC6a3Piely4aMuMVjOuoPnsirBf7EzWYyZOG1U
uVw4jccC24//keRUMVLMUI0EybhK7PVza5iZTf7Nl8jQTMacfjAuWw+FRfiFzVVm
Yl3EF8DK4nlsFjliCKS1JaIOPEtsNyTWILOvw2nPIZDFakPpn1f33m/SN/ox/SYo
Cqj759HcF3O2AKCKETF6ATvyUnG3Xz1S6+LK0HDyvyaG8LejRU5bJrKY6DUaqYGI
RWyrn9P5ECIrVULONXVqN6pzKWcKn0bpNBUcwO5IS5PDn/FTHoJI8Dx1ejpd/PII
Rh10mthIUdfWHizFTB8h7C7w1CWVa5fDc8m6hIn2ZktLMuYUVINFYo2R5rXce025
z2pPFDD2H8wXLXX3pFriOgZj6zblpRmNhI9ScDYSOIJemudz+XOEecVH9SQydM8s
gmCKzQpUSCtvcsV2Vo4R1W0/g2Eu9pwsHyJ/nic4lYXtcrdR4IDAxVI8QqXIuK0k
nJR5J6Fa2xmXrCrGWtuT1ZmdecxlXw186HLs4ZymMiCiyIG40IAk29BPu5LHx3wk
KbKh41Y7kGptmhcuXgX2emwOQxfd3ql7ZTTfaWflG2XzyBGBxOa2swA8uZAn/27h
+OK8CdiUkcmr6JZ4N0q6fQpSVeZKwazDU4f9Z946dCTj77Ko+wjGkl77+XKEEHeT
GqkLR9jaySsqtmbhDv/P05zpTeqLW3orVHDaYnOhw0Un3zwuX0lGYk3SV7HNuRAo
LF/zP02YmJlQxzm8TKVIfg5hbk+9sCY/hAO6q9yYRhiEvp3jJOUqfCsjXsNy5JTT
sMxSnIg5zpyzF69o0i+v+Efxgv/PFPdkoMN3/kIlo6awqfhEFpk1lxu+gcSX5vgG
PNGCfuYbZRQiqQaqjwrPeAnyuie+oWAI6abGzIldIxVc1m6l3RM3lpZ6kaIZlk5f
G+c2AdRs9OZeFMccNAkw6fUCq7jU1o2xS6KWwsKcRV6gs1OWsvEfEZWBPaOf5K1J
7DvRXjAWQQaxH9S9uSURpLpquCYN32OLPZG62gep5Y8cj5hSlcWCj7rYxkEBaFvf
9YK2f5xFBHycUqHIr81QSPsAq05jOcApYHKzozAfY6H9uv8dLBQLLbLEzRZt+OZW
+OpmoTLoaiWsBlzWCxUohc0PDej46Mo6Z8Te7tL0TQv68to3I5qHoeC+paR0XgFH
Gz+6EveQtIqhkKZIpWPPsyZPUlX1bgO8bwhpDdShlr7XGVKoLfOcWHF1B2b1Up/b
Fl6kf5JWMLtDG7NRAfCTEuYYL8IpJc6vb4T/hTVPgjeY5graIOtz61W+P0TW0f+F
iH6Uu5aB/82jytKkXVX6eK0QTISSRKDW2ed/1fERg39B98oz/WOfIXJZ/FwnxLdU
qTL5yd2ndvh31gJq4lCrhREr7rwtMbHuCAbhaILL4WMDpz3n+z4wv+rqp30nOOSY
k9BsPHuJ8X9Hw9WewD43kfIZjlkRmcuH/zdzpqo73bfZCejvqHyzCPAakYwCc6gv
LWDITrq0T8NznlUsvD79EeJAEy2LnbmmbCpGbYUMZWWJ8zDnZcYg69Ub5PQ6c1Zg
2zpjY33BdYr3hwyopd5Aphta/Rs79RmpB6Tub7YFJcC21CN/GHuahvJ8FPmDVTGm
QNAj3O12306stWObgVcEtA==
`protect END_PROTECTED
