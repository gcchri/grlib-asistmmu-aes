`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
33ffodtTGEewArKRWakthd0CLMo5nquCscbmjriZj+aIN5qbVUPI4CzyIulbtFNE
aXmdIqB8AnWN1fUZho16Sxcc9OfgPG2oE6Y9njXqUIXtIHTdLvqDXWS+8tzwYtGr
N4zWFDe3fhpu1OZg3zELe2oUQkWohtTabhKtUtY8c6uE8LKgxkYHFrcEc/jlMn6V
gYIDjE2pi+DMCAc5p4wqWGc5Cu1kCM2Edj/tEHD+ZVwrqo6iWHfjokkACi3ozfwQ
JcQfSIQCzFJ74WbnlmiJBqzH2FPGpvXKeqL1mbP3GDj25Bo/25VF4jwXg6TFXhUR
y0XH3q9Go3D4e7lYy4xUYDHQa6XPBNzMWKcUOdyxlyuB9yjdWn3Yl2+7qmz2Mggw
QeFdyYT78eKGJ0X5fuiqTBxM6q6uZhrl8RHDhCXe+onkU5bhyA7uE9UBrlkLX3ml
EcLodHez0L/50vGfe446UVlWEfbQItC8qBRNK8YiQkyy/FZgSKPI/NM5pZTjibuS
`protect END_PROTECTED
