`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQArr3oKkgZJgTtJT5lL+h7UeShQdVITQtX77+oRTEpBIO6dMgNPh+Q1fk6TnMWH
bTn7NtfUUP9InqjND6MmVzIxHF2UPbkyXodV7DmtZWeq7trQF240chEJ9TyA4Eaj
5pW915OBScmP8ONBooCECdzeHK3zatOr9qEilYn+aCRHAoshMUkBMQGsO2KaWwfQ
bAfK/fBJ+iaw9Xyxqnv7NBbj09JwDhAd9V/NwTONPizU++HqXbEXTY8rRUHUWvzd
6y9sq07UAaqAmou7dsTyC4FMN+pSbGoGoePCOW9ooVSz848X02pJReXalvbrTJ/o
ta5Xy/Nz52m2pc6NDfds/56pCNEDyq7VQgY2U2CiMNwNbd3cSJKG+ArQ6nrlwO1C
MgRxlQYcpp/mGNQP2u+exg==
`protect END_PROTECTED
