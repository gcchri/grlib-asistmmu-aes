`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GRZsJqsx94YXy9cr/KGcl+wXqnddewr22WsV902wA/IkDyfcA9PrlYt8QQBC57WU
upKsDvS3Jan/Yh5Ow65eBrrU6bJvJxj+3htPh7YZV0n/bEAM9PdvPvXk977SF8sS
Fs1nm/p3dTyYe2H2JOivaZM3BzSwr+B1+b9pYq32Gii/UeTghwBycoXcgIN1N6r7
yWK6xP/Mu3C88sWYTNqtverMVzthWnCA7bM/V/LWnrRZtkw/TUJlzK4sVbgAeMn7
SvZSmggo4HuwGmIb78Eoc9yLN0rtu0vXZ+mP1nzb++6rqX8YPzVX30j7758DYtLr
KkzZkZXVuJtq5YJsiJ2ozD2zGCnjAtA9rqIIQW0myIpYRCzbbwzCJpg5pDi0by4s
fhENKJKJyUqMOa4jArHzIuTuzbKfn1YkkX7RFbgO2ymvOc+GOf/af34sl8iqcTxY
+EKKyjw/Utj8jWjiltUjr8ePAJpCnpCC+7iv40Sf63I1QK+ybVdI+S/G5RkdPQGg
jkthnhik/jfrUU4082dWy9e7VrpWPyRnfmLYcE9X/5nWWSXNSDEVvMHm2prwbBLk
6mJttwJxXVIm4IFkMQlP+xx/qQnimLxbQNc258VyGRF0K52s6FcxoqvYgfS0qIAE
68ANw0RkEPpGhQNtLjy8xdDNxijfjh3WSmV1GWJKgW8=
`protect END_PROTECTED
