`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jyuN6rfqET7RxYo2fE+Q1l7L+LcQLxZiJvZdVBgZTAEB6kuZyjN9Chm2brGvxvpl
K/rXVJayN1vZLx2qm91UgXMU/s4DCrQcshjE2noYK+Ubd8j+w5ge4GKzPrGPs6Tw
DqL05PvI+BXrtWHr43ko2bDz4D/QadLZchIfj9Pfw2vwabu0pkPq6rS5V0iUrD14
XrRz2Ti64ARRj+bNZ90xX2flgNL/IfUqwphEo3XbShK7KdhjYJKRHZcBxF+OI7XR
gdhiXJ/e4eQ649RUJDS6iTFAXrQySVgDFPHk7A7bjYoFvIP9yl+h3+44GlfQLM32
AdEJNjLHkV5z4b66se+KOHAJ36N6NeUePvGYQAFApsE0o16hMKsBBzJNihRftJFh
3S7MRJwhjMBJVgOGT3CuqnKkkS4FpBu4ZnXlbBZfvwZMlzrYwtY1d74Qmz0NnTDH
2V8fxBAjIltqRR96oDxAsyS082NphZYvj+3h5god0cg=
`protect END_PROTECTED
