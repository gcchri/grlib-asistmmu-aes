`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
waSzp5duREYmOp+NlpMI6g+ZQq9zrnWhkPCJc62pXiHSnUNf5vjfOx3JKKGnKh60
V6i0TM+mm3+WQN0YUp+Lh0sRL46Ko55u3bGrx7Qp6CqSAUS0MYLK05FS19Z6A5RQ
hP32Feuv7Xf2h1DP2TIxR1ifI1hulat/cqfMXErHJ4pjwtovJm0910DZvSQ73Mmu
9S/T/NIIlhSnulZXT03phW/wt9LUePKKveZFEGMex7PODlJRl98W+kyGDYlmOyfY
ZNpwSzdIPRvWv3Wnwvymv/AUTvHU73aBxH1Mbr1cTxVWadGy4gJa7BFqJ1ODDxUa
D6gVLySHfl7H0+8MS1e2YJWjwODhEDwPXH49bYMux38Xr4lH68t4/ADo4cC30KJ8
EW8FyDsK1zyJ4oIO8ARQPRIaMjk7/zsapr/ucvEmBa2b8d9IGRLJ2x7JAD3i7nmZ
l8gvfLruqMh3cP0iQ3f2NH9ZmHQcTEEQ+Msf7ErbyiNCsbWoK+M+whPs8nbD+a3u
`protect END_PROTECTED
