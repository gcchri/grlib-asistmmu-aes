`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
re9usal1F1YWCZkmKHrwPEYHEb0ParGGsV3TNzVBNgdgcfnqNRQ0v1vPOOhFH/Id
zaoZ1Xv0ggftE1+JO7NMoC3rFlAmsIvbNwmmcPRL7+22Z+0uXl0lX1CZHxC6MPeX
vYonHiKuKnnj5v+ZtMRb3JZG6YyQ3COmhLOOQ0r5Ey9HEZXckTwDNiyX4AkwYA2L
Ct+Ha8b+NRnFnmE5RWi2JpYSUUJGZFE4Ktt7LhqC5LyPSmM5beIzB/E9eHBi6PeR
AtlO4c+2Cr+h9IPzw+pbnQ5u/nVWhNbfF+adqRydUEUAVZ1id/UkGi0l0lz1OuJK
c4Jsq1ejhXTYkoVSzuPROE2SkqKqrRXW/QaDlchKqW3AWwuy6bvrUXZBk+nTmKns
b9JOZWRIHEwUyv/+ZpsDjSEOhsVJn9drZWgj37NoBsdViJiZk1YxrNJ8aD488TQr
PT3pL22FoecI0UBbuGmld322081RP1z2zznzn7GhfYqwoBabdGCo0nRyC0dwAL9j
vsYgmBwUpqY4JvWp6Lp3MHODEdEw+uM725OVui+8jVJ+lvZoiJI0jTWRtAwVajRi
4Ya+q3GR+tMFCGl4/lpvrHR/ew4reCl5vgMiKf31N71IBK4/9mWtWvhJ4yp3/rwU
m1RqrW97IBviguubpi84QNbr70eJMtYmxwSnnbi5a1FeLR778T+sFd0710fSnIyp
Yrw1sedNUd70kACS5OYTAI+A+ZeMCsHUMYxZzOhNTfLKfVfz5ADGAwIA2d2RI9Ht
JDr4q5WCQtxBIGlLalmYBgKiyQ3i0wHg72UXu9ZpLLpq3e1mM+BX0361Xg8LHd/A
e+ZMT7TbLMFSRf2Wc2OUhwrYHztXkUSa/S6eYMiORPUVhj5VMgeAZ9Gc7tQexRHu
2z8+JKwzkouTOl0WYGftTXcZcdvObQ6VW6G855n1ya8P3Mg5C2SHlRZgHpaxyiuz
t+tgRhmcg4UtNtcOcrMxpi2AP+CWOvLk7qFTNEgz/Ws6uAft92XNryWaiZ8Uk+I4
lKrOJcAzQA25lLacPpwc9oCeolNxUcW9LDRVDt80N9zTXnlnwVVInirEC3VZSJIi
4n4L6br4C9UkPLMxMIx/C+F8i2S2uRq8Ns21jcz10fGH0k4AU2452tbX6I5dZSGz
`protect END_PROTECTED
