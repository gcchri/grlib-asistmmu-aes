`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OYzTPTy1FjxTVz4+CyKl58faXKPUGFM8pAz8rJVcIa68IbFhgVYPOwp2PTZR/1OB
v3b28CdWkFjKhr0vi0gVKVsrLL/sUS5G+vlZiblVZZkT+13XWjNvLH3EKTBv5Bfh
ZEAMvezqwbKEGcsw4CiQtnWd0qxNMfv6vKpQCc18n0qOepmwYaYZF4HXOxTHOJSj
sWG/IiYUbshT8sPXuTgQWkkVuCDdkGoiY5S5zusw8Oo4ZjlNcFeVsB9TAYdGZav7
gla8EK+ZaOYZ8YP86hyS340iI4K1Nqa/BeOD7bN5yvxijJ9e+0VQDP2VSFHOUO5c
GHKUETySb3To9vPCPslwDw==
`protect END_PROTECTED
