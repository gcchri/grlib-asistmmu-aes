`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NgmV8h/bpPXGJy1GbFtNEqm+SBdFyR2LNy5OEzWcRA4SpkoYhsyG3LvDbMGzSy1C
4CJkWFVFlgGRNEs+PC6b3brnuuY3D9rlYfNQDHXV0LF872D7NiaAa/IW32qIfrua
RocTPOABiHvdwWbx2NQmafSjXdPW9oOQ6A7yD8kzHzkmruwn1bAWf3BIbeihHgbE
Dqn3cfp8IW8zmO0fQwGZDDCiF/weSHYj3Y0r2vB+ad5SANJLNfT2dnXkAZ3evC5f
syZGfKnDyb09ZCEw3semRZa3JfxKbz9x1XbfD9/i40KBBzf3sldqcuWiRPZkOJAw
AuFrWncDSgqafO4f7UVqRWI31B3ODLC7L2Eb4tMomV3q0E0kkauT0I1UG2l7wtOZ
zSSZUZBmkKMToPkOGQUJnnTXMVeYD2yu0sbiiD0ay8k+fa0Yf0XVeDiNSBAQEuav
`protect END_PROTECTED
