`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j3jgv2+2NCCB5p5ZPagljkIQAsN/PoaFwPEpoXnf8DyxER7a6pdYu6ZYl60JzjQA
G/GTITBY3q9y2OHM8GwmLVoof9TmesBh8b5mtrmVxLp4+9/C1UwXFSfSU7z7JeCZ
V4xhvg1F+cge9DiOWzdcVlqGaIXoIDSKALe69YpzNdGsibWYc8DlXQhpg3cBUmAh
hUrRGFqYdwqzwvDqH3z3xh04wo3SnKIVgCwbioFwsrI7Aega6Pufe5SsP0LpwfuU
q2aB4tTayhrcTkINtgn/BVIuAFPzg2Ih2lHxBhENnyzMS36BhiR7Gfa4N6CiBldO
/HNvkyppFccQ4lUZ5szNDQ==
`protect END_PROTECTED
