`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iqFW/UCZ7TwWpmSJJ6/RL3M8nH4WKfebYtuoAIPft7uWqNcEEP4vLhfVbGXxagNn
figKx88NlOusp0yS8+eLum8DnzX/1fTi6p9tKcf+0LjvqtVyEDa0dUWHXdqt3GOR
9MlPvIg2GFRuJsCzkRqRcsTOvjcFsbYlwMDMbRnWfbEoKmtaxAkDVASLwWKbBSQJ
mqmhQInjLB7+r8l5e1oqNq9eclVwee4ylnIa6j+Fir8JRLF5mdBEEBqWmBem1mjJ
p0P9C697HewJrcbM5ekoFAcAx2YAYHt2FDV+bx2mDctawBRm068WF6P6hE5q11r3
AWbClTv4qjzNDg8uw6qzdYrojeH7EwWPvz413dVioJvbbOxE8mBSR3S90pyKBt8H
iq9cemX6JXF/W6HT9NeAsB9+qFh239PBt0NoHyXBOKX7WskxJjdUcZNabcGgDTKZ
gtHpo8/0iE8NZLd2HBZLndyqZippZo5l98L4zPDXzag9aPGYd74U2Z/IvIdc5erx
nAO0UISQ/6fOn4yqlwnWNkrGD9g8T2qhxH9x5lXWrJI6rPgafjuGQse0K84Esp3P
`protect END_PROTECTED
