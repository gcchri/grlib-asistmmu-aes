`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bhV317a7z1k6rDA2bajCi+RU3IBeDjD4KNR+ZQFPnUML4SdMpUg2qOt9pHH8zTiE
h0l6JCK9t15jILSoNYAVmCdqPDYaR4rP8tLrOe6/biaGwSE/yvY5YIiE1i+/vsQD
ky1VkwN5Stw9UnL5DmuRz9R8nJGyXbvBSnCciVB2QcyHKhLAnCpPcdmpfw7ry4FX
z++mx9Hm21EF+wAsK4d7Uob0mvNe2DBVt0JxZ35l95+8GDHwaCJXeqYk0ET4SkKe
/ylisI9OyQSBbB17n7qOGB+ibNaBQAN0O9THmP6EffUS63BWrn5VcOqhdF3t2MnF
7tbmzE0ynOw/p2SlcQBnyCqVs3KRuT6HTnm8WPmsQnh2L7bwVL2S6OV+T08N03Do
2WkPGzjCYqam3keS3Q7sQ0GWUX42gt9Ar31ebqF950c=
`protect END_PROTECTED
