`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pAeUQ1vtrc/5gbN6KIVWy5zkGuzW9pbbZJ4MJR+/qGl/rGaWTh3vZjmncqrjeX3F
8adOHyaKMHl6y/BigS7N1Fv41IB/O8cyrhSv8v7D7ay9UsOIszTXk7OukIOEq/AV
PIXLxxtx+U5NdV8zLGD/7x4ky47ylp6BsqU9X5GoLSeOHT8pIHg7d/Wmf8z21IQk
/MncCICYdCBpev4ms23rA9kanj+Nvyu16NmrpGuMJBykVPgK+Y4lUtQLbH+VOqT1
Ryh5G0RZnrifkpyKQfx4cN5uE8RtSlALkPFQEDlqhEiLwZYAM7YD5c+KhCvtNzrh
Q1AM2GwxFIcL2mEd+qaEF6up4CfoRnSf1WSYXq3q5V3UcozYXjwQ0KkcmBmupmXV
ZTM/NcKUtQqaJkP/We1tCWT0RccF2o+veVAWpf2AJGib+eSBILGKq1ER/aaaBxJH
vuayC8Yv1bEN9hvRpzi0G2TgBq3Shtx+/B5cvvn/1faYGcp6HANkskYQfZkH3EIH
1FpsxMR93XopGGzIOaA392pKuYE1PXpzRrwiir6vRQjW54ICbHFx4GNGNjsB/Uho
GaVBTtsLBpqDK8oK+UCgs2P04QrR4Ltk0fTn0zfknjl6DbP/0KzgpIi2Dfn8ebSA
mX78PJy6VZD7t3v9LLY/i+6vkr/pemsE4L9q8IuJBfgNdcoX8Co+o5VbQDU65/C5
2DXR1Ga+XW5GQAC82P2UGwkQ+gbLE27+j2zrVqY5tH94vM4t0yDR+ait0F2/aP/S
jDONAvA2VLXbpmE7Q8dMuV1+F5j1B2I1MG+SwjJd+u1ve6aC5jCwXCLHQvnbvtFO
PyBS0Vo85sFNv7/BihhiQ0rs21xmuPJlVV4UfO3uI002uxpSiRhdBXDch/+10FH+
Rt3X/kxw5AZViMZWdxPWEiL5FgbzO9rWX9mlj2GwvAk2jpKgY47VZd5GI9UwkkzD
`protect END_PROTECTED
