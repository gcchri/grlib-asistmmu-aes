`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DadIlM4uPSPoaS9ZpCJMlY13sHSH2FQFbdjbSUYvnKjf9cCYERwRMAGMUAnGxae5
lyBGqYj4Y06p0HRC6VDsx61jwAjkAiQDp9Y8lrf3uZisda4sn+6tBIzzXc5oWWAQ
tFWEi+DzJRM5ZlE59DJBh8bvDx/rmfMkwJx4EBlvu6MvIigYHuLa/O/+t2HkPOF7
Bp3SV2EB9m4KTvrZDIuV1gLKUZEfuO1F/qzW7zeohYZ4+pZzVIvAnMT8KlH+wXgS
o67vDwLgQ+mRBbSj+mJ2Bg==
`protect END_PROTECTED
