`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RfNi3bBbfOGV+KFjmZ65a7nZR2D/ey7Be8leizZ/x+AUbbE8DVAL3HERg9u1asHr
FgjEhx+ZY1wtzEIl+KKXvONbuazJGCk4OnM46Avxte8fHGIr4ujDvPR+DhlLRN7p
ptEFimKq8dVBbPIs3NuaGowBJ2ixt0IRa7fAj96JSq2lcXe5e2si1DTosAHPX9qN
XgWWNKTK6mBzL6trtA3p81Y9xYRgTFB6D1KVDiBpYxITe1jVu5rpNynyWgD9bBs1
DRfevnHb1xsqXOF4Dr1FucYNDG9dOLPSirN8S6Y1IwrZsSuCDsrvXMGfW5dLsic1
+wAg62/H8oXzlKDtmluuoH3GHnWP0wOLGoRW8ENetPAkg0p4zM5ww/fndI54AK1q
UXvFLY79ZGBybDh00YQ67ujoRLkiWbQDZNTBShtOD3rcOIOoZDWU7jCsIxTjUTEF
FLXUyJf15hElbwRZjkLeY0c8PLXdkTGCwraN/asEpIh1wvyKDQLpPlz1K0JN7rbo
NWffm3shOBPpZSbDpHzKpjjE4PAZ55OV6hC/NYjb4LgSXOmimORHw1cerbSQBVzG
mUqagR8zleAAFg76VC6KzapRo9+HL1eaMO7tQF0Kh+ShMJFlR1V0m90q4reHLfbI
wlQgHztx4X/2Z4cxGSCkxa7/BuPfpcqX9iDR9kqA5eOEWTkBMG0KjQD8+EeKqSSc
MJN1f/7V1eMQ7qtHvj5KGUoWLYhkd3Jy/YJbCNhglBuYWf4e6hTS7qwfCwBuQ+oa
ndQVF2VXEhTWlLC9zf6aAw==
`protect END_PROTECTED
