`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8i2Q1bxWUhtQOiO6x9/CXaxXMFWJrdLU0blmGLpZcx/PGl5Z+EQCeZOVZYTmxlpB
9daruSdjUeIJ4dya6dwbbMfh7YyYJfPmB0P3ZdTxjTBJbNjGBPOGk5TQty5hGFCc
weA0KIhJxYlEZE/XsW5Gw4Ymw6BErZzzOy0nHYjqxvzyyCB1ahBqTWaKB816gGD/
vXv3CBlYs6vGy8FJf0xDglJk4napvu4qb4UvMWdu7JE8uQ6siSKBAFd5D+I9B8+H
HubKCNb5WRpYVRBjydeOCTZey2JjVHXdYcFGZ7wB5TDFR5WrzW968BzSFWI7vUw4
7lGLCMitVlv3v3N6SS94DHAaHOQIUueMVevKok2Jbv+Wl9lMhor9VhZxJDbNjzZC
Cik0VJcq3C8smoKIZFblEOvfA6iRVynUDiEtgPT9HbJXGDrFBrwLZTvGKgZW8wDP
pBFv2cLQvFW20HRBQfme/blMTpRkiB2JH/C13cuqpHKsoPbelbkL9OHUyEyzrOX7
LbD26Z/SMyHoXH8UOMeK6rbPX/860OVSBREvBOJhNCKbkuTAAsscxRh6PP8VARo3
E9bNI0anvg8hWwa1ZDEK9S8kMsmjbYjsAwhjc0hqWO5+sLcNiGKy9ErGyK3kkCGL
NtFm+BQhd9QdpVqIZmMGcv5LAvA5+HyGroGfDomyH8EM0VSUMKNJRkn41x8KL6Jh
UwuDSYDgzJMTksS7hFf5YNHFYlv6ucuQJ3UMpGSjqZD748LFFetIbkSNMhJpZfEt
QDLbDsOVZklZhZxo2N4Fa7kO2NyQ37LnVw81JeDGe+fqwJQD6VS+b6m2yfrIoEwZ
WVRVIdTRJxGf/i73gxUxQlGA3MltXXyq2YIry9aSA9BgctgI96rNtZb2eLzH15Q6
yhBzGj4h4XDmqtK5xgzeLlMt+NcpGXujZJQN73uPi8Uyz6//HD92Bi602HUwKEwx
43E6/wQ1OhljgwzdTO3P8dZpqHvYwa1hb4HKWSzJWm/iQYrCAEuQ3xoQO7UJnPx9
ebH2gjE0P8IxdPQa5z71ptkbWeJYfsV6jALumpIj3dJsssAmBMzSBocgMy+XNl5A
d9Ky7Vn1EVewlKkCH5p0zm4EJe5LtmIgYMtGfJ1UnmwqqtK0BZ37hI5Vz68Btg3Q
hxy31GUP6Sm3hdTWwu9Bq+jOpA5SyuU42TMlMxp+QMFIX18HDfuVrxCRyQNHR5EN
e62g/uu4NAqMW0de37Y+bas+nTRCRGOBclT8QKbnx1rvRuND+twylFicRJ1hdwA0
aN02ZDXFoIId+gnJUQLQW3YlOfmiFd4Kama/vyJe318OHG9EGWwfrB4xKQXFAjR2
CDTXIvdM/ZmC8dYOolhH5f2Nfsm01dmjQ69Bt8XyH3AN4Z/tEXOC6/Pxt88kRolW
FbgSJBttcndQBvpY6qE+OAGysXfkJFDGdd8gpkZ6uLfuw1qR/cVvQPgNaExdOzYI
JXVhmlIDiLr/H5YKLcDGcd11Pe+suOT7GvUiwpV8EmsPTOZB8+SufLEk6EgIbZ6V
Xu9R/a6ZE7U/AcUaJ1n7o3biPf9zSYKI3p7BzftiVzDYF1tlGNHmUgIdNYTihgm7
29zgL4COjD/bhBf7igATCsdH9RwrB/kDMGBjfyMc3u1LpBRITT5V25DscXZvkJTb
BGXTLv1sbAKJsysOlEEKsbFcQpjud9DN9C+KS+uZ+j4XeTviAVjdCfM9ZBinqx9f
RggU1lfES7lXlSbyPlC2q3jTKpL6uHcWFQtDVQ6XoD3niz1gA82ECTnMNg5pCbqV
CHa7bA+5ynPgt6zze5Q9dzlZg9k0ObZNgRTXDiVYohGAcqe1r6TJAoOdP6G+1yht
IC3XIkw6IoE2BBysuZcRFOCPKq0+WFHxP9WndX9yIqE0AnrcfUWHNpZ3rSUO1Vza
2N/7E3ie4bPMa2JsGYZuEq6IgmjhCGgBYevXNJ8LwgOJd5Um8W5UNR2hv3iHaNzs
0nKHgEPzB22KpS40DOBpZ5DHdrRhopSidDb6AeK8/xnwQ/OERU4CvayyRrHTl9D1
oaTeVLc8oOCAhZ2QzPlq07tfaJjk5dssNq11YhVdXi7TSWKf3yzJE0t0lyB0gS0z
o6fdexc3YE+pMN8acP6ycXdJ9B3daCKqaNdTDxCyhKSBKb+tsspoMpYkfFfEiobO
`protect END_PROTECTED
