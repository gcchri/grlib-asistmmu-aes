`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f4tOT0coqV40C1uPSBdtex84hH8XYD4NW3+e69qd8F1rtT8BCkUo1J6aIj1uXij8
rggJ5yqlelkdApelrVVkVvDuD4MRXsF0bH0j1/mNequXOqGx1AtytXwFVWYhGTei
h3w3nKGanh0tLl0RJr+0jTzsP+zoU5Z4kz0V/xryC5wT9RPwA8EehSjMYRTkzrjT
DdTe3C45kcF53B6cbVawKf8AeCMS8vP3xbMdJkWzJVwt0Ggkr0yEQfVpqGCOnYbu
yFMvrowrCa43//T9G2hiCwSyy2F6acbqQq9vhIyHmyO8Q6thpkMaabWJvnopUT/d
3joHvcmIf0rqGLRhdpbtYtizunyM2792nqfSH7lffU+uAyvoJCiyEYVQaOZFYa3s
pijIO7r2DjYOlZ2sU/PgXngLW011+63aH42Lm2NkvCsOGfcvWAKkwkb/b1Y9Me3K
zhtHA18jhrWiudxh90xKUSii0syzEkxnX/+pZMFUf8Ls5GaE3b6vW/EyGVn5wt/9
oVsIq9qYHRNgYvxHiKB0i2BJDHTXsgf22+LJ8uzzbNYKVgj22EVjN4fw8ty84H+M
uzH5WLQfYfAfH6z2eG1ARpN0RXgegfktBmi3jPYRj9pvoRpLl8lCkbDbgBWehqOX
rskjb6tvApmoRPvuYK2xvljwZmqNNmfIeP2XymtjfGl4x7NSYApBcSqcQxYIG5m5
I6FCGbGjXHuH/HDSqC9sPE9mN5s63fulvn0Aqo1jB98=
`protect END_PROTECTED
