`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QdLBa8vC9jhCUrOXCGs6HiczqcogI2VAb37JQLiZ48G5+SjiAPdlCIAClYCJ1rJ8
Je9UquNcUcC5wmnMNbmxyRkiMCuSFk7lfvvfhoxC1JOckTuTTrUUZUK5d7rgc3xK
MmI1DRr4z3tyXLM3thDMbJ8Rd1Q1/VTI2VobIZIiG4cadQjZr+OU46nN1ucbI4HW
9s27m5Ok5T+GLtmo9pbeV938Znh8Xp3gocQP2Jt6w7x6SLdLupOXldXGfHIfDSnX
ciiQZYszJorQxOoc14YpPLAf9xxvPml4FMN4au6H9lkNSBa9RGH+MBa86CJDMmxm
b080gor+pvA20HRZcMioEnXZ4oJN8KlXzeOwF6k77azZEVDfVPadKgybGHMI/uco
wcOPXiGZK6C6HZ6yfs39xGHBzjYSojqbVBG+lIoFecGTokjUDHMcvWDXleUg6YuS
eYq0btSdlYFmEx9lyjc56GmVZdYq4OGPts3RFeO3KMXWg0RhFMeinhRTPJEonaqJ
5z4zcyWvye6ijDjTLl7P5Hhd9mtXT5oDA2IxcLcRaVmU0rSX8si8QpT/Kbr3ZWEq
`protect END_PROTECTED
