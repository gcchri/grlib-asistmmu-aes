`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xk34DMfSv+nEx6YS5/LG2SsWHe6W0CDBRNqPS6vo4nw5xI88DIE1FSyE+v3K7ebV
SeuX57j+lMaTlAVJoQNRSp3sfxs7N7nCF+EQgGPhHvg14MeHxHtyFzHrCKk8zmh0
kjEIxMoWu/lAEtcOHluFF35cPvu6TNbQzp9vjF2SwNiYANTYZ+u8LBiHk9lPx2v0
yalJMqqaSKwsgY1mp3PnH/6KWXx6v2fPqLGiPzyxT2UcZ2854tWO1kRzFFtHG4a6
mzbKxyWeh0EY+zi0Ts70hFj3LtXiAdZZVbJFtwUDirHYRHUScxvKiJu7FmC9s0Sk
qskxXzzLT9GgnowKCNi62w==
`protect END_PROTECTED
