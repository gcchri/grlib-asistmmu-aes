`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xo9AjfhIcVMvq63egt/fEkUPwVSbNPPUvdAbTyjv2SmxgvqwW4VLnIa391KfQIYm
NaA+cokqeovZpWv3NSgbGT8mGvAonqOQTwNVGJTcjgqoCAw7Nn30E/zp92Hryp2g
Q6oTISSfLQXmepdRLOkR4g2wEvE3SysbB2g6omPV7E9pswrZXjihtJFtX7bEcWs+
V5+7h2yP3NRoBnhD6+QxPeojeN9ROux+0iZlRkGAkSlh52az96qg5rhQAdnI7Cdi
z2KcGw7gbLIL4sG77jo1skTBc4UWW23yUWlBCf8gkv+fHfJ4bYvyeeRzeDyRMhKj
poD+mx9ziJFR721xEuHaj4sgvAbEABUfsMmIKj0Oe6D+ETyrjF0TICt1D8IPPTBG
v4PalVkGev+YMtC5ev8nE7HRGfO8hCNjp6VJ3szhkWI=
`protect END_PROTECTED
