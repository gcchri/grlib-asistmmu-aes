`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5+QYXlJdTmyhcZa4ufqLt0BVAKeOtaVa+HiDHk5BoRe6RYxPXYrcHLqT2kOlfuKC
GbnBZIn8A8pXFgij94zuX6i+Bnxtp5DjdQldUAnPAh3R3ZsFoKlxDPTYLfv5QCOj
TJbyB75c40MeOfQT3BwVYZmR+hh+0UrjeVauBFPLk13Ve7++XG5C6YeaAy+7pFZR
ofPvsLkpglq7FvfHl3/PSGCNfpAlEpNmk8hjAQCwqvuSWl1KMm9qtsIPvAo9bPm1
tsHdzfBjYa/8YhMfexS95wJPrKtcmFd9vCYR69Bgn9Bc3j5uca6I+/2EaDW/m8Vi
KMvtHwlP68wJi60vHnP84sNuW0M6JknXbgj88HVkIsReyr/qbCPGxPA2JiFtGJnq
iwLz32kC1B+gvZbHDJ/Wu1oGw4TD2ublTfeiAyAU4N5UTd1565jUNYgwYWe1DACi
v7S14Rk1YYmA36vBggPlPQ==
`protect END_PROTECTED
