`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lKdZuM9GBXzoO53ww0x9ricbqcxp7dqZy6gH0jyPhSVBZ6OY5xQc2Z6LS2OLKG6t
gCOfBzoAh7huH2p1DyY1pTwLbNR8S+4w9t/BkjG+WeA5iZzOG+44AHUHFbQ9dLNo
Al7OTubLCG1+WW5v+bPQBL8LOthU/luGJMW6CPcoJOhxSVF3zjgZf2ilK70LgsIR
2/VTxTJe4OBoupd1clGvQ90YpRbl/XnfHNtmPlR7Pul6a4cdjLwoPh8AEQo2hRyz
cNwe6WYiEMY4jvZR7WNwofFdIPE+gudu7gMBF1+ZCu9Q0LI8DBG5QZu/pV6LjI5g
6p7vxFs/M5wQEjh15VeDPeiz3zaYTf/uPb+uMObptvhBX09Sc/t3yDS/s+4rIAbq
CguAQ0X22/hG63ZBY0I8JHzVVgNgWs5/ggL5OBsT408Gqm4BKILdM68Yw0rx7mgc
FVz5MvdjScMpfi4/P/Tui4ITPXL0s3E6ooEXRFC/HU+5issZue/fKSk1tVI631Aq
iZy5Yq5vefquo6ysQvR8QegKy6+El0pPq5ABmA9tvMAn4cdAeMc5YEO9I37tKyK1
yQjGsJy58ecvfsgzEdTukNfPYT75vMv4BlP+/A2eWtzJ0gioGPsFjqIo6SHjCl8S
/2YqE1AD867CCFN54VRAJCvhlxdRRVuvmV/p2X1WNr/OnwOEKNGEIxVb4c9L/sV3
gX88jhfI80e3EHcItME3Hf5AVlU8RYA0Wpm7/6p3pvf3MryFyjIj6hToWNy/Mjyr
EQq8R0y7pu04okeGp+4CrtHFRw68bUGGWrLZiCN5YzFftkQ2VLycfCI1fL6fQmsJ
sdDjZjFzyTlRikal4cWYd3XCbzSK3mIeesfGtoBTAYZApjVxKD4s46gA7cbL4ng7
OEvASbt9Q2B4C8b7UYnsETVH7dfMpCmVH/uyATdCVZ8Aaabu/SqrcJcvry9kPDSP
XV0xw5Piqqu8RWL2Wg6gPMdzOxVlvbTiZSB3tz/yaK/JnMCPZw7uIpw7n3z8FEwX
THNFADKhHFwSoOvLXuPp0ZLUwhL5zYGlQKGXKxsCLTqHnHxqVTAYLOS02s7cak9k
vx9a7ijfNx3HOi+WRA6brK13EFqsTwl1WU5Skxu40/ApNFMP4eGGpjHvBd2X/RyP
vRo+xZGmqqKr26G5TyAiDDQsMfR7alPKgvZjDqJln7YaAAByAXDevFYNh6wbkC3P
6mjmsyHMUqiM+2hliFBSOl+R5g+BzPp+EAqAyz+lxYqrYj1IVG6wxMmMXw+Q9sgy
k2wZfk2t18MRoT0oMFyiF3dAY5hgQqF7InCLuu17V6B50tK4uahUdhusM3/G7eS/
d741rP/+WhIByJitqB0LthU79zf5nPwfYWJpXQa+2cnGUlSan94OPdsfMn3V/FnC
C5oYF2aru6sZ4vp9Aq/kdsoVGCYbFpoTeaooey7f63FWFiIDB6oBxYOyRmD7VJCa
SXmDpbun9P5Z28sx7tN5q2wh+Cwte6X1ghmFoevBWyqzzgR3bNGIFH7jmmdrG212
VEWWwabgh18wchQejqFzxIaLwuywqMNkNIdld1rc956Plaz1MPi3IsOmH3ZdUDLG
8JBVdxH7G6Vy42vMzvhmibyafI5JwrjDcZM24JX6rXqRn1OpJ5tsQQWli6hM6oaY
8nntAAclqZHuygaAAYl+3d+KpOSSTIBHu8hYacOyeKpnQSq+WfSrXynYQMmgpy4i
Ldt8Bxfn+FJE2N5zLCrX1uOHPytqMGL5G96qhScWbpy49Llc8jb9ACXbgMngqrWI
xY7D0OOCcWpb1xxxksGhTxDkNimg98EIXD440aBzLAIph4nX498Ff7iSOXhebU2R
EBIOxhCvqgQ9cVfT131eXqPjwEq5A1XCDR9v3UJkeTVXsCZpiNPgFSEIiNQWwtNX
9+l1SB+rX6DemDC5ObrFj9i8zK6Z0C2Jdzcp8ZXkK98onZz70cCUyC48q9IbyUA3
3jIrUWkclWRgrAAR56VARpSOll0e+6z8RcLhAzpM1oW8TBrJVLbhuM1us4+Q2uvM
L5sr1CzBvKc6INOwnv9AEmI72Hlxjl0RzRIklgkCNYfNZ+NY92KYuC3LdIYs0EqK
A86m6/7il8b/Kx4mamdkbVFMhONPB+24hOLmjIsA148=
`protect END_PROTECTED
