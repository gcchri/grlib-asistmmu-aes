`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
neE0QJQm2hIPf+ASkoGCi9IKlocTLz9V0kEzgfUSMUtdR2p1CQg5sE+1WFAvAaDm
ONr03UGcQnAQyKCozu7NPPskqRvBL9o+tpqsYYfwdR4tiM5mVHNaAMwAXZ80Yhux
CPfAJkdtXQxvNaqC4Ujbk6YXSHT7C+b14Laa2x+3IcI3T7O4ESgwnLg6eUeM8psJ
QU8lNjcFiILHY27xRN7VYrwnGWXdNrJssKZzpssOXY8QcV+488dgm+M04SsNeG3k
khtHJmTtNxd9LI624PP0+QOYWbIzuNqLc+mCoZE9yNTOSGW3p9I2/mpWMPAXZvZU
tuAYLzCkvVf1FJGYl2pNof3dQf2+8phuO53aDlhzyGJP/Z/ol7mein73+sh6X4C3
0+qxSDV6ADgDo3DTD9VLzlwZXxjOYQKxhUm93s6yGWl0Apglj1h6NYqGB3ZE4rEE
o3HJRohkLYHyqsFnPrcZs6Xh8VRf/goEun9rOzP+eh4D2Y9K73teo+2tAGdsK6nF
2HWq+5RDrDVhNmb6IDafApQBfWUG3mJ5L93x1iN+86MG/AA7hA8fv4Gs3Ro64mIR
R3uQ9IjSXcMtJShoLrofpcCXNJwA+oZfTuXh1aca+UHaMkzEWdPLP0SVGELDK7XF
kMqjTf1x7s7pNLlMfv2915u61jSAhSCB0QpTIbIDJqsL1K0nyMTAu8bX34qWyaxg
Q0NvBcA4lAd0suMB3wLUhBk8UoNs58wbaSBCfDiS8BbWhLZtgEQCyZYpDjdi6GHH
ETVDn0VfFSILqBfPdurE8zuZy2Ghq0tqqCFIAtcMKCeQJym34Mkkq6qH6BDiMQ4H
vcz7wRpFGg01w35yBDAag/3YciTdPLrZSe+4PZA7AOal8bgFyGSXnqqRvBR1G1tl
XunPUZ1pGYNlkEm8uRP/GY/xpqv48oWGewpjIpeU+O0yxECHwa9Uov00APH0cf2h
kNV/aGn7zbYQ/4BFJh9w75j+LEl9eUJB6NiHcWXmsmNkxqizVDYKZM2fjZu3rONW
pIQSsIx/myqJWKReKqg56HbqRtBirJbGNS7ncnc/9nstHvw/kk+WwfSYdH6/3Xmj
UDZXlYMK1+0rV4YLkLXCBL0agTKeOGpP2czZQWyJyNzKmhLigt6di97tMoEhP21E
nEenrLdq7soFpJRzoPY0HakmBTw7aMLjbMxLampMDEY2XfCyNGQg9IUztxWsaNDK
Ii4Ib93JILLpFKWZkUzPkPum5UUdVfzgQiUmwsguSA7KruaHVJiCon8K8HhlRjEB
lIojfQ47s/sJEdPS+I7gNIYS15cTjdWtSrXJdHknGpO8Zrp+KYOk9ecz5Fv1hVTG
D2xRvZxoAkjnJM1eqY0fog==
`protect END_PROTECTED
