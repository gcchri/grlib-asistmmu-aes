`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uqKw48cJHdi99zaZ/Ojq8Hs2/Ya7X374SRdQ6yij4UeU9QwzZRwrHk6toL9ok08r
PYXZv1wI+oWTbxs+xkzVKh0v09hzoqQ2O3UBCyJTaR4cu1TqKSdIcD9QBE9n9mzE
aT0DZ6XZA893QjTOg9leG1USX9JDvpZ+J4heMt7lUTk2545XHqYp4mavI4lgoryV
1b9G1c8TGQe9aGomtqeQTXWO4Z9kmJ7naHMyjF1ZQx+mIpyFUp2AXwV6kusIDu+1
qLJUjSjDz9GjzevgMZ2jAqSMgAHcSBs6eE7Yc77KmAr3JZpotIaDthrV4BAuBexW
eRutH25DHoFWh8+SBb9pEzoMq/LDqeoXJlIX/pP/VnyJLbLvCLeaNEnyDpMqm/96
WWv9GrlV87w/dSshQ7beZd4f3cn2mMiE+5eTy10S7kY=
`protect END_PROTECTED
