`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EcFEJuK9PY9iRzEVsMXjJ40QxDZdnArY5tCg0iGpmdahjjlgZSTOzH5jGWWWdUNB
/KIT64xo+BS8SIG5MqhsZCWiJjK0bLO8LD+vvLvKq/DkB1RUVeY0yRpYiTDqxU/5
xhmhC6+b7S89cIetr/QQPfM6VyAGdkjybDYPJFoA0OVHtyBPKTe2Pd5YQ21Up38J
/TwHhPabb3HzrvdMJ85idUfAzZl2ZCEhzpMKQX/I9SJIJYh3EiheJXIfxOA0QAFm
fYu++BjjZfKp2C8gp2fp0thxK93zNx04RlCCecO2Jzb+1fhOUXT/7pwJhbDTrlqv
piaLNZF6qFE4mEyEEsw78jGwAZi0RErjBRSFTDh0u6lBM3bMXiXEkkb4ckWwiatR
g9sLH2Zg8FLW8lLDi3NL249E4ARFLOd0U4F8HaploeGDB8ZqbpSQSv6upVWskgGQ
zJpGqhXh0Yn9fcx6VCkceo+nbhz2CrgSNHLtd0afy58Zl7xVZXi8hRO8ZJbUNJy4
1cYJW6skNLX0ymwYxF1/IqBia4VUT1zaTY3z5AY0ch97RHJIu24SPUoBjjOR6ZL2
ZiUSxn5ePvQ/s6BTa1s5Cg==
`protect END_PROTECTED
