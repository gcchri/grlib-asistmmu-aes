`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0jMsG/D39+H/7d1sy7WK206tN7jc1n0jOSRQln7Ij8/wVlRF9+rqSnYNirrPQTG0
7PbiQLWRUePM5w21ovVoqy2ZFFf3Ywwj6/XNfk93QASRG3I82S5udEOyal7tMJ6L
coVu0UCkinZZN/jJcat11a/yZ1XxUW17h19HgXFpfjH5baOYWJqDYjiqS96vEP+q
u+bMmDsHyrpRPWaweEBKdfCnl+AA2CLLe+tLObnxN2PUQuKixTALSvWtj+m/voT8
zB3Dyk3TKVvvuk51ChlKujJQbo1k8yDP0bHGcglZPOrTl+ErTFnA6sYhLW2QcCLf
5J0Rt1uUMvzXoTg84JWttqjavW5mMX5KX1VisJkPFnEz0aGrHE3GCYkdcTYU7Tnj
NlNuBsfydGAtl2TVFnGOUdr0dFv6XKlHLxrq+fiyVc8cb4p8H1NOqjhBsZJa04B5
BS9i6qMteZtyBTbhzv9jl38dR/hApRJj0khxesEp8yRXSk4IFUXUQuVNAM35osDq
Oqgrxj0E8Q4c+r/4JMAGb7p71JxvCBpGNZlneINMQR4d3SGl1coYwTfRfHlKXKKs
FK+F3cLi1TvtjP2kg7pFuh8ASO7uFMo4rjcwYe0yMZeIudimTZlk4ZuFdjEgmbG/
Ex1+jwD0JihiTXiOTcPaXcGEUoH2iTTSjymIXDzrO/szpFT8YYpucWapWEM0kHem
5mBMWGxtlEnzWsHO87wDREsv6g1rbW7gRpZd1n8imQXo94ZRJRDMLVeUOh45TgB3
bab1Q7Q8XUDkVUqWz6Fyq/8tTe/cWT4elOwR8LZlpskUQscAPKOdLDw0bcAgTgyE
e43eajiG896TUTckWZ2VQsk9schV6SeQF/Mq8U2i2JOvyGaLrDV6imgI6ClsQD3L
1bQtgR095vKtXPPOxGMKOKUuwKRMfp7Nd68h2BPaZYhTp4EAIAR96JM9yIcO56/n
sTUjTCG/9GPB6fJ86kl1d0s+5GkW3UqpDovqadhJEhPFMk2dcdTsPkRhUEKer7uM
i1vTBZYA0ArxtQgpU50ISJN76FPlrGzx7t+t4BJD9nHlhABCzsx7VHTtEqe1dePW
ZkOQ5BfvJOlpp7hP/Nat+00E0nhpghGcAUKtNlx96O8oROYxENpUE/0pgCcGyhXk
EikVDBCJIPavs2zIH2p7CILUWpSe0LqIjkPZ7YKm2oPb2ZswNsWeeUMRy/rOHyuf
CPjerPRRniXiJv0fSpMo+G+3K/k5NBe+M1ho0ql1R/me1MYZCsHai6YXKsgu0KqI
ysztm0tKpqZpGW6pY1PJl+GY+LeWF9DlVvOyFrkPm6pdHm7vbgXT9eyWi54/iyYD
gaH/eDK+kphXogrUfBFjUvdkpbas9tUIelftvAcbeDevsAVtuZqDBHx714OG8DCI
n0m8Hdsy/31Pvo9w7Ppp/oCR/TgtKMcUL5fbgojSkqijdgRm8EHTJjv7aO9zcO3W
qc4DgDt6iZ3TZya5nmiBRbRRNAxPGABLMyW+o5nt6OZ/WFZHFr18f3UUwT9RYxJ4
szuSlduVbj3d8sZEcXNQmQPt6rPGrIHf5oN1U2tRMYHHkzEVIqHk3rHsUTtNsOC5
X4jzHeAwDJoRf3YgRMxhMpi1U72vgdRjaRdcKGt3CuhpN/+TOthET9cVPja4UYOV
RFE/zAeu880vq6WzwuE/yiwHF+C3xBXboDMsxjWJ+0PJJAt5EdMonC3B/OKTPSD9
jUjlHYpfu69F5ieV0k95Y+bVcO+2mvuce0IzPczzSNaEpD9RFKwxdSuRGz7P1HdR
OQIOv8ouXcACzsBtNVOLQFp/IqchiRG7BGJLtAUhr1iFPKKzSVha16CIkr5kwUvM
2G1q9Xkmcm8TOFYPNJAajXrwiCqdRXpbbojYkIh7p+E=
`protect END_PROTECTED
