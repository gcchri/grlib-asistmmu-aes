`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ZtujuTWMapO/1WKvdD+hIJqLg1DztsYX9ixpEsXMNNbEM9MjBpEBy2hcGX61Vzw
aNB9WeHBZpNIYbw3kQR7Q8wfQ5C+fRsPDG+0Ci1pZqg7Y8aeZQllRvguyXQh/uMn
MsmojCf/SCn6REfC78UIWuovv3y2BgoCP+s8o4BeOp+u2Zm4gImkbYyE8dPDD+B6
GZasz3g1SMOjw7kNirScA6uJfq6Ptlt0hR1Sh0m4pO77lussrH8R+J3BXwsTez+p
ULl5UPZ/TxF4ROwdrx7/TND4o9S59ZwUm0/W60p9XMF01R1zwEI8aGHNqmceg6R5
uxebmEHNKGyizlWAQ2u8agXV10IlipYpTUj7I5hzp+bN9KNGMw8JnPbD/Ob8V4lU
Ps0ANp2dKY4AZRc3C+mmZ3D2ZNMkbX6xGwfcJdu62YC8ocPFg0Ownv85Xg2vYsP1
XlCmH9Yyr8RUXZX765e6T4ekvd4qMet74rNX9JrS6734CIhCojDBAMQnmk8gaydA
ICmrQLAikNgV34r1w4XTn34BGizohyJJhiHe0m+Pw+rCSQehJUVFBVEOTpSO+Rx3
Ii2F/jBTQQNcGj/tV/4M+FAesYbI/MM96kkLDpZWR2k=
`protect END_PROTECTED
