`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M+v8q+l7UFaZWfTGEtTO0m0AaUtRp096Fbf0UIcyS1psP919qpX2kElKgjcA9iwg
nPSi3AcaGjH6doE0kreZrT38iACMoAO9KeUqnxmPHY5andUj+1hMCY7fv6JjUPf3
lTh7jUyIasR5ezCxqzNKaPGrVLhTP6LrcMtodtoz/mrOewnpAkQ8LMhd+SRPYo6W
tozUCFFnq6JIq55s7weU0M75n6M50yj697fAbB6GXe47BL4t8QfHAbMyz25wckyh
WCZFfE+To43ANJm9yV8aJ74YuPm+W9U9yM6B7PlC/1HAo2szi6Bb3WPeZ+lYR9Tn
rv7DUH8baPJVO3L+2TrkXt0Rq4j/DYfVmFsm/MBafzgrwT/pZOYYCHDyIKmFaZjo
wgb9bojb6cboAQRyqZ8l5bTfj/Wq0akU7MObsPjlLJTIt5y+qWcnOJoQo/TmYhZv
JKFfojhalCYnFKNHI9mpO5nAlUKj/4vRD0vhHLzpwy9N2g1lqy7F24+Wr+OcqmBx
R+fU83Knk4n1FHH50p1gKM0BqcfhGZNFoJHIOBIFnR41z2FIdFPoxtS+3/By/FUX
sPWsXErcV8MXDnnrNsVqT6neF+nDqWWsEfY3sZX5LuV/pGmS0rBP6A1c99RYjUzS
wHQpGSkJlEgmhmL3MeezOSeAkuMeAxtELtMaVcSml0M1E4bBphm2lNUWQoRGnMbG
/6bQwaAsVcArUri8OShY2w58Yew3BKhe3QS8bOjDSXzts7SIKkhsk5AIn6WV3Gp0
hFodjLRCcH0KO4tDQThKuKNaSUBJmjWvIsTBUgwT0gvL3qxa/vBiqySGlD2HzEjZ
7ym8pXvDH3UkhrcPeY0bg1frRPmw+tMeCmabiNzqbKTWuyhGAnakCsODQZqmgzTM
kzCkI8nRwd+sxuh+hDHzM5Et+OEygNul29RgPkToFb6UruEGIa7/o0TKeYhzXgvv
IJxnoqeoZmZ8i0RdtVKVNLwmpI2HiIaSsaWBox8X+ehXUw1IcBepviJY40dtYvtY
kZAVJiApBmjQXLg3nE2/YFXQSiw735q/mAtuOMepXX/Z8h66zMBtZKHcPfNEE+yg
8iMWM6TYXa/o7/+GeERs0x1o8irksCNmKlMvUD7NLjd1u/v8yROJG/cJZ+SOfPng
iaGFRiBPYit8t34dbHT2xefMImEsC2hYy+rhqcb/Vu6VNrVUvwttB9C4ctDT5hd7
N7nrBvKg3FQaIP7FfD2VlH1bOTmnkCKBHv3ttk185q8oT7oyMmQcoTCHWjo/yI+R
FofWWbVmxyxhVq/Es4braAU9/Ei2G6/tomI7sbAyrIxuaSO5wlcWmd0QmGHsDxUU
6PKv1ompZZWb7WTuQjQ61mufZvsTeI9WqMcAST7wmrxrIlV5Xp8Z7o13qpw9fAit
dO7ZEJETlosw6UL9y6k/Kz1xcXuMs5qEk46GzQJ6eGLSLQJnUGKVEDVNsr2eoqzV
rvfTzKB8CgAeJFnEoFEd7VKUf3UU5XmYMiKs44RZgeB59+l4q9tcC1MuoRydPW+Z
gX7dSJbfzS/eEru7lola4Wda2N6RjM3mQwIaxHoUMSxAmxRFx3WT7D7lY0UImdx6
HK6W6sDd7RneoMXwjXqQ72stIym3tVKVuQgpaymFeZ27TBLP7lGXUPy+PO5a//j9
uhM6j7ESlRiY5bQjxWPzdsD0xSYgzdIlvbaNMopR/YlaPWueGG9qnmaoVElV1kdk
SCbiZYIi5+gnI7daK74I2RXeYx1dm9KkC056wiyYTAMCLp5ZV++6/ShFVAK6Hx6d
qIcgf26JG1cT6luaOuA2TVsSiYhJIMtTfJ1CtmsYkSipJvYC5uqoJC1Lw/iu6n7H
CwgSkWFwwcMnyCM89zwo6/D4OElFctnOR1dAAbpMwg1j7W1HwT8K/QIZipII9+Az
gnH7mPS/rHIEcqJjDjGXdDSEOIeIjqIELwjaThfSMJX15t4oRt7xROeBpo01ofmV
CKPdedom6DVwVg4nE277Dx2KOeJVnnthmFY/QxAm52/kZv3fO/jjHEqqTQXe0gOt
5wt0xIWBdmQzLqKggrmmcU9dUPYPegqxu/iltfmFMKtiWv9WG+dfYMR8PY0SY1dL
5SG80Fy4VYHCjNWSEZCFB6vP9IarSfyMuEBq6cDX7RZdZLtsVRzrA41V9BmnC19q
GlWdqVYf56wIByJReBonBG2zk9hQWVpcE76eNTc2v8oJWLtKU/SO18dT9QFh1gzE
qJVKpA+OJs+uUTZn4Tc7y9BLpQ6Iu4KZdlgoV5pf5TgQAPD2zjxp+gHNzUyaVXbv
EZjtKbNTeR4XTNjU+tAmYHW28zsgELTRGaxmrImtxRDIOBVqeodMGg0ZxA9ZFg8V
sEaQr1Z04+GMbZS6QCgGhn0Vr19dfdIGZHgx2hGxvYiWB+j9oQmSwM9NovxIx1Nn
47gxLwUv6nW/LJdzWmP1dDeMpSJHb8jRphDpj7pvu8/ipXiRbncMmCTZ7gyoQMnf
T3KPxItPNKx4VTujCP/JaVqi3huc1jqbaMN3cemCAFX4pobhiSVsKZsGa5go3ZY/
oxTDZ0eJeRj0a39ZIWBxIYwbyP3Mtv8yufIlU3NuH4InteCkujaBsb8+5CFttTW4
d11qWnqNm0WTIbdlEQpjXSZ4rKS1bRkFM6sdnSI9LbH473CHR++STMY6l5RyRLH1
QkJnPntfMl3W5GdVHSDsNiOEv/u1UN4rAd6n9XSAZ1E=
`protect END_PROTECTED
