`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dzDaXkq33WpMfDCacFbY6edkl43bZjolFTtqcXJ0Ko469Ld709ET5maIMBaMzTaD
k5hNtzYXdjgTtWPPF3BmARpY60GJOpZDWDD0sducCUWyLZ++cjjfyjFcfdlqBb4a
xN4glXLEzsjutJo5GYSXm54eTuggpMGrdwjWTFi+SbJkFg3ujcwP7c97vI00GMGR
YkBUmKFrzaLDvoAoPMwbfyK/gEqoIDc3aMAtrt663Kkj9Umhjv9FfAxCFL+esH8c
z7oCX0TxdYq2t6UWxFMChtXAd8Ea9eZeZznXYqmj9HOcLCl5qS9S2CC9GTKnTVLv
MAe6rsXA6yXHMT5/tLTliIr/oVTrSBDEeOgsigsZtrzwjwa/+IOe+8Ib3Bel4SNL
TNYJsMcbtT+HJ239+pEPXA==
`protect END_PROTECTED
