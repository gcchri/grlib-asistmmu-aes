`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pYe57c8LZMbMhmCjJHVOY1sfNUG+IdF/hj6THQRKGgd4vBPawiRRYVW/3viZ7n8n
p7BUZ33Fekq0RJg/ec7PMO+WyLbar+yc2yLF0rwgqLQ94z4kX8U30wYsMyvb+tqu
5YnQMi7hPDWUTaeefUkFTR0XKm5WMsMb+nsm9A2sm7OCLgRlEnwbodi3fFsUGo8O
jN6zVNWMELxt8eQZLWUG/U6mWwnQyL/E4L4ktOP7hbPKc0onvthqC/l/8v482yB9
6PUYvwgTS4nk4RnTYK0HlNX+8hLyqJxKXplMc1uYZwehtZZp7naPEPv9diGjg0C/
abQ01EcPhhERHEWnl0SPdMl+cMdz/yty7x5JXagR+LRf1HtcSsJhOpScKHluD0Mh
2EBvnmHBk7KIpTwrr97UxEfKzrQhrdDS2e7QPuxSK3Uxq52DqrxEaMDh5drmlV28
wFha0WSbb4tXtw1AouJGEAHVURJwvuQegzRZaZnTYqaEYHJNES7r7ga0aK9Zvvpe
w8I1wNQkS5hngvDWvMdDOjPKaUlXcqw8Rg0ceLiM0jjr6rGDzJvpi2ko1J7EwxQO
yTzL2qVIe86wtjiOx1sL4DlTl/1MPyiq3p8hn9aRwTzQOfwngKg9hpALXmcCuTXw
H5yGcQAlzOKHgRhyvWEfmA==
`protect END_PROTECTED
