`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T10Xg8s5Y1mofMrR7nQIsN5i37gqcs4HI8vwGQa1AaEYcdTkgZcLYnCuhqXhSk/b
Udx+ONChXsaqBx1VjFEu3NSTVvy5ESdv6FuH5GgiAKpuAfOqmDSVDi7ylUv1AlNo
7Be+BqQJVPrfOv1jv+w9bceIZNlzYsvLLta1CzshSkK7WADvUSIPQ/QYlRJCMqWc
dc9cMg++d0GyY4hMAQ8Vix71BbhEvCmpTn0Y6LuMXnuvmw6+OzLM1TZ10WE5Sld5
J6udy8FDPVrOcElpdX20efRZ94i4J5HoUobcc8eE30A=
`protect END_PROTECTED
