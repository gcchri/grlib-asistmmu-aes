`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MKaLIbRqdwGL3TTXTObw62/wR+WYBXSY43miz/jks2btb+qe53m39r0k0ejn2wq8
NFl4ygfjtiVqCQSWfjfWJOFoJcfnSItYLKMYHgmmWkHiP6R0XJVpeMcW1w0LzHf1
RkwAcF2MCvWvVheuY7fQFdAKg3l+SkYYaPszBNptEoyt4OHkI1eQyGM39u7aSqnX
+K4MoB/QNSG3JANozeZhdxOiRFSIpWd2BVRqJvh7eKaiK6elUGJzYB95lakF0Z6i
p1WkX3e4G6u5bqWA4cf0Dfth6HPzgQxiFIy+pJsod6wqjTrVByOEopAxPg9Asbwr
QSjR5Gmye2O9/mysSwo98BvpRnnzUj4Oojhm24eckNURPdlTCYZhyYnTHLziRc8w
OkdISVaMFq7WQIosfGxzZRCyqFf08fI+gSWo/WQQYnulMwuuVl0W/UXfcFMgKUiY
12nZYpholsN4osDnjRgUjGL73iLpkC/L9OvDp5P7bSU=
`protect END_PROTECTED
