`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+LB047l0J04PX16TCUwQeYOq+sz9wWrv8EyVV+z69QvgNg5qzO4S1d7GSxr2/Aoj
5tVNe4wb76hIFJKLk5zoKruLMfcQg9Hypd51bO7e1v3kYVA6aXi1vagc519fEogL
MWscUDGKB7ScS2/zyD8PIu0JYuygN6UDGMpwVkt9qpIpmZ3NStMlozCflCcr2nyX
Y+dPpyMljHUSoIMLy7XyNyFG+Oe95VnPY9N7c3goXYppyhGsH0V9X8+5M7AUfGd4
eO22F29rfcShCQH+zR1s2VeRJWy4gfhgc1Kdc6/mb99VgQ3KbocHMPtCOZoY8LEL
7OvYvPAp4J+DzR1bR+eOW0maimMcQsTer6savI0D3RkTCKB7VStMo3sg156rHwfS
xwCF5ilblQVMCNA8gyWDbulAUdtzaXvwavUkjsHTuwCcj/ZucyHg/zYixJbsxDFI
2B7bhcPX30zFcw1/DiRGH2c/AXEpxmcintQRu/sZeCNjsyHvr/sW+jqez1TPjC0l
ZXGNmhfcgfK/Kt/m58R1Bcia5NrlQN/bYzVj6JsoJvJmW3EC7TCSpz5H1oKr1OW3
s8tgpYBUY9BE17dF1QbD+U7GdBuAez5NYcGQ1ADfsVlQANfGvOHxrfkx0T5BkqAY
sSEfhjHhNtYhQFkrQQu/14YLvwvVqZFSHKc0rTocgCyFYXfg1J5MGMwXS8TLUF5d
vOLpxAKTWY2FUSJtTRt81OYrpNxWZOOaLGgYzZUfLGL5nSqZrvFZ0JJnCjc0XQLI
jaQD+BMexnQv1482vDkqm3IOKnHgx1tl3kkmmr5GwfrPyihWgy1Oab2fZLM3aIKA
L2edjYGY7QKacHoLNhW5m+O5lnWYIlMJsUce2TSGmZ9/fQ4+t0J+ifl4tUDqxvNu
+4g4Uk3a3W+AtMlP2FU/5wGm5iHBVHhvzF8sJviQxNWoYLdi+dcMryU4vwWuKnHQ
`protect END_PROTECTED
