`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qpUymOnXcs34bNvp+ZGy4zohckYnNJo2NVR6xovtZEmYznSBveMWEu4xFi6N+vG7
8q81Ix2U+PPnQxM8iQQPfN0pCRCjI/UF/WSw1vHozpmLQ+URMuw7FBGJW9hT9CVK
ppoHQ8TsVr0J//5JkUrv69FXHsT2Pt9BQLo13PblYt1/hdHbpiygCvm0PuDurvy8
hus1nZv/gGT1+xcGkwtB9aV/a15OWQMwAUzWacFk4foHyZe0cgyI8Dm/LPMJM2la
32G6pRldINgfmEUkMvi5XaFIA5wzDMJFzdju+xltqV18tCYdLVXNBE8YWtiliQv9
KUFQ0F8YS/ovjiiC0CphK6AoK1nImID3/CPGg8WrwGeQhXsJ41c3CtWbmTIYWZlt
5UUAkBuNw3DkhGMKg+6J015JvqRVsFq2b/43P7JOFZbyYRXuvIY9VGLWctl+MFq0
4V3oTjpZqjFb5hCMEMrGBHr3I2CU1QnaecrdWsORyvNrgRJFDgkOQ9I6TrO2hBdX
TCRXCfpDRjGolHFTUwqKIeKJKMjkZwDSTzTk+aEwVuOnK5ethtkzB+SsxkBU2SwR
XLRgIt2O3YvA6BOPdp0UOgA5/eh9ynmzTAhpaqSv3EKmiPy3aDzhgARXZxw+A+fg
E1S/AVeDyT/w5+LDZktG6zTfqwsGyeSnwvTjlnv1T3qjmsLVscoGgOOs49edsCVc
HiSI62WCY4oiX72vNbtswdgthl95B04kPpbhaqyqxBSGMYpAxRV4KPUyoKJuUj/3
FVkWIrFUOVqrb8Q9/38kKtIyI1LOgdc166IFXFbU6V96hOhZM1GYse5lZJeh+BO+
03QLdiA3+HXwFPKtTSNHUnJCkXSHLd3UNcTVqIBjkzH683SCnoYyWifW36eKgmuD
9WNzV0nM6GOYMBtoA7bSlu83agLZ1kk6qUyIGWe4cWuTCuAsYnbLQSJ37PMLoBmp
9LEMhWfBlzvX17TxX3eTKqFiCgQCqj2LjYX+MRS56tQFiGYOHX3pQNZivT2ONopz
5dLM50DCaq5ioL1qh1iDCRx9LzxXPcWz8xai4pgqvk0NJiqc+/52937BeeNN5DsF
ZhlqIgmxPshnG/my5e00mgK8dV5iQpYN2DZizD8Bz+8D+RgpNBBi3ztcp+PjMbZA
w5sbjPm9001Ac3EFo2/F5g78469eM3yyVvmy5CFUIqM5yu4veu2b5oW3fB3KZVXX
gIT529blvD5MKy9E8PSiJMQfz7KLJdUZf0Vn/aZMAsxmYLz2CWVXIGg39VqLA1JA
QTyFxyjrzLcF4fOIe90pnPFDB1bAES/CqzRL8fr9E8gsJeHLEfFE9msI2G1fsCp6
jeBG6oXt6zwmKsEB0cei+lb3PgWR1WAJzgDgWsKx/4DeF62B/Zg8nRQ5Us+aWagh
`protect END_PROTECTED
