`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dlZte1p8ruG1I5arHPpkNFrhp7FMj+SJmTkcWRh1GiDhJPMVxz063Y4l9QYHlQIm
0eB9LM0TrU5jBglERneuIGkC0TyUa5IOxxPnD5/OZ5j+CtLW2Zo/76Z245E8eWNn
HQmiEk9aF54gBThs6WCWAt7SpfRpwE/0CumJdQ9FDgVxgiaTo0BwsyUkS25Z+oT8
U+RZFe6GSWqn2tjC5gDGwv0ov0Usrg0B2gGQZDrhsJMIY2HDAp4pFHCoL0yZUJ+i
2lTJGVciVxJnI8pT0c3uLfjbyT7KqtGWMIN8jVEMTBrj2EeP/212g2gAYIhjprMP
jE4Fk8x9iXXTA3UosaBEc761aMqica0JN3NfEjvyMKvjLa8VDgmwFd/b1HdoPJyG
THZnCtTqf87AvuPS69RVuEyLVzW0cfiPf/55w8U84cKQxLezrGpS0wZTPlHNK3/r
9TaN1Q6JcbAnqdJaoxAt2pX4LpzN+ZbBkP9ZzwU8sFAPLzRXiSffx9eVQHIoTMRb
TkyXMJmHjUaVYWUAbSbCBOnPtp25REeXowigWcoudeRmdHS3LdVoRQ0QKm1hmkSZ
nHv71r1V4rHc2BqiF87wihNaZoytRnw7b+saptLZZwlUlSSraEkhOu+R//egULCm
`protect END_PROTECTED
