`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PkYwjGQj/BDMubrF46RuBobphO/40E/YhrLmOOpDCX7+xJlcYeAXq7zbMwIONWG3
YVB+BoDgXudYc8P0e8YLcPGZ3R+JZQj3wzCOgP1JzboafN6QcmUK5+QcOJQT0HdQ
xyg5g0lsUppQ/VfKyn56yLuUkq2dZrH+LE8eOT4ZGhgUroVaYzLCqPuTMAiUvzEb
v2V63qpWlj34cp4f8eSbz5SUzOcwhSZUfcm8egmkBeI99GqBV8XnSxQbu6AZLhrX
m8fUrSdQ34/rsLrRWCB/PPf9CgJl4lQaRkDizjC9F35QGEXICpVgzTK+0cNlTmFt
scBAOX3sK283oz8YMigfEQ==
`protect END_PROTECTED
