`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZAzSHl+1RKL4XBa4XwPYA9v14KiVMbFLLabpsikvkq0VzFjS/0g653LHLfPyX9rW
GpOKgM06M8sBDafub7TrQqAFfl/BD6rXFFRZUg9N4i5juxcVCXuPYYAhX0ovJ3Qt
PkxXMoCq0NaU6jm6Ahud7ggDDTQSYWCnJKLxyF5vXMwB8mw7TRjsadQnUX9jx1/G
QaKgmXQsXQd5RFLpvsxm0YZKBUn1OaKskUzLHiAM5s8ox/rU0mOJui4KDy52IaCT
RjYqZYzsS4yNyCrbhhuGeA==
`protect END_PROTECTED
