`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kJriTBSVs9OQgv9agQPBfghnScNQn0xMCLi0j2yXJSCKpCgmhX4s2XSOeOSy+H5X
qmbGtfXc1eJ8Z6Ps5Gx4hru9tScWRIj90eAVHOEZGSn8L5OR6We+x8pcRay65yxS
9PQt9eKuEUkXxEJ5GdHBjLKfFljYuUU5Cb905BCfHS0L5mz2/hXR56sis9AHcLIG
e5jasJcr0i7/faqDht/fkdbpmMuCiMFy74fHPpt005hz/MnYBcm6Gh3qVr0ekYSX
OV8EtHPoB+T/dQlnoeVeIZElTlbgg/qZ0u+G6ud6xueOrf+xqUl6q8cgsR9oNR+2
OancN1C0kBy/PSynsJmnLg==
`protect END_PROTECTED
