`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MfwoC7+3pGv73B2bUyVVTLR3bSpidRFhpF2hx5kSOktvDhMQWZ2WNsB5VnvbQUb5
uOrwkgzOffyy6JiRQOvO1Y5cAvVZpWss46kfOFbUtLkH9p0kd76pXsqA5OZX7cF3
4aK9zP99LT3pXoOUfGH4nK15GrxWSRNfFr3cWm+hvNvGDf1QFRiCndf6i+4JuRGp
gE46IWJmT1+kwX01dtkM60WMao4XTzU5BSk11g2wJkjtt2uyYdJmLLixQBmrno5g
qD8MZOMpLDwEqGhSx4mMYkkK/LcdRs2eJKl+kx4oXY2gYj0gizWw8/NjQxvL5lPP
cekId+pqxe8GGsXPGz3nH45rpEyWe9FxG4vkCV2gW05lZoxt535zWMqKbTlqg/aI
up0MvbIdxSCT68Bf26MEQTCQP+p6ra+QI+F+AauBcOY=
`protect END_PROTECTED
