`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fy3xBQ4SdL25BAML2p+qFMGJaekA8GeHadVEMIOhLiPer1Hkg6/HkH82/Op/86Jp
AjzUhGpuOwNTUDo2WT1ezA8Kax14e6qp9f0UyYH7uWF2F72OKA0xJJyxywbBgJfW
cYHv5zm6BG3c1+uSy3t/2ZbbCB2b9PP6HZN1rEIhGHRHbHAh3hjkbX3eo9b2Q1EO
AW4Uxq4YpDBopUCLBqt/GANWWifTDIwMNCqe/nX/MRTTr6Arg4MoWdZrxedAluZA
SSmySTc2mpTvO0PbrApqn5iZuw1607U3PHvaYEpkNYeFQSmV1bDVcDWD0Dz3aAzA
7Tl7aCzRz6wsdJ/UUBAG+0RSZ38RJPt8YYnoCa8kimfzGgHRsqCvjIzQ5wCDPaeA
td8kJRpYKXuIsuseZBkNnNq8XQosbInQ+YQZki5zpHAjtsVqK1qZL8Eyt2eZbtr5
faE8cWY1S6+N1M3Xlu+MBKIElWoVR9uDE+6z1QSOZFTfSSb3RkBL7xW4v30LZSfK
+0xE1vpDVw+kH+12Wkv36mQrRJ9We0cc6bUDFHsi59W3bvCcl3zbaATKV/QihD+K
+wlQFlbq1ArqlEfghcGXbHu6XQBIAEsXmrxAbCMWDiNVyuS6xvKRWn0H9Oxs4O5N
HeCR+sxDF2mX+XCne5iAGsRvxce7O99Bq9nu7MYx/jj22iKQo0iyOrTT7RwuHihx
ObAXV6ajm54os/dWqnB2KfKt/BTQWPtYNNB2UHgm2KHPt+r6m3F0AHJifNMqmrnB
8hpx8d/LCCeGsrxfPjIDa7dcEbHxvdvFwTpSG6jQI5d6fEqTKv9EJgz0s8/uXzjF
HH1AfsjBan50G7IHZW2vskluyuMM21iBc4uq130NZfXdrPhB3Yr3vlH8b+QZT4/R
wugmMhVcpcg2Hoj5I4ICX9AEJBvLROiX4Q61xgusl6JvXuud+Yzk4rBOs+dY1ZQt
ChQXQfzxe03iSAC2dKsHbMNXenmuSoKZFTQTL/eAiQs=
`protect END_PROTECTED
