`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cmf1Q8UpXmfbqSa6qTIqATsqwZuOE+70wGhGRQnEqa6Ef2CIvMRf/fLddMS3L8DP
7mvzzOj6mpw7Vj0XISqDXJd3uQOOd0rvjoTwUpPh4Cf14cpAn+hchhBIV65sqHdi
ceCU3KlkejjzKad+E+fu2x7/FHZqkRWPit6/4AfK0sn35w0cqxiGRCE7z+wKKDIp
5jRv7ZZe+NEsfdLtt6qWTfCzbdOPhEKbq+iRF15nu7xD/GIAATuyXq9yyYaQQQHa
J+NMq51sO986UhgGxxfenqNQFuwDVQMElcfaV4qWT8Dvax5AVE5OrHU8H4WfMBtv
7OBfZeUfkHcFhhlSeiPX612pTh4PV2dj/DxJyyrwbF8xFqzZFfXZnh1GDQTdnc0r
3gE1UWp9bmgU0WKEivxR34eIVPMfYMUHynMEukacU45iMDgY42F+LLB4QXIqsmd/
MvmmTNQm07IqLegeMvuSH+s9815K+8BL1+WBM3KGUBQJSr55ETtnaS2zYm0TqiV8
`protect END_PROTECTED
