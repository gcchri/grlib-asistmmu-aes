`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zLPu1+SYtEw39bspyx2jh6vlrkEiFuiiqaNG2fT/0jR7fXurdte7fCnm1kqYPfQR
JTdX8Qv3mGivFWqEzorZn0f88klSAPI76dxPnBc4oXl90e7oJv9peesiEtz0zwJz
OgzpQxe5Z8/5/3VildVa48/zq6rhpgr+v61x0jBdyc/BcfRfDu6+tqnWJaw35adf
miA/oXJUV+pUCMJlDI4Uh2BGVdRQGzMyr4tUHE80JrsCUnx9PYE1BpkU5RJ3a9vq
Znjth8+qW304SEd/oeC3ePGbFSXPkpC99juqqb+0I5usb1gnnsCpM5UqnKK6HYjl
ITzCLnsz5wjXd0jH4gpXvg==
`protect END_PROTECTED
