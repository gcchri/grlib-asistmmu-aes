`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m0oT8ho/eEFGZKP8GVf2dqoTUxcWwta98O2YM9Opll4YLYb/YDvTPM9Dkwt7VPs/
gKprB9zlSg93EZJ6novGV49YpJpZZwf2XPt0vR+2ogPbx5LY5YMt9CBfFlyVvfWL
Jer+H6MBfXZdffAEbUSg8pqZO1j3SfPylBU378AaoyCSWehPGBEmL2EIGIDyCSLQ
Cl7leW3MzXfaPkzHu0zEbXgvw2k1X4ZmdOS2hUuTl/R4KPOkYAB16llNgDe/y2Uu
WaHRFtnvVQf9vycAKoviYAf22YDG/SfCeTqIfRrNG1MAQPRHfsP4xZYQ7X9GM7Tt
KtG8HHJLOtKmk2aLiivpCMM8WN/aWRT5ibXhQEVybGr3CdkO5cej4SL9GZ1UGgbF
FdQszyO+T6PokFWs9LPqwp/guZRi6oDFbR/91cxjvohbyG9a4NE2bteQdiuTOBTr
jzogL9DST3d8bNdGKjygSA==
`protect END_PROTECTED
