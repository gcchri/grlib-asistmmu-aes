`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oerPoRbmu4+kq6ibbvDJtJaYl5xi0PxbenWIUwKTWUcV68KwrDAONnWoA2CjefIN
P3jGAIrq73AavI0pqGWBUskRGirlXH3zEZjkmQX+MZOutsVeBX8la2mlk2tYVRAs
5wGagngvsnnmVkRUFD5n+eO/yfLvZbzAZJXwXUIF8bVD81Dne1wOVK5vLQXAszf9
5LQ8gWCt9URJQQyyQ9Ed8qzcCsJDQ59C99sCF4qplsXK/YERvYDWvnhxH7+Z41kr
D2c9mkz0iYPBYOkKnT10E9EdQ0a8Yic2OJ8jyMdBQpfpMN9wTbltZERz0mkCa92U
lJUjYt8LjJMjgltn6bHVipzB9aQM2u0BnWRiFgeUASL0393tfcpJrbEHH5FvZxxe
AKU2tU1dVThH2ToMKUzVSdkb8OdwSCfKzvkJQtwUnK8tOB6MXPoD+gFO6MY1NOlf
cRzv24K7FxkkrZVsaNBX9Q==
`protect END_PROTECTED
