`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GBI62xVczWQPQNPKhj/OuULdyLyJQ8b6Mzwozv2wg/ATDknFX3bo2xDt4QOUjSf3
/mStvwap1/t+SJpeUO2TgjAitIKbuqpVL0vVDnFp+xxqnB2c8Xp47NxzfKUZAz/i
rKE1LOb/zVxwp2moivqS6onYruKDkuwckzoqi5tFzZNres0BBgZIV7ZPVTPaVr3a
L6glNPKq8EUEmW8mTwZnoZwRIk8++bVWQgfOlw+DWExEpzCnri/c9rpz12ThpZVd
rDQLmOO1Y9HtS4e3hoDjuF9JqH73ebX7g5fypGKPDdeTzgq9LR++2QxpIRyzpV0K
`protect END_PROTECTED
