`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ng/IR8y/ZZnlDk2Q6TKNKNVQ3TfyC/FAVbQ7lBsvBkuGlHexcI9iKTNgbUyvQSbn
26yDgd7TmxVoeOTwvk//IJNDWaser6AjIy+iZbT/DUuoXVbPlZtPmKm1Vki2OWC4
MQzCDreGDhzanITjNdJ+IicVP6AAhfWgpKPPMeiGYfGGCMg7LBqy1polEgQ6ZZv6
kPUxmBFucB2i3QlmgMiVy5DfYifT2nb38QiKXONwy7KVssaJHykGsysq3XAS690u
DC2NEaznzAnaWEhSS1zTWPBS0nyIp0tkqNCO66WT7qf3xMx326fDiW91tVi97t7J
ADefzRt0nM2dg5ZTNProX5IIniYtw4b7fyJ/tszU6RbIlHzfkYRk3sqQ+W8+tOtJ
qSCGGt/7W4QS6P7wR02eab7Sn9iXYIajNr66nj4Zm2DN9M5PHAr8YtvFtiKy4eIu
Y4OTY/B0/3AcE60NordY9F1QxD21L4iJVmmBANe/demAsTUmIFvAL95sWcvQ4hOf
SxLIszHBYuB5OTNE+BtNV/onWlH1N3JWFTSRsJyt0PSNlxYdqDyT54CyvbHRXEDn
AFQ1ALieZZEjOcOx7mWM9VSu/qj1+bXz7kgOa6Z6+suauJOROB611XANRsvzIBAB
lf5XTAh5sCwEO1Om2dzEjGVVnFVHouzu3yX84Vx65yxPrTU5/HX3SKQxeaMzI02U
ONXQVlwtqsLV467JBgrYI93vDdv/b9jfyyM5JdcJlP39N39qAd2L5mSe3NXJ2Ck8
+uVXygIIM4n6BYymgdALibeG9pjIeefwDQPHy/iZBKUaKcHwKv0EJO1VmI1Prjtb
gMvX4xCenDc9wdhBj5ygRifY7qWJ+R80HU9484DtMKhWA3gwQGPiRKoLnhTST9yC
pGCDXww0iZ1iBdANlkH9zEW7LDxaDtThF4pwnKrV6OhOHBAnOQ0IBXWbMueQa6uD
V31SuIe3/g11gYUeL5Gbwwi9ukV+nca16QJxt8T2Hzglgjy1fxrnFCvGl6XkIvfO
RLrFc0logDq95aNM7aboNoCg/qUoPpzOOB11rimwiRxT67u8Sg9DAN8vR5RdhdDL
chohiuW35voWfo6PhV1dhXYMudsG6xmwwP6PKxQmzS5HMKRbMGYafXfxKVR7KxJo
I5m/CpbjOPcXbBQE+LR/oOztZiZzdp/CLbfrp6P/Xf0iSdFmqY6ndbv9gVyW7WBs
pz6YVX0O6k4KSL0P+25d15wkz3LcksIhoXU+2eCpiqbBERvh44C6wCfAft2EZnm+
9Hv0VGdWhm1i3XacQ3DC1DKUbJ0NukL2YuGMXiljhMHOj2TQomzXz0Xfz0xnGOlD
k3qTF7gDWTr8dNtsuaw40HTo/EGVQWfpCzahgklpQCaEeRELFF0sx25eFmddrStz
5vTg64QjAFO1I/Ba0QcfVJq8IDD8hfCs4ZQF+514amWnxIEhcp2QsA3HXnDWGhep
ghpnc+UHAcxxUe9Egc5FRJNtCILGrZn0Il4ABWhdljNNVzOcej03pfy6oTAHaFuG
uzpF28tNqq41LQuBkzt+e8z+O1I+dVHFFL01loeIFhTUobWOAQJcnEKg4a+hxJxE
qOskfAiQFjTWyof17S0WDDXdSdkhnOBWdYxVe4iSK/lo14U8uZdlDe9t8g6VTB97
LaWeqPW/r55i5E+TLOiMHhBjHYC7jDGjjM8XEjk3dd/2CPnMLDPu/P+pO+azfXfH
4YQYSziGd9Yx6jUP2MZXBnR5LoHdtx5ddPRcXIKxeYcjbwWKVKMfvvGhgkFL9Jg9
b5qbQuBm6KiqIS4gfUread9iBZ9IdluAlT+XoLCrEdt29F3w3DI3ImKlv4Zpqlvz
a5mMWmVvfRJ0qxlKklItlt1gz5MDsH0dwoR7Dji0rTWBjtW3UVTa2fS4/ogEXSHi
0b9TBKCHmtFi75R9x45d81bTwhZF9IWmHvHujD0G32QWXILWzv0QfFkKZI02qmHX
tBiy4ULQ2HQ8L6kRzDuBZJ9TeG16DcSWF1U/SprGkdHCpyx8MrSyOv+O0TpmvOg7
aW085Nf4/fM13lA5QXrxJDoDx87m2QQBx5RCsAxG7PQpX3sAHktsUhrNKAYfUl3+
AvBFsRVSYAMfIeG/R9jBF+DrWIV/nxDPraHj2Rn/n/D4xWk/0IH2sBy1NuLnVK4T
aPkZsvVY74rX2M3M0HkFg1+ekSLImgZeGyKLm5a8cuxjJWIDaEU3401P8Vl/zkQX
oAMRU7ITAYX6WADH+V3jTn4/ybCBMLDToBA9vC8NSfpajvtu4y46K8areWWdReia
6PqIr00tSJBgaLRiYoeoW8t4+szmRnb7KJtpFfzWrwvEh2H6hc+/rmaxvBh/KXox
WkPBiar1pIlvxSjP3oHF+ELifVep5kOCg9tiwIqeM/97pxZNt9AQO9P+aDM4d9+N
RCS+gZnNVZVfbVl94OT5Clwp8YvGgRPmRsfz4Dw3rGYN/Zp0VLFSGa3Gc/DG2w78
JZwIZ5zhKYDaNhEfGnBS71P2WHwAwuvz3WvUCbbjc256xY32OVJ3S9s2Ldj8i+qv
/evNBIQfd6dtnl1kHCJ0/ziZUrpBMTWnVjoOvU1GSeBO6t7HV9v1dF2LVJxbAYW5
wmF4o/+sYYtDQ8TMVDxBzWk2JV3HNbM29ossur/zgFB8ucSmqyhrP8NzCkxUk2TO
nWP07MbBCXXonQKlUZxpmnWfcHX8d5WSSQ7+Eom8Xkk4UcGmEfvFGNaP3Nas19Lx
MHb3gNaK1eSAN9/bae0d+eVpK3NmOLCepHpusDj5KyVhTiihz82GOhQQ0SEMHi2K
N28uW9FFTrcld25QthnWlXczlN2A38gQGDfYwZ8zpXtpJMasggNK5HCb541oqGIY
XHgUJbMolhqEKoFaouGMr4UnhcsChvfHIII8mwnxCQe7yTsYDAJZ+fTMFIG3BlmR
ZeGjI/16uLdOEpMWJIIENX8WlVh71O6rwChxqgEcu7sbSdihZlTTpMwS03LdmriP
4AK6FH32x0Wi/T8LV2AVLcqUbIT5xn3LoUAllMq7+O+yw5VkQgOagjr/5knbB66z
boO+LAV6UP6xYak+gkIQfscE5LA7c/wbbqwDUAzsb8aAiz844HpKm0vtwgWyccje
qqQKSC9PHcfTKEW7LuOeUnRW7gcfTJ1dOY26UWbiWIcIaataOoi1P4uRdjp1wUs/
bl8QX1r8TJklaeBQbWBUksqMSxydwjVO0AZBoRgog3uoBvurnzLYAcWt182PVdAo
5PmVyzxQoj+9PicHJZ4QIynKYJQ2rqQJfcrO8uuJ9uhsSBvuWA59mE5Y7BBQbW5H
cOX4Lt0BJFt8sPnw8EAMJDwIZyJmwGMGxLgsSfO6PqfwOOlSJ5sc4jJZzT/Q1C2Q
nbEKO5c7pOVpyzvX8p+rrenEQtSqS8KLNRbfIGXLV9GMt1Mn6icOxugj3m1wRq8I
g6d7U+360XQv323ma5nsxK1+Kl/BIupmBTeyVvusQ8zR0D3FImc2bmV99Tbk1uu1
QbP/3GvVzDU8NSjkc9rAQPiEXjYzrBJy7WId4el2nNFJjrKhLGj4T2aE6lxVr0x5
iSJ9YTqfVuMEDtw116e1vLoCli+2nlJjzavcLvrjik4MCzMb6Vx+VR5RZNm8UmGY
7q3GPr4ZXtb2TEaaW0jjrjgEUvCYfAmYGyhS098vb7MezR6Bm9MdX64vvXsthUfl
OgVSG8vfYzKg0cz4hNxvqiA5LWxhDI3BSz5628z3Hs+L2synI0mrMxouLqyBtrRr
MDPWgrmZRTgKm5a7DSDwb/pT+I0+WylfXs18T3pxUHgJC9igqjKc+5qO+/cU9eW0
mMCoXaMpgHJF2X95ThoGnwgkr9TtDBrcbhsvJUIzo3ol/kAwe+z0W+7WJ9D+nWuA
O8rmfaJwNCKKcNCIgz1paedhU1y6ixzHJXmNnrqqvrRvY2W/TBHNAJFMjEXQ/uqT
o39OxvByKzRg2kzQ+b+MzLA7SlwRYwaXXwHmAZiH/CNcu682w6JMRFNFVOg3XILu
iGLRY2zctF6e0qJIa1jlkziC1gDA9cnEhCB4S7727u8N9ECCU9bdQidPamQT5il3
z20RvtLrPj48kgz26HlzGAMJwHqNF398gwoOAUQFhlEBIg1KNbRZRFE4E3g92dZf
dUWauIqwPBDYTXa4ShmIoGYoan2NWPsEPMqiFoGY+e9e/Fc5grVgTstVTeSKSg/0
P1vPfevDlY/mLMj9yL7w+cF7IurK8NDe0GliJvFbrU/kx9cazdf+zWQsIcg3EqRe
IzkgXdh5bnOPSUev0OnWGCFJGyq8QCqED1P8wxzxifiKoQ/D2CzA5Zlv+ha4Pc+j
T4FAJ1bQhYNgrVsUgnW6gGrxrNfjMb4JIt+4WA3UemMotSAzdZMGtHUfzpysNnum
LVjvSZYfebzBZU0SX4o9FOihVgIrFCHYIZ7El9pyOasp/Unv193XZ0eXV/T2xMRA
lV1WP5yEaelL1aKMcoK7eJXK1nXjc9ebKQ4o4SsT28VPN8NFCEheYV9o34BthgLs
0EiorZnPVnwYQSEjm//2GYyE98Wz3jWrWeihdvyAXq/o8/MUygFmi4h2Srmc8bNl
0HqDiNNMPt4HjZMOyq47KTt6fhgLhY8YVP8KpU4QH/8TXR0yi38kBwYMewP0wedx
I9arqQSR1CAEnHPgHm5xU5jt/4CXpVp5obgDVBzK0DqjiXGXcs0vGa3sHCAdO7LM
GcSiPVeNz5gEcaszqZ457LxPi1L+8mzrl/cOaSc5BbzhC5ARK3/1JZ/2LQnSn2U9
CXm3QXrvee6Rs/IUrF2rjqfhnOu0tnYonFVlUz9Lqpe3J2q+vMweMojpqpH+CAiy
3OOGTOKx4xrRvGJp8WpzyS4PyAciYAtWvMR8ENJ0mEoOaN9XYryn+XxYW24GQwJv
3j5LfXlYUaEq5J2+/EPheBWGR8l8g5O20FLcOBCP7AUCt/zK7CduREj2JeJZgUIQ
MeKKWDMd0dyy1NXiocTE/s8ZG3sUUuQscwQtJxYxkmkoeVKelTxmOUhWFNmwqXUx
gr8vwwO7TrTpYoC8VNVPMqTHmQ8k47msD+SWwgtliF37VEkdqxU6Faaq12fI8nPW
v6o0FfvoMphO4/VZe+AqYMAbZ+eFEsh/N+IeWwclSHFs2VTHD3FYHiCtT3aRoNh4
iythnP12oHL6R9ooQ+WpsRR46BgTlv4+a6uxXeH8UOrcH7t76zOPB6yX4FM0OPe6
J/76Tz4aeYQ9quwgwFpnkaEs2QPAihJocxs04CFHRY6Amsyui4MPKFUjWKkMSAEh
4x2X7UidkFGIHt6yDnP7dv4ynevU3aAVkzucu3IiLjpqQ4X8Gw+pBAgD6PEv4jS6
0bPXZl6laJcNNYngUxSC37rNbtNThlhfdcBU7Go1CzmeSFrO0uB7eXrXyHvi12RK
WrboSlx48r/l42xdho/3x0GF3a/ocNkyHlaq0qztL4zlbsWlMeI3yqKi29K7OrRD
kPVqh2morvW3+15fq8mfnLNMTdgtlfpPzHOE7yVeWjlhqZmKfoxGJgn3mrydav1y
jVbINO/VZiJtmTIkHeeBgdsramQdcmV4uSBji25PEnb7/KP94NbpChE/jwPXAmV3
JXHTx0u6tPc/HPr5jnfDsy3nDiRMKeVVltoJ587bpjc7sPacKzDianLvcnM5nh8B
ciNRSPfOSUdNOVjiXwpOpQF/ANAj9TCODjU7i98Qygj6FLujiIg5/PB5DH5eovij
D9As/ZcUHtQ4JoKu9V1+tnAPEC78BQpoj4zg1f28PeSiMZx3Oku/lG5nV8Eqqti4
8mp9oK4UvE0fJbPWAMc5XIo8xJ13ASgGXEHaxSJAVCH6hTOkLoP3n5VM5dbh+Qie
imzpl0ok7Gcut4tMELjrsxPt9FuHjHyjnHjMEW+GYYwyuqKs1hOmClF8wp8VsSQs
re5MOufvW2o+svIE6E6ohIr4zKIbkT0/5+rPptXm+zqkS1hU3gkCQ54cmprQwvGF
tr+TgkYvNbohGEyqKqfzmPcLtzIdUsyOpjvfS7DKDdwmOHDvt9i+ShG4IthZgNVx
EZuvQNITr1kUwPsBlV6IWrED6GkwC1RSYR9ihlh306IxjNwvkGrIqS1+FIQtIQ5d
rP7oDhwyccbhMlkrvTgpUGgOzmTwnTxJPvkV+su5C6WOYBd4VxfearM5tKh4kpzh
L1955tyUGzMYdYAvThXous3kuI00ZzIUoNm7rJQ8WLRDGoP+lOBLPnOJka8JVyMJ
3zlaIA0nqCBaTHgMq8JDk0xNnr5ydWt302p1s8CUCiYD5g1SareyWvQoBKmbwhcK
oFCTGTzWYG3arMHGdm2yNa1lEYbc6XXTYWaf5NUDw0atbHc6JZrBeov2YEPpqMgA
9KlWHVPpsM+Zlixlid+wcTPXJbrkquq66aG+w0YOQDbGhLnFaD/hkM6H0yqQdBdc
85leL06nf5oZajHWj2eyecrMOw7c31Vz6Q1Y1AbTS9rat0+xwBFKkSN6yj4A3W/f
ardpo4+gRcOXd081YO4FlxGlcXkK4H5opV6jTWLqGB5SKQXqsV4q/xmYkUOsJmWB
6rZXmLiAvz6gTO+Nf4W8h/1d0zSGnckxvfkMVbVfWJbKiSRNnFunVQCTpFFlynMS
DWOjDcJoEWDgQs1U0r0hgwjPZIoRWBLQsBRxmhmIJx0uKzwtbLCcS6tUTCuAuHad
I6qZkkBzPjQ1cqd2XHTxSTIFyWl9Aw5cw/lPDq5jmer7y9tt2FoLqDW+Bk5WELgW
q0SZZgHpaexpBgaHOATTaILx294fL67yFBd4fOL5QF0/oBw97+xzeHuFa9CNkEUc
8Be+TrP66j9zmoU3YE5aWcbeDH05+zXn1aCKnzusm7dzkx6ajik75NYWPP0toOW1
jGg7DlnmBqv3s/wn0H0KuWBiyws83F8vXijR+u249L1YHm87PSxz13hejmch/X0C
mvctAPEvZ++ki2skQEWdnkfPvl7TTER378QmB5oj2g0AKkyHM+i8NweTJAlsGhfE
LqMcx3fQYPrq4GxMrPZN37yh3PlKFz0AZLyTxlhFOtmcCdVf3x4PIRm1ofB9Msif
nnxhQSqS0E32d2rz01+GrpTWVjFYVfrbix4FFlnom5pzOm6mhCjQ/MUgNMBtT7hT
P6v/GFeNWg7zH02X23thjnW6jI8wSUfavtBvi2yQ4HMN12ycE4A0NvLg/oNq/wSx
f94xxPraUms6SJLuL3Iig7fvjytfwF/Jz2j9TUqzhLrAjKe5ABO9RQ7+882qK8gi
Hjs+JjY6bi54hd+ahLVbIFcwB1OBVKSZLKJGaH9z7bYCPWf2qygRoLiBX8W+WbHo
06isr5tbCa6V+Xz6enA2AcaAsT3NNROegIaJ8Y+V8FYsgDXfkdxI1aEHNBGEj5tB
akXExKQhMQks1jNlW8FfsammxqwRSVgqHgTiglwvs5vHLVi8VdBQiktdVWoXL136
f9EOpEmVFzbEYTzwC723A8o7RTloVKj1lU1Blt374JgNJb7czZly3pWqL9wk3InK
gJLZvs1kPUTiWVBtIYJMqrVCaF8/T040pzELOxsR8qjumME3GL+/G+yhCGNxhLmd
phG6tf5DIVnAv13LvcBJdnuAzaH7bYiC2BXi6QGI79Ns65UoHHFuwZbEKO3AVDz5
mgc+yCsXL+1rXl1j7EMUVwWcQaTDc1YqybXgqBiwbHyI2yiYtXWW3jVTVSe5aS29
d6YYqa+vdn3a/mtNatqViEzYCr3G8Mo+X6XrTKcKsuF6WH+cHiWWsvxcwIfRBp7Y
P3G1iEb0ruxs7kMJzLEcLLzfkMSNjhdDjb1Kn8KPaMB62XC1dRn0CzjD7AT6efEm
00d6A4XDhfONJjsCDNg5OCsPK3PE3EaIt2WhO+YUHGyNIWW/zGQIXkBVVIik4NyI
19nw7/5bXD31HTim7tiyprZS1woeFc7hXkExqt+5nmvRMV1qiO0YUoJK9z6iTLTL
3PjfsT8JwPjuG9ObFPyDz/6Txprd9kjOTqhHUYqQnFu90FiaUd7I1uBgfEu03iuw
m76QAtmj4nQhO5wxI2BNOco9fQlhPw5Ob+iCVSkArR35K5u6D3SIdCwNGJLa9yIs
wkT5IXkJEhlk/YIK4cPON/zVNTk7s2ubHvRwrEDbX4qYPFI2wJ2JM+Vpj+uxsho2
UiSiW4bvPNi+qAfLseynb92bGW/FTU0ZeXohtdfpOq/eicNQEPhIe/swmDCMKDmT
Plz33Hsg+EArpFLnTvafuCsDya//58UkVukjdNdzjcHR5kDDfHnvZ7qfhY+QKNtY
o8YkVhCPJssa31xgFVGiOa6yorzFJEJFQv6a6iap4FDGaqTF2mXWBNSc8KnAGDzC
oi10SAlBlkQ9BnAxTKmRIutfSfROGGA5Tn87Ln7xKVj6PqjmnpTso6hZb0LTyDJf
l5n9q5JnTuHsxdq9yg70fE0OiedIFh8t8U45GCrfmhck2cbu/3NnK//2aT74jHun
vr12YKNrsBVgtj6jUPwaQ/C3cIL84iDAVTy60M6vgQvG15MLQCDsGuiQDAeFLOIo
z3QhFxvfUHeHsIhbX/610YSkA2KMBorU793zCz9Fc1mS+sl1R0RLPWwuea07fH8+
bnot8kbfYkpNrQXso8YH0ujwj6n3/1LEP5uj1ui57N/r9p5vTgCWGnwgJYt2qToo
W6v2UbCn6VrowkXOkjw1YKF5MFB+jECwn4XM9Ivo4PPlYRHuGOS9/2gNagOunoJ7
YIsOzKgj8YlhdstGeBrD1zp6ZDinaunbwJ9ITtYjlN1BiEY3vWEs3LvrzBmbgFC3
gVRDKGePkH92uKT8mhcI9ELkTK4Gq+oVSMsyo9TIDPxD7A0MRfSCL7U5GlO9RX24
o8fZoBvo40cGntjhqVoqIR3i/zNdOsgJfqYAWtUJRdY6O1uK4kn5ZtlEqyoZRXSp
/L6boedXfZidTUP6jQ0Bga8huRpNuRo8wV7U/5Ti8cGBtXZWNktZcKcN25rB1r24
gkMAerqDnL0SgKp3LtXgiEYEgUxjNpkR9/sxOPITgPM3Ypt5NZUQpnGvAKCTWj0m
rtaVmFQyQM/YeGUQz/fyOj6tJEG0MPVX46RRZ85sn4M=
`protect END_PROTECTED
