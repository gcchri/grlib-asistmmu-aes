`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rwk/T3oJ8PkXLTgObSBXYPwGk+ZwiK5o+1PpwhLwkQ+pQmCjxws2C/y8CjfeFCME
uGDpAqKPhJDxLo6SuKi89s7g/RSgeeTuTWwSdHZ2n8EOR8aiGl4UPR52WtWlhP+d
iFtuMe+0G7u6BG3Cs4AnGSARD17dE31gweaKkek3+mzwgslABFJCL93vR5KHfKnp
FFUskQxioI20KSrchbzNXYdLcx6Y+AtV+G6JM3TH+g9bjhgNd62XFkxLWWp/HWzq
atJMwOoUIMd1s2obGpmyq9sTBAXxhQwsdvdgatq3MQlx6XCINjJ7x0PYcmlkZATW
bWxKblE6NDH/zaZC2xlXwkSwnhwwg5SCeOP3tvqdEvbg2jYN5vvk6NnadjZ3o9Ep
xUaInUdS86ni7wVyQewqKu/QThMyGvPlCqRGBX1AVg8LscT+6ty3GjeQY2ICTJsO
FoaRX/zD+P4Cl/h6QdiyJysaoXgOsFpl3dUi5IooR/KxpLd2sQUQ0n4qMlhxFcGg
dgeFUdQaLb3YgVx7bnQNruyNsYFmsKJiCMGEupSGJvXPJjHpiIFS2IobPPfYMMKD
7tm129cWj+Xu51W72Qx+jg==
`protect END_PROTECTED
