`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2rsFpIApopDtRNbQafNwRQBNui8vqtdw34hbl67SPOeLoyu8KZ5jS5IJkF3lbmbO
MCJHIyEKUG6+gZ5abm4yBke2g3L3rlPbL6ufsmVVUqf2MKW73MgI6jmAqi65jju4
uCNOIvYvUjifL8rPCH49rzOWntoKOfuUDXz9QVqEfBzBwPplHeZlOACvnljsx6cA
P+/h5BS+5LBcPD3tEiLRoO7ri6Kp1SSse8pYQWm1TbVc2qP5/eDv+FZZavqLlJvw
v8iyM/m5ZtcuK0P7qHUzSOVoZc31/pduM1R4o2LdmH16sh9jH1I+vo8Q/kbuqueX
U0x/QA4Do3WEc2MSvlqzaNQAuYljp/AVP/9OvphXBURg20h0ltP5aYhGPL7ecyqW
Q+mY53d6Dwh43d13uiSO4gC7b1YCVkJvYRJAWYUyMA445sXojb3Q2uZ0d2ptU+qB
hXyAoIfwY9mtXgguf9oJVMy5gcgZS3JHn6gS8Txqw33AK/4f9AD+nNGGg3/wGwlP
6qwMrbQ1toleyDBiKK+sXaelvqArS4VrMh8sMnIYp+hQQj8OOHiJ0t7shAt7MviM
+dro2Qyy5g7F9wJN1VXnQgQas3jzHjJnf4hZ1MKPffewlDS20x+W/GfUbl8h75BX
U4WzyniyZ4ffeejkH/KyLDGLMNQchjXKQLcbJEUJkkFDNEWrZKTM2nyk8T6+jvhV
q6MvvERabLuaelPYfifiky3kFOS6VfQAqGGoxL0ihGAJ/PPL3CcXVIXHblzZso6P
lFdzJDKl3NJzLDCErddqXY4Th82KbnoYVX0aoFJ17wdgeolamafZsf69Wk4TOtW6
1XMo4xphly16wr6EPOGpm4ccGJn3WF/eNdb/Ugh2BU/OSBqu6GDRwL/7gf8rVkgJ
6IhcQ4EPrJz9CX9KcolfcBrjHgEdkC6sZ7yWrkUhdbKQWBx1s6wcXk4HRmHC4D/y
LREJrYjyGfyllAa+BuUR118bY0JyQeKWl/LZotdWUwUTxQEecY0+beHGExed1Tt7
KQdFWGbLPubdJJG3qTGqRbQ004ZHibU0eUqKlE/YdVvsmKGejytBikXnX3fZB/8t
pOmxm/L2hD1altEGr3XK3DAqcUbLP3WOb8jekzV9zuauGr8lpULbAd1wSJoOXIst
CAjGNnpUP6dlPCEngNJ+hLQtfiFr/zfn2DcJUAQw2JC3NHQShxAFrKFyY9/jIw0t
lO1ynbw3iIR3QyCJnvevnfzxtxVCiHz+1dI2rgNtsus3BMibT2ARlc8z/crQKN0h
3QdSrzWMeEWj5qK729mriJnyrO1IeCjOP++HCMkaImp5GEauRAzIwRF68Lnjls4g
yNiMhHsrX4UCbk45jH2u9lcrrcnz1oWTPw5hEx00eKmKZLk4Idpuq2601wGNm0Ty
t1BNzt/BTK+UWN+PlUImP92kczLE89HiOEtNFWW4HH4/i6W7Zsp+rbm16mj4DS/x
FOhqt77vq3ApxdBLyyPZDT+lofFFGu14CDpUBy1gZ8CI8ukHQ67QyDEk3KnwccFY
rWu6vOOhfu5cbVwso6+y1OCTWj3t52D5DQZUE+p24acX2hCARUh6ffL1UF8IG6gB
QejnfxBaWBKGgnoIP6M1gCbpMwQQ0GsOput+RcvXsnK/5g075sHyCBpo6QRg0J0W
1B4ueQ58Wme/dYxtNfJRaaxjmKy80jSxvqNvrC/DEePf7hsR8JsGYSgMkgBzj8Xv
Qpaio44GEc0TarErydN+7mtHfNO1PtYHcUVyQ4eq+4TZfzjdGnCxgqqDbAXkKIry
q8sQXPL9LNvnTvmecdwkG91mg0AKulQsVS2HizQd9fsM7MJKYw+m/9jXE6QDqI2T
73iJYKZ6Qa1kaBZ8LFCkqI2KXUvagcdXzZuMcwi8SIZYq1GXf33q6eNj6LR7dIs2
bQiGQZsXS6kvvhYPOW5REPxuJpIfDoL9yt3XUjEFr7CWpSwxChwvXOf570tyfR/6
xPtP8ReP0NI+NvDJ05o//7KNp5SeiAOrwxPbTgweSDJ7TLhnTH5Q+Z8lCQwhxfky
ofJOLAnpdSytgePV9ED98oHodB4mXLUpki955lgtrTJY699rmote/fLcWeJc0y8a
BBHYVlee8UXFN89iE4HIXW3ThbrVUDSUbZduJVmAGPqUCpyRlHf31qt/rdPz9EXT
7xuokCRT0GYay/EgLB56oQ0yVLm1qneC48JhkK1xzQfS0L8CImbIvIPPD5AfOx3u
iXnwkqZ2E9a6noe5cb81HnnF9xrbLUisDT6gH0pSAT5JezJFolew1KohLquk5f34
ZCDfPJERRZGlszgFyMj/HIUwjXknjhEybeX7sRYUclMk8UVm/cQzuRH9/oyXSQbT
/hU4TdRlZ0IXZrlZ54XmViDBvfDzazhmXPJ4h2WHiyvypC8Ru+Q1gFBSK0Yt+k+w
jUZhgLYYWvdJdLuh+okj8ZFiEzP6xXdho5h/++CKyg6012oSRN015/s3PAggTO3o
SzWPJWS2fSvphfO3wEoxbZYkLoAFh6iA/SDfC763syJSjLeXg6PqHdKnEYlMz3/q
6wy3+5q7rIM9MyZnQHoyPOVDtxk6YWIWKjDX/S64IB4f7Fsysuy0uHcaqw6U1bBy
tgP1xTojo4dxX3WQ/rK7l74Z0DZ1YIqV/yGoufFbth3di2lSxi1TDUbX91XLgB2D
YbXz79B7C+agsec3+FqJOTjcsmx/yfjz7Pk7gPXq4HM=
`protect END_PROTECTED
