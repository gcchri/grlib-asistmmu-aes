`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3c+9CIRBNO8UYsTOLEF+rvgO9ua/1nZOz8efTuZwwRp0jd3N1avRmAAeuaKdpg3Z
+UJDa5d+MHGzURrJ2dowlBfASTle/G8m6rvqXQ9rlMz0gei1mH1Cez/R6eZvyd6g
ekuRBs8MYKnF9ZzHAvsCxZ8bx/FpN++Cw4v4Lbc5CaZ+grKvNJl+uNWvVKRhsLO0
JoGu6b54ehl06g5FFNH/mE6KAShsZHhlmGK+ZFDLxLvhee95IqXO3W9XlR9gtZqP
75rGZsOAKSljeP0h6ihy2M17sf97YyachIb+8pAPrGfrslgI3PfRLBkt2pUrRX3x
LmqnlfpE9OWEIGnKX4QwGO219z+jT8/TmrFpt6cgSOqWKYZQmM51wiT4I8vOUxrI
Sewk+EWOjcQJkhCn8SFBuQ==
`protect END_PROTECTED
