`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UHXDj3B00WHp9pwEzO/aHSKLBJgo7c34r1Chihan8n8qJuYpWxCY1SAWN2ZCa33b
EEfokSQ9F4uXR8RHCRsmCoUWxHIZIHETrk0PV5AxheU3bPR8uq9QV0cpYnkw84Sr
5opnLIoyIP7KWgIyoOt0tAE1fNToDxLlnpHDMIUTCy/opGINg5BpIeDQ+PxP8nvB
EWUYSqewXUdcxx5sMJ/tl9Fh6RI+fgvbGpIF1WSBYgGGgeNfBZYOzZiaI+//GMTV
okHgPxM4CDS6G3xbq7qBFJLIVUNw1QlMlqYAYVjdPvklNYZqlbT+MUChmsKy3Fh3
kZBvL83xG+iUqTngn5Jf7EjlwfR3DsWufVzsaUKSqZMu44ZtwjJmNKqioLBItBZg
UGkrhXwYutMOmL8ZyZiOnjb6QmiTp6Vh3H81CIpy719ghaThtbJ68hX3Ygj7UfqV
485Daij/I/SUxE8biNgqpqUP8ZcKNoHbmjAkIdwE65jTJ8WmeyJ+BXmg/0KoOys8
zHVjbm3H3IPqBTpcTDDE7zhYX+fdftiz0UytlnpYnKpzPMN96BTv0U7zzNQ0FZR+
zIqbgCqQDdVeOD9/6GvOgQrzJpsNqL6sY8I2Ds/y9Ab7W2SJeCgFnfStzk8HB9Hs
LWVJnhQKRI5L3KKu7s11pjJu+UJ59f4h1vlCezk7yVF5gIJnippGmLwHc9XRwwrm
l2gumXz40cg5xCIIZQlOsgMCIklvuwdDHL3+YczJKjTJMr7otfxIcSzQ8zIbFUhK
LbMMqegBZzhykxxEKhlRU8ZpR1n9pr6Elu+MTeLLXwzAEYEIrWBlJKQM6DEqHMgT
C5EuOm742v9hM6o7xhC+OPsal6NRtAsohEz3wrbxm+Ss0N0YHo33qOi/AtSyWp1o
yBWa3bfh2rXONh+X5sqaunuUdzMpRUuQZ9z4QDDsaUX20Aj+K00kCdIDyuD6dtbz
GWbiyDPVgBZfEcU/IBEBNoA5e9Bhd2sGv9twAdjC7p0MQaeQ6aNDwcxGhecOhGIQ
6/u2DM5GnMIBkyVl+gFbkL99OGJtyZk6Ly9zh5aH/CRc49SZaiRBr2zhUKaTLypn
u8/0/RO2IeFUv95L5g29+Wcjs8H5McFNAQhhiEhnkKWzFPzpyPne4yEjJfX1uObd
RPtcjaxUoyAoDO0vp3SYGdJbeg1PWFkoCXdbk3iMhIbLEoc3YgqBxikh8lpVp+Fm
9jb3f8kcywq2ZZXLPJ978P4ag7bOFUVKED6jk7UogoSx64Kh8Livs1O8w+yzCRWC
FAZLOv6Ty45sdqA4N0xSCAiaSXCkys7K16kETgLO8r7M9h8pVpYme7XXHXSyNk/F
TJPSmmQWgH5guBPQQvOvOp/JxZQcEm9pWkoPoq/8rZVYelQTd9dULcroDB0N4ktj
K8mgVZ0Z49K5xcwmQw5LqaglVTT3RXK/jHDLbxYUDzioO8KFe+Gk5K5HiHu9hU0b
LoYSXyD7a3Q9zc6OkDhVltDe/5Fo2+cUR28MqtqafRX0HPt1jBrLnzAC8qgr93Vf
g9FiSgtM6+I/FKc5CAAPjk2fbjta8VGGKuUPJ+O5r573g2VJbzwnazuEEceSwzNx
PmR0YrhH5hvByWkxXot08f02IRug0yyX4q5WFTTzZwekbhJJvA8YjsB7qVubjgTZ
GW7nV9rMOYTlc1KTQF2C74vUbbUmbU7vOMDkXrmUBe/jdJROt48yiGR/mpUQLglG
pN3w4TDLy3s8HDSHGdfX6ca4NBIQFy/YdRRNbSAMJY3Scn5PtmDjpla9w1EQCHdb
EvOjCr7yIuuX1SKVnrrN2uLVLNkj6JClM6GrfBnKnpt8JgwTLK/VVCpjj9BYx90b
GDEGlf7xvsNkO1RpiNzDszU6QTKoW97ppcQGzX9/GyEXKcTBJW28+uNoOm3VsaFl
NfN9YUkuVuMPSdQMaV3ukYsGmfxbVZ8A/vJ1RFSg8DhZ1mX+lb6oUBYtRuJhQvj5
52Ty4kuBTU/CJPruL+QzNqof8nx15tkHwKFBeDtciLczXnsS/i8Z9semN77X9phn
hwz/6SC6YD2AbPXZa83IVgEk1CeUH8y3pAWX7rrQ6ngVCuzqHvfBChM2GIWx0s5W
pvQUA3iVejlUpL+F+0Olxwg/HMGfwnGRQ+/mkV4xqv9vARREMITTrZhBKRJVysB+
5wdPDNSGSgQXoN1YEcqyKOmOq5RzWCTnkzN7xmJ7jfrZWLppEO6PNu4kKfrMIoNv
Aq+TbQtAjRKE+Z21WyuHraop9frtS8CE8ESFYEd7ZLOjJhQuby162yo4WlKgHTnI
8R74A/HXAc6b2zA+m33w0FxZBu0yyTASOo+VjqmBktSBbceojJ4WczUUF/83wUpT
Rr42bRoZI/ipuPEfp47BXz1i0xqJi6xy9BkjsAblfp7DaJQGKGRADzHcPlYv3Pf6
lOcy0HjNr9xw3sHNF2F0BAVzzaGDeFThiikU4ztNvA6R0Vy+Xfci+4URUuiC2Rd5
LnlvrCmFoO68OjInpQEslPYurMykF6ECCHzplM+22dlHJMJV0mppRPzs4opZ/4AH
E0ArbhyDx6fuvDmPG51yLTO6owLAZkm48i3YGWRrqPmcv54PpOQaCG8kjMkhvZ1q
NOCMmbwLjxvLkEm9GBe3cnmk6FFmjyaf7Y1ujBXF98WNcrE9zfie98QafpihkCtg
cJPGOLYl/VoykAVIJv5W1PtFUMF80u6WiQmaOmt/qh9LzvsupinHPufrg++hOA0U
LO5lZ6iFZwzRicxWMw8MozW+Ktf+G6f6aG4XY48MeELiFWtStpbWEVE9nBTp6ugU
ORp8gnskrgWnw2Rrh6p0qCEvJM0uiueYU5gl/aN6Zw/b7W8K+r2bxgQFfRyDn4TD
9RNOVyrhuH/px24iT4XIOnyEEh/EsYyqN9SyH36YL1F42NszgbdhJ0Eby8J0MRPy
Ib+7yCu1ZqbgK2YBuhd9Vf8f79GRDnsUWX3S3hJzJxOQoszcSjvB+Jb45d3Kq0zi
45yyZM/pMrnaPw6mVTB6fLRh9UHXdu4haU1yFcldL4hUK1UDPT6kyvpvnymKv+Ui
gd/UlOjjIMNWTp0ZzIruWdZ+3ahns2VTgluoPeXAGzBTO6E//cmXVJxZp1tkWKOb
A3WVs/spMtsXI0yISRBO7r1D4utxN4QVYTdxEN9uEpR1Y5LCgUQldO6CHCvBAIMA
+5SL7vWUViU67+peSn4HpbTHhgVPtJTljL5g7bKL/F9/0cyBKze+T3O7qPo6YmkT
4GSmcBU/TBK6fGxRtyc80eRBUqATjoii4YB1DulZTunMWfDHxYaiJhVWR+OcKNM/
7HM9e5rCIcDk0D5j1eEs+HTKrYaLjtD8CnKhS2kmH3PGFXTwEutEc8CB+Q4lIpfE
gowQpeQhH7SAwWFyS3rpRTILILQRQ7765SLWecGO0HuMu0ZBqHcwVPI6K1+eVBGb
awG6xL13INLBhcgMdyFbX6iH1TfiIWbORQ1HaGsx/s7JuSBZmABFFOoX6N61c72y
DJKPHF4OdHyR5Bx4JmDABaMi62Gm14UlxEnQr+F35BDBQOJ9m3OoU3c2UPUn1e63
yOjuX+wqeETJwrMvtRonaHL9e/UXUzqTe7y0cmCQCLUv0KP6IH5jYh3rDyrcmvB3
euR81X60NWR2U3ShIbO2J4t3xi4i3aqkpgQUCHhn3muS7Zg+KSBS4mjhD4qeuIXI
N00HqKOgvvCi68a0B23IV8l2ifskRcyOgi2yf1EwI6qABL97BAVCjtjdwoYt760E
RjzaF42Qat9EnjAMDDnjYC9xKugGftoJjIOrMdnkyA/XLpFsxAbgKA5k9vFYh1W5
P69BAOku0fomFF7lT4Y/pdD4yYLgn+3bz95Xk7pzgw5dA1xTywCFY7LudLAdwo1D
keoIs4mJdcRUDH+RaUY2yDtrIcqHLEVbgfNita+nW+De8JeViIa0UIPSsx20OeuW
sUCVBhRSnVBgDhsElfgRJzbfbJ9vSULqxu/pa1DeUevz72WPQuAZ/TmCF3bobBJ7
P3hchIr7+0Y84ub5MD2illPre3aa3Zjjs+v9Khi8lhk6H8/GONJqxK003NCAzs15
kVnsJnBH5zlEaAkCMJeyyo4YVQ5IlcBhIP5Q+KCsztanlFyiuDWvTunF0vwgfDGc
bDgc55O+c0xEPSwXfZrsqUpb8yh3xvsd9CSLcQxFqGfVA1wAPA6VgSvYLu4dpe04
eCBu/j4m+aMeaXCo9iZbXkNwXrUPiXNNRxI/rifV5fk6BX0ikMHxBnkW45sPwjOD
qVin/sDZ3c4oZagr/dfcD6miXN9e9ZBUSEVDDOj8AHvBApAG2Gxx/30HcbeIEjHf
ZcuanOTPQ+IKBT8cfCPLMEnG5MED5OYuHA9qinkhudaXikxFeRYtVA8PyNq6U3T9
yjO8Nq2aVd1dLnNatwEMf8QHDJOTaWmUO4G4FzlesihDIznUWoocJ2LupyhIzBFA
Yj0OztLRGPs2gahLR9dgq7BXWWhRPwuOT0pgg5U7DX7IRi4Xo5xQsn/OOwFGQaKw
uIusSmDryjlS2s4JPbtwxKly/h0EhD5EkBn0I2J8HxsfP5HHJ91taaV/eTX9lwnp
M7zqO8VPIV17xdyZx8f2rgbEg5Vbg3Klkgko3w2hT5fVfueSsNef11lnhQfHakQQ
90JWZzxyRNPR5ijqY/RT2z8dZBUv1+gYcHr5LKU1wqO3mxZQ7HcGPRV8wBuqZykQ
SX59a0ukAG/bVRf6aZS43o6nICh5RLarytQdof/AU+yGYvfYVLTRF8Q+UkzdSGNs
Z74lrMVBImlytiyAvfWlvBi4BLVltDd+orvX9uRuIz/r7AOase4Zqek/QFM9HD8W
gAEC9HVF+MJnxKUDgpmsPhJgdCKx+J95CqvjqBJ3dnSl3TDcB6SgT0RUkmNcfpxJ
RlycJsIX6P+XeyCV4K5Z5m2mOUm47pv3mjphX9D3jqMjR7Ejw2aSuPhwq7prmWkT
dKnGefQLwfLeNf8TJhItgGeYLr37fEeYC5W4q0jI64j1+AZJiOzY08nyZirEa0AQ
2V6Dy4D3WR/HMPR9ZqQ//AyKuQm50hBhoXfQkPLLe36Mz6FnMAoE21T8IPB3H8Qx
BYFRSehr0+x+6CTVwTxFTmFnZNmMeJjUcc8FUqQ6aLauxCO8DLtXdO/iOb0nsDlK
hQnImXsE6LV5t5OnyE5Ilz0njWBAG2fScqTNNmnlsPpEdjDBZSpzhpi1ssJ/06oI
8KAPIRwkulSf2Pmm9PrRjRo9vqOP3m8P4+y6/8yoKI8S7DiZxrTjLOoXD7hzc8yj
IsCfx3DpUvSqAaAxihUS9nURZZrmHnrbsAdXpBExaJia8SxNhKVwLD643qDl3J8b
/FqzOqRny6+mmO4bCYSS7kBuANEaYbXwQrJ3iPS83akN75XqR2qNyTnru2nAUFvz
78Yc50JLCRxC/Zbn7WAsoZ71k86f2pu0GA0Hq/z64ZHVc0BQoG2Trk0Qaumkxrmt
evFAlAIsih2izdNPYXqbg6Q1UPr2LAEXWeTkOZKA63E9mPPWOE8cvQQ8JPy80dSN
eoVEj7zssEtTL5Z6D0jfoNwCfTTQlhjzmmnsbnTao8Ein9HfSN+Bo2cu77/TM6MK
hQSXcg/822jP6KSbXnYPJczQb3yxSFmdy9WiEmR1TGZm/Cgeme2YaVo7xZBW66Uq
8X5cVuh9NcwQ7bACRKivpWw92WUNNMsmE4h1ToVkPDrJ0vBfPycj8B6+4UsAWVqX
kxiwPgkxVkfrrmFRuTTXfvvPzv+J8xJRCL3HsQ1B7cuTJu2/c8RTjV7+VTK2/Wvb
vXWKbQBN0CUUvJ2BlETQ+Ac1vrYp6m++Qu3v/Jl218nMzQOlxfgLKpzPyqJrbKmc
1pp9wOg6fic4fOREcC9NqIZ3gK/YED3Se1P57bX4hPLGJYF2KmnjGGsIH2CKMMkN
8lSM0QQwspyWfsmvZkWd0hv981gA035w4Qu6PCiKah0cID9lyK0PYFrmIDXTuQZP
D5LWQIZBf296vFEbbGXrLahS81rHj2ZqYwfDgRgMQ7Q5KAm0U4BhNzIRF0wOPqAQ
Cz+8f8LAS7DOh71d9/7p5fW9TVO+RCyf+qO7r9rD5VhMEVBa/gQ6jI3RLMUp25ji
bEvQBD+swqWkMdMR1/HYQ2gntfZeUeaBNFcvCGfxO/Tx1vynnPvekWTj3JtamRMF
KLUdx0im4iK7r+YrUG+dodzobUOj+9YhEG0dw/xPP8OX7SlD8MRMI0hlJS5Iw8O9
prSOQCa663O0Kz7JFqHpNXVnOPAZlVh4jwCAjB9EsP027q7NNLYuP1EIOXPZorhp
G04sy5SJOPbl2gb/izM+GzMmtAfpE/KdpvM1UKM3A4+h/U/lnTzIv4GhTWCWoREW
KCc5ZoIoGPjdF6CJkf6+2jG+mA7S4+fAmDCXuV5hv2RLYI74Ro3YAdw7YMUEwoP4
JbfWOgmGI6O9CveFyBHS8CD10CO9ShobNGR7LXUN7fOu0hbjfwI84XaYqY6rRGzO
0gUa8+Vo4BLozN6hn7cpQokm02w0QCHCd4EsofzrRGz5aKWhpEZNVgUJk9rOlvXS
tGNI14jqXez1Oq9xiNjWfCh1jSCer7kay0jV62H/HPb91gCvv9sV0S/RjaRA1sHX
4QOsZsoc1fowAs658M1gK8i0EfAlDK3Ur1vOFl1WdLoYtPKdD0MZqlmo+NLNZkYD
HbZS0K/EAmPrVLPmDPO771V+G/XXgtJDG3rkkn0SOwg+/joYvL0ZLWsgT1Ue73FX
kXMdy0j+TT7ociWlWFKRBvrIp/ezBeumQbcXIfmXPKzvu4iExEkIxNzBqeGsCmsU
cRw5bRLN6Xc6HhKX3eLGYFLxjyw4/LxPpYnuID+CbX7OvPMUQBC3jnMNEcmJzuuF
tA1mdnJRJziruNUmNR0JnA5r9KjEPUbSo/3PZ6EMeZYqlTphkSNN3rjaQhca8n+L
/3IQMlt+jtGEvlHvqRWjyx8yCqewix2CmwwzfWrDvf10D2OtlbJ2C0dVSwGxX0Nk
XMyHaAqfwda3LSoSaQxvcOTKM2Bo7rbyz+mfgvBodjq6g7/OuSp3cD1vVF0HrNAR
bSUrnVKBAyw9Pfwrnl/97RYeGRWBi7QkXBgnH/z8R36lCcy0i7YaHRi/Y825j+DW
k2n4Fq1epoD7enRft2w0IVja8Hdjx6YNbXs5iIq+pgqPdNDZvgAtDOTJlTUfEJHj
DpwMKhLNepQzybBCY2l52h6DCoNzCXPf/d9ek6UQymOAeyWobKYaAr31WSP9D91r
dREkPKfRwGxl/ZsyoVp8aQDdh+G8LKdX8WO/rdJOxgrUADSHTardC1x+kSqURNkh
Jesle+l3Cd1r2EH+ymvV13UbJNtvr8b4hOLzKBMGKFRMXbzJcC8JjHx/jefP8CqB
v1fL7hd8zJj6Q4UVEIX/a4CSnD5L3P1hXB3ggvqFzmGu5/vfOzAYkpMRzexB3HiZ
uQQ5V76GuATLqYLMn4l2RPbw/WIqWWojzP+oPwyK/Ge8XaN/O7vnnglyPfvfk71b
D7aCa+ad6QFG1lS4UxYMG1IzcW+HwEQwP3xnNWrIMK7A0wFnFC+eyEDzNnWvYdpd
nKOoQqh0WoAutTYLLXvei7GWQWMYsjT5t3j+sKUTGdz7K3sr9zCwJ0ZJ5d9JQrFE
1hB4OflZbOLraWLHtabZrTNklI7aDEiNz3ZB+aCMrEfWUj+EyuEk5iFcrbfX/kNp
sIUDlxwLUpe/SzCisdH6uDtMbEmboiOjqMaCk5/jwJMNysemIrhbm/nQm4OGvK+y
1sbeixzt4BeD+2bVqutA9FHpq0T+X4m9mt/DaqfwvCczmTgBpFEON21tmn8eYjeI
jHYVgvo/Zqj46yWOI7iqVHMexY2BIrT+6W49mZg2etWqF3uPgtQviHorY14qGUSm
cf4aJz1vcH8sNXQ6AxC+FLlpsFoQE7uqxntg0E4CvEWizNl8PRoNWzLN5u7s1fW2
WNkBHckmtoHWxqpfYA9P7qu1zbEOaVDCRCHcAoMrlCgWJ5w3uFebW3gvr3+7OLFQ
0VhlKQXUWo/gIWEFaB6KPN1JYZvt/atyOB9Vba0nnVyQ6RK6HMoacb0oOwuD3zlT
EHxNoXDwn1ExhjbRWnwJ5Yt9XFiriG7POtTy9Mm4WQm/HQxRdpQ2iyqYEyP1yHvt
+6WeYvTrFEDbyE9OQ/AN8u3bMauZ0v/jY+/blGq6wPA10YnMTTJ5ZWUnqOaGNnfm
6aIEtKQyNdNe93z5n0JBRqT23eoGTHYt5LHr/ouAKRdMx94kzbtfHEHIXhXtlk2v
3/MqGAkQomFZOLLR91zj97LTwDC5rL22MR0Yknm0pd+puqNabN3XmvjTa+OdnxUZ
fvXZm9D7tm+aLMot8CicV5MLsb2VlsCQVDKqgm+iTrhuvLBg50M+valNjuBOsGrZ
PSF3Yd55+wQt7zE4YcbHtlD9gKl8p5+va9LeYW4FB+GMoljYoq9venEbhtzGi6I9
AF29PfAycWc+bADJ90pwdu+U/6z4L6aw1LTY3itHGJB7ZlwKdQdXksdK3og8M3Rr
CmBCNo+bKL3X6ZPUcpyDovZOwWSk+Kb8vLK5eq8JIALnty0hbqqVI2vu3ZAD3tNb
YillaOyD/2Jypz5ExB73Vj1lseGotFDqzTN3wE7rM2V7lrdK+ayEkxk2hJ6C3f+m
cEqqhLP+eVqx4qocM8lwVjc19+kltfS4fgCQqwaeurgo3qqvE+NWdxdanyH3IkL7
p4LYnuh+GLWpHeVWpEKI9q2/1wpJFpruze9THoDNo9O6+6abTT6jLsCWpKwC9BSN
5ClMu3+Om149ILzu27PbIzZSJ4/6DfTlGX86ouQ+6VkUvAiZGs/8dC/tB1hfa2hE
y+MHfjlu25k1WDE1tuVItQ+BilCOR1wFAkwOHwxHiY/UWTIs2cZOAG9twbi+q7nx
yjKcoxenLCWYDxUnG3t5PsNCtHozZ42I/J/XIpAtAjkV/OrI9UM/WLZCCmHORFOI
pGlKY8r/oAK6RvAhyW0zlEBanmNjlTw53yW8VurI1O22/kEhiurlrtMgOrY2F28X
oBfft5EdCPBiCiEUfE5AhbM2GtW5vtY7k0rsAfAA1pW2Mx5W2z+fUwMTWaeSuLjg
3xH9vEPB7nraiK9ev8BcDyQFfp103Y6cBNy+pnmD232Pnw/8C4okoI/keEPnz0Me
t3jqNtyKkPIPbxwBX+u8khUU3o/3w5jD32B8WV+CgaYdAZw0MzFsJYBetWI83j07
73p+v7dr3g+T5Mtmn/sChHhmibfBDFaay030jdXmRAbpg8sSGWVSXyCZpjNmyTy6
U3CnskEbPeeb2kKr0vTMmhGcNW4TZTv5C38wvcyPuoWWxz1chqnSzyIBVP2kjSja
AwGJXWVj7r6gmH4OHRmI2j2HpvWaTF4xibEQBEAHpiJyVMMvcYYCXsToQ2294Qh+
XZSjsbYD1ky7gbpus+xWOeNzp/3dTrClJ/SCf4GmayOGKf6kQfSh5IXumm8Kkftg
mdEU1W/jpMWbvvgpUC+292HhEsOgYqb0Pu7+m8KdFZrIm8dmGxf3peLLWVGsbToB
XT3KD7yeyReFttnJbiqoEDFteR46Z8nuKa4hZz8qv+ZfjutRw1YkrtJFpwhau1Qb
8t/w1V+IkZVk+w/ogD1RBGLYytQY0VuvKRBpZvlqLqc22iR7ZrKmo44ER2DtoXlX
UPtjQun7zlfyA2tTbz+Yl8VVsDFzaXFhcog+z2HvgDI+nr7SBNc8yJdMJlhVLYZY
3dAaW+/E4RS5DQmkyXXefcgFfA35y6PvplJ0+jVaIclyE4fgIXS8hRm0AjWgnTPl
NfnJvdx96GeXl1Ffy/luCqglOBkI8vJF8bctzI664eeSgq/LLIyzhMrRoHFYfFwQ
hOERFu3oc9b76kaj2p5OZY0sFWmZQW9npdg9T2vwPeZf53b9WZzZx0A0XORnhLdt
yru8rl7lzpirV6E26mm24H/41Gjj50MtVskeZCN2XarHUW4l/mEiHhaCNZh9el+y
fNosBdHjNHWzfMmKaFKNSYSWN5ce8CRE3sNKBMwjjBb6BEmAiaghe1R9zCERPWAS
Z2DqoQel/IYzy/IsF1F4men11i7WhgAGIj9ywmjgSGFh01hJptbNAxU6ISuFrtOB
cXnhIfB9XDXBz+lJPouIl8euFQ5cIJm9CgZJ+JOhKlfguf03ssqkcbeBAvq5URre
gh6fKsuAYEzSELFNHRCMQaQw0ZlBC/8jkbKYmLtRMtPexvdwNOdOAVzsEMH7+pXL
PZs0+Oyl1glwR+SktjiHGnbYzymFbDfgR2J3NrF32BFcp9soEmQFXVd4Mf7k66S0
zwI47P0w2+ugiaxbbQcCtQSHFe4zIAl6YrlYutLHygJ0NEX/Bax1wd5rIA6rRbKo
NaGZHav2PkX82UxoH0+dUU5H4B53AABxaVJqmdkAR7/ayqkkfEKloVQxEJfA9AnS
8QASH/fXcE/IrPx7oa45ZpN8xyFU+yy0i8U3c/UErafvZ3GvwIilVBZWebVQP5Se
MegEnn+X1TKdsM+6Gkk86Xh7rGRsPWQKmV0+jaSpdTbcHF67Wuf+YgH7rSvf3bEt
+HbZnZrCTEIwbg84rB2kY2ENienSG5+jJPrkMvtLiYF51A1tXUYDZ8WBYGaNdf/D
/zDWVgJ5CXLYXnHR+kbixVUt+j7osNSF+H5osVXYFgxdtFUmyR4BIBjQZELiI5rS
MPhWU0UWV1fAu61AIYpcIyAwrfIkx986lpCyL4amOtWGLoyQ8ogLzoM9hNPMzH2h
7JewzFOq3GfSaKIlQ+/AT2I879qPCufm8zmfkTXQhYnwseBgBoCoKiMtC7I5c5jW
az6rBRqmgIe6J+IbK1rIr10CZpBKYDfKRL04kTqjXT2gIt+MiFZjur5U+Dur4ztM
ocFrgExqWFjwYyZwGdVV0enhParQG75OSpv+N8vHNAWPdahjCZvCYGNWqXu7i3Lt
LG43Gdkwa2PLfUD3UBTQ2q4QquhOqoWdkZ6FwEIhhfsIY26HX5QgSpCDPmNUKFvA
E9LuUDV4PqqYXfMWhFTHy8aFul4RHnOaEwThx6EwaAEH22HAqcDGuiBF2Gi0WX91
Pr/kXqisLuGaA46VkPQWtzfjHsClEilb+EFw2QEWPWnyLCtE/gGEP054isWoVsgk
Aamq+wdVzsoBd1SlgnenynScT8rFrTx2pcGTcyOTkibJiWwajIcEUZUL2zSfIj6p
fsP9CbLraphyfSiWvg6DZkOhNC+W+DoVCpASkwDH8ncwtmLJSrr3bbSI9RT+9/2v
4COvTtRqF1sXMZ48NyZoiNKnm1Lw7pu2GOBdmWgTgxd3S9iivxEhMSe1/pip4eGs
iQJrpEuraf4Cml56IkKGCNPmRO/jCUAmJYs9tHYY9Qb5sN4dBTvi4NWGOYOYqBzh
LygZL5IK4hYUH0CY65aXGKQHcSufVuwHcogxdzpGRJU5NOrMXqIC6i2S7mj6X2qH
yOpWu3k7GgNRK0KQCnQViiC/vGkcLT2JiiGYEeNSctjN76nOQlOGy+YT/Bn+dZ/B
q4DF77Yqg8owCfWzoSWEZRIBL0Zq0Vy+qPiqQ/1FtsyzhHlMPmxvXep8/Tsdq1LY
8BJ2rbccl/Q6bLMLX3A9Cc5VBlyeJ/RgIC75KRElTob0lqr77KP7N9om7K9+92qm
EEZr9A1RQsNhuEljmuQkuvBrat7aLY1KO/zjPFnDRWuvly7qsUamwsJlk66pID/9
50vKn17Oyv3rZclhdhwhCeCmRens/m0DKoK+zqIWW0SYRVi0UvCfCyGvR99Kt/sZ
g1LtKqdxKMpwHE5nqK5AIlqZDdvSRcHPmCB7RywI9ZxEVl3fH2mvQN93Sg7tfeEH
Ubei25AvExFrrVNnyH/fB14zyoMxPwqzh1LAczaCdfwdI+DduLdDZekfAvDR/ofg
YFrYza4uz0t2+IG2/xYVm3m2LisjGlc5G8x+LFPtsuRlqsuNWDVwU37sdqtV2XXP
NvHVli1HbphWhO9MMUCghVsA7EqSByPRvU00eXDIHXnfS69lU/cuRMTfzBjeXd/N
MmHwsF+VSZH51ZBt2ke2FoT4PIj2ejWu9UPmIAawz0gRBZri79ox0y+PIFh22KFd
P7me+k3GLMe7uBYbgoThXVzAntV7x5rysxq7MRjadCpZaMhJc7P45NNWjd7qh3G5
BQjcjCezo34n0fidRS3FSzEfOyCwrompYh0enu4wLZ95rZNDzUq2zLZa5zVODLF3
S7k040C22mGtBfusJ7PJwVetOqpbg4JRHZTDET9C+JkpfqSCzitBH+xQuXQMtBlj
5+Q+WwxIbapgHgsL9IqF1dCEVmhSFvwLirZMC15iqat6x8Z7RID04ii+AqQlmZxP
ZOvnQN2h3Y3oY0Ls01hRp0ImwpL/tnRXLNB3Ar2LoBYDV/IkNc/risCiXGtgPrCc
6ctKzu5aifODrs/c7k7Ult5/+fMLLYDFb2k0A2OXtQOr3Jsg7p+IlzB4NFYUh7uX
fMUc7PM/CX1mDDP9n8vplSxiwy1qvbPolbM8sAyD+D8c5kW8B/iMmhVvsIZNWgqU
TiN2lHJEKrYxATYb6jzVJ0Tcn21nZdt1SGBEF6ulZgElT09B91wTRD3aXSQN2CRM
2bIuFjl8Fk68HJSsKgh2L+hiy5kqYvRRqSnjAQKVnMJAbni7cOarYv2LcJ0vkxBR
fAlg0JVkDOJdjSZu0Upq0HneWYe3Rndl8p2/pPonguet+IZH2TppyWFaNRAcVV2t
uiIictjQh3HUint7N5vnb8anO+Ywrs4ZoaMr8udD2Lctb8SKazu9ttRHBRfypG4j
RoHKC7oxQzFmchYPu4q86NA4NMuYAO3maocDszMav2w48qgtTEjwfeiVHifDgm3h
BSIpuQYDMnGKNh78mHNAnsEaf/n32AsnZ7aNOTPPz4zREivYkYgmqGHUHKD+DZ2r
OWHOlWrldnFrn/skE7Ljd4avPZGhyelgK/uqQURaXipebxnTRItcW4xly+CNVBlZ
aXG1TE0AZnYRWtsfZbdRw5oXSQ5QZWBWVhAGj39dYFqVFEhd6QWlkv9aj9SmYv4L
Arc4yDwC/6wNaCovGh5WSD0Ne6Djh6IKzbjbvIolRJTI5Zz2OZNlk6Vl0A+GFu9c
L0UpQXdd2EvLw0xCz3m4qubKN1XZV3ecuWTn99ELmC2Dun0wr2lMf1OH5QSes8rg
syNoM1KRjy78jiUROax3q0KzF8JRJFnESYmUzrk4U9eTiGEFSpCvDa/wzdGV/rBW
5aJ5OlGrgieYIJfNfO49156RMeDTjfaO/1I4fXD/aCE9EEFzJ4g9vnRV5bqK/WKU
tChsBYh6NZkH1wFONqsq3vryVpOol3g+Fig7cJWcCkuCcDmcApXPpj+64bt0SsEp
bOx/FhxlXXS8LyUDejsJ/zWSYR6AsJuv6NSx4KNEVDrOVTOtD/2lh451tXpXq9Me
Ege2AseotUz6GTYEfYH8v37lyiU1DNsuZLTb3loNNxLSrVEZuNZTGPnAnPun+Gp8
Eou54Gue7uzE02WfzXgEifwJyHx5D3il1osMMw0M+hfHMjAbCB44Cuw79Su+TGEG
z3JbUuq8uXKL2oveFyWVEBcAJR8iSE0a68dUOm/snu3fvjFe4JAu8oH8PWg//8bC
XOGamiE28tFrCjHlcF+HKi7tUimDMhRvS7PxFiI4nzoKty3eXRLWCXkpAJjJ15z1
CFQrQDc5Gfs3+HKgF6+70Hhl98GYy5QFF+UOZN8U2hVPdeNpyxdZVhNgY63RNL+z
KoTw4KNR8izT3aJMJiOgQnkNzKzWNfED+tjcku+wwmu7s415m1BoKXs3XfR0kKjD
Izg0LlxEuVce8zP6IR96djW7TuR65CCEJ0vVUG8UN2INqVfb+mfqF/e8JPOAfWN2
yFnlkmAaPBtCVFIDNnWuuQZfZsrmdpC17rUJiKr2GtDtthmb1wiTo4mGJWkPF8Ew
ljWlPoCoKHFj513NIGllHgRTWbVDoOohnIlgzU0eRD1I01XlGRFnMdlpnpMwd6Gv
+gl5yCAGJfttrpIWFjx/895LHaavJ6vO5h5AsIu+VO3P91MAeY4IrqgWbcU96hmg
TEKe/zEGTu6FuYprlHLLoagQyJKjHKI1di6QGEbi3xluUuUxEKsrrnR4bzNI7REI
H6SCKEn9r1Vd5fCOXU0U9CfkyqaxJIbIBN5cVOXePfjNBeLldXvFDKilLng4T/96
M7ShaSBPIBOV1wSOZuZdC8mtBE+mrPAKPG+2LFKOsnPxm4g87vP+175MM6TjyJZZ
pbovcJ4HcR01qKTyA74G389KgkEnDxNnvrkptaBPDMJF3UikU9ECr9YsGX7tKiCm
5XDtdGNhIKUeux19yOa15xSArnoQlmM4zT02tSt7MOns/dWSKTxfKJnpHlo3OAWu
hc7c2LbAOmjIQu4+CJPsxhCZigkKoe/DfC0QWN9uQM0mdgaIQqdpSPGHSlHAHTMf
S4BFRQ2z1T2nwHIAMefOAL3KA6Ubaw5BYWlseWY4e50gcvFfe8z1SOn1RfqhP93x
Yik/5YrCkvqLjD48+rxLe/92fnR2cTv9LnkqwzwM9BLoShpTIqYFdRKaa5610pR7
RyhOONh42SjkRm1NAyoU/maUbUQmEJpp4RSGuS14eiG3On/4Wj7z4kmyu2wRijQY
lzXVGQnKjXQuBxof+Vm8Mp2LIjdMBJidgFhN05Xo2sCC6tL7RvLGoMuK6wvii2ix
Q5vXn3nCOw4CdNlTlb73t1AyZbkYpTSEub/1ZIG8zcIgogE2PQ60nQDUx2vuUqVH
t16zy6r1+O0amDFmOYLeyWTEyh+IyqqWal7wR7hPZpZOsBG3DUGluOYmqgSmS+gH
V+dzxtT+O3RD+H+G6JUdDKC+W1h0jN/SVZxc1E14ewDy1STOyGPGwkN0gTi27aGM
Ybd6Cu0c87pI11wyVEaqVVxm3KuebkfLdQBCpyOxv7NPWqFe4l5FwDLDArPoUnoZ
swj4scLpVIWwrxJoXwY5ITOW+Xf1UMC8T3MK0FXmlX00PltMzptWZstR90+90WCs
P5RGW+a5LkQaYenKZGnP1THUjolzeWVBvJmOnogdc7urrQHhX1zWz+FcQ+qADdb5
XJUIVkRSPXP6d8iqZjL6TFDuC0f6y5q0GPd3eNs1CqxcIc09EgHdLT71mAa4qh92
aziqF/OU1owVy5sfK9L4s48V9qZbUSxEZEGgNfrcxSxtxR0b32yMtHRQVuDyHZur
1DmtwG+kWymH3h8XD0T8FblejADSDCITjlYGdWjCJB6xEp5fkCfsRkuD++gcmZCy
lKSYE9bVyvnS3KKo5H+Q9TWvd00FaqIBoLeKhyF8096AQ5DCn0agS0/KVN6dIjZt
e/gai338XhD1XvFTtvhca1lWWunY0Kj99mSdU+YJyFal25gNi7CDoLmmftlgl8c1
gXB95pEqSxpxLuv4QRoGmmTNbNiBIvy9vMvwbAQ/e4Uj4MjngJJTI6FCq/IbGH6G
IN3EXsGvAS8QFg6asLHwllDhmdCrQxMZqaElcyeB3bATSypVkyD+eEEVYLYnzUs3
bwSXWsv4XEaUei3qwvcM8z173u5ondKMZoJ+35EDnjp+W6iyXzG3eDxSbw+v/q1w
xSsGav0A0KzObUvIJNu18ji4HovyUxG6WbamrQvmHhFlYe1pLfIsVSKJKWR/GDsW
wt59aRph7ScHrV9HhNuss00LlKuB4Hcbwhketul7xXNjd5qlGV6HAByaYrtHR7U2
dwvlHEKFX0tsSQirutag/p174XKVMEG4LTDDdPbSODwJIrS+4PGePjQn3vqTI0yX
sc2M5El9riwJfcbyfCac1Ls8mEQcTAcDBcG4b/NYrFJ8OMYolNQov58/FbjrKVUk
04qeUKC+KG3XS+Hw57R+8twyRrw9Iy39taxshhbG6oSgRfZLpCFRkF+aiRmFjqkY
jrbPWxgAj17JKg2rJ6Fiq+YVT6FwMTu3BZdF4OBsLKDubzaCAz8yAeeff/lgU9aN
TF+jfy5dOB7pM1Q2mmIBqkXLiWB2OBB/4TSkw8p+xhSDGCih7ZTFSoii+xMw8tW5
gPiHZItkwCOl8Wha5q7GFMLbbUFlcQm/pXQXzXiWoaGR0r8tqv+TDB2YUKS42mdo
3RrCHxESGtfeqklyz4hnCNA3OlHP0LiZ5kz1ctzyNS9RirbF/5qwZZ6A1Xpa6lfg
T82p3GL7LQv37FpcR9bPRJABfWHZJGmGAWAiKKgeJqSfLVr38tIo++g4kYoGMJmI
L8eR7sG9Ge64w92fcbqZd3f1+P3oDMnjcKPZwHRHwd52f0D4CHbQ5YI+dBxl0Aos
bw/3rh7DolIDcmaVnZGfso3HdsyYxrqQJmM2/OBE7AMB8rMovz3jlHXhKcBBx/ev
xONtc/OhpDf8OI/w/jRFseToB4ehY/i21ranbhIUl0MMsj7SUA6+b6dcPoA0nE4f
sfa7yqezbyJMfBrLcF+MCNbjcD/Ir7SJfpKrQdt1oN1caBAooU7/mgSNHHgCpPWI
khTAyA01kOq19KcAhdevffRg2VNgU1s4AWSIw6FEqQOV2qzfQtKXpXjH9wuBFoG1
cL9+uShmkjd79DB2sqUliSELCvz1mEvMf979slXVr4jBb10UuRvuohCI1ChGsJlv
1L6EJIA8Lolrxjj3pay5wGeAw/rh9RW7lEHB45Mp5dxOWugpYlFjREk824JAVnqZ
BRTSh2UVk3YRqRSOMOQXSHPe3BvNsz8iBNf8GwlbNM3ftoQtI/BBY12bh5DIXrb5
kJB319biP56u9uH7QmsWv/4bpVfYfq4aVXQyBgowvmUaLLk8uXS9WUbE1XBD0h+G
8bvLvcZWddw/dB/xymALmPco1ozrTk8xFYjcAH/3ipQRXP5LUUt0H2nl9qToftzW
D+uZYSGcpG92t8XWHFFG1UQdbd3i6N/tz3Y2HMKTV1p6fjq6y2uqMQhcAF8kpZ7x
+SL9og5eyi7cSpNGAOXVTFHL7p1kZJoV+fhPBEcDDwSv7z/cCx/mHYDVMCs5oIIO
G/ZF7h1pFbDuSyTlrcAuBAwG2wVY2FeFgCnJfEDVOZw9Tw9eoMmO3KetarguXJHP
gct3AdZURszZ7JEhA7QSd0pAWg+wNLatNCIwlDsTr/skT7+NEFb4CWPXdEjhH2kk
ZDd6F2DYS99IwX8GU4+0Cr0RrNtqv7VCHqbEWYBoKLdEKuFapzRJuQk6JGVqIrrR
VM6qUH1WVScA543RoHziQVHFf6KWB7L5/HFtmsofwvGArYTXT1d2MZYJSCuZj73d
L1jT17hKlbSunqdvZlths34qa2eP8cKst1Mde7cQeBhxh/SogxEfK0iyNNdhHlom
N8dE2Lmwm8NeKZwd3KdIRzbYN5oBV0fS/gNe/ydjPKP03R1lbbV0eCkWKFIyaC/0
L3N/7dpTKmR6/i+vrSe5kqSbRBRh7M0IDddTSjHuSSGoxzyXeOkxHFIi3y+OFNTH
kZDZqgG7HGC5TYclguEwSz6cTkPjJo8j2vmYY+AUAGQlMuaRHbI4KahWhKuORCtl
UmtQMUpoKV2jP5TY9vKlYQSmehBOaYN1WvKe/TIk/RVFjUcxlPKc+8m/8t5WrDb+
Xe7zMZm6Q0HIacPVrZT2Mm1ruas7Hbwz7wHLrF1xJqgXFQWNaDqUPS4MDo6FnBLh
9Xzl29HELqFNnX6IgzHJ5stPCrsadfhGyeh0v22OunTHIk0Sx46wBSo0D50lYqB+
/xYUdPAlz69BYZpguCCEvNKkcfVkPUITVcGefexeI90rVr9bedmsuTpCxjxrz+tL
+AQ5gb7t14W0XTwqUWaEJhdJz28XhRq/MlNe8CkmpVakiWLnFyZzD0xakn2FyD8X
uPQVnlXcFKIXrviAzuQvfJGAqdhzZiXwleeZeJRYK43wjAvcllyIbSCHmFFDski0
vdtvYKrM/ZrVF3hjFV6S6fzqmTq8v+t35sYDn+sDMKXBxt1R9l7vKZERdbp1clE7
Qu693PQsWYn7czUN4wIhqspKyZUcvSLKsMedggNsZBlirD7cBijibPokyk3X6gx9
pSIvQiBfprqsctrkSmT+SiPRnwzAFCcQR2cXlnVdqM7npL86tu+o8W691uc8jHol
/f5DUwVQ1p95MOzGeQwkRBqrpJ4qk3by67JAYoH/sfOy+ae3qUBEbNHinnd3pUjf
xhNsJTLvw8nJygHWfOgqj5sQZ51XLYM6uh7pI2s7y5P4nGnknSEEgBkP34yYIhFu
1fPBAW4qLdN/Tyr7vwzfhr8lmmdUrNkY8OnFq686tdPzMp98ZkEk1l7w8ePaMqO3
TalSf739UrBO5JaOMrkmDqvZsbkaPTtYCQeq7zkgpre9uVFgS84mrv9PV6V6B1M8
OntCvF1OXihzg3lXcD7pWC5WTOQVCFyv2dMtRTp/QYB5iYWgXDF21iWtHnAPqwcV
F066vFMcYjol81pK0q6M7HCGGn5lW3HiUD7tGcJRNMDivFh2IsM7TmFVSHBg8FQI
FvSSJAyZFRw0IgWxcHN0HYK1FulsVup8HyK8lLlKjumOqDcMwTJ3goj2FgF57faA
xJzJzwiu59IIwlwKs2y9XOG9UBxeHx+zLeJ40aXHSAZtvjnJPUlVwabnBxzeYfpx
k+Em/2ZA+cBkSHwjcxB6GKpF9hI7sD92dSIsnWpxRlD5sKYWlpzvxpKuGEP5edIK
yvMaQYz+dTzieodwO1CuNEY4ivxWiQ6edbMr0iGOFfaB1yuuOYuO4M2kGM3ZUeoC
XyAdpYwSCfcZnzZue+cg4MNE3MaM+o0n8KAybWr3hlAYiX5l9UwkmoNyf13yCuli
llXJ1sdE9I4mWUREaNPt/TFGPDCU1bDqvI7wcDsUhO/qU0FnHHaRAjWk7zWUNg0s
8M/Bw92OnBcx1mb2lfbgyHNgS4YDVb+PgNU3jKhc1yfdyj4jm3/xj1g+iwsB04S0
nDD8jymX7/P11Cd9nJ41y+NcTV4x7IC4Wfeeqqi8yHgm6nQZUt95AObMCCZO3AfW
dZw5XifTRVxwaJ6n4FGK+u6aIV6C4Ls3kviTfW657gZhLqcEXzw1n927fwKE2r0T
MR2umgdmJpo+Kkd1lY/cCLdUx4hVVfuJmgFIgRa4J1F/8EBzk9OqVGuMvR/9h6eN
G8g+LEpOqcxQmPhQZyuvFHUsorcbpz8k2DqHgDKbvDg9H1aPFukSR769hEIVGEkW
1zMK/H4JiK3tPpjIU7H3l5OEh5t6j1BwzcR1ZU1EX6S0mHxrkJDe/dI/qAVF6fzK
dHxd5pnLz8He8GyWqxPEwhg4QxFfzBfmEzu/OLsuN+gNUm85uOp/aj0iex7/DdAR
VFTUprVos2n/MTVq/qfTojPauDTnVNhApBpuHG2SXmwm03zkjOXhkSD7fxRKkslU
gQCj9qAZsRrXHszTjL7GbLrK6n20bv6X3mh2G0yh2XlYv7WM9dfBubzfr74E7Yfc
MmOvRYPDE9dSldfSlMhbm3LXt+L4gxf0BKyJMQUJv4w6W/z4t4HsXx0fmvoGz4Mz
MfKgyfnzPurIYrv3ryMhh74YxpUDzzm1vLtS26dEeH/FGI2vi0YF4Ev0Ix3m9hVY
hQPGQ9et+rx6AJAgUtrR6/RbA4NC7GKmumaS8tVI+J/2PnmC6BzCpcESLNHsQDtf
jJd9+XyaqEyZb+PfUkFYmp8oorWQez4vzdPB5ByZ6GIp/P1qPq2zaSRFuft3/LyF
ovSTGwhA/NBpVNg0Z9vDvdqs+7leizj+TAWr191rC2xK5AkmQCeWZEIF91/IFLMF
oNn3zu0Nus2XTO0mSb2kA38jt93Twm9drV7nCwaHbP79gp95OKXKeh6qmW7oPVSG
4HE0WsHj+Qv5Zgg9Fo8B4omfVybSGaORx30LFMzTKr3a2JF5WNEA7wRFfaEjNNf6
18bdA1Mg/lK3hp2aCORR0eBbenUh+tffR7CAIGQbfRUKnFrzfamhp7kHXlxVQgDn
VHJWwNrShGmDvnK6eUtBg747B3XrrtEj+eBpcXR7ZjCef6E+SdYnoPr2qol6UsMN
6jn1J04Rcr0tuyD9W9I6UokZV5UEh5MRMBOvvHn57p7UBh/aAYr5X7fih8/XfOqt
vgHywUt9KYZR3uVKWSuyoRUtUrs9a6+ywMkvlJg/OGQSDNK53q2i58B56257MWPt
Yk20y2k+HGLEMuo47kwkM2fckqcxA3AczKdDANOjLMqUVjxo97Plp9aEZc6GxFi/
KjO8+IXF2GyohrbNqgm8aguJkRnctKhnztDTisCPcdPjalt1JEBMXQWMu0xfWQyS
QKJPqwnBTTVLTkFb1kszbw6bfMoAkD6B1M6MI9rtdkvhgohAgj2oshIhwwJizhUK
eTdrRnE0mCVZrikdcYHpk5AUe02XX6RJXos/8M4jkfbvxFFw/Fx7c0RGIFur+3cR
8JsSo8/8JDy7/yPQGslYpF/gujVs+q+gEQU9Hn2XFr2irYvS6aV6X/wGaSXRSECq
agYDuoY8mpcSKxlA+3HWk7cX6r5kCM4NuBqHvO/6KkVNZA/DqLl+HX3yg2WAGXRX
qgn44snXsteUlkRP2caK4IU9ZiS4hv8n/AOjp8cOVBPFF3tZMUrzhqamMZxsPOS1
wXiD1A3pQLceWpcVTkexq6+YAwfGGYgQQY/wVQws33Ey5S/6BoRehY9vXQXEMwkA
W0mw/LBeY6p2fnaP05WMX5liqeuCDXrlM1NV4E9DwN8tqdY3A1UgjFe6PwA5IXfl
g5mvDWuc5ZxAiBIZzw2eV50bZTzECx4LReMtnI1FbKD2KKJgv9qRCdGSBP1VDc/t
hnG9xxdxsOced2P9CXtPZgwBGkcFR9SoRJx9L0yTPQAhabfblmwIX/7n0gV9B3/t
zZpmNnzG0ez9/Qm8sUlAq9AyQc3Q51MPpex9pR7p+xL4sWVqvVOqYkIpII9dVR93
ESPfSKercx1MEN3vGqmNX/l29DMpUUfMOiBDao9MYOvDHR+3o8Xv4Grd7QakGXBo
zjtHApQBcQQMfGt+c6bmFIFF4xq5CtlGaK0k1/aVTDF1DCXRqxRx5TFNR15ABfIh
FM+OiRmKwJn7ETqzpYVQv6dMKlIDce5MANjrWRroi3Sd/6sCQNd0yOE4AJJXGtWI
4kpd2bjd6uZrgYN3CkpNUPF2LJ1dWINI4rGrEdgYPInvSzbnxhhjV5VMTKvVd7pK
eK4neDxIaMA+Dor3D7TqHw7/7IpHgODnVwEOt6BB3Y6Si7xmaOebJCx2MvWvFwU5
1dP9sAMyxEOegwhwIPfNs3kPdClFpAhfdRPgxIDYIq0l2ev7lxNcHqguQ5GNCI5C
lYs9DoMogs9O20wnKxQnb/Q3VSHxnZzWL0DFTcbfX3TN8mY6r7i8mmlctUHVTzWM
gZ9ys4ACkqHEPuRKk5kuq+WI5NDDmGwqzHJ3VTUWhbLolF2MxZWJlEBJYJCPw+LM
mxaELPxj42jvBYFisixsIU7d+mVAmbuPnPeDDzBd6gQmjwv1+A8byU2ZIvigAHrV
g5/LswJifq20ADjSgS30alwpF97l+idvcinLQmOrcgZ7fjRkOc8lKHmuyXx4W3xz
Vauym46ZbBwuPTvBjzvqoD2hFSOtdy+D9Go1uV1yjIKA1TyoaKgtgC1KSambm2x1
rEBkhlr8Lh/+q9GE1O3wIgwy1tzIsLzyjybsC9rURDgLmMcxuO8NuuAfVnyLSqDc
ZNnQt80NbVA7XqXkyZHlH21jo0zao/tkg34LNgMB64ar7Dx8TmFsHdihle6EN+Q2
C77hjp92dnia+Sdnl/Sj/+KfqQh3iBBioQwTCmE3IMPRW7tMts7rLuG9/GMNDC70
8nFGsEufW4m/BUK+HD4YakrqDUNyWV+MSyPE58Yw0btJ7S622b64E/TF3nQrD6gN
NpuiU7SMzuxDMETKQsAfKvP4W6dxcPmtJilhJGdsrUyVzDustXL1bLHgVUrog0hl
zw41nRYXPp7QU007kf2EGLqynkbbMIgOk+2eME/x2ldSQLHnDLwbay8M+W7gdUoR
f7M451MNgXHlnloTAiMHyFyR17tyJiI10n7mdHBJglqLsyJ9RphY0pxes3FiwIWG
X8lJEmHDLVfNJszNXwI7QexJ+q2JGl+eUcKjJaLOQO52peLqpgzRKA+Oc7h26T4u
/1OYGRNj3Pdl8D7Ma82IQETdq4Xfz8G7lV2pxgHPX2tSw7YHrjfqUs4zGHUOhjaS
IJI5jg1MS1oBMeKDDjLCc+qzasWQha0oPlI4pezMnwfLHhmnn/Y8LJLA+0eblz05
EVy916FTxTM4aWnFWejfTMRhDj8ycU3ifvfnHpd4ArWzJT4/6T6bo/SiYRQpqk6t
fs22NGhwRvUJFXHGTYakDDmnINq/U0yVY71T3vGPso9KgRm8KZBr9Of6qehXLe6g
E0vee1nSyEzPyVIIYGy6d0oGQjbxAWYVEW2dZR/xHdQutlPJYrfMbdbmuyTFxLaP
ZWHZQ6t5cuh56fYuqDAEWAZVyx98cfAJ4PpcWrwxkSH3utuoOgAHUFbWshAnntOf
UXGindvRx+fwsMNlNAdo3PXzk40815Lug5wtVhyOenV6RxNsV4gRFHe8VPdaI8Mv
9yR7TiP3l63nfmqWx1K3l+5jgcrp2PscjkynJt6xW2Kgd7T6Sybsc2K7t3UyATd9
rsS0LmGLt6lWBXZejSLZe5GK59ndNEfTZdZvIKiJGOQU2ZNoMlzGrmK8gCzjoDcM
aGQRo7Xai9v/E4mfDJemgpZUirshSb0/KYPyLKKYZuAMnambRZppx0E6PKSezgie
DJuAaEth2mH9T31UjQ2w3FHlMZ6sSRTGcQvq0iNRyruNw3XSDZou9MbYKsOsFZo6
jlXAydn80E+B+nEv0O2h+e8TWzKhHQVm1mHLBwTCGNvs649ZdXuUp0FMyGOtTChr
s+A6VtbPuzDTR9j0D3eO1BUk2xhuwK1Xw3GgCsaAxAUXpT+uBQYk5CyaDc0VnneG
o1RSH8vOOlHMz4EMfaFcFovbUuULVWOGurU3uiXugCP5fsFQrbM4KGXGI6ZEaMJI
EpC3AzyklJjA1l9U5s/ST3ia0Z5501fDhg6+j2VuskRSeyl9MXkX8NNQiExvFgQL
pyuzmTqvoc9b/d1p8RVj3CXMiL5h/wbzAlx1nQDPew3Saa77yc2QbqGypLqdG7RD
AnhjKwAN9n91SP53+FhHxesTgYv2Bdi9HO6MiJK1Zk77xql0KpJ2ckRBDyOEnY3J
Ug95VUX+nhZ5CcobvIJ3Kak/8+OGOM/zro8rhxUTD9jbjoKXrOnrqFM5jQ8xoPw1
iRZwdURyctU+l50quxE+TnZLbVn4z+wCgwEIHp2UzV2RxB7ioZYUpLm42IQYxbT0
+6RFlxpwB6gBNBJrsS7XWCW+lKQbCGcFQyV66Dof7znXtQ/5eSRAu3fhrmg8R0Fb
hx4y8Xmgg87yGk1UnYy2p20tCSNCV6YWTWSzsCU2gjwnT/ntqQHicGSb0KeDw/Sp
FSfAgkdMjQCRKMs34dd/wtuU7udFeCln+xn/OwdRX3YTTmsZasHhY81KY9mSHfz2
bmGuwfpyWfl4AcsvIsO7JPSYVEGfX8JWfDa0HVzxGaCTKYunpaYXvpAM+iPxJ+sw
LHyvSaNuvXF41t0uDSupME/kYGMlfHRMd3dnDOe0lTMQFhxIsQbcKkBoCveuN96T
vv9tFvVakZHyR5tmfwF8bt/TWqf0Pdbo37xxZ23REsWp0dDpWv8H1SobmlMUvyFb
6tTiPFqdkSs2BjIldfH2O7hLPc3LpSbUXBkhDF+MQAm07W2bxqwOT86uR6dupoG4
4qJ6h9OhbOYDrjRplrcxuqnljn0qwTHLPs+7o0AUTrvI9k2IhImSdGq3ZvodEyRF
pI1VPnKlbTdDTMgjBbdbRXO3BzSVpoBxxJDKZIhIEOcvBskNSuwhm+vjQTk4amdB
wW1nThTmPhypny5xXfC8Xm7kedAfodcdUjXrMp4X8yWqliE0Pvru/h1Rhmt9i81v
D/hChh/hOV0vrf6zEJBYm/n8PhuKPZUAEEIs7Y+ZE6kLtmoYGrTGMiu3ZU1yZXe9
pd6rJu4scVZtyPLG5WPKVqJApY/Q45+bW7/XYnKIRD3i4NZskg2oI7btnKtFGoqQ
MdbPlTLo0qmXTVY6w8llBjaop31BSIQrdeE3vElkE8WiKLu3GwOlLzsM6sznIb1A
YsWA5vbjPqXZEcSE2PAmGnktfhdM+okLbmAw7OHdQxX09EV6b/hgXwW//aBCjYKV
xSJEFJt6Upk5QsuAsHkvrkNj9oGGgRLBh5aVgyZWK3c2Vt7GJqcbAR81FN9v7o+r
cVainh5fBrb8vg3ANGcPHy4c02bENg1UuTJmG0dlvlatAGqncsB8s6J8q85dc4sS
k5XHgdZvt75hsdKckJ9oCsOBUNEE0nTrt+nba+tRk/qaU6PomB1FPdfgtYQ/1NIP
egcsiPwRKkMqaWjGARApysU3ytS+scI/R4V62kB71oVpM0VXeWH1QHyscAqsx+Pb
eX/QdGGVlsUVbXkRKnnIa1HdTk7K9QKV2o5nW6HgU0x5Ij9ozf/E+taoyxtjyPCX
gpktZVCnDHu5Unr7pYN2evveRwTHmB+4QiB3sQUrtIuElHFK9yHhSmI5+ZzBRu9L
ppJ4eLzfONuqUoRkg0SwqxpKKYKr4/Mj9K9UsHkiYADBihL5SSlYrx6Tc3QAwAG4
6poti9e5DGycQxTM/n170r5se07IXcQWzD1yOlRLjT7OZdTdvEm9BLKAT9/VXtgm
nMh5wQfvMPjSKSQAVDf2hPfHtUWRA3m48IbnpLT/+5Nki+ktxWZ5auLnyxHT2OUH
e+nFLzVcsrqa9gB7OykakVDjhWDtZcEItGQjSqJeIN7AkhYYXmj6i+PUqDtknzRX
CKbvWjYO39TQT0yTW1ZEAe4slyXuXH3PwHXh0EP6tq5ObduBL/vGyYL5KUQG/fh0
1LBkgevKR68s6NAoNMxfp2Dok+El4Wgmt7uIeaevyWbCpqqQkrjjcQbZXUCnBYAF
okdcThbBMupoUqQ5L/IhISZcQxNSFE2ysi4Lv2D5sf20Hj3uOZvyRPhXpuD279DU
lIBB61V8wL4vCA+lG3TRIIucRhYowCKJGs1cKR+q4quWvLSdwPXCYpH7eiFUmB8s
uyjoNqJe0fricZXo7KFKDHo+GhnYefdNUcXV2jvcebBxR/swbDP1bCx8UVVfCU9H
9ybQfgV+lIxGPve0vAt/C+C0ylxTR4nd+Air0IxR9id9wghhb+q7E8poYQVsYksy
s7VdGF9ur7LZjzqi6Qei/ObFPOvbmpt6ORivFbmNQg0I8T0kj51X2ZrtcXu8PRX5
o4n9r8Y2EcQN5vXgUPhomTsponOnKyGcZHAKDzh4hf9w6JdT8LcCEO7rMVAX1bv+
71USsJcmRnyJJ6fphcrW1LuT9zDUFU4v+VGGy0fPJI+LeW2oxUu1/7NGoY7iAjAj
yhZHix3z7MUT3QkYNjyU6uGE1rO6mHyxtx0J7T3PETinAM1IhjPpkSc9N7SYMbXH
ajYMp2e0kDcBRtIyrfIOwv6Vw2NyhlYkg2gVhEnY3IaaAKhRzo+lTNmZKiN9b0vH
sS+g3cPrOVPqd292MbDBtPJjC0fWZ9o6qEEVOJn29cuyN2Ckeu9mu116nMehXn7S
jCq+3V5ZICmatz1UPFSvXD4rUeVniCCIRedFkqXMWtkuRDwpid2wtF821ymploLz
xZwJB6iSmQ3JSZHKS0Eg1bZmItDYGvzYqVdape5LiyJSvWSXkF+0FSrhvBzjhB6H
OHTd/FaObTYAoTg3yqz+7ECSPdDYfMnwOgB+5zZknPiUc8eG6zqjPiFfp6eg2X68
jksK4RyFyfk08684ldpzv20vaE5vNpBRa5e7JEnnk66R3Ub80CYvsunpFSgwu+fh
2rkiy/U3A+pEfBiET+pQITcV/GoBQmqq2lir0oILuhIRLDYaeUJsRmJwu5fBm0LA
CR1rmUdCEtoTsMP6ZD+pImLwNqaEzLMcffhrkCIN+7S555e5RTRHr4nBhp+XH0Iy
dj9xZYdp/ELrDq4pQ7j0D0n/+6G5puv3TnatuKZfeZ26l0lhnRNSJBz1GLZR2lBI
qhxmezvmfWPJ5OH3hGYDkwpGTAV2kwq7PgMHpVQx00rM07dDeOnTBbunGtBduZwy
L3/oEkvr+1g25jJtUTxVQMvxtKDM4wNUVvB7SM1nONtpQUq8sbOIMzSz5rUIsRiZ
rVnno6wIMeVXCZuqomiOSpRzQ5m+HeK+RdFc8U1KcXGHoCU7vcEV7dptdVj2TWra
Mn7hlwiX3wKbFqzwhGNwF2a60CbwyaMLxsMKbooexcTXlLxf22R4PFu9tzL2xZhd
6lASUe5a22lU9LD3MwPsBGbm1xiz/0cFll4ZtpcRWUI6l5NfaUYmKmI4+rhjxsX/
esJ+UICpgPOXsR2zSCjdFKD8SAmj8U0EfFHcz+pyz0w5gJXzdvFd/hgUShiiz9Fz
g2r5YU8Du8Mbu77pRe5dQ613cWTLKJvvgIyBQQmiGL+7fHmIlWe5Xk2jEmwzaXrL
dFIxmnPylxidL3+qkO1W4kjFuZKioFtXls4xgggtgBSsH1odl82iGkPlUTRA79Au
3xVdkC6pI3B1eFpO8JfTkQm5f9NPBCo6QlMeDoa6dIHN+TfvKBeSn/h2pggV7Wvj
dLYuqa2orHXzSP/R3s6K5qGa5RLHFeQKCAyvk8+l4UZYmVXBsgEX7xcLC7M41OPY
BiqJp2u4W1RdOlXrJzKdNTUtHT6LLhEzLw7LjHP1DhzXFhRTYUzWp11CzSOlfowz
/7ztuYD/s3GQsVSwqdEygKHCA/Q/wVgduAnyaxzdp8XxYx0FzCoKxbJ6UXHS5myh
QhKIUP9Qw9HW+3y/YsYHczRaQK3rjr8BBjUg3QVtfgg4+ATLcbgQyM0uyvRV44ig
IO3IVPbAUC8ny7rMlJvo3PunT0kDFRFCMSzDu27dXR6t1fTh4vl8xObGFaY/P446
RMzAFX0Y62ra+L8uCTP0d23bak7WAcXnay157qIrgYDYN1d+5Z76/TZnWfjpjIA0
kpHDt7rnAQMviacrQZkZu2/0IYXyHvddgMwvuoZtNfHDcnKp0z7vzIhA8IELy1Pr
TQ3W3MLSpoceqXInt8zSBX98NGJTuwRobRE3WYGq1FzPfSvBbzz6U1rIlNViTuji
EuqJYewDbPn55EzQ1dVX9bLG7KX54FN/T6Vvmu5Xad+vyBh8477G7GcftLwr9E58
1m9GKLVQYlSF1YusBU/YP0z2iwvrdAaHf/PpkCbfPCBm4/MU/Laav7jZZyNwG/dj
tM7o1nhWPF4f/DpT63jtPU918AvliTc65sQYizF27BJegob73D+et3CoFC3bM4g7
5Cg1gw+S+KnM4Z6SPZzVT7jnzpzd0g5Sb/t6/fA3xhjKzhfpY+yMYiO/PGEi0vWc
cjXUEYlOGy6+9OtUYWpE/zTBrwoPxW7N1oNOt8mKOf2uk8p2JgSXAho0R8YM1yui
ZvCbanRmPxf9esmg/EYyG13qShbq8fo8pkkBJsxqnKsm3kVzBpdXjG2nj3yYgQXu
95Qt58rq7j5tOlXcfS8sWr/GB9cVgg+EJ/nyTrTF1IEhQ2NNCryko59P7rG4YVaU
Qrdx5xXbKvshsK/67I5VrtKqBBYP9OEbSCd5sW6inK/TIY60yp/qiX67jHwsnXRv
aioVs6oruKRfsSt8vPo/mNbHX3/k/RLiJlZV6atlaMAjZhz4rZ0NE+nvN4NpKgMT
WyyGdslBt1P/tggk0kR/UqH8lS2fSVEDBpwOyXZjJMExmaj5sHLzJnsukWP+kkOm
tBRMMDpcWvgi5ijXH260NF5xI/ST+ra8W3Qld0cy6SVY72ZUDG6zwuD2AwH9k9Z4
pEWztHIck9HscU8uWd2oEfE6tqftYVy+w8Ael/v54Xess7nZas6LWGXffnhem5xY
h9hCOihN4KA5NlOS8WgpigrA+aNIeHrezB6fGLLz6sFSnfGVrqwKSzNwW3O09UVW
AJdzy9q0JEraFIxsfy3HLJWoGpOGDwJre8+c+tfzKsKlzrh9lhO4yNYIkIiFZ23T
qdzOCK2RrcwU7lWn8NeQ8I8BU6jyRGoUx7bb+LXz8dWesoPxRivlo/xYx1pZ2g0z
De4x+lrfzxIrsYlnagcdckveohN7Oz0Gkwr2QmI+sGWf1iQ64U8+IrozuLcEtZGG
YDH5z1VwjqluaPKVvrknKsSXF5JJtNYcZTGvG3EeZSHg329pdfQGJ5/Xu6i/2UbV
rLhKQrleclIW6iUOlvhrDkrJ1JJRemDD8jPXWqslFha+28bC1Ns4jjKOt9nY1snq
T95rNNfqZUCeyquAYVvPl3THRFttTDNTMqd+HQZwJOwTy25D3GtRuBet+uB3cnYW
4Lj4/hrdUy/80qBK0yZ0RWCjHjAwGvGJXS9kZeUZOuvjCvxSusZE+J4KiVwIBHT7
yOeyTlWUysRYaXwj5BZm2Fr7azsWcq8Zy+5GhAYZH4A6YIIYHFSnh/1COURF51jr
05of3Mu+uYKXwdnv9v4qc87ssbgj2jxYqT2bI8ekYunhX2A3H6PvZBXBmDNjWXQo
n+tqydx6YiTdo2u2eVWPGJt1i3BG4dqVyx8fPtmrrkFZ+aEq8JaU20NW2bpGfovJ
0Xi4/1h4cqSRAGQgmNKni8RNJLn2ZExRdQLvyo27T6X3NGFeJtIyOokBF+/WHJuR
TmYyoT7heL25L7dpY0H0KWECvMlTCHHMy/SrGq0sZs5fs7WMP/F51SYNWru4a692
iyc+FthKIS5lZHWVZuzudr30qFJ/J8W8Xg+nkDQGb98nK1NCeNrvSObej0udHDC/
7zkNHHDNpb1ox8RLIDMhZFS2Q6Z3a0NQR13qo6zC5wVFVVh56iwAXDV9rekjOobm
nftvVIp7XYo17Ns0NJN8w+2dWucanIDcQt7ZgxHNRL4sHCwnhz65CabpffUiomG5
4E9xU2Xjw9SwhODeHegE5WCc3PvH6YfHa8IorOOPXEwcTO+SUNJtKeH/yPEzBRB5
ucOCOawJWmTtTB9z4562tCgJvBzYxb98r/wFRA1RU2/mDW0w28xjqv88lWY19LQI
qMY2tHiob67ZWLays4ORlbJfVdQ52kcewkzTCfS9odOHaGJf9/zI3IhIsc/Uf2NJ
t3xC5h9E5s8f+cX5t9wn8my9HJaXTB5cV+DKjo5+2aPoM3LzN9u4BO2mO7zdSp4t
qbrogoPCYxx3KgD0REdfyK471PxE+b0auxREOSmz32u4hE4hOny8cMP8XBW3Hjb1
tFqiAdMzUty8p+6blB5b1FPn8xgXlmFXlojWHrAAWbT+/l7KFPvQYy7g1DY4pLZr
Vf/QUJd99QKilJ4w1nRwMlQ9D+MR/TxBgadg5GNKUDnbXv0I53CFlpvOObtbgo+c
ksOl6KW/Z4EwNqDFi7h+S7pK4BEEK6isbI0ITZDXJv1PRBT1R754Z41PGWTQ4By1
ywpsfiESF4GplmofhdpFDAwOEwRju+lk+5/fqdMaSfNNoppurxUPmJ8jeax8bUPE
TBhkGSzsXRKcjx9Ofn5uQyQo1rGWXpShHfSLXawKJGPtTIZTnEVmkdXbap3KvhRH
TGWLLHvxBiX5+0LwiQjgLihNmQMh3gvaydK/fp8NbP2jpNKFo0jzLN87yKyxM6LE
8kvmOfQUpBKwQddvFjXKNApCcfEB8Hj7Eb754Vu/p7AvQxKkbQg9ZIjccgR+sO2a
Hfemnmd4HwRY7nw3aawgbx6JL07zhFN6dX0Q3wgN7EyIjRBFigJQ7poP3S2KeewF
WjQq8CAEUMIAM/1V6nw7eLUZfgM7H1MnwLA9b9HbZ4BjTp9lEN/rETQ22XxW2PTz
ulx4EI+/7vmCmIw6KSI8p1ODNE+Tq1+0eIGKi3zWt0zEMnAgcUPzMGHBG7q51AuD
A2xk0iYploSgDcPFrpPRnb7ReVc36FKvvR8LYTPqv2HFWQioFR+6D0tPFecdKK/+
xg/6K/q+sgjySeSoA/Moqqzzux8CiHHqRrXbJTPBaZ0SaeMPs3V+HsxoWn2l/YYn
f8NhIQRNarpiQT3086a/C1PntOYjXEYo7F3jhH5VrXnQO7LCcM1y3nB+QTuFYOcM
3snT2Cy1UgG8oUHO9q5RvZOWRYUuDAVnWHwUaC0yBTg2udGGz3Gd2gLpK90e/uTl
FOmR8jz4/MsrJK6zjMBnVCNHJ7rAPYBap1bNVVFqowR6F9cHmujTRKMdH7PolLgJ
EN/NQNlhISAsArkEQsh/Gm1LbHfcy1Y2Smt0KG+ju0QatIkx2wIzVTXrcogkv//n
n0ssUsY3Ef0pAApwKjPZeGjg+csBWgCYuqrrgPPztmqltKIsbL2qapsl+U1ptDff
yVnZl7p7WW+YyT9V2a3PaqO0eIfLZC3opP7gSRAmrOtf6DuwWBL5qjV1rlUxcOX3
WRj5CKYzbhhqhf4L0K0Zp1qslqtJEJPVG8DK/pAeijnjN5VUoa905rWPrgLWANwG
O5EOFxF8U0BeuEEwUqMT071fNT1/3yZcbnh21+OenQbq2aeOxkI5nV/9LH7THYMe
rZGX4aQ3Dm3tURp2ssbNtt0C0rmNh9KWrQYKEr26EFZwhZ9hKA5tw+nprtalM/q8
pknHep1yOdEXJMEdrlN9cnWLL8fXrsyKVWG+Si50qcZvicm9gZND3DfNewJvvCrZ
bTLKQHshNnFocW+3u4zhVw3NzxQqBYwCOGOg3/7IxOMe0tTLFM304mM8ln6PiUT2
sb2Lc30J1F4i3BNpAtCAlY/UFQ4s5tiZuRMXpqLtpegaYfa1H7Sxs1kX3lebjfOF
OQ3fm3pOTGUUEplrv+n4/VzV7i2J3j9cYTtyzp7Mr5xZP8uxt/w6C3QajvHSqUiv
JNhIbrzeQhXEIgajKgpcXNX+0jzWfSIaUua0uOo4RiYZvv7NLQOfLBZEhUMu4mlm
VzEiS0t/b27iaOls2iMzRAcpRWAtEA57Aie4MlLfYJXEHWRwUBOXNnfinXr4lHui
WAf/XzlRjY7r6wuQt0WspbDQbBsQvp+YN6vim8F6bBvTaAxnHjVtBAaj9bNwpO2b
RJq4O0WB+waov+sq5oVDhaFvFEnH9oZzw8Q6HBUPWIo80Bv2RvXkuYyHEfeTjS1T
HGv8Ts8OibI3H++zjrzwnwHUHkAnOtxQHR/YDD+BEjdkZbC9p85O64ogtDDXjFKR
ySFC1jS+7P/R4x0BSg1LGu4a2AeQ1QukenaWSq3AQO0eRu8CUNyuxa+dF4mqIih3
3Hu6i5a2PsPCLmCdKGybb1nm4M27Fbih+kVziRnYKxDJS9dVwusuKChOwB+e6kLf
ZHhv2S59RDQ5giNDlHBDfq/9g3dvL14siBdjQIcSt4EboBU5s6FGET4bhb38nrWa
rahtwSXPLeIHD0lk54kVy28aAMZTbwl0Ib/QT8BFMl6jjUi41jR4mGsHakOEd5hK
gFlWsIzFHeTcx/0w3d/QDh4jw8c/gfesQYyQqmuapfTXxmQiuxYgdMJgaQVawKAJ
QvfyJX2mjnzee8fqSe6LtJeLV1OKzabNWAr+QwVrEmpGA9PJO5438HGa07GioyHA
URQIcPf8MitSDLTldPHdFpZ/Cay67HVH1KiG01yTNkg1FwlcIgg/qSQpIpwDUf1S
pUUUO05uNW8mUEfH8Ce2UqaVPaNEU+6OmarRkZXwqu2o8SMuszHy744xi1MwUw9W
Mk2vvt2AV4OsjW3EAkJJSBkZif70r9L5VPTuKGbjnrag+QSqJ0J6tmooAAQZ6arZ
KeOivw6M6oNDKozqUPCLayrYjKdHg7Zs4FnoPbqPZ9VDMemkrQb/roLJZqq13/0g
V7hFr9/hxDYNWxLTThUdB1TXUc0AAJAv/CGUbs7nivmJdg1AR1+uYvniPFlhkE0c
gAZtXGbhaMJjPx8WVoHpI2oZj0E6oE7wfF24EaDWAWwgswLjg2U2fd45gTdQ4+RY
yy5ARCq97dR3hXEpIMLQ8MVuiaCCtkSBcKiwwOJ1+VKdO+W21/ldgVcFgqgKwTjI
LspiA0RmdKSvouaHxPFGeTKR3AN/q9zhIIFghabPm9bCgYtNYIquJ+DvBTE2mC4m
UA+Q8B2d012WuEkPR2JkGap56t9UG+eihr4X40V5FAuu1IRuz6vIfA3P+lxSUtuM
iyTTXDlcNWaZIIs0TYvcHJ2ZvFJuj4iTNETzJaYeX0kjuyUrhQcsP27x2UAXkoNT
J4F4lhlQAcrBGok21S5vaDIgMurH0U5tivFUNiTPwJmtecnnnEwfJ+J2eMu1gTCW
16uCuGQJf02RaGRgCXtWEchlutP6Zx8r67O4tRf8jxDwt4Ls8XtNwSqBdyissRnh
USLvOJ7/nSMlDVgu+4A4HOpoeXIILfHu0wnS+DL4T5vwqfqIlixrkUClcNZ1Iy2d
25txSEWlznMgy3v+eDd5iiWItJ0d/icMAtASKTgz9c3fPoAE/SrmTUJpYT8B+r7U
sJueWisCMS/4x/ilyesLwZY6MCZFzLIion/g0LpWXXmo5D7yKhjusXihbeBuCneI
9tFRnhBSj4z5D4Wpv65Ro3XLrllkSeGBJp1XSsxixEG7ZGDGc2vePPJh85WYK804
nl3xNeNZuzUPDq05EHxkQzAVNFXDugfb+xBchfSAHk4fapEkKs44verwkSjQsk3g
7UX6FsfEbXvZRT/T1Pc8LDxqXcxhDNC4u52SFMjed449k4zyj3SUgfN9wKoQt5Be
ZbyjDAflU56sIHdMZUXQx+721OZLRskYaGE42Gsp2B9HEnloj6fZ+bbeEnXEQJhW
STAibZeL4qWhJzIe3+K2LrVGIS9I8RzP6KvZrU3mhjiwsoVRUJirixWO9gEjtWOV
LelcHC0eBWHcZnms5RQYzUvXKCbHD70N33hWwADWQ/CJDREaU4hVzVDUeNgrhvc4
wGWzCKlAcOnZTk1SLzo2qOPX0Jsj1LaSnx/Ph+KNB7W3FKrvbHH8n6qksgNW2KIG
hsiij8TIrk4k9aYdN6FN9ZOJ2eh77o58VVRW6dZjCH+OL8/ZaDaBW6KhrV9ZHEJU
S6gtuVkm/qjzZMFEh8wq9ctiTIhUqAgn8CTY/D/Il2sV1ukz1rj06fy6IaDC+kTg
4S6J7PVPM8FZc+HzeAtKipYSLYpvwuUTmnf+Fqjg0zOZGGu7ytFmMUuuisOG2ysJ
OWM2x77IWCrQ7/RykW1cGakL8VP9ItA0zA/N7aayRznJSsG2C6HEdgJj6YB8je1C
KFmOw3bhN4Ivx2h0avmcPzzBZWH8xcQ8zWcl3Lk0b0iH5pGdy1JXx89TkTPw86k/
l1u1/6MQ0psc31QNOzUUdW0XHUIfcuulLy2Uxsx1swota8KbUxxF0osrRW2IDrny
xFhELchFq7P1jBjuuu+5m4vW9WS6Y6fYVPlpPJhhFwDAJ1NejITtaTbOBU5oW8MH
AuMmqnaSZb0KkEAwTTv7wFdxsqughcWCKYOkZH3mZos8U9UBYzAUJfT4I0ifiFle
3jjP1HSeEOkBwZmO6dnMNoP1WjZ+ZjWCG+oBU404ODWpYHuPwEUVnQueWU9R6s6Z
RKaKABepwEekHtS8drGf7pIbqJEQhbXXHeND540mwNA4MAIrLvpGS25uWxZjm7Xy
NAXN7gVGN3um7qwvwAryBVtB2pdLiwUvl1gxxfLCKRUqGKpfya+Znc534qicWqxk
o9Uc8ZVB//113cPdGLyaTltFUrUXuQoep2PzeMFwoBTqMf26VehUFsV9w7jKKRAy
ix/Uv9qRju1aX6ioFEhHEmaJ0CI0wLnskZwsyxSMyBDM86xYbAxp8Iu6jCA0nqGc
AVDi7kAAPFAzka9IS1snM28fAr0fxrUqgXUY6H57EVKfmZ3SPA9jLpfw8SoMbtz2
dfey2Dn3xfxmC5rYYNb7p5+5Y00jOVNTv+v1KeFoJrFjc6JjxYzRXo/k3+DVkXCV
mis/wy8/k3ALV4YH9e/3wPW737py3vFcU5qphU5RhqeYzfMdGRDEw65V6uxJQ9fN
ulgC3WqRKRbXUWyaj1Ai8elcw9CrCxDGQVvYcJjpAKVCOXeHLu+MhWnsgK/2xLEJ
inWm6Gdj+Ps5voyD9qKbU0e77SXxLTYmvllxQWteeO87d51Fwj220eoEe36vyK2o
49JrS6kpGOWEZ1ikwkguOmvbUrDgiEZvNf2WhSyFEFRZnqcRodyH+L5aa98klieB
P2cOvlsmkr/X421/ebkAG2JrYT+Qxu6pgxTF8JpQ3k3YxWEFbeKOWWN8/TuDVnl6
7qiyS2GeFCQhsKJm+nrHMw2xSo3T4mbqg6uRCsS1Dkfk2x4wkSXgNgHHd+8LfydD
chYFCimkMTtJUA8CAoy4YExo9mFcsn7SHLrDUPO3P+zKkft6lPQCqZodykheumpz
POd1sDgNCgzgyrs8V7d+seN5LYp7kRL4n8lsVQcD3FdIu+mIXIrdfFzzq5GQw9i0
Uyg6PAtasSbqM+QyrqeF4o9XAr9OHC5kD8c9PcjM/V3/69jW3KDJwY5CF2g3fzx7
fCGJl9ZBkjGmqkAWoLWNYtUZ1foGWD2/tLN/CPl7gqRAi35Q0WEoPLN3YT5aZa+3
09s4tLAuWs9jH/A1IUN9MZWvjt2EhIEpfZy/KaUi47RSVzdVAIwOEJM2RhWvM7Az
MWrZ9rZtFDyKiMnY9pr/tW9JaYGTFLbytRdvXauE9E1O3+ShGQQLr1jKIl4bWH2g
32LsVFvy4Pmu5MBT4wh3j0iDYGMCv9qpfX3raKPO6hMeGJlPd5Q8lfX7VgbSWp/F
8Dt3ENWxda0kUMmfEFRi0JPR739S/pni2O/RmVtRvq7hf2VPMybw319lBPmwkwLf
xnxomxQxe0cNBgy1/XGzavWTd/pfVOYnQ9SLQA1oRzxCsoa5XKAY/CX81Xxmz4wy
pKs0Z0BkxseheGXzrNpgXD4BfBYjxqvE7A17hsWeXo7htb+jpcS51m7sfbzps1Z5
G32BVqRwa8DZnfV/EH0Hi0b98hs4E0ildTbQiGTraghJLhvqIoTAx9oTAbmdjlJo
sOmYMyLh8KTJsLE1QDTCd8Vr2e+5Tq0byyIsWA83f82BnW5dmOFHI/n4BzJIoI0g
8WdyGuMY7HJc123SWvv6TfkM3LHuQiIl4lVrfLHZ21wbgnvg5bq2VFB6KEVxJTjy
kGGMDF+ND5kVL7rMpHHefpGd3iRffvl3UA4j7C/eqkiY9pInkQPysbM09a/Me9fP
Ni8mp6k+Q73lQ2u7x/NsS0UgKnev0SefE+feCsC53xzKxsnpAFK1cfp2E5/RYh2x
kBexXo1vvbXqeEfzYSqr4c2XTvKeNpbjHNc+QBT9zzVkssI7/igvX6fh5TGUkBTK
pgKhuv1rEURGCzjavyhhFHjiVV0HpDlQCQj5JYU24W1JaH7pNDhn1Zo6tdQ+1tA0
w+OrRShkgFUIz+A1BcKzcnrdjXayfx1r4GozdT+4ryyhbVPfJPlmGo4YKOz1RmgF
glrXxvs/9teTHMCnL/x6tecr9tTffqd8X05cKpHLu+/FgpU845CCYEMFxxHTPF8B
EHB0skvq3DoE39+iJejz6zCmZIw3nBFnxWGueLY2XP41LkuxKuyN1dM0PK/17nBP
WIltyXp/4y1q4PZWNOXHgP75dZ5PHgXGrBRp/5ZOAVCZJjnYiFCkdv+kleBB5bTk
/ZgbL9uMPrzwAegAyab6QDrTO+sBFwQPwbsnvQP4wMj+M8kF+wcU2Ulpgd23KJUg
MYuwyjaWPMjxzi+2zCbjfgJfN3oCq+WW+AMSD8Pxx7AP1ZcqrRCsJzaHgFJsK1KU
/MXtHuWlFU63ZwMm9LmVR29Sjrt5PHz3ufD3GFR7EWWgoFGU44UDkMIPMMkJa/La
Xl+vNmy2pAbs8/a91X563PyE3xpyfPZ2ntGKoIJaGbRJLwGkkkXzpGJVVqwSw9z4
hMBD0m6Ou0hYtbx/P9nFcHTMdUHkGWN5M9k/lqfOpBrxUFatLqILYyxpK/sV2Zy1
W5v5HeDf3wHd9feSUDoLWFKY7+h5xZEXU/Spr4l6jENsX24nyMpZ5decpMGMeyvv
uQtOIQpTHVvNhd7zvrKz4isQ+PKsT4g/vMhb0vFseEWgAKhFIynecv2gbCWuXrEP
bDNVmI/Qqo5FcScxqT3A5iOfjICoW9OE+0wJIanJzh97XD46DtRHKI/27+meyWmd
Ne2f30G/rj0vgZs21qEDwZ/Hg5KMWd/BWEo0Y+3t3VMPRfoAhdu7E4qWsn/FoBym
5wl5m0icMDnYkvA6OvTikGA0rclduSHZATE+VdtiQ8sROq7xL5yXEQeVqEcc8Ps6
Cbj6KNqCDBgTRuNJL86h5e4BuRRi+/7eojL0hmBqlhCj2upjdJsSi51r+/7or/QV
5HNIX457Ldga8/mA/DTEzEUJrPaaAUgc18AyFOUNul6KpNdwkvkYHUMTo1AUMTik
Y8sTYksWG7DNSvytCdYtbuBKDQpHvBX+6Q1UZX/4m1zSbUMj3T7xYePx39AUiY6q
`protect END_PROTECTED
