`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6EVoFg4ZOQKClQPUFxTfk+u6+OICm+peA++1LLGtvrv9+ev+zhpynUxLb9EMtopc
fortyavLCBK/6N8hAZnhdYB5Ekw9FKAnfVPvuk2Xvvry0XDjbqxecjLMrvVbRzyg
IUF+2IAvPOjX5DB0ngKyN4WmXq7NnerEnQdMtqKWcufNQQlNgg0Gpe25Kizdu2NS
DIfPUpAjLc/XtmKeOUFB/Qa4cS0LQmOhpiqqUCCZDIih3oDwxSPRMfZKMbvZjLf/
Rm7Lc7vAIJySrdXxKtIQ7DsXRdVjVO4Gc7qvMjWzfccqswSz5e8Oa5jStITOILmt
0KumIBNSKtK1B6cNMCPCzy3xm8fM6NPf+/Wg2QcaIaIyUDFLLG6L4HjTGGOtulVQ
zWxqPSlUkt9Ea9GuQuN5IeRHLatGmBRrb8Xn8MslVwnpNlY3xZvJRru2TK04wNP6
w4RBDzyGhuW1DlS/qYg9+kuzrKqLk9NjcR9zsHeYMJ+iJ6rJwSqjadMr2110V+YT
mk1cILftLHu12qcSCsWROc6y7Zk9Y8R8qumD9aRsVTw4ZBm9v3xJERv4eBic9zbc
iwQOh0r55jQNxTJ9KEyXxQ==
`protect END_PROTECTED
