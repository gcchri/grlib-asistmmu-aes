`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ip2zWyU7BcBfv0LYCaJAQTEHShULI36y4kKBgJhVD61io2WkSeHgUbdJAXr8m9zf
yPi+y2zmU8qJmXOFqojoREiW5tS1HbqXXEKvC0Ja7btU6RMCFJutVbjg6aWue+7f
qYMTG4jBaOvKIbVq2IxYk7+A0pEd4zsfmm+Hu3SCuTUZZ60l/JIeJOJGnzTaoqhF
8SzBGxco2YVwEOclamgG9pBIGpStr+g/Ta5zBqwU34ktrW18KX/7MoDE9xWhtAty
LONq5aSRV7LWfvAOzXsSEqsEr8jpcp7kUBXAsiDPHySoVHMIK4wG7HaZ3lCRP8gl
kd4BXX2keQRntNuUVfH8kpAZJAInU1QfJ/muQR0/0IPEaJ6AwrwqyIL3fjpat2K0
rPaY/Sw4Ka4aiGOhDh66nrwS9N8re3XqAbXgYin4pNunrxb3X1d3wtD1601YUmjP
oVKjOqX8dL/G6Cng7hu4725G+GMqkIRkIFbwrL18Xy153QmuMK1KwINPxaldiaFp
CLz3mIOEfdXTkZfpKbut4IcT+EHSMlk7Xn3LQZZvTyG2Od8keFZp8R/C6NJUPBeE
KqOyf5m7ho9Q7eqiKIdEJGupS7PlIAg9ZXGiB/tRvM1HFtSfb+u8J1KcMg6SC5lk
jG7EivvlfSLc8WhF8KMJo9jLNlmkvHs800BCbbBYVWGqCCnmd5BHnV4umVYZZUuw
JfY8c+V6fM+mm0VBjrzt/1ReDfokjxMyyz4jSKRhgpfuU9XhMQ3LRu+gzDmBQYxP
2kq/8Vvt484CnwWR1Uo2Jq85Q8hKCB98C9jRWvOkC7cqccKFevYKXT9wXqKO874y
CXoyuTMzLPHHaoGcZuXZsLbfwB1vW/cTjeRiTFhCP6MvWJLybUJ7o2R6LB0F+80g
uI0vM5PgWAVKq1nlomUKnQhFC8cAE5GltC9Xxkk+5IxsCvYs6FQgzrHb5bdIbkoX
WMs6gzibqDB+mDE0i7UrwAFwqvj3QfqY3zBez3VOQNpMEKO28LyG1IzTPiIc1H7h
hA7ii9lmkprN5fAjx4OzuJQhWpX2LiWdbNjRwgwAA3L7Uv295lidugkyEZbm8a8V
nGEDEspJjIB2MjzB7WY2YJw3/a/qJGageYUCl82oP7AmHkv/lYGXHgXOMZpyG0sz
CgOn+oS3yRAccgogq5EmriKmO9GxATcOyaJyiLn6NFhvf4XAhEgZnG2ZbmLIg8gN
ggnCP8/Sft4FM5gdoOfcbIwkAB/3a9/92q0rxU5JQNZxsCt04Vz5GRQFmZ+lpptT
tebUo2O3cg/STRiiBz6jYeP8lN5k1i95FQG1Gj5E6cSMu4CDGjsAUkRpbsvuTB9g
kZBNADLmRlPG7MzlxYr6PQ==
`protect END_PROTECTED
