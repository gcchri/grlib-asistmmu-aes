`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uKOEHTswwoQSR3D24RX/1E3d0adzFxg9AqQwwAMMZEql7g4HBzkqqS/Is/OSTDHp
5ufuDZMHC1PBBsy6pyJGeTFLgVhKENPqXI9cwSVT10Qkg8oti/a7IWFxOhGUtL1s
h9mtngKmk0S6bAxrY8jIfVsOlGtpzKHCq5xcWTx2s8gLvy/oOASmlYN03V6Exnb8
d8Z9YNViR9MWnLYLWFCe2VRgrp6xHGGlaFjebPy1i+QhxVqBPPBuJ3t46GLBtKGt
24m9fyk1Jx4zhFotVUxKy87AeAx8M1kPeTVQkhjoQWCZgFSP2DsfuacE81GaOuLH
Zjj0154AtpKF6wxWzosvTjBMiP0YOEzMflMCNh+bbQPkYyCwzEaHjqI8Y2dlhqyo
EX9yf8YMjBTigG39hmEKZuLLfWOzxlM/v2lIXIWvqdVch/pbLNFYv7onqoOlrjlU
`protect END_PROTECTED
