`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zIyhdExUuhkP0UAlxXb9ckYgbxGtO/ztARzoFldHoOatTaNJbMrdhjglqSkTqW+L
AnzwgqEACfdX82E1G3rUNbpSSPF5yXwT3SamSafd5rbO7D/xukcUkRBLr7XkKyIp
U9eE5b+Jxmh30SciW7hOgdAJCgNOpize0RL1lXqD/DkFBbjW1v0W4eQnQvhhEJbV
lPw36UgqAJrJ0ehMN1t9mak9wNJJ5vtH79yqfhP3LSU9QFV0Y7Dqmi+GD+7S0YYN
OTgls8LrRmEoEKASoCfKG3MmFV4AigOy6QXx/o5C+1oVLBWBHFmzEY3xGEaqr/wE
Ojicr1ESs1y3mAuiEGqlyzaIQicVraZdjFQRZwtCtiGhy5MjZA4J7BR+i+xqDqve
Ha6D9o3g8Fnlw6xJVG/b0tSlDaVTFa6uRZzn5guICUbV4YKy1AeSP48Jr/82GYu7
ifQG6sMdT6X1TRtSVJ3+DZSJ1ECKZAy0QHdWa3PfjEJoH8Nb4JCzx3xmp9bS63Vr
oWrsqbUF8S+YjwOi7vOSDsV8E0er0zhU1hMHwLBbD3Z2lKd2OGjNNIoJx3qoDiCk
`protect END_PROTECTED
