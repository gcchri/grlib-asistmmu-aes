`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nyB2GsPx/SkEzpB4ntyMwk5aFqX0L6lDu8hiUxhOf18M+VfQC7d0GLUW+ee65FZy
iQD7EAXSSrTwrEEzT5Xv3ZMX8pQWK6w6bIAhbR7be7eDmrcPJcVEexrNSO04p4YA
FWRkzEI4v0YAFV6OkKqSTjqnvX7F6KpGZyd9XEXW7WM/qNn5D6Fb1PofZWdJuw7/
1PSL+PPP4PXetJEwQJOOI6xy1N5FH0nux3Am1AGmnDSYtJyJuVargCL8E/03zrTg
zh2pDkhNLPJq9NOhVvMvFbRiksJ87fJmCVIWLWMyz1iycCSEdxf7285e1F6Hryhx
GQiTcV1OPSqGGz2v8QQi9n3eYoOU/j3xRSXf4g022PYV0oNAUQycoS+AeVeDKo96
VegeI9ul/AGdAWIhaSlsSm3kZnifWVz/U2thnJXz4VwaEco3dgAzPYZE57SIOsRg
PxYoF97MViywN9OhPUJuJZtpT3Lt91ErEFlttRPpUK0o+qCUkI5KDas2KcXVAyMT
9Zb/sR2SFmGIzMvUKSaTOt11CyLdP5JbcgFCmMaKo0mtje+rjNTcCYvEguqhMHLI
raCXm8izTH1HLi2bAB+1Zbkltcbb48Y74vC5JBSbAUUO3jacMb4xMFCjUpKM5q8p
WD8Bd4TAc3mMosPYeiKxug7ZXrmB/O/dP8EZ5mMp6ZFN3DmwVFMvziM70b+bXeq8
CPnGhO0C3vaHB7gxc588kNEPJ/xOTSQ0zFuWFvSXfU04zId4ZmWrBxO0WURUoYgo
SJ3oS1ClUQBW6dL8CHJvmN77AA6CVR+O5VRDBShMGXT7vqjKkOmF6XLzhlVKBisx
4jXorKNYeFxssFX+HvYB7JBF/XbVxxe2VuEr4ghhmTl55aHWcC9GgoykhTvZ5khh
9vo2TadOsKcILdG5/nBf99OU6lPYqtqhjvKxNVJx4LO28lhdxgQ0lYjGiVjsN/nf
CrhdRiEpZ4WdClGjuTW+BPLW2onQ4tr4oTqvZDHVOmWPCu85bqaa7JRVDjxshDrZ
p4MF7yP4J6OgkSU7qkYGLpK79iTFliVKAql7CIDx2XWe6LQbJ/QyVEERsFurbbHh
`protect END_PROTECTED
