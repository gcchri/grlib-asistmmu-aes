`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v9di1VYQgAMkr+yQ5lLT/dUlJfA6O5NanyPsV68RA94NxO9RmfI1CySMMPJJxucQ
aJOBLmGZep/Ubk/2vdHo6j6HCeJyIDIvR/GpKhrV8PtVFC/ZTeogWs5LjJIgdQd4
VmkBrBRrPGxEZdjqcz0Ecx4w9P7O0TekGrnxSTe2EEKTUWjOxRvub7CsWefaa2N5
cSLuHdbUxMQawQsB4fX6/nAv2HjHU0nCXyUKTFv+FrZPGAVR3F5y/Lb+1H0v6ha9
1k6XkqL8amlHHqvJzvDYgSGUJe7Oypa5yVst6MEunj/3NR9L5t7m8qDTXuhVgiyR
8GUZ3LfcTEwSMzGaygVM8WhjL5b8DSVWX/UQ8BKYQdcnZW+MZnNnq/AdtdQprsz+
ClEZkCcgxmMaEPnW0S7gkrvz8CeXkhdPP3IATQ+bw91x4salgU4A+nLRtXGnSNAM
GSH51hkiZhF5L8MI2HY+tBayJ/EYmdM4VrTedYfzNNcDoCbXLvQ9g+2tuDA9H/Jf
auY0zxrdIgiYEjb7DntRm1mDODf+bCW4rW0aMeokLzB79otPoB8sj0fpAIdAR+0E
atfzLDIERdbECJjB/VmW6FPEjjuJjtUzeIv199nEQvqWo2RAbBSy2nFet0w5etOC
qEYmWbGOBHNZe4MiiK9kbGyzdLRVmbVEl87aNC7CW+0B/wUr+PoYDlZOxT6rqJvB
SfEcmGwBgfdt0u4xXe/2SMsqnsZR74LRczWgiGgiTjOG9T2UpfyqxmehTKy6HH0q
m2C//I0L/rxmSX+hgjdhVukZrDuqNxXzdjfa6/BFMT7ZTL6/NVO4aMqN9yH4uMa2
QW+68G6dkIuPf9E0JHdoE5nk5fZvJkOm/DOYGRT1441jV3trKChnkMBp1j8sUO+5
meY6FILGHkRfsjOhUoAZUe2M5ep4SAqlU6d1SFE+B9xYTSkrWi7QX/NIlwOdlTsf
Er5+qqj2whww0g6yILAtZ8v9ZB0rHX3l8+FGaP85e082j1P+HcKSrAphEsljy8w7
`protect END_PROTECTED
