`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1kWM/5FmgY7CAnKc92jILBcwnVwKwTq4mkXdwVAw5y9DR4ke84RCOQsIt6euvTLE
/5ey9kU3JED2rFDnyDeLF3/Cd2yBjxKxz9RXDOCRsrCxwGhu5YUNO8WLmUuBLkQF
Nktd/gaU8hDvDRJi75koAXb/KAsodo24uG3Jf4szIEcxJASRfEsFrD7tqnoHhpu4
gRrOjDKhZxJSEm5P+6RnoFmRfZkTop49SarlqU0PlUxBJR2/v3a1ba1wo8iQruLt
4Eo9Ib9+W1osH7bUJ1uRmg==
`protect END_PROTECTED
