`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UvFZUXyZTx9kPFfTWMmlqH8ecIGT/zmU5NU0wOsOurgMAOrapze8RTgvAaY9uN9I
Z+ZckexQf+/9kcfmciNfq/HyLdf2FrDJsmVQcHimJfiJWCHxbDxGsc7Kem7Wntce
2tT1WqdEx/dr1uUYpRtL5+DK+A/+NF98Z4+asRzE5LCEptW6FqUnEoQvp2ZzOLq2
gI+a2dbMwk7W4rF4zk2PNC06pKgiAgBRj4qHS4v0tIc1hMVzetcP02nqGd5MxVY7
KuTtt6OWNtzSdes2gRJ08ra4jMdf8f93iPIze0VPIdEnkWafeG4InBCTFYfPlMHA
01AVIaGxMZciumcwgn2y445rTWS8hEIgHbY2SxWs/bbsgyIYdFokVIZV3dsKI6mR
NdT3DMi9yaOE+VCkD7+4Ma5fscudUdFXgmBBuYB/vVkqt3SIRBtZFswywcFuWlf3
zJuJgGUuV5ZzQX/X3eOZrrXrTLb9HlkczZCiOCn6jKAIkj8t/EIZXfK2y2/ZT3l9
61Q6VHyiKevGh0PX+LYMmQe3GPMW+Aqc4Fa2niyooSJW+/PV1O3yQYwJ6fV9o8qv
ai6YieQrfqeWXZVkJ7/EbjFvokH0IHN+t+oEnrmaO3h1TfSlcVH0pHcJVh5t6gCZ
Ne9iBzumlgGP4MctGofmDaKRHMhM1qEjIZoTE+cY9G4r6heMyWv6PIcDt8csWSPq
+ht64T6dMi+mC1b2TWnwg2n1x/TUdCqCUwBa8QhiiqKXVvmzThGZ4dO6lczFhEpE
FPS1SYnL0J62i2sfMO064T3uoo2hIFSmcT4BdXLO0e+UJoBE4I8fjWLrl8glOQzG
FTO9k81wCJZe1NX3PY0gaFR71/flKXBPtM/FaC03IpFkagni0XxRzPD8A+W88Ykj
ACAN/XvFkfr38yDaN+Zr/mfV/Cq4Gcbbr6km4yuyIuHmxadB2AljNv3tIouHWD0S
golqmQskwzh4it/GGks4dcqW/28zx3BKSyxO5kdVjoEgqGR6dHIY53yRHOGbGosY
T6RAxSnd9YeK2vOcanZch02wgra1WfsqAlxcC41bbIPEk3RWU/ihluCOS2UxWaRC
06zOEaH1NinXxwYUODCoryGVgU8UacgZd3nOdstKqZWfP6qasHH+qyifOWN92Sds
pTivJjmq4dYgAbldBCOOFV/3Ple6wm+cRld8cDyVYkfzePS/ugW5LLD8QOASjPVz
UkbKznKZLzkTNe7BM506bkhLVraMDzcUQki31JDqsRPzCxUJ9kLxa2DxWJl9nE3L
3hptfGrH1InsSmrNoRyPSCFRPLDRfG9mYJCexHsfyEVK2uysymn5p+U+sp9zlGBZ
ZHT5oyA1B+/qCqQyNppsuiZwJUNqCYsnJLBepPRVWpb1m71sR0y7dtVElPl88is/
ZKGrepGFW7D41fYdeNbQbhfibgKS2+IfdMhUmrnyKz4NSi1+nP2jDOZa3YQR2bQC
4j/S5DA6pTZ6V3C8qa+ILcBYjzRFJFeIsqGhwVD8QhU+AR3Y1NTrw2djleBON1GX
4XKPmdjLN/N22TDTTD33eNRxckXg17v5YBBAD7ZqhNsJS/WEeMBcElIe1Ik7HI50
33WwtlkksBguXO4VBwGzOysOEQJzWn2FnRyzWqLj5RfBKmMl7M3KI/JdL0xQ6klx
Zp7ltpg8HlsaehPpHwRGyBagxZjyzLUOOwQMDecSt74xXk7OhKpoi7WMNEs45BeS
Eyqm/m2x/aQZlGmw6xRkEbCROWQql47CZ3mQ/kK98IiZn4QnVKqXHL9oAmI6sgdy
UyNbUX5eh1mC4pmCVtXWUpFdwECnkNh1rDbVo0UOOp8+qX9Xk5acNzxkn4GTqxon
RnkWp00PeR7PxFHhhKcmzdNJ+G5WKs1ImOiRnnk0NuJNv75k4v92e4SJYLdKt4dg
j6zZcm8vI65KuIJHmboPtbjVkmdfE8wQeId2wWPaK45G76xt/bqiejlbuVMRkQY5
LnBceGJqFxbhVufTBgG1lWcqGjXgEI37fXASoqRSMSFeYKgvfetHS3E+iclcxJFJ
P2vqtuVnqnDBeSXZuY9WQ8kA1MmTWeP/jnLLqGTU3l5h8+/G6fvxbkPkxXXsBJLq
wSYVG/iq6YYI4+S6hpatNv+0b4MY6qq/K8K4Fn/5OyDHOnsXiplXyvgwtoiixHGz
BNy2ZyD5zo8trEVSPyBsfpv3wekwwpjf1jVty4sjyms+djtPsu9n1PSkvcoxQZxh
Wcj/wSclJgXojEW0RfzUgfNCi1Sw2aHfzWs9UZx5HR3TBCgSLeK//79LCFcjtz7K
0JKE+asxMP2PnzZpHsdcdMLrNRdoCsOkS7V46FHkeWFqIoR+K7KLkFeXBgEAF0/5
5DhC8OjtwVi/DAmnRV7xcfax+KOOphB5sgkqiF3PG1ioR/l+bd4pINbPjUcWD3Ca
ThO6gtVVmy7AiHMcosM9jOxh1RNy3KIm79zpT/WWjrf8m37BI7M5c5WtsDZu3Nlp
E+uAdcwG7LLm/hf1ZC9ClRuguWlzTxhvnFdTiOTlovNa0QbaY5uiPjStj7Uqu9Vc
J6RUIQ/FTe0Ym16OwQk3ThkQVAOUM2QY6gjOWSb10z0TmCqbR/7oYPdX83kIIBJh
LKNvSifxevwrGc2YtdA0bx5siHi7Qu8FO5QAR2LjQuN1my59k/lLtCioA+o9ZAdE
fII/BYlLH7NCD9l3iOZq5DWIw/xnUSQaBWLzwEeTWj0vUiOP10j++v2VfvKFf4AM
J+fMuORrHvBQyit9W3hgDkUIhuEjQjRxLGQShuTIs6/D5qjW41lUvQ/+6IvsJA1v
7YLbIu4ceCKYO3P0s/kxX6Mmxdyl/DEBuosAMTm11qZZnaLMVk0FTkZzcy3oWiVY
GOIDGVMc0hFgsz4ti034JAxqkurZ+ssd8+krGGD8RelQ02d3g2gIdugG/vS+mAPW
X+qQOOi3OYl9D6BLLeAtEz4/pmWtU9P79PYizMS2GtQThVeald7Pqlr1KCVbLN6r
tDQHmrRndw/3xWEzjfM+6IwmhJMIniuHY8A2EJwft/g/elJ+5Gez/tcmgRAOpEUQ
7lSSW0ZJViPzytUuuKs2dCi/kczPChkk7RaYQDsLuTqCjYZ+1jPlM4EpNfX+3Yyt
RgZiBmHcQdBj9KtrpPOYzEBcnRmgPKbr/T5+MWxIO7pSyNIvmW8v8zoE1FyK+lYF
sXGoLNMrHyICA2SmPvYjvRzm7qm0FFVoG5D5U1nLStA+5wikdzT4UMzWIXueBmd5
r7hBhpOcwy3aVf1y2rR+Pj+Agfbe7+TG8NOwuzHw+nAZ9cYlrnOaxRWf9z5B5Y4B
TmHit/tiGBzkWV+dd96Kq5pe/bYCo/1tE1Q17ocoFCxR0xIgeTvg0wO7wbRkoQC4
GM/HUc1AqOBNS0mXTynaPmyBJQU/xxLllSYTjq/sF5Qyqk0o9A+ixmMGs+zo5Gta
XT6JwC7NXnb7iEhibgZT0iv4esashkeLZcLtjmScTlvhQvfAODJ5JFQUEGxFsTBY
EDFCT0JZweJywIjHFXXsPifuvtyFvAZRH8bqJRIfkp7FNjiCj4f96ZwgBfD64q8B
eZzQWmpJ6IJDOWBH7XEfzGVZ3aZGiA0jAPbGs1ZPUQhHsUUkFqn3mBMpDCz0EwLI
2NI6nE0J0tVWhQhZq91lLExCCDgWET6QImKPw3OnvQ9Mm9Rj+gSDq+d5OjwkkHH0
OaUXKQq8gnH6mKGbTpj6lnhVz0VOg/2ZgQPsiEhiBtS/0GsLpN3kJfchpEo+RdwF
mtauhjwX5q+K/5bUnNN+7qPUbbJg2H6ifgclwy1xBwEXdVD5altFZ9VTyg3jxwPO
D50ZLe8Z3yTRsGZz+HkvLV/kUHwb+R/crlQrHZTLV42ErelWCOOL53neu3/iIQD/
XBtWWWBWYeGMBGvqttSxUQKHHTWr02XiLgOOgwRrp9SjF2D4NkErTG10JFHFWZHI
dwi8PU5U9BrMktIqZdT1uE7NCa9TZsODAsHbH0xsu9VWzgMiLQfhEGJXXmT5Rtrp
84S0eWf/HYmUfxb4M8pzco1bHbUYN4FMpELzUd80ZGcBM+ttCExrXDETcTHJdjJv
Q1SrFluOS1Pl7O/WwXcUgAGVRTLIG4V4FdMDdQRZA3aH12KJrEoP1HAwwgQZzqc+
G5jgprVFONsM9U4eiseVQ7s3NT57MCxKWlPj1Kw82hX5+pEkDVEJz9LvJyLybDTi
0st4L05bibbfqOUimvF9IZyjO4bxuWYfnOAMgEViahfeijrRPcFMt5+rDwwdfbaA
HjEnna6ij9jhKL/zwrdIdwl57IfPZV5VaGSfRihScV9cU3TThkdw9P2zAYSe530k
IJcrV4oYUdxx2A4dpzjC8xdG5fn0wGudNtnb+H6yZIJ3O6VkYFHnz0xoUDEDRXyl
OovKV+HQKRp9zHpAGG2FU1/P0xwQHF+YLnCHMkD8Dck5hxH4/RtAKHl1cIneWSpM
YwtjfPQwY6vWmkpBK9IPjnFwLPdux7FQYbyODWWWKeQsFr6Q7VR5P4kOyORN78Yr
wRKXrk75jD5wRdwpgS4cY651nF0lRKYtiCxM3RlHjfTZ+oZN4jIg2lQMXHhxko9m
V8943rU3fZnLg0mVG/ZYbh6KVfwGNWqG5LEFF5PRachaQGQuV4VSleQ3QjYL0DDA
RSVZoBuioEZnHvCC+9Rf6iu7Kc3oYwgoWcshpL7EjBspzkKru4CVEhfVx4VwsWi8
uxxF12muE+qTBwDw6l/ycngsPhqqa1lmiTSnP+zdfMmIKN+BXGtNfacqUaUKJr2j
vntVBpt0iXiQfF+2+w9sWGrDUcskrWXUgWCy09A4Nlcihdm1vhZyBMXmubcWqNbq
vWDDO0WVieNx28CHfQnX/XRAN0TqmH6gtcBv99CJFY5zCZ3aRDB2M2PHFVFkXzWC
GqYgvLEqhhjoPVF+r23Ls+LAuvvNWDCVMINnJkVzTzJnv1R9i63R9WbWK/BTEkK5
OszVrOzni14lnUmsJERVkLA8Eb+SGnJRpTBt6Zm0O6VfNT/YMywKlFvaBnd1feMl
h41HiS7ARTDLFbPNBeQjbVIs0AMNe4gYt9tXkqf+sZsKV0ia9/i7C66vGUgTQ+QN
3hE4p70rFcXN8dE3Sr37cxPurOaG7Lp52Ie5pff+TjHc680BRhs+2Fa6ZDfSGRS8
T5TLqpE8TBvTb0MxS+i+peSRSbTBkgyEsZTZ5y6RzAsGQsntQRNEpvkRjHlLvvyF
AAJJjx/EOREXTEQwNdzUJdAxidgb7+iNdjQ+/E9ksarAYw7bKLvmMZychnJDZ+mt
I6sQJLFTrbU5Z7C7qebZf99Li/dVy45sHJctjUw09lRs021lyX0hSI5aEutaDDYY
iSlTtc2dnxRktSxEmFfdYHSr7fyVRiwCkECq+qye2ezYWni4JpFIhbRWwbOlO+Z1
zKS5Mklp3pARtnssY8N+3ob3juBCsBuOWN4BRhZDcsycp/FRlH+/ofXwXIwpcXw7
nf4wB3AeCDHhYNtYbjnnuK+jSMfw+/CJ01q1dgYrMX6rFQcwbXP5Acv+tLKYTgVY
YbmhMoHV2CL2fiMSXCNFxrm33IgHbiXRpNtupdyc/EUXZUh7ClwmuLmNIRUWYAgR
B5uaiAJgN1rugzJaTM7sP2wmSxVMJxMXysJ0lAIMoFbA9Mg2LPx3DsUTr4l8rbss
n7DEm8CZebzyvqxN5bVYr4Gis4fw5+pn8A0w0FmoW9mm09JL6bdcy2dDE4XKW7co
7xiSR3NZqmt03+VsXf696zN8cVrmOxAEyWMoURG3VOuPASDNYuj8FlLMyhrIKivT
QLjJsNSZKNnc3udWjfiwILRszaEI5J5DLJjYv3lSEwNuJ9BLY+jdHBctb0mw9U1x
bU3p5/7hQOnwpIS8R3DnfeId5uJ+rpW6GYGIXq5+NO1+qw/Bsh4FRGsp3yeTR9CJ
xe/VvimwEKSMUfz9qdEBj+wHbt5X+daa96YEVX5FC3uPKlxzbZoT6+CzOMkHxhrb
88Da1SIscNdCLy09hpUik5yOm9vFYW9q+GhU0whOuJWeozAUdwfw/wpavhL/5q2Z
T0XNMwBZ3oEY+2/qyg5efg8suebCFO8/TR88EVRND232aNC+uHkNAbx/Ce33sI67
bVc+fBem4423ZqdelvgGj2ZEf9uSIE7qnu5v2LRNiRSL9uFeIXTj7+X86I902ZzS
DU/gXQXCi0T6QOmyI8tsfgDyNiV/HofMK3oNp+Pe/d2GBpuDXGEAlDypVt3/chru
OEGZ3IcUSSumw7Rl1Z4VkflS/tv/SIPIbHPEUhnu7F4ILtUo2xNRBa+j9ar5tl3w
44ijF9uTIFNNB6CTvGjb+R6/kh3YUa14ueSmlwE1132sexzXEvoWg/dy8xDTnvvE
+hXzjTkiJ5M/Eu5UrY+Z9F7bn9QRgM+6ML3cdVQtRtlu1FrpVpo0dR4R4d+yH6sq
1I2COG7ev5F8xAYvnOPNFyVtxnvZUW9dv2xEk+CauCcGZ8i0H14gzvAMr/GVdreV
KGJOuOOTJNEGXvs+0hlhlgjk8M3L+M5psYNc11N5daUmXEZvKPL3jQJhYzcRYm0p
Ze82KOoKvCGk9p5mrAN7Z93BTmUB5dHCPMGid1Tl3x15UD1cq7rqDgVJF72Ox5DF
IOKGbx9jLvTlzwl3Vf+zqBtDWer064UPNE0rL0ZnLGuxr5sQnzL4JkjIELDPoRIB
euwwj9cJUrgFq/8RlT2jsoKcMBdA+Qf4+Z7oE5BvxNNtMCNzhGhMVuxOEIrftvHl
9mImHHUKxs+vPYSe9tj7uHkRlTKSQMtOG2nSBqGVD9BmpOl2Rn70mVTg0iBX6zIH
SCvPm1i+FOYsz9sbE7FwRlGI0hbvsKhusCQ93P1NTWqoSTgE2bHFLGZkK31es2ht
T0hnHSHI7hLbXNMph2Wvi3x14XnxrQyLo98TAJeXFXcS5kf/hllohqF7NPvastjW
UrCkLnUNxSe4OS8JWX77njUVx3m7NwtWiOL/DnNA2FAMjjd7PmL1QaNUC943l0om
/PdNMcjvcn5vvPCwEdasVws0gMUu6pdJ8hpIaY0rBDxbv16sEzziCcAueIooee2E
LhLh4uB7RmagqqwUvk/wh84g0qUTl9v+C1sofvTfK3JW1++WeShpsN1BU0Q8m8QZ
8/dc3dz55AurFOYLMS9S8hLHIQNoQuZ8orIutskcl7eEiY/y0AIhN/r2dFqMGPBr
2DqTWlpvZhffKhpMv8a5lG70goP8V5LbPuU4lcW6xia73pOpJEnvy4S3AymoJxJy
4ZslsywGROVJVISMLI105lYv+dUm4hz+Xu544CPosL2GzE7ABIMsC5mU7BMITYBc
IXIrjnencmHwHdVh4cuW0qHAGhd9W2CQqH31OGxVyCYrfhYMIA0ooV53CNHJmflh
g36flDVzA7K1UOTYwb5NkV3nv5oluz+dTXS470TCsJX/TNOFHlv4PPdtt9p/uXhx
nfAgsVTsBZL7Xt1iRL7BvCBPThnvVYHYxWmnk3ZazLKwAYfYN6Mb8zNU4n90fLJ3
udCtuAuT+/k5qA5wzUCp6XxjGsHcaNoltUEiL5XgV3rbfRmvvJdy15rS0L0OHSSP
k3yRfV3PWL2JIK83obhvkraXUE2Ns5Kbec8fJFx1NrCnzgdSQ6/cCKsUeja0mOq2
SG7wUkeZ4G7+Y3JgFVtJ1gla4WsToVdiyf7dQSPP/kZrzV33/X1A9nNv+YYbmofV
LJA68gnM5p2npR7XualeTv5ZncKOSEaUeRSYAbcy8q45j4juQu0EjkWIuB1B4zFn
G5Es7j0kCb28UdOv/ayf0tJSlWUHUzJj32eXj/fmHUhFqeqGA3uXcR6RccxAGyI8
42NdkPZud9pMhAyz4h/ytvXkNqkIucY+81sTPFCXOzXyuhnaFuzPfw3uMlcYJJ+a
MCyg8kuHRwWEVOsdMBoderkmtuDlYzvrak8DkQ2fOX+UggD3/vCWGEUzTxiHbsoT
VAWXLrhLTpAVWv+Pm6JW9B1gITC8pIimn+Eds2b1e+oE4fHUECPOKdk6LD51yUPB
TrI3USnyIQN4V9DbamaWD1RlgpGrDj7awMNCXnrj6K+SCACUjg7vxPGS9M7vSg3N
R5/j0NHPwzKnYqrmDPf/8xdjQrRfKf94MOdTjIr+nwbHdkhKp2gHUQCnnvxb5u7w
onymW/4i4Xs8Uv1ww5xBOuIkF+21mwmVZkr8mzcoFEPJEo+1yv74UEAc9qTEOZPG
pLJsSVTwLDaXfMZ/CDQjEE09LQUrcl82Qvf5fp/C0ZYFUhKP0kvceR+MrHsaue+o
UwDW3XRI3dzuV0GLtNlNVTXW8K+3qbvFKJeav+LoDBxHvXZIIJSDYmFxxESrIej2
MDaMY7lzb7V7cB/095PE/8OrBYz6r37WVMH9Qmm3k+1ySETTWnhmgFGOvLV7Cip3
bpQgIXf7FUbPZjQrUDP2lBIHJ9GLdrgkQ7iAo+aL44qK1+S1zas81dWN9VYAr9Ob
924gB7HpLsMq7MSTB+fG/qJVTBOywuzcZavd1EYNe/YhqZQA/X6W0tutEtob7O3o
luBJl7n/gW7+lVQgoUVA6u8q6WQ9G/L1yk3nwr7eeA9S5/Cs59p399lx6/RcfZTx
Wp7dxzJPwsuY9sVtbnql3+XFkBQvUYS/gJH4gME2BEusiwge3xGiqB4HVg0GEelu
KJj7JbCl6DhoZptqm9NaxnMId+P0aQKLWZzkpz4fR8+YpXMtayH2gFUy55TYfNyW
AZl0J3kD4H9ek3WZ7vD6jQgVDOqOgC/j1wBWNTyCat4a28FEXGUTnqvhZeQtt6rn
NFVBsMOGe0Y0ZrdFM6OkYWlPCrVJJVqswrgUNKHDun35JHvZz3Fv4sPs9KAtl9gh
aldiJgjXU7319gZOTBKINj7yCWFX+iqlMGdbeHq6miKKzP63n4s14OCXc3xIww+0
Nn0rYnTcpi/gJ58HaBUfCwx8zXWXdmAbD9xyi2mAxSfe6CRFGptdCbrmMM4e78HA
gw78Nx+GXuoOBl9btuxnIAbfXlglB4xUuP/SHv3dRVbyotnM55wtB0oRTJVp9hQa
vy6thusb/BB3X4FG5tP6YdrP9Jv5XNRO+9jOuK5iRG8zgud+2GzJIaB+GmPp014o
qiEgk2WLjppBzfY3sHtuaBhe/jyGI5DPf0YlZakDz0xJHl60Qo0cGaoJGHc0gW+Z
qPQHKPDdmluqPjuu96ON2qernJmTany40GgSDiu08lyxFXmdpnvCiX8WqqECi0U7
gMuwl7v9SCVKN8hxQGwVgxMCnlT0ICBFFUfNBOjHvxdsF/fmUoGsyd4mXW2gY0Ut
de6GZhoGUTjaw4eNFrJat4UZXVu9vm6kRahtcvEkCTwNCxt265DGgWLsZI9c1xdR
fcNbeovhEwVW+EHu37GXnlZP33JM5EgQn3Sb3Nkf9zyyxFceTPBL+fMOvth4E3cu
sKj1C93//w830EZ1Rd1geC5f1HrxrHkIAJ6Kawo9957Wksj75XZvMszRc1y+eCTh
UDIXkelgbCIu/9tZMdEErbJlH3yNNyEDRT7j0/sJVOoHiereHj0Z5iiFiCvpIdG8
fMqP9vm6b4/y1N/AXIZ+WRocbHMbpw7wei0oRdzEzsAy2NlyQqbrDgEtIGeoktpW
hKuIMypHSi0OgLAolVKkSJPTt3Rl1y5FBFZlAXO7wkavMPHj2XAd/9uORmPkTcN8
OmyxanaT4P8wBxJ4p6uGbHbJ5E1stJxX6UWvWSuedUJXT8SMus07kR3yxXcBsrZ4
95JMypOhKElf2jlzYnD11TSHNLoDDZWMLiz3uEGm8861gSr1zrixEk3a7lmjtaUO
P8BW1e7tNVnchYLciqKVOtELdgilGamL3VJimYWK2ZERQ3eu84AFXADjpill0lU3
C9Eamjyy6XciD2gpkmhnZanyjA12eipyEe0phyStqhT1bDhKDVbJ3yqxuchqbe9c
DHvFu2Z6UavEGBTDSARAnWLCttB9pE+CbK+yEGLk3Uo8VJ4AOQwZXxLC10iTG092
xBxiyZoTlCyYgAt5ve1KM2oDizfKqvkCJ5YZ5AeMdAabN2InkvrdO9LfuppveSaZ
cKVzYwXumiPwCUDMdBpz/T0taqWO3dWeIBRdKA8kAqFUGi9x0fXp2mRB8JbpZrTn
uiocS+a82w9uEDVxJpPaM2h30SweKNIxPLWeBPxmDeIbtu6tPKS4BN6pQsMXtGGF
ocs5VnjXUk8ziULhQIeHaP7wX/iZ1Rnm8MIYkdoy2FgKKJ5m2m1q2mwfs21okmbl
cf2sHwedWPfyXUkcxxzpBBZPb7H9/fBlYMFTHj8nhD98G5U5Wxs+jK4K+YM1SpBK
prWzjoqMWHodrl4WL8TRXms6GgOoP2QMyerJ03B13ErUJHS/47tq2jS0qrxa00Uh
QnoHSlwmTP4oPyvz6/cxrbSNmqa4KQAOQu+lcR2Fgv/aafcwcdnNc12k4CjOp9TE
bUWLrsSO9O121UNTL5jIuDhIsH8ryxV/m2XKR0Sf04m/Yyz8FOy75TzKVMMIFkQu
x0sOYMykMYpQ90fV0XHBk6U1vG5w24rRbjVzHJovdUoabUDoFYqGyZgY6LYEvrC1
Az6d9Pm4PhzykTbNTAsT9QXFu2giBItC6Glqu3toNh2bRcHo0PQqgC581cbTgKlB
yt5XlB8czQV65fDm9MldUoUp1sIF3OSMqQd4DgobZv1E/Q1FoOvgBV685kB+Jiwx
IEDIWIqCc1FY/osgmPZNvpZymL6TCGn29ncXfOBUi7aupy2g7UJFtQ9W8ALJmbDc
AAv3dDUZmeap/dUiyUROykJQKt27QvvddemZ1obTnkfkvt+OwXUk1duaMwZ6aMzp
tfts0qc1EjQVQHsVSfjn4wwqDA+scpCbu3gQcohgCsJb1X4N6r4h3IrexIzRniJq
iMieRyJ9AsuFhutUrw4cgJTNHg38NwCX2s9yDO6cYei7Smt8Ut1i2RBhJd0XvMuZ
6dG515f4Mk+3KvIk2+j751lwUSY/pfCf2CLj4LkrdgzCfzuYKyE+fB33KdR5HiLo
DpTfs9rO4PxzJoWEBlTbB3J8PJLwietjZAobcN89ztGilH/kbd4pyY2a89iwaRwn
wRBZOL9wWZK6YV39f5SI+Q2/1COPAwTG+TG1bD2kcPRM30figyh193Rg994UT8vs
DVvK8XZe4FAbo6VDfUmeFBLu3TzQhvg62Q18PcOe/h/PB+C/bYWo1a4xPAVNXQ2G
FOtzb2T/P7un5z1A33qCLIvW4GcQgu2EOv4WTwEWdF8kgyvzDb3q9LLRYC5oZ+bB
LckPBnNjYznVIOiGzhMo6CqwCd03Tu811TkaGpnCP4HNPg8HlyftfjA7rZpu+sij
qtL7uzT0ahczA7HhQeyUnGIeDVMO/unhz60BefpiJBb7DGQ/l/FWot+NAiZB9Kxr
EeJ2turwKFeJER20TKPEVo9GMORyYT+1RvvRxiDLMWmKXx/lOIzPNS4Wb0gIork0
hySvwOQ8CLa4jRJZ6uC8M5wT3eIgw1WKfUKbNXcEBji93kgBtnSqQ9BBmWFPxgVu
jwx8xW68l9AWHI/xde48wmvceWM8V/0voS9lFxnCnnW37DWR74w4A1A3lUXRPbSE
1/Ia5V9x0NpYqrpta+jYoyKl6AGNtjqv4ulFD7pzz5wwVuwDV3LsDPcT6817vWjf
BEQi+CBg7/3dO0cWChR8NbVpvi73bdK0EzcEyeaEwZghDzXWTvnKTUWWgQqF3PDo
snqfg3gcDNMnlfnaFLcQm5buKjvmxJGq1KMfB0ILQKF8rVTATjcuZ1BvmJYGK4My
D0Hj30zXSjreKQpoCy82/ltowYACiIFuaP6vKsQwBDpCC7duzYJta45ShmOv8YZc
EUl3PGTIv7CIyb9UHfQn2UzqGR42pZ9Re+Clrn8OsLseREQckSXrJWfp3qbxrrao
sHb5icgL0OEsVa9+1n8cbPnJKshhEmVGffzw88wtAbnTROvskyTYgWETOOHc9rQD
+V8ekYl+MtqtXUSM/rq94lrkFkhwz9FlyAjUlGp4FASshMcEalzj60dvF8JY75Ev
4JPE6DrVyADCf/2trj67otqO0Sr8+mLGKZ1xzg1HXl3M6oc3yPCtV30F4d1ghWYr
NB4HtepupzM4di6c3YirFqBbtb7vF/NUg7iovW4jyhGy/R4tRAA2KLjkLwtL+kCk
7BjBx5FE6ix+ONkwzzRDzQ91BAlANbUl4c/69uH6O/2tMz1KtyU4XyWYNBNhBz5Y
U42RNmpbLi3/dyYxANMu3ufl3PI+QVUvDbQMpqnJeis7kdfGy9/qqTegkO3VerkP
o2WIIYSGqBeCRw9UCifDVE/OKBdG5tKjvedEe0uRkMAvhxHvFEplbmip5XSgDCQM
gEDZSohZ0ynJ2kU1vJ3mOS1wZ5IK6UcrL+IMjlPqasjMeQhXeCvupTnlmjYtPihs
1Cmcsk60DWhL7e5yASc7o5c6xi1D7epkghJn8XqszZTnKBi0t7u+ox3E5ev7G7KU
Otit2mKA2NIARIBO7tcCBRRGwK4jWkuBnqki8Vh9GqscmyhxAmyjDUdrGZ3Grg5y
MVAGbH9KuI/TBJekMuMxlubvGNFqIO9LFbTTo+djCeY7e187F+7uqizQNuMvIzeP
gk8rCO+tiseJkWPX3VqEowe+SPeSAny18TK2yym5fA1CkJSnLM96VXvw9aHRU0yK
XQha/Qwlc5DQ/LJyq8J4pYlc3++T/EDKPj4h1hhM+evBajd8d6UDgHKtuJAKmZKd
YOsBu11k75n+KGtN6Q5GOyEAO4W+VjjAw4g/ODgOAQnFJFTMT2DXVpEu+IFNhJ3e
IxRP+R7ABsKg8egJrzkY1yZ9U0jp2yjSHSsEzrawhQjRC0X9KwVfHiA/8AHZhIYt
K63rOV66u1/vb/ssVyL54vnEFADWhYgaZftqdYfqV8G/MuwPW37QkWywrchqnc9T
HnGAVf/9uzaDnQN2B1J6OzaYBIZYOAJonjC0mnVgAvSRjw6vO7fxOzqwnemg/ZO6
FnZS9TU+XtYfbWOIDgiEoXLOCzIpQmapZuLOfpU0xYBpMSwEDJBMSFVnCFvi0CXs
ZFiOXa6IoMtCmRItCtr9LlgrPlBqeH4PMhXgdMGHkkEhzMxFcKNHLBS+ahZkEU90
CEQpVIbjTLpGbdK8C4HMQcioq1Vz4bvgSrceWqsMwx98W3kJ80I4zPjzqvffOP6a
QGMrMFn+gazN22VE5ATTAZeqmKSPpvoSRiylsQtUqAxs6ncL0WE+RpokvpgQtdt9
Gvy8LWJLehO4Wc8nZvQ13pgEKSAG3KMZNHPczQrS0BnSe5AA+1D+d0GnlArGoLr6
nuXKFAATUQcNGx/T1wob5xv3jddBoR0/VyM/EzEUG4JDyqZ3FYN+QQjqjxHoTmuy
oAHY/xj7r7UbJyL28aFjp7q1aniWTROonz2/M+Wz15EOH/vGHVfsDgTopSFcA7FB
ViKriHRw4/X7cYwuiHPd+aUeE88CTE4ShNp5R3oTJY3R948YzW/N3uzIMdDSJKOw
y/lOBsJFL+5ie0uuIbThQuAVO2GLzdGt6pCoUSphWzKth841uemKKfj/E7Qhb+nK
1VeLbFerD5PrkCnsRTveFGViCmXiDXzXI1w6Gzgx6koqesJHBt4LLSlR23dbEXRf
1sNywaBmnHUwMUyma8JML6FZ0ySH2Cg2aNPWYyXzbER2LxfUJPxFuMtqsUs700ik
OVzBH1FtQG8Srs3Iug1MHlwX9JRpNKYRxkEsfOV6H3DxYUwLCuqCr+wQF3dxa1SB
XhyqmMmBQizJaxIHgtyLYAfuCtiQIIgPfV+Lf9+2fY0/Kp716FAn4JHZq7wzKgbi
PatRKXPaDxIUnVMAC4BmWc9+yEU5aJd56ST0S/tiWVQBXIx2hzpTouh0Sp/gyZL2
5dUQXyPnYCwtqJD6ELw/rBtLg3db9RWm6NV+3pwiVy+Tw23l6+RqA+U+zw+eR87s
2kCs/Qw+VJRNff5kTiRqq3EQyruFsV8o99EBk5HsaDE1lyP/n3IDJ+qbfKkUZ6GK
QQ0Pb3EDRGA36CsxyazDnnpVs6QTyyxp3YemjNSWOdkp4cQ7bXCjfoH/gL+exPIt
HAIQrOxge/8Ao3fSYV/i4l5BLdcifsg0asqjZmgqBCcmNhHcDumcDKBbVT0AjelF
7T+2AvLw8Py8dOWW6u7sWHXjTRtsy1Sms02mSVn27+I94VOvqcOYg3Lm+i3ZN4hJ
tBBzYxWLEuAhj89eN+FDdMOFAWO2T+vxh97BuIHks8YxW3khTf8Bsw26VIlTvkNf
U5nKTU1uVamQ5lcGY0YMEuJVEfYs/oB9YSRBwGT3/47zHu3SyVxRG0cD3nvcqzO+
vsvE0jQ+kvM/3lz90BaCLnzrJYgnw+HSw9hVyKy6XbBIgm6/3zPonoC6mdWtUmGt
UluZKJvUGVGg1463YquALjEY5COPoSDzmwRAkRHHsHOOG784/AvrDaJRQATPqswY
dZ/ON1CAF4t8+x1gu8H+ubP2XIPLdAn4qcQFRs0Y7HCj/MUOgV8kjEwNC6mN9k0Q
Glnbxp3gnV/Fj7Z/glZvCmDX2ZkH/wXKA69pd60Eovp3G9ujBakH2yJ/UhvCSP8j
4KjFkSAlN6jo7i7/UeAodpDNMG1796XMp7ngg3NE9h6H1BNaB8G59arT/z5q5/yS
I0U+N+FZzwv6v8303qn9zmBIGMVrh3YD+i9yrlTX5ikHgRAJeBQ6lSABMPSm/Mdj
iwuwEFK9q3reYzAI37yFGeSsip0luRyMbQU4BMJruxVweIoIqnykev9/Vymm/TLQ
szJNMXXVzVOvyoPgZbS449VySIx0KkR+k4MrAokR/rtp2r1BClrf6/v4V7siQshu
XyBVIG5I21wUcMVsQvV5pA4K2strEEvwR5gKG/u2OR+MPdszUybNO+Hcmj+xO9Pn
sAyGZ/p/xhM1CZ4BYc8ILZxVb0wFRzAnTBWDQvPNewm2PEcDXBx4usCx9L5/+wbS
5dd81Gn9pjnx1uKc/DaAc7zFHsNkYJMdoDB/v6sJD6jNbtPW0CWO0va1psFknoMR
95VY8EccXxP4CuNFWMRDSuNJQax8mZEoIyLzdLyuWzjiLf34coOaqD1k+M0LlpUz
9wAeXnDGTqhLFPjVUtyA3rhiqwBBpj9X1bTBgqp2ww6gVl1PtOrXrpIKXb0LHAUn
G5bpBXASRXtYz2QBwTxAoCGlaFgTxw4MTtWHjw6E4CQ2OiJ6VU+IQ8BJ9EZvb8uk
o/7h9C15CEJ/SJyhEtXs04ngmx3iPWaftW/Vo73/z891u6eMt0xVVA5ibLe0HBbB
aUB4BHgeLQE4wgW8b3dAZcnVG29N64r8kukPDALiIimUsUElIBGZ4ofghHmJ4XAn
phua33tfJQx6qY4rmxYKqE24i+EW29Ocb/iykWDaTcEFjgd1nSWrR9Ok5SJQQAB5
pcQmzYjEXYzdKCWKNXefMZ1P9NJ3HWE7hDgVVq3X4fF8f9d4JBJI2FTtB+w93ryO
K+zTjiV5+Ko3QA7lfgafm8ftypQsqQutS+UOP3wEPf/11Ww/qaeBM9dXpOOybBP7
SUQE/MI8X65BoOh6IhMrEtbwbW8KBw5Ep7aRSp4AJjI6kJnV6fsFxnUU1pgLOWow
g6GRpgnNoYPMcUL/8YRTlmLyUwAtKB/jMaiDCH7ur8bVQiHha6ye/hGVD45FWxTp
yRbOjvOxrN9A+7nPk6KrGElpIhJmeIlTnTjTZGDXVQfWFIvhvt1jRzIS5cS4mo6a
maex9XUjlfDajIbiIEGM0NthtpM0dJ4I7BcsF6HavHeQAiNAW4WQNxqr+nbOpNbH
nYVYApov4Nh58nQM2PbbNnxQFwRUKIOjYqxQOne5CnXdJdl5fRk+PVJKz6EbYAQf
x5xbVJZN6runp6oo+aUQs1VVtLv2G99HZepxio55WZUuB5GxpDm/g2yd9Inhyvip
MOQL4p4eeChdDnFeSaY7pInL0jeljbsJ6ixkSD0fwm0pmnFngvzztDGavgtQPB7i
gh06d6QEMGVmVxDNLADoIGHZLkLC+DVv+crGlMtAICw1CTuHx9ufA+bs0nH+2czJ
6pdVn2sEwClebA2sS1B2GV1aFIp5+oqwJO4MK+GsDvzgPiTtX942alzasuW/9aqG
7s8JwbCgyIL6hFmhIAwXJ3kRXGJGvljcPGPB7fT8p3zkkmxnQKBvP3PIfefiqA5w
xIVeKtAppBqrAxC6w2mxiRqcq8ANtZomuOzeMzN20sccz2VdVd/mb/Y9pNV9Zy0q
zoXemkrQSzWb0qCk9fRB/0ApGM7AUn3S8zJNBDzTESLWrwFtx1Wl8XGKf7cYRrR/
wU62tZlsykcGqZcZkFumuh3iavAeB1J7D+NAeUhsEZ+Lxd86dTNVrIpfHJoxkOU8
XpPRv4sz+ddJhaRicm4ppukN/HfMxivw1TjhHZfNk+zAudhrhZLdaoQXQhzT1UMC
eXwTxTVLnMfxhpD+N+Hm2HuRg/fID6xf5sC+JmEPrFYK9zEr0OAVSmmP/mbvwFC5
ZsRKQS//m5ekP0P07wh62x7Mr3O/BVwmFs6mEP0RLWOBWm+7SCo2dpVU8OgvUvqq
F4IvBJiD8htEmajDY2emKJewMkawvLMz9W9JeLcB1ehmrPJrodiCFRuSLq8Cu99b
h21NvovqbkUGDo2Xw9LgU+sg/fKXUWgldpWkK67OAPv9qF/zkn36mfKX9baRsLwy
NUKdldoCNWswyHiUJj2fw+L+Ql97dfyaRRTWk6y10+DxzncRTOrjqeXxJdgxciQF
ehRmlV91L254kjhW+Mz/AD0bNdLjP0gQPyGS6o7wtm4=
`protect END_PROTECTED
