`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aX6xszik1eVlanwb1i0E0eP0O/F6LcfjQT8+kvfzN+SBlCk6n4fFTkjEFYL9baqF
hgb2f+WskewLIqgn7L6FCkgGr2scT6xLRZCIXqR+TLWE4iBF+CaSHeyiaVQkXeox
KC8RoSIL2Af+RGvZGZSMum1z9c8O7Q6PBJEWa5E8aqeoMIePK6NUQc5ybWz3Vpbs
a5V827v5Qie80OG1xglAgMDu8m584hVcPWEhbatbcmeyNIeg6DX7RLHa4C/OhtX9
yf61AsDC0gV1kihiAIVcsFuoU3ODasi+ZoplrTPyU08nOrJ/9Orhxvgar+F59etX
bmd73U6+4rvvgp7SyQVgv4JwuQxtsfMxY1SV+8onaXH2y+O+Ydgyc6XahGCG+DK9
bTstjaFTqoIZgiCVdPRtfOiKvtApW/7HIrCktNuBuRPh4Ck7Pbum9jV8aRWuO8Ea
qkioQE6eEOatcE1ezhlPEwDBRT88VeKZ4wxIFpzKUz3N3yw5w/ODdur6SAw27a62
RufaPLe/huVRyS5UsKi4xHEhMALNNj/LSNp09yDCfMuC4Ymob7sw8tA1duo7MI/X
QbEIV314EqymalVcTfQacA==
`protect END_PROTECTED
