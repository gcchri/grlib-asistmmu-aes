`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dWKso5lAnAEFvfGAMsAsttEdaJYeY3JUiXdKLyC5vL8yWzIsMd6nKXwnzOpwgzo9
cy4srVt7BhOHudayqE5I/6wzzuK4YiQan9BDwKZFBlBwwNQs7VX/UO0fmX/afC3f
VbZ+e6LatTIofNNrKmyYFUnPtnA/VfwzyjNtmzWdrfv+9AaaARRQhuAv+fkn9vr6
H96vZjFHvdPM13KvaARCdBBO/sbylFF0cGhS0HWAulBje/C/talpReSngE9qpHY0
f7iie/Itc3/p8I8GG7/oPjlf6P6JV2Pm03qGt+KrCNLQOEY7vRU0QEpPiWiDnJBG
OUD8v3lvd56Nh+SHgelrIUl9eLUz1hjqZxFXU2cIiqe46cp8pOl0tEs8SuAFfEgF
9sengYQIJiHT0RjXl9HtfcaqWYlydBYwgVCnMINuDNJGvfX04osuX11gmgAxtewS
GkLidmmdi78tH0eAJ9I+hpwAXBT2UCNFq0YjXtifBkVYyLqPervY8w52YcSwCjQz
fRU8sziHNqN+JEhwv4tNmWUlM0x2DFqqED9wZiZQlBCqTKMVJYOgEKFJE+YT50VQ
fhv73pCdxcXZoU7wmQKt/tlSRux7NotAfdYSPVDI5ripoyauAs5kFI9cWcQj+6Ih
2zythltzeZNFbxQpMTRpKJO5eRBmSc8jGVesQwgKr+a4lrO44ZAHJ9wZBdH6WbAj
dAg8AApFHV6tM98/S50OIMlYx9QtzrgHUH9OT09Tksgui1QyVyQUlhulMVLoEj9T
A0VlcOun7lCJc4AOmXv8O+6TeW987IOpyv5LEyMyzisJpGPXvTIXo5z+itn+UsZM
TEV7fKrrDBDQO0PWhcBsGt35GKtE0Tsw03Rh1OGpOf4QmdOiVqdVkwata2AFdC9r
yaENUoK2ydjpzovxwgU0kaMc/hnWpjrUBD8lUvpWUKIpLugqt+MKzoEdzqCnVWbV
TyFe1k97TRIA7qpNKL/oMsPcZKnTrdWLLFamOyLzWw+WEXN0C4jI1Tk2gSrzgFtC
ObYqbuTniRV+m+J7g5izk5htaky/aXzjgiL3Kus4Nf3GCONw9giXGsXLRKQAHcgY
QwuZ+5VvjJwHTbJExs2Vdeci+QWQ2kjP9n5J6ljRJyTL0IStuzObGT5Wtk9CUw9t
ysnBherF1ex5YcqPvq2pMqmEZNzYU0Ugx/FbvRunwQDtYiDhHVQMQPoGH6Jt/y2B
hjJekIKjFR1DlzWfVWF0PTr8C+3jKiiIeCoFoYHpkmkzRmnBv5eZaO3jew3+DL6p
6jsg9zHZCDDKGBfWwZhy5beyhiZTaCLXuL+lhnV0DRA=
`protect END_PROTECTED
