`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1HaTz7k08GTnIeF44eNdHsGLNMV/5msm8W2QSUt5zWcJNugXlFpLL23+/SLxv5SM
uCM1AGpih5WPeYyrEQjA9CegKqAnAmj2M9ujF0KH+grnklDRGGGI6wwxXYmLTmaI
mlbUPpeHvoq5tT3oY3LHiTVB+erFsMlvBfUBRJXK77Br2f4sxPhMWYzR/jKnJYC0
HdtrJradu6Wx7GZ+rNsYhFvvGFhelPMFax21s++s8WNVWbLYEpTpEyZA422APhj5
B+6ADwvGfGg5by7OzPd3piKyY1pxNUWgZQTYfcDcj9E=
`protect END_PROTECTED
