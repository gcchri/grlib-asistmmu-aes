`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5MChPxlgPPVxotH8B/lAFwWdVneeRlCvTfyPx1xXsEDR2H8nDflAufx7PaH7zaVH
/D5/5MJTrzx3ocd9xPMP2NgKmVzRKjdQxYw9kG5uQGMJQbBnuLG03t/xasEsK4US
aRhYp41MWEVkG6i2J7932qLF468ppqOKklobf/IM4Fq/v7Umj1YtzWImHkDyGW6s
0zeP7fi/wxHtj3jo3/Y4LnNhXdlk1P9wttZtqQn99i7PNnmZpXQGr9VRazEbsHhQ
EzvGrTwoXcsiJ2+XW71O9/d8MaxPYoRQM8uHjYU4boBNcjPZiXB8MublZ1OXciZC
M8N+GOG3PqDEdb5LBkvFDOWLZF5QPHGYNtYbC63ntjV0j+n6BPGDRxIVNDeenWxc
cdN/BzwTwLBHu1OKPqCBswGQ0UGADgZxn67xSfFgSWH3muZCo+kIiFhFeEhXxdqW
eoXvlOQBdGDuG+L+13c9IASLx9KNeRwP+G2mctnjQcnhF1o2eb2xBQFbJMX8P+EA
kIO1P7gU69A5GtJMEZz5i7igOklxqDFWXuG8NzILj1OlNmT+BY8QdqMd6umCnd5d
Fgb4hVkbQD4Iuwi/wwGkTo369roSud0I75Is4vNbKsVWXj8Q47Hz3P0c5C8hWVTO
`protect END_PROTECTED
