`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
soY1ou1QA9OJ4QhQZiwuCVgT+hwoCz6BC6ZFAoDZaaWCVFhvFb5oS6zg3huBjBVF
wS8gSVedi6jyVROIueVcp+778AWS/gHmnoK94RBvUEr0ojJrKT2L3BUS1SLhLMbt
CJ4aRC3lWWTotQ5M2T5V0PGu0izA0vKkHhbUpCH/G+PaymgtciEz1jodPXmbuvTK
LWyK1b2rt7hfaRG1OTfGRH2qZygMNtnaPZVKyopk1wOUVWs/SavG4w/cXsrSoPLD
liEbLOpstO5ex/+Kibq4+eTlm6HZGO8OUoe9PItmaE8Q5YQ1T3PZ7q4ujB9AUMFN
l8Ztqf15S23BmRBS2dpNDNpWnxJlN9dN0RV9VpYix7aF/wGMe1UgW5hnibkkvAF7
JSNoC+PFKhAvEdGSpdeEyqHGmiGuv49isA4nRMTlJBRpjPo9FcEnJ0vJOeOwcUJw
age6FeRdODEXpMpFtQ0V6Um88BBuNZu6keEnM+5b64F8hl/FarOHBTxzQ9xqTFvm
DwOIapSvND98lnIxjad1wleZ7Pmd6HdAdq1CIzMi31jLLefYra3gjtBzvQJK5aqQ
YtA/LpO5Sxn629S9cudUU2nt6DpYpEwOeCWWPmzPm4j43gPCU0n0mui9EwfQRPQl
6zaGCCqeeIE68p2jZMmCVA==
`protect END_PROTECTED
