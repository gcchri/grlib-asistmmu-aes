`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vBQlL2sjoOsQrJWqJIcbVr0t1L+ZTHSEFGJFbysKqEwUkINVhTIVGMIrFVuqArg0
fiRNBio1K+7VbZ7YimhO6UBlXJkjNsO5MbvpvsrbdLn839HsrS3HQ5xDumNlh49A
pLRXsOrZbRM0fPovDYIYp7ASvEshzjuvVspY1J+16VfJxu/a6J0fSoGXnjKLwryn
wZt6CWyVZMilulp+wL55Wqj3AmI2f/Qq3P1Tc4WU3gI0Du6TtmzC6WJMNbBqznOT
m2hRXXcFfWQjmYD5urVI7W22FRSMKXcBS+0lsikkp1OI2H3PWSE4OX3QOR26xJmU
41xOphPww68hLa6fmXgawDcKFxUVwSEeoIrznUMzyQ02a/alkr/xzMsLCN0I4kga
ST+Tcqa5kiOABmECMmQ67ETY7xdAzMCcPZILY/gYI7BvNULCc7t3B1YZpgKerOe/
EFt5wsmUBkFkBHez/tPTivND9CzfRuXPjCI5Z99SFz1kQtFS38Y5Svhu164HPKre
OH+Pwcf9uOjZSFyYUcLJRftB6cDARTyQJ2KACueyCUq1GKiejkmWf1y8FReWwdCm
nWvHsRNGYEAm5EWzaj7lT0pjjg2AK7cgj2Nxw7eOWXyYRNtInv1SzLh8EcXv0a1z
5O2Ixsmg+gU6UY7Wxf0YvUIdztT+FTszPxdb5A1UvKAsk130LZRz4Q3mpKEyDRKt
RsYLgZsHb3hVHnqfoy7PdX/Km58sfZtPdTEW9AiFwh17VxXZJwvN6x/oKceHeoeh
bJLfUBxPDAm/Lz5p92MM0JxMcDbTfIaZ08mI/dNMp/javULclNWAmKKV++DkpmsF
EiAj9kdlRGD1dgOuWzo62Njgv2tLg4EjBZm/5xSKpbXv5xVs131iqvZFSc6hWmge
pvMYo6NwiOuzQBjASwmiT9qI/Hqgx463PJUUjtSpk0lPWeLmq+odU64wsPgb/Z9d
yqwkAmJNEdBXAwVg4ucdVtGOQWP9UbZDjMWyGj2EMbwDinuVGJQNb+nCiNS6ZKNQ
2gi1Mt7uw0ej8+TL7sTr+0M68AXrbSM6d7dGj6eoeCTBEN9gTUMtd23L0lD2E+OW
4zFrMdNMZUaUQsb49EZUf9sVQCXU9JjX3nuzzOP7WZZnqmmsGSLvpoChWle1dZA2
YA5+Hy7hBaXHRMSCEVA+iulImMP//PphgZiTYnk2SSUnna/PuxwN2OxEQsMSU8AM
VM7xAKQzGMdTpN2fGPOSaMhaVFYN44GvF0CxrhTOdoFvHO2bKK+WRRtFSguhPM7C
i4zhkSd8BBcgNQ+4+E8N7bgBa5bliXzF+S84LAdw7kWfoayll41yzLjMfpe4cklo
QNSYs/Cu9ZO4WjXRax8+mA1gyEwBGSa9dib0d1UoizKWtm/M1SM/9paU3XFFjbYE
l63TvdrEkTulbSGnahHjE8afNSW/JgIT1g+5WNGDx1O2dBCb0RT43mtLom7DfwxH
9DYp6RWhaYNXQbaGd8AZzaRS06L0fUW6kTLnrWrjAR3ZCyybbRF4hg0fdQtKW/St
fJfOW5+237twln1At/Q3KxaJZkGnSVCFzwMN/NWKY6JXc8B1xQ9QH5zoFgIO7/Dd
PXRQYBFn6IvXcylZn9HZvgD8mfHzKUuQTVtWEhCOBcgwLoYMpSWZTtuKPkZEJpe8
AniOC396la7RyJ20+Tg8G/J8KcsKjqd/liOU8xGsa3q3ENesgJQNbqYNuH+GrrbA
2IkEuFvs+CaaTPMDiot9daJED3iqKc3W2XsLzClXYTxXoKZ88N01Tjw7av4B4LG7
qsr+c1SS9vCiloGWg370VGL3yXTFFZyefpZigQiCK/H/1Ic+85/nh4qpEJGUbXIL
4FETyGnQ7y6EO4WM4w+OEJPZZJuLThul8iVvVMpKLHqc3YMurSjFvGic670c6pEB
eNgRyB+SfNCpyfmcF/ZOOkC9lji4OctWjFP6kX4SAxM=
`protect END_PROTECTED
