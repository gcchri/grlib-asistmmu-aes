`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n/jvakfUkXNI4MjmULgXQfMLAHTfC1CDCnj2D17Wy5Kj3sEodJnxvSKWODUyF1kx
nGV0waf8UF85Kn4ZPxHFtkUkcdChwL1E87jQvxNtrNcVyDrMOUb6jnw5aP4htIlK
EcuIyiQtp+HJy8L/6r8emIN8hRu82+zLnhNYiHlDrcosr9GJp9Iq60JTYmTOM/2N
r5vmF1VyoqQ7XxcLQ9ezQFdGR7m3HjGxVjPzLyf5kTMrpv3UwZs24VULERKBA0bq
LX3OkrLnnlZIMGppKDGYYYvgHm+bFN4PGGnPK14rviEFhsqX25LnvArn/2kAqGIp
hGZyQSXq+TZguqfRULBtBBx/s5ofHOtSeoBw01Txhf5bHoPKpcx8P44spXTB04hN
dHQIU9qF20UC11JbJRIQKQvawK+Ol3S2XI/XUZJP+oaVgijYbn8owAmb+iRjnexW
Jurr7MaPNKxabbKlhd2tzclL3L4w+BJFiW7jaPHSgL6ykuVOKno4XYQodVb2bgF/
`protect END_PROTECTED
