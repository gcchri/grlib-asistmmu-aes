`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AHAFZDdGmWCd4CwNZoIuta3umlb2wg8iQw7RHbP/gW6KJEilTC5cfVe67YS9XN54
FN4SRJGVWhXWWQvyH+RnhGVEFsycuvgNQaeqT7s84T2T+CmAwzxCbvnkPtFmedWe
JGbNCbMFGUNdlfLxrVYvthZGAwv+ZJgy/MJF9I3vQTczlmOT4LUGAvr3KQANxRg4
IlRYZVD+/kdQQA2b9RT9/rSMJb9wdfhSkY+ZWFpBxAEQurorKmYPOP+/zjFBTWye
LP2j5KIRhOvR5slToMvEuqipIX6U1WtRIqj8icmw8NLbRrVNas31pcIlJKfZzoDD
w8CNrKRYzZ15D7u5FxvQk5BVN0/4GB2ciL7u5tfgcoWXPwLQFH0euHYIv57od99r
TootEo5RrnfsRWSzBtrRqAkidt+ISzS8oUHaOlrUOiuBFmKekLfFJxQd65V/iUkL
ee2c26cPbn2UABoC6fq3zHoZVqlJlDiER0Kx90J1Pc/gjKB9S2q0NCAcokzXIS/9
sxMO1OZbGgAofKEZ7/B+p4uCEiWgr8UCEcWGPTGjGC8+sp9EuqJqNx08RbUK7drY
6FvRBpVphTeAZ8ORCgr+8JLZZ1jB+vIDMp9lycT86DTblPDCStnPq8kq6G3X4Hhi
pFtYUI45gmP9J2NznUkE0az8s7xi1YBdMrw5ze3Ua9Y=
`protect END_PROTECTED
