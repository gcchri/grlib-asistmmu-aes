`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WVa2M5G17cPSG3WMQtf7BzKdXBDsMGSaHzYiNbW3Oanu1UEKNsLTwwumXG52TgYe
B0qRGEoPGUXNGrbUYMXVwhaGSb6rJGWZPIy6fLBnmn+AYH4kRViJlirJS8bQ8QIB
xOglbqZsaSu/14e+IO51QybdEOGqUJhx5R76jDCnGJinE35N7rhKIPx1Ob7onAyh
t9pJvuEnhLP23gFIMQYvJFJhEPBjnxdjXUGlJY7O6TDyFJPD5RIhp5E4s99XDEYi
5DylbTkFY/s5ZpVR8nfpPSHLpQarCm3UE77aMXpALpFWP6DYzpHNgnOQ8TsuK8gE
wjo6tUd3rnGje/d7IlO4pRFGkZCIDumYEUs8IeZIBA09GryiV8fumAbGQn0YWeLl
R3YFcdnRt2MAvLOt+tHOQMm+5NA+2a2gL7QL7k/gb54=
`protect END_PROTECTED
