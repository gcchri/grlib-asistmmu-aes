`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A43yJw5UdfAmbDMlGWQglYO3OLigbqAMM5ZtUGwUiW5JoizyNBu9XhqoshW4kJ7g
0o4v4m+xoEo8rV9zB38fBNWrxMynDt/zGN851sHH99SSYH3jz/pRZqBlqiaim72l
KjAosxaDdWZV+nqjXWNvp5taCMTveFyj0xeyiScAgi2E/9Bj1X1iRUEiaiM4TyY/
aJHU77xV/tFAFXFk4k1qx2DY2Dr1lKWGVJtOW/PP6jUlDpemfFmHEORS6IXx4Jk8
L7edIXJOQL0aku+MFEDIbBi1qj8zm4n8xYhqb9ySLnsoK8RzapNTWAyQTv6JLjR+
VLouvvjC1HiEpyYyP64TkrRt1muW69eAtPTcPWdSecw4If/mZqlZRAc5v6hOaEyz
LeDikZ5DETvVSSQCWLD+HoFPvWpYtWPliN7dsWE0LdCR7BefR1Bf9MzV/828qr9f
hiKwSC4Al9nB2p78c1AyaueJBzPmlMAVmZMDEzwLqlnqXtpCUq0oa2afF9LIFVKG
Ge+n/8AzuIwAgGdq6MHEWT6PinIw+UiZEvqcXELopknYxywcP4xP1ydNWWMWEYqE
Meuf6sJSRyDiRvPfCDvv/C3sbt+TrT6YUO0tac2TTGZxL5kx07imwDT42ohv3hGx
FrMzGQUNNPeCA0jDVo3ZkUx7spckyHP8cntN2pbz94mRE2B9e3ZAYwJlalUNYAVa
6ol+2MuT4tznOqv11bVxdMS+0L0A5HcJ+b6BbB94BVtbDyQcC7MDXxxvu2XzLRxH
7lLTMBa2qlGg0NyB6qR/z2jwADHrI8auPgFdd2By6uNFWLau3VtuGpsxrjVqucN1
gUwIChIkqQ4b1xqCJKn6xXaiaQDqEnuYWzS6CLFTMNuGJPbITQ8qBGtmZHEsGUt2
qRBiUI349gM6bfiRQn0o5n7VRleSPU5P8Q6JQuymJLK2Hi+XZ3P4HMiE6ycA4mqq
5io6a+CCUJdXc8N313rkdxoWOk6V3HZMDFY4i0Dls7+yao3OGa9cnc3V27PpSMGf
yaz0o81sGNHgXhzrLvOk2Z7NzodVALTzYqXVOb53ZqFgXueB8p5Qlpdmk/9JrES4
XR+9sAUeLlWNyG5/BcquK/siV7KAgNTVSAIcBRNc+tPFJNGznPwtNlVfC2Oy4fKD
puzCZfBpKNRIAF1VwnDtTSxdDbU9PS06DTOShCwIeg/MOaADabGgp9UFTDuoj6Sd
kk7dpKmezeVQmg9FluW0h1NJmTG9UFDvTsiWLpkmjsupFSvzUA3CYD9FG5ObdMmd
+EmM1cs64J2Rr/2JOmToR5lUicJHQR2tlbsWmfCh5vuD3eG3shiT9VTFvBzA6i04
VW6zfL7U0N8n4AhGzgEucXj4vv8eFDA94wUMNNC6X9CJokn/n6ZaLjRK61SpdW5T
+6AEfPEryLCKgMDquxOrLvyg9HP9Kfg4tbqgcVfOZlhcSoYVKnYEwlxpY0yigfI8
mj5DXq5FmeMv45k6I7VW9tw4d36Eo9O4zF/l1AkMLsHIXxo3fI4jOBQfyMXOvAzK
3Uz49OXuU5m5+bZZXTzFGGXXMmqkW/ZpUtBTtSzsQdC88Q3K3MilWUdE2YmJB2IB
a0sh0ANQf4gYbK7KrMur+rfqWY64d7ZEzIxhvxFUsRSaBHqYyvPXqMa0y5Gf+OD7
m0BRt9sujpOSnAbTBKOYI60EE4lDjU+EjyK1Z3SdNzexFqq7bVQDEjbE1j0cY0qv
i72C3tw1jqtvw8zhdXUm/k2O3gmoVkUqvENu5fGQsmmzBqCo3tcD4lcChyv+LuAc
6J8KczmCLX7A3Skci0Aq9dvYURJtBtmjOSj82Jl8Xx9GTEtfXKoeVO1i3PzuY/s0
Y8d9FgjTiQ0HpvJ8GxfGH1F+WVzdkRA3GAYyK0KGAchwEJOMcYMmS5jmkuzYOv8X
mEMWb1CC/qzwo3Rxd3PUawpH9+K/aQWYiNMFIPMFqtL75/oIaKgEFYxuX4OzDMqK
i9RNYVzehYLrUfwWTGMr4kfpPIPveGtwWhSnTN2NBNtwT++rpKFV6SKM7F9uMbGa
57NZ7q9rVfhaPC4pDWsgAWHmg7xmqW/s5Bq6l4NdKswAduT6WdpxyxMISWN6w40i
rvW6T+7NUgexjnxh7aXCIHCWfx7+qeYbg7YXUAJfHDf3SclNV8rsWg/8acobDuYM
tYdWK7MmaRyTRrTS6exS+fhj45qqI/io1HIqcSZoWXUbOc8jETJJGEy3j2nnIuv/
nCw51fliVqh6SrdpM6HJ4l2+JZk9l0C3N6amaOedJagaT6RaDSbm1VnckDqMCydG
lucYtHmDUpCF3MNBZltYZfSvraUmB/ZXKksdLf7VVhgPr6yIrL8ARfeGlhKc61yr
wnHbSXx2oeXdwpDWIAeW9pXH7uV8Wa9ko8cst2wx5UJ1xrUAHgXZEpCnYW46tMzK
i/2lWUvCQpl8Aiit1qGglOjYgRlXyzYi3ePhzkYr2cn03V6/ZwCKzgtkaSm8I13L
Z/An/hy4QUOMXTYGsp9/ddtkv24EtYd1qNBeiuR2Ymx7Ha8Ajkzk3TYLbZgkBSI4
5plyBSQoZyo3D10HYUGY8BYxslA9iXxPYYMr7OK1Y6ohanb46QFthoVsFtosSwb+
+u5GwcuZ3zd1X5DNslq9rvj/pZuUSVcEeeQ9rObizRLOQ3l/GeouZzW/3G6TWwzj
SOuZyf28WcOhvisila+4ql4RNt1WGQiJ2X5ABpqAtgYFBugIqEqjxa1PtgXTfpKT
`protect END_PROTECTED
