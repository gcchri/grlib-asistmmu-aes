`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y1WsUne7RzPiEJOcPm9w7E0skLdSLv6kVwBLUf7EEEhfZOD8wKLJyw5Xrd875dAn
PvuGzaBl94xZJFF/CTkh+1XfwewBPmh0eBo45ezrshjoRcOeHRFTTcip1r+eBTS6
onj9f6TybbBFuvA4bbLbV9a1T23l/cEQCc3Mgao/pG7gNOl4a/hKvUSZAb6AndIR
8Nesmq6VPoZpykR7jP1a4jZw4Z1frtgmRbdRZco9WEIOrcgLiPM3Vli98/+4ZhIO
HR0F4x/nSrZ/Bnr8UKEAsVJVH83WZ13pU5nzzYnJGSRlnlAG50pBfxSi+T7HIyF0
YljwF8XqjFIDx/ttlvGrkA==
`protect END_PROTECTED
