`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MOi7N2JJSYhFikmC5MD7vdU1yf+F/LN9p/6TWXTecJbpBkzO2u7quBcZ+/t6QcIG
vQtDmMiQw/cPgYZ/TdkvfHKYYsv+JbVeUc6n1g8qI6ng4wdsPJdOPJHsRWJU4j9E
744JV1js19Am1artj16ztdswfXZAIRi4pqoWVrkPYsEQ9GK6OUeAuwQPbKABTaHM
uh+yAxukGcHFUhP5aIybcttuYZzy9+kiPfm61RixwsAFslolZCp6idyFv/8aSvef
79zRBYVvRGlqk0tH1Uuw1xtkq3lT3WTJ1yNN1EaimAznAUTNlasIiEt+UF7ARHnF
gvVLnZRfGpUhNhJC1pKSLE3pNKUGIuZ1jO54KYilWSaLNxhlNDH7Vxb+h55lzzVQ
73TVmLZduGJBg7JoS13ImKCrxBEgU2gJAaqg/+R3HRcQmIzGckv7D7Qldv1AnKgX
f9PNtjDNW2iYUAToSp3c81X9BMPN8fjPP5C/dwwsSPEzL05+ZNX4hLmePwh186RT
mlkWgphOJMfBzjgSdRoTkQ8M5aiiQB4fr9XlyM+xa92mzD7FVSkvsFlTQ1R3+dTo
sDmZI0PHhfGwfqWiV8BgoJD5Hw/B1HDcctsmDwQEbkKng67c5LMUyugLWvCquP9f
Z/IURx/g94aHZJaM2z/2wh5nZmp60bKY3gKhOGD4W5dRb84WMSIhP6j6/ACil4v8
yGRMszZRovvF09AbIaqHW/bMScTxt5YO6k0EjMdTs715Vw+edchXZn841aXTd/kp
j/j+RuqjR+j2jXm4w9AGKtbMnOC9bbLhKu2c7EfPaucobA0wUuplkrRv25UYblZJ
3UN69xhnCSU7W4iNLYhLeasTbB5k+3bB7akjwxKm/AKL0jiKxaWAQUxcVdNy9YTX
HIkmffCqZJvdaT207D2MsJlvNBkAHxUidvav5EAH576U1zS3feiNvM/9nEnj9UrN
NJbf/InGxQjZZKPyAwTQ2QsOq5odSMaV5Wv4u9/C15FJmmHuS1guKLOEFdimFACb
A2T4JJhx5S5IcWIBl5Ff9AQJN1woDjW6gk9vbZW+Zxcvli+PLuk9kqNQEjZlGofs
klyQ9enle5blkOGs+1p8ODhCdF1EaeKR+fFvMHM8Xi1+UpOqN3n3rTJe70VdK82I
xCMMgpENEqhZHiVk51ht8maarHt6DMOBE3HtWHNMo1GQecF9JpROjDd7dsyj7/q8
GzbryH/XsTrDsLwTzWVWWy4Rtj1Jfp8cXkqqA2X7YCszEDRhaCoA5gDExBBrgNM2
yBmDzsiUvzbHPMtpAIRk303K72QsFISTmOX21P5KRcIX45+rcyD5p3udU9/kPh4V
hSoPrLTp1AWzyXqX7jr+VFys6C0f2QGzuaqytF3mVly1POHOARnLmgniRlO2tLPs
/YsCKmpIS63k6m5Hlng6oXP2uJMB3oYILfDZNFhQb7bIWUo7nswQQ+n4KKAoptI3
k/wAFYceT2wt/KC0Iivj+QY2jq1GcsHnZ9r45ZMj0huos7qNjWe6x19NCJLPqDuk
mdgrLpWooCputgiwL5R6yfukMyOGvfqQahPb9tyiOgUGq9T6jWHwq4Te84fj9I0j
p1vulpSRLQ0LO3dYuaTV7R7cdlo3XIxaQFmWhyRXu8QgYR+oGd2EvPjQOy0+/anq
4SkuNS/MxPpBb6YQoMsiolQgYPwgJJaN9ST02BExLlt+/Lryyo5INu03Hz2wGb90
Azo9o4Lv77OO7oyT8kgblnkEsvo/tW6c/bocVJQhZwjaYnb+IFtu3tiVS/ceub5A
NMmVJgxk62vRYCsZbLgAOwez+f64kOO64kSZpG0HIxAB5Tdq45Hw97eOaFX5l2Ra
dsXRvKFxywkfZSxoCKtWDR4mqyMDf8lotrbFRo0zjv29MzTIKTVJMgWidVfRbQd/
zn2npSkhAQ+k35TBLGMIfE1wQ77yzWzlzjlOpK9ZjlYiK9o4Y8hRZS4ZVgHVTOc9
LHkILukiE/cLTfrv3T9MdZKzrbefQcdAvyOI3MP4+d3FQ5VWHhCwlnH1fTgvLpeC
P5O/fJHF5MLkIa2m05g/YWaFC6ZHxhGXKff2WQnBDnTgiE81XXB5l5ko7yOQiQcL
Mcs/kFpg2Ay+4c7xHooH5nwEAFUE2xv22oi/TeWkszg3w8EOETZkhSLvlVwaqKtU
VGWHoSIfzNkqO+bxOyan4SzwIa7TxXEEZcAzY+OO7VYqrVhmIrq9zzVSd2wGaIUU
vNeFmkOFedJWVEy4+JsejV9wlBhPFpkT3Xgg/4jGmHQgQxk8ZvbLkseK/ta6pyT5
rdI1BQaxoc+ZBtJfh70eWugoUmyYWgZgTKffgfghUiKQPjIleVuQw3DwmBJsQ9Nn
JPQNyCpe54zMWvL0swkQaHoX87Xdz8us4IhSqxiRw9PFCozyjGLUC6ZUQgpjTZ8Z
KPAt/s7AxgkClrvyDynOAgg35gRcsVGvzmdjkjtFHR19ZPCgllF7oTvJzk31+Mxf
`protect END_PROTECTED
