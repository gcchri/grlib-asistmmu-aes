`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N0IXlrkCJeeKu9bZfECtWaRsGUA5YwCYAml0eiqTZ225Nn4dOEZZYFomMSU2MxBS
LXxEHBggvxDdz9QN/+ZNZgaBm1A9GuD3Ra6Jc2Z9yize8YGestLJBhF4Ht2tVDBa
FDUAss3FWU6IykBZyNLquU2MqoqcWdtHM7Q6G/IN4XYuTk4X1m/FKJtY25aXiE9d
TUKM8X47J25+S7G08xlCyOqJjYBj0lPa51y+A07LVzux4ZkAXNjtv2vQm+OMvAKi
9rGId+QgV9q2tqyxiL7nXEBLz0se0r82XZZkNgWzCVGVKVRRqaQ7LZ/+GsdnztAm
hWDfAFqBQS9doDFhzj4ZSPsJdfOzpChSlZ/ldfxNbLcF68MeAiVNh66m0Ouh0b5G
L2bSKGgQS0JP82+2fQroiEguNz2wbEm0tLYymrAXDggQ9eyFrkXwsBaLB3mnMnXn
`protect END_PROTECTED
