`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vVKLqlWx8riq0E/P2g2esk022TnCJEvrJvMJFexXV46FPUbetfhIJsH+m528cqCu
j4qPVrhy75Jh8EVQzD/hsb9R25t0GQ+cL5lN5X2lyu2uLmG4yFENppHje8d73S6b
2ToGQVmaXHOev+UJF3Y7wlZjnJiyIi6xnWe4QTrILZpBwUqONfoGQOYnPABx4A2d
PEysMKZqSdlc44pdHPp8UeZMu/SKcN682+ZGh+Kn2NjJdcOLYQzl52IjMY5PlD5R
Q0dRcSS9+uDrIu1cdN4LqhsnBSLuK/Swzll4YAVgI+mX2ty6VQri1IQyC5QWwT5Y
P65kjmB16GJO444ElKQx2799t/A/NUjzX5oYMInvpUYrNAefAIdlKfkcP7uQNo1B
mOoFKUUbV1dxxl88aVXrpvlFGBKlSRem92blFVJuBapOPRwclDgXyYjndjSMokW/
vNwjnaGvreFB+jnzDRRs6/4800dAD+24YU/jgS+uN5nVq3MjZLBwQ1TzuxhzLlct
`protect END_PROTECTED
