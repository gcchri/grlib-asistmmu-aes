`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U+wwFA9kDQkYWyPXnbzf+M/uGDkBH09UJUkOLpV9+qgmPxtmTEbhcZwH45VgP2WN
D58CqUKFrpEFQFn9TrPpiqwBx9ZfaJP+IX3CLpz6uaXSLzhg1hN9lTzeEn4J+KVt
31sQ+8fJiEUZP+3wBCreB7cyslOKwAKpya8rYnOuJvsJkjDtEGUqOz0wP4zBtFh7
wKrSQvrVv2IEv5mgZnfG2KesY98T+h2x8UmeGH5sjcJGeHvB5adm2d/MBHcG+e8J
uZcJNlp9z+1qSWUzfu8bCXyA6QvAsWPSiSJ+QRpoGPnxdOac7KWd/UzPwpBaXBTq
0omVUz4288BTgeosI63lgWHtCmx+Kfdl9zrCShzIvrv2ihr5IsA/IL7FzFtJfCcX
D5ZL7v6FUU5lcEE2FBMtBMORzV9AzvLC5ARQLi9NguRmGsxOPEBY6as8ZjW9Ff1+
PZ4fcJltQNC+f1CGfX63Kll6pwJy2yRVQ4SDmy73OMM=
`protect END_PROTECTED
