`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rKjqzBUGmuLNpoMB9E9uCwsNPOZa5Uuoja05gBRj7zwRT6h/1xYceVo66gWRARa8
ZM3SaaSEnFfQQBiIAASjLRhEaxhd/85LayH/7+lpdyo7QpliUbyLuPqNo8RIT0mE
2AfcsLbNsSGtS6amrZS4HSVM89FVQaoulH+9LLrnQCHUPR323WGCuXNVzit4GIvY
LYSmL5nOjnMOmMk0KDKnFr2ncehiNsswPh13jMAuEq+eG8mst4pRk5cUkG6Xnomq
VRSrmaHa/N/v7WXiD4aD0x1gsLA2ikFRfCyFcxwU1kz0RLO8liBSg6Chy0InGcpO
qDxHeggtkW9rUGRGxLSxSvmGwMeBK1nL2GJdWyC4+PgqNHsQmCBJfR460d+1a0hE
39EFGXccjWeo8+1SdBgtz2Vtqsi3qDSXZyY9sgGIFrw=
`protect END_PROTECTED
