`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YCuz69B1PkLI/YKZOxo1Gp8eeY4Tmd/2SUC3N4lNf4qHB4NxUZaYITp95qBJpjEj
inH64xV4hlsPjVsy69tKbzpmcQitX7b/D1i9DJK8RE69jBWWsJDAh7N/dgE4AAST
63jbIAxGRWG+w0X3eApMnRfqv7w0ZC60dZDmBDcyeE6IkZzw3FCJXuPca0f6Da+m
crnMQEONSxMXWFjpP6AObihPtj7VH/EkwNDndHfKZS8ehs6XFr1U5zfcf+RzArfi
FROZdxoXdoGWcoK7p7BZj+Y1aGr6bASZM7xVE10vFXa/Ik2JNfAwBtoTCKNaEMXX
VWQ7L+XsWv1y8i1iNQNgOcmwkDe50pMwC+ir+49V4RVxkhzX3V/GH9WNTwO9NzHu
2gpqf0hWj4iqf/saHr+I1iidGr1Bp53Bzk1xUC7rSgW9vn4fdZPo/lHxeod9YDdx
sfkHwEfPnoFdC23S16+TqMmhD1+VaiY1d4iZPUHPoovJiYXufrky4J4pdWgx4QeW
xouLJnpTw+9DwA0MCcPLylsdZKjpr74cchAN3eIBTlLhSndFagAd8V6uZynl+mQm
RsEG4mBXnfgfcGmNL8XaxL6Ipvw6mAZrGCTLfcOZPRvA1ZYTs70X9wyPDryBWTf6
gUdloKaKehq8KYqw6EGSAsVzb5NpW+i77TaaOE7YoV7LnH251+8gwCT3cEs9Z4Yj
4IckiMio0mQArBslJk1FCJQ7Mi57DTmDPi/e5dZM7dtmeJz9Wy5dR+d7pFsHm73F
6mzL3hFKG4C9Ag8dfIvC3BkZ6MMdYoZLKq3dTW9R8ykILnOsXmu0pn/5UvA7Ydyi
KnWYT8rU798kYg1LSDrzcH59iRhC7wjxsiyG+XRN1W+WuXU0uIcWydOxK/ocXSSP
hRUZ4DFbHxyPZlmP0Pdh06MYA8WPVaYmT+x0R0MRxfIU2UkCJoKb9Tm5vaZ6mB3Z
Y6RQisS8lCIbEw7aZAW/AfsEUlUrpXej2ktd4qk8+OpdDueFbfPUCU1b3rY3ZoWV
gQ9FGDZgM1GpyLoxkJfrn9jeNQvOFJV0+HNKvvrTB3GZXyeHix+1FyDM6qawVy7O
r02gSFXbHy1uACiDP8Tj/W4ASYwuUJ1LBXsfhqy3c+BZlIshtVQbwyUhMxg2rk/q
CiCZjs2geir8izpKm1ihyQMJxQ6urCIHy0iShZ6JRCx/GiCNhCXfuAeWvsM57zvf
jXOgDBHFRU3I49aaJ8GQDk9bzQWCj173fNH7gKi8mi0Zs73XRvbA+AEI4dSKc1z5
BNjTfDMwlS02ZO9VS4inNKw8dXE/wbN7Dg4q9CmYSgNltvgHuBEmvBP0Sl4LgMlJ
8JJOjAPEgArhfnO+TjtitXyVJyQTyzI64FyeNud+gBEsWNkUB4gJKiHpBxgZA0F5
sF03+ISbvf11mtH+WyaxQ7utKOJgBBFUrp9m40G4MXggb8S951QMnuA0n/95bgBO
/mglNLtdFdqL155mBCHP7RDz8NpLuDcZCb+ZgH7lCSLWOLyhJ1JrRTAP92pJgtcS
tTYSY3uhfz1K4BT80uTmHmpBmut9vOzcB5T8LZuCkltSXjpW+7eQM4zmQxjkHkDQ
Y2cGEkwCO3y0K3aW2mlsFSTALKvvNLbGbM5jTBHMZqCv+9Btw1wLnmkmUMU0U/O0
bxovLQjYwxhuRAfxZt6UaJiA+BuuB0/RzHditaMV3P7PXmuhrluZ2Xd3TeOwHwvu
LPbNYrpgebttm4DHo4ltfQ7o7fhxwscqLNu4LHuUacIM48JlJVwW9v2mqc4/BJO6
Q17hmlCQIAy6caEi0cE/NryfmI97o1woQ81HcJrqPhPOHlx0RTSniYxyh1trhJsm
/aBIz/jnQP8ZkArAE7YYeoZ6j4Hq5jcf22F/LLJE9Pf/Sbc2dD4dAQPRL2djohzt
HPELbmLIvOJ/wY25ApNOB9LY3Tf8TKDJ6WVvfPiNm4+lojuIPNAXgKTyVKYFTqWQ
vGBY4JFJKC8cCbBmko+jbaKHjrN397DuF8EjAzIAQ7BhqqaVDF9M2ovdHiz+a3CK
y4XQV7GTQmEDTTB97tfZSQSJpZEK7nL/nGT+8yP2QmDr4NJ0QkmEiwwL+Yh3cAC7
S4b3ML6mxEAotDS9Z5y5dmFIiC6/C6CPORonfdkFWf3TUN+GSGXCgYyeUc9JxhkD
vDzuRn3eUF6cdBGvvsoujYZbmoGtok3sNqkirNVSyzvPoX++DywwasfdocIpF5mV
B4unNvY540RSLTg/ogUbDRKeg/MLxe+GMHZgmHrTTRxr8t6n56ooAHTdGMsf28Tu
XZTjPyVr1Cssg2zdDc1zvB+vATHJbC4YHJMX56j97jK3prP6OrmkRExlxZqaz5KY
/beNgMFADyK+tSmsO7VwruvV3cs+Hlx7DVWXnBK78zoC4kp6LMLW8hmlyRtzFGYJ
0+tIjSg0jVQWAENJUNsXnApzqAvUNa7YT2e39SdGRFrkB6ujQAQ4gUsGK6BY5ADB
opV050ahCsrZHJoHdZA/uINxfCHQWn8gcwRfSbHHkuZK6H43uInx9k95JzsIUje8
hM4c58CmrsfEaIK1W4cbotus0Z79anYW3AcsLJT4PSJCmGGUmO6E9J8S7iPpcy56
+qfUIqQQrgBFnHypqgz2n0rJwf/2Rghx35mN3/gtlg2b8ESQ7Iyg1JZbJ5ZAlqlz
ykuDGlIZFOTOuNXt7AdmmNvFGDIBO/xlrKy6BpR7F+3Trq6+n0TqrHsotMoanVLG
vqlxSY8Wc0zXadRPkcj1rGB5bBsxFVMy62LXSSRBjNqdOQyC+ev3oieiZrzuGOJm
Zii6+9QRJjEwKd9AzCULdf66FlG1M96IWNyZSlVju+zMy/kiZXAT9shE2BGAgeF+
AxAeDzveNUo6lzW/k0CG//QISt11y4LgZ++64YpttmgMJMmVHHY3CEVC7rKm1jIt
nYl5m9I3m5XLA5c3/DpdoWMjWdFMy/85U6ymUGiuhusrk0+KrfSRdWMMqNlOJhld
0ezhzeYcqtarLxzYie+0gT+VjLeTCd8th7xsRbAj7nc0rwg53mBAdDzOeKV3IBzb
MAI8bd/JxFgIi3ANpGhOx0aZ/RCKNJ7jqGCd2ZpVH0ev7W6y6NZp5bZf6QWeugrS
Tu3zuIH3o8fC3ocHHrAilqgrg1I09fKIT4J5nYLdNY3sDkxeVKwBbhUWMuV+M881
Or/vB0226uW6gr7RWJQyS0kl2CEV7IzYqPN7di2Cs+Ck1WK3hZXfKK2zn22JFA6C
`protect END_PROTECTED
