`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I/GqFg5/XucqYnv0QRvEs2SI94r/mgzIfZa5TNVDmQkU6FPRtOgSs0mJQOyvd+hy
5i53bnDzk8yq5SOdwVmWrFq+KTuVpp/beX7oiqMLo0LSAlBHV8h56PW5giZI/27k
8xUSmhfFfsoFsvti0QLznDZJNdNjE4OeHvLm2+hewHxXLL4HYzAo81YMVM/yhyIY
KEI6MU6YGU6fv6ApjvNwePlkoLgOCgKQD7+cmPd8vobDm8GIVwFI1NDriPp/AyQ1
Tpi5POJ5LTG5cLEQEJuIe1/y7hvCAdcoOvZUfF/g6jb55t7s4unG/RWJG7z4iUrC
m2Zmve6lQM6ckPwhTgCe3qeSWrZJocHy8KQENWFZfMP/OisEWMEG4D0dvnxa4Pvh
tWB3xLUrhbut8GTM+o/pbUa7T1KosOovBHtlbBKvh/jgiBu4CHudaz+WwsPl4+th
Wnou5Dz8yFy29lk+PM92bHsIDf9IEng1HssxNSycT+MNI7+/upckc5Qy3TUiSgao
HPctJiRXLBuCqgAp25XnhDNQsRqtP6KnEAL0wJicdjTiTSTNUcUcIEAmpjfXX5MF
M5nUyjKFVLtFQOtWWoLtL+Tg+Y1m9Q/JoqVqoFxaqhPGV8qqA94fcHzw4SnuhYUn
rvv6gnHhLTyiKzb0Mqbn9HmNnifaA6ilYhXtva8qHmmveCHRypBkY+1cPxq+1lD8
qB36/vbH36eWST9kt0V9571IdLKe9BpawrGjBWSUQO5enqUrqlu2xYUzl92iSpQj
6UAgJ1vTwI/ITqsW5v96SvXUt76jtmEkIFyTNu0Vd16l2Qfkm6f/U5zTzHwzTmGb
Qk2I/GSxZRUK1ksrItRoCjriAHBiD6eZbSemfA43S7QiCouQUiFCagA9FEkQwa17
ldT5yDSXiRi5lMVdG4TJML9fkqt62Lt9H+MT2iVOGgyjDJNzbZf1tEV/GXTZaARm
`protect END_PROTECTED
