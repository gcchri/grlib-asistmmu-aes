`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ysBmbmCJfPdOTaeBZ8kSDM+mNjEYQI9LLEP55Ut5neBd/YJR+axhtgmwDv6+BTzi
JrGVHEEVnV2I6Wf0eXHVf27Q1MtjRPb78kV6uBR5W8gfmBeXXkhhAj5zK0EwjGxT
tOS40VXDEnqhwUht/gti/G0fxpWF3Mlp0G2kXKJDBNii6PBlw5HC7Vmygd+VdpbT
Da05LQJJ4PUbBbcLkCbxbHeS0HRvL1ODeZIIcUH6cRsUQUMVRwPHh/hItTXSa62T
Tynw4yrAIB45K5kTLJNbGA==
`protect END_PROTECTED
