`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b4CFsYbmHow0NHocv/dYl6Dymr8GI8rDIs0EetQ4dwdCnAc9tMQYDW0WG0xL/ZO+
khXAENebxbYHM4Rw64FhIKF6XM/PfGSg9ivWu02u+6AJYxO3YJ4r05bqFo5Z4Cws
ZXfvBk4/dhEe5jC3WN9ZbtQhMAkYx7JmXuZHMU2RInZsp8uop3k0U3u5UdP5TxAe
2GwTbthb7oDPvNKydygzFsmxw1PtrPB/+11lkVS3OQ3MNTPF+hCmcDlSDOhVRHwx
0FwLQe2F54xOw6nSrTA2lMo4X9wit1xfgIRql6G+O2WvfN7/hs7j6OQMn5paYoM6
gjtM6wg6JNJKvpZaBLp0F7nRCzMhCVSZS/R2TXzNYSjoSDyOLX6DWyDm0ynX3f2T
9BCU8RobZuYkddgzy+b+yoAosOhfJf0+SFLF+tVxcqP2DHxhWa6KU2XcVBhlurDr
ddOQX5POkKeeiOgIERenWksxvhdAxbeyxHxAhUl5dAOQb+nbR0kwO13AM76iRSHl
IIpLYeWhF6Va3FFPBkKO5g==
`protect END_PROTECTED
