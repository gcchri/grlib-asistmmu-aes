`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lW66e8UQfw3B1C49rvv8CAPwaXF338LNFQhn2ICCKnBT3dnkIbL7FSbCyXihJQuz
z9z5Da2Gd6HCqDqa2mK4rIews5d0xpd9v6JuF9axuumHEp+edjkH/HWQgrfU7ktW
SYXlA9gDAQl1c8b8tOMFqaHoxc053i7imMQPj7zZy+auWamrKOLBMW6L0458MVp7
K/TFxEsA7jzvCvLDVUBwmdYMb+si3FL71b5OQ6U30bmsEuzJw4vfF6vMFKvngvxx
1Z8A/+8KXHzAoH/0tbUFv0dVpNs2TFcokC87aXQa5mCWu8GY+PnykUqUdKo0Rd+m
N/0uBObmdq1eUti95sN6rg==
`protect END_PROTECTED
