`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vQ5rpuKPz45fRfXLoN7OsxsClReG+ZKf13NHkhy7vUz5FmBlnGkjUR/Pghbjh5Tu
i1CMVzK4+OrX8L1aImO+bHP6N9Nd3tFciXUEwckK0Mti+ZSVdJT6Nh4mjgeBaHk5
5Uw3HXsWaXzK9jNgD4GgglYSWiYpnP+uFyrqZ1XA5Y3go0gPyGdaaJMZT2P7gfGb
XNRf6TegNRwns2ax7/1x5VSc2dKdMZPUgggZgFBdrBe70m80Oxmu5WIy4GJHd/b+
MVjXO/AEQ6I34Bc0e/kf1Wn4YmXRd+8WxuZ9jFvBVEesg78yrynUENk/Z/cRPHi4
iXxi03vHq6whmQkdvYe/DvZCSFgQjgWxd8ZmHq9wmomSaAffxEd/yGK/yqC7SRmD
r+NKIAo388kCa5pM5sXRP5Y7aFTamiV0I+hvEx7MSMuJS9yGsar+C8PoVdtWp5GL
VrNOeUiYP8VrQPX6k21JqhpFW+u1rl1qqUXyC+fH1+O9hEhps85ipOBeldZYAf3R
O66e/BQbI9Jf9MsGPRB7F4UxA97XzC9Y+loxytT8Ud4cL4TIWrlfx2ADRXuKlQTn
r36jS5X4u19unmGU+0devK21esCiAANBNSty6gO50Jk=
`protect END_PROTECTED
