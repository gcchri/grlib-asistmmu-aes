`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2OY6d+y8gH9AD8jyK1pG5aTSoG8pNRcLq6nW6hO0p9PGTTFoRMaejl9AuVmOvzsW
b0bwnBWXN6wbIgjTtxpOOncOiV9L5HVd8o7tOnYtMzz6Ndv4COeSsuZwxea5WkWY
0Y34cHfTJfZrFbjVBNwyWcgsWiv4Kf66lXlRqWs8LvPZtlqC75G9SNjUoA95mtjz
FSsrgvDQc4FWQGJh7bAmlPqY5ji1LmAhdTb/U9l7Q9oK2QNYwB+z5pxOyKOPzgp1
TyRv2OjZqlyeMuxqlpAx/tkHnVeliOMtSeM+PeTO1IlXDvlxV+eFkKYNme0n0wPQ
blDPZoT6q28aUn2eXuUF1J0T8pd41yzZ0i0e9eoQA7vMs70jV4oRkHWZ9NKwjyCo
qijzGj+pcy+Pohnwt6x+oNWH9egV3zeroWQLGVZAKEGT0vk6GSdpKzCUs+BjwoRx
`protect END_PROTECTED
