`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oolW8WXWYIK1BNbGUIjMwowcFiaAirIWPOFmZ1jh4/1F630haFKgywClyqpqpObn
FVLvkXJ585k+2eadSoMP9Ko/Z5krnpmY4JBhmxGSrFufgu5ZqqVRqbuD/ZYq4AdF
9RHEIfNFaF6BfqY/h7escFAQYpmeY4DQKc+pXUqOoXtlJsJUQ9Mt096ZwDVIWbmD
+MH36OjsjzrJjOCVyY0pTSvXF09s52coz/gd3hF+xYtUJiHtQRTIUjGzuxToglhA
XxCRxFoS4eA3cHY4Lj4+H1gAVFKhmWnZsvOdR4Rd9rXmqoNm4FpD6ITITpdaVrEP
OAK4+dTdLu23rc5Hi9Nkk+rmTfdxUYs0ISqoFJNpaIWA1mkTvWuSXA+NyV9J8+x7
tQob4o5jiSfvSlmZ2XsX82I2RYwTB4UyfelI/E2KgpvVkSttJewlpdKLLvdGDCuh
Nsau23x0xF9TYIkVyxrpCkvJAaksl8vmIOH+mODLEGftpf+MmuUSsSu3WoKo/ag1
`protect END_PROTECTED
