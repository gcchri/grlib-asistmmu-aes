`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K48mjd781lDJlR/II2SVusC1FrIl2idkcuG4rwlpT/j33npNB76BWQdSAmXYdVEk
3dBhfwlkBNJ2QaLMDNyxgSP9yR9IuhMpjNcOI+hecNenzBRYYiZcyN6XGSjfmIcv
rGzhjrI7jCI6XO/UuTp/hhuO2aVqG7i4cRWTdNqAuSE6cjM6cClmDnfc05QFmOPm
meepbH8BiNjBoHdUbQSnLwDfnUxv5HThSKdYb+4qJDPAiDxE2hiXupm5vfw0XC0i
0fKt6Md8GbE8g4pNndAFpb4qKSYwBfNBBQvxgIjN9PEjWlY8/CSQfuhJ7w67bZvw
35IE5aWYY+CS12uL3IWwV8TJPvF0Bed570zhQUaWe8psP/BlmIsGQ1ufMJ/uVTvT
ia6WJvGUHBXOtwBXGQw898Ial8VcFoP57LyVEe8EaMBQUzU7+3Q6GoTLMKGdAsPX
FYtZffw+PseNH2QJGoLzQMm2bACvXzRRfPcw/d2dji7vtoekWapmWShl7XcGkmlx
2TdtyydPWFrKcNciQewFj9QGAxora4tr/BuwKGk/XZ50QZ/UAMgV80Gf+GVKbM0m
PxkabBs0n1T45uFozOBSS96eYgTEWxoTkt8EGWn98+5bw12rw60DF2SUP2wZ6XNd
/wboEe6uQSH8Olu6Rsn46RmFYT+eVzNNdhw1k0LQS6Vx2BCrzzxq0kqt/eOsoF+Z
suVamHTcW5hEVY9MpbVhnxDABun+et/0h/TtVTxqotA6fB9Kivjk03DloMsw4ZXk
Ifhr4z8eNneeQofOxh/fJZcyhG9SYqE7sWZbpzBrpY4gpppZWSTSq1GZFKUlZPC6
gLEfRZe9Qb1PCbYfmMeqLimONIS3ytDrbq8YZ114TwrVf2h/Y0zMdagiZiyo64O3
6AxCaVjKrKaqwh5RrvSPwQlLKcVStB0bH/TZxaIREy+G2i+KIdOPTyqQ3anh3Gu2
Nk5BfmE8DqUhVDv2sk6Z1wn0ItZLZhVnOPTzZfgd/LM=
`protect END_PROTECTED
