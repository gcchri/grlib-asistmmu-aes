`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jC3zgDuf0U0FqPmtNoC4ijHMPjtoqcxXffXu/mnD5OdLnuRvNipy/aw68vhWyXAg
KEIRi2CLXY8Px1rt8pRznJbLqbKhKepQZEUtw1QCNfp6fhwFdXiLjyTxM6iVpgcS
chmLkYdmPvU3GIY70xzP9yqKlGFCoLe462jpHVAUFJAQ3oJSMto7h0NCCvZ2q3PB
N9tDHPvxWE6zsrBHFBBLd/TV9xOrvTMfWD7ELPMQABCLzwWHuW3HA1YdQlUiddyu
YHo0snmIcdsA5rbjn+zZV18xG6MnuLVdWfMLX/wEk/IIuR6HZY+WCLxF7AqtahBC
NgXvq+h4g0YPk2MQcDoUPSOf3TndUhDF3mcfAgL23Mr114JL9b2uGrLG8wH4f2wY
xyvHlnPud3h2mCvpmuf3w7e7A+TemGswGouixT++It3HJQUB1hn2RxPQTqMVQG3t
INGpUwX24eY5usme7UdcjO5aFwhqxptEWjaE1j5Q7Y+02PCv2QCI27C92BQNrAbx
`protect END_PROTECTED
