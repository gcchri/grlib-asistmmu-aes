`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LWLKW6CRmai6p2XUvBzRVLH5zwr6nHUVzaLiIgDVveHJGeF1bFNBHJ3r1MNuTjUr
OBBAQpza2u7sVlj/+cpDqaeZS0MNMrNnMvm2O7tal+Q43tltDDarB8fqSbS4JvmF
y20RBOT/CY3yP/xKg28KSAm4LGVfdLVWFHFlBSUgD3rZCoo1n3QAdo+d/amB0bbC
+kfIrpXRX9pq4uANCk7PPERGUM313Sz3wlTYrb+HgwHOOSIE3V8fWiJWksK74S7o
WPwdVY/91OurkyXjth2H28QtzklqOMskeQsuN6JpqaSEdzd3/Ko+Qb5DrytTU7gf
TiLGlYj5f2z4Da6nl4EhfIMsdc1bdFmDKDO34gBQLqLBZHE4ngmgziqFnloqttHI
myznHMlxDsesH03QEgFkiILT2ehgD0GLu8T7pxNE2+r+XXrPkwfnc1pc+hxNnta/
BcHqUnMltdyRF5esmmS+YRKTZ37SyQl4mTvgGqLjal6wHM9O+2bO3zsyA+pAQjH6
x8pN2JGUwUOM2eUiXxhS4NEVQ7UPJjv+lm2SBfIsx8hum5PFuXnReVAWdy6uVyf0
`protect END_PROTECTED
