`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RuvX89UA3DYyHdAxSJ0Q8jxGVnsm/VWXcejstc/R1noVpijvXePHniHkHDBdGbv3
6vDeK+UWTL60uUPjH5gYh8PdOKD6b2zgdf7Fb9zd4uRTeMeK6bRLQqTOdMl5NkI5
cUsdZsE6iVwaoNcyor2GCHOzLEsTjCy00wJFp7cFjQvnrE9xZUgpHagTYh0JwlDD
s/PR8vlTOSXu2sw8ZCICCCP0Z1w7TLQnif+2OsrNz3j20r9mYKw2efEIUmd1D+df
`protect END_PROTECTED
