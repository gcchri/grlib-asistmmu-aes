`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qTnDyXE/g2cholxjyEwxIpYEUeyyTwAx6PQmcODDkBLdie6S9gaVdeRHq0X8wok0
i+oLnDsjQYxmzvXmFLUApHnSbIPS/b3AOZ2aORvzno5arc2w2Ave75SDbQT1TIiF
bAAGK3ZXDKBbnAPKGzXdQKGoXZwPdDG/p3p3uIKs/jP6OjU5SoDL38dvB1Zo/sKF
zsrsvtNhEGwEIBYZ+qPqWkCfLyODj0SFnZkGnr5aDNxx81xMQXa3rBNc31kzJIYp
WmQ6SvxAZeQkepXT+ceSnSIW+l4OGQjG/RQ/bYcqtwA97OZILSflAyNFe/tYVGm1
+BYM1yQVZ1Icgr9EGbFFhef8GR7qEnK31LE7Ct+X/im5vA+6Kt8H2Wd3GNCm2fM9
rwV/hYW0Xrs/JkXJfj3BD7SZN506CWXWQzeGB+0bCv879fdMt7Bd17c200BPeqK6
eEUS972j5SJZBvdxUM9oFBVGGAY+fUUgjhS0gBEXLqI=
`protect END_PROTECTED
