`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7fwIOQ/CKxp8QmhpHUosUELD57O9TMIV+kXn7DE8kWWfYvPbPNadH75h3MuI37RQ
k9If8iDZjOLSMmtPLQf4OSaTEHyW/YWbMBovQrhgdPyCAQPTpvNtgyZoEvgQdVZN
bsiCQEJticRWd/HJq0xBXSIZ8ErpGNNKPiTuPCkZ1aEpgdJ2eN2PwKeTNUwZ1LhC
vW3C6nVad7t5Hq/ngSPvs9t9HKA+eSwMBVzfLBtSBs1qPRhYCmwnWqU5skYAH8ZC
bW2wycW/sCaa5rLCK8J1SVWB5OOdiQyS1uwDYRSE49wSKJzpUPQsL1s5mZ56gWd4
ytyrZE09BTbrvAzwvmvXvw48nOmwBd9u7wNijpkaJqEQktamQc1YOyJ++o83OOrt
Qfel4lo+O1+cBNvjeKE11yQL7/iy8XZ2hVIQCrPEBM1fukavAbJMdx9KPWzl6m9S
0ahicujN1xb2vgp7YTkgWt06FKaaRl5JSnn6z6wr2uEWE9zK3/C8d3abSWROucJW
1YJAx4/K6gFRVvkrQh5C2VZ0Wm5QFYfZeDZbwGz1eTzaiZiZQXt2YnInzUotdTpC
4wg1LZCgQLwOigdJ4Nfz5TZMbYcPx6JjxfIynPYluSI9bo7yryeASX0evHkU9cj5
uJ6YT9sSyRa+Z+X3d/Xa+B2UuyZ7vqynJgoFVaeW7oiLDdWea7Xo+UDhLQMCCx7H
Pk404dDNS7HsTc6nANMmQx1QSRrHEVE7hR3k6uQm/9Q4yw1lJzWygWW+PZbamzTH
xk46xv4vw+CniCVb4hptzvzj1BXgwdlzHlp0CGWtjwk6hFF/VJvtTt4Vu/PLo9zS
qeDbTkjvA621oxjHlgX1fqtLhSwpMJpqb+V+BxzSwI/ZPgAme6GM+dz6jL/rOW4d
gqBB9WHWnmKiHJMNY5guIcYmhRZBj8U4onIu3xVfAbXxeDxPgeO9H8rhbYRxZ3Pe
OeZesyQw7mSDidJPYg7pXlcsChAM+3tqCEZKNebAxBhu0fmro99vD4O2mvKMvpp0
bVLEW7ixpjqGxvMZ4viCJwyx9dMi4dABgutBntx7VHL/QBTqmLsqLuKtIEMPT+YL
wJw0VLkd/IUjgz1v9FAu4dgHCdW5w5cQm3kWlGz02MhU9E9xFO+FiuTQUjI5rB5L
bVlJtLZeu90EYVQWUu1PJ7fYcX5MtuW3zoEQTJjjFRFhI3jY6sE+BBgRSojBBsE5
p38LINe40oHqXsq674y8Pp1AfYWt6IsikE2I12OHSKcLgFH5w88KHe138vlV7XXg
42bSQ6HAf25v4TU8u3Qco/6lwpbcGA0U9d03ey6nk4DZmaz8wq52j+VUm4JegMH0
PpMe78UvEG6q4IdTiRYKpe5JQK0mK+6De5o//WTX5XwT5pqpXlbyS5Lq95QXtPPq
jvEcuKeHq8VWIcT0JoO4YVprTePDuY25jwnQTpvfCpkGw7JU3SrzTCoH77tuNxSM
wOlIwiUBCfWpe80/1CGoyN82rmpZh7PWJBnVTFK3t6UFYnAk+sqYCq/tXC7siJSB
zk1PZD8Hkun6whk/5cTK5akYnMIQUlnN4B1+HVGdeFJY9/GW7aDMEV6944PgdSJ+
v/XuGSeFpLTLt1h3eE5I1lPF58yQlyr9SugN5tZM6IOyuDSkeIbTLkB/QFQKcwyT
`protect END_PROTECTED
