`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0yZgfzM+IR56eEc/4yNPHter6iIXHG8qszVfCm1f5Uw9bzpHg4KHaJ+KvY0h3yhD
rCaMlnaPw4Wbhs14HH6r8AoGp25/bOpBPvgHaseGmiESReIRetMQ9fQTSYG0hUEV
rBznH9B4mnjlYulojTL4vcFPWqrihGlrLe9nV2oQwCUDpdm0S3mVjQi/U5VvjKpl
AjAFdJ/XU4Quh18CRTaxQ56N0E+llhhFw2Zu3AgEJt32IwczEvqGHYjL11bRb7QT
RnBro2YQ9Hkf6WPfZHmKNWtIWuLFXOJfJuhUd5Ds/xUlcYo8JI3QG/wT6uriEzRp
dxROup0cRC1IJeRw2kQM1Lu5KcK6AhBmcFe88kgRHrOeflkkZsm4iwuGTGEfN5Xa
UxbWP3OmujuhqqsH3/+H5W/jG0jIhIlb3kl25clceOUHNvcfDfVpYDXbaeWcrhiS
CrPv0Ki62bEot+aw/lh945bNeRTnnJFLtCb5WigOpSr020rVuMG3EfTP1njSAnIG
kP+wKJvqeOdEMxwxuEE74dT0MMHHmy5OKKkk6tBix9q+w8bIlbR72m5wCMrMOv6X
TFv+8T6Fl5trEoYeFjRPqRSFe3pkX7Sqxa8Yv5iZxymtZxbU365YDyN3QHYdLs8Y
xbmFcm5DMuuVaseFrAl0e8oPqqkm+ngLpoSsWEUbsTWe5+JP7+lHr2gg1eiTWW/F
j+TJNyZSts+y/HUi3jzWViPhRnkyMK5AFUw5aR0YZKPEXTsq3J151APLVdSslUas
JwMgiEl1oKMVLLLvqFNIw5/tqPrU7g2f4kMMUhlq4DtXQ83mHoTv6SjI9tFEoKPf
P+vgZloxL3/GkIxEX++F09oLFirq8Jx57NT6sl1c72LvLKkY6bfiKOvVh22e7Yuc
NnNKHTfiFy6tYqXyvF2LPF1258zMYnd9NobtqBAwfcw=
`protect END_PROTECTED
