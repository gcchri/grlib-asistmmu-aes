`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
03qb5VPfdSZa1+PUsdQ8ARr2bwvQuiYTtXargmBhGE/aPNMn1BEvCbPF6MhDSpyL
ULuGV/B5p44fAlHUzamijSBm124rl23Q6lRa0/fBglxochuOk/k/FfaAk2WgMh8E
sxZ2WOGjbp7IThoGXGnY0gWrRPAFHLi0afVPXi0ii8tvDh1Y3Gu7ML8wG71RjHHf
XmwvIsCFFacFd6bM7PzvcfPoHS7qiEZvFVMziOV63JCyqWHgumvliIT0K0HXHiTE
1QNrrMdHvDT/CAfjYq8cEAvoHWNZPOxZirGAoydoDB7Qc5qbpXjJ/hAI4nTD/nJu
z9+hbrBDCNTo2Vhxqa4rg4pvMv/WFz+H/8k4CtP37sZxmOA4+ZIpfEq/VqCbU7fX
joQuHDk6ZTW5rPoTuCyTmkN7BYx6/YRYKvaBPME+kUBn2FInFr8iF2HARhyH/tR8
1/UMcd5/tkJoy0ZsMDo3RPh5L0tBw05oWkWjhQDaX/8=
`protect END_PROTECTED
