`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hBs4UilHkhWhXgmWanYcr1gkT0D9EIPYKpyv5TF6WUjt9rg5bTEMh+n9geVabjFP
rl7SJcoP7F1/7UiTVC2z5T6HcpgipufiuhNT7gzFEl9VoUFVMsddxZ3JlZpthzdS
TC7j+Lt7Btj/5fhePpRW5LvWdEcw+nTAPQZdK8+V8ibAWL8vyYCgalOEkZyDa6pv
Nxf8wjdwe97JGYpiAHi6rVofOphH+IJUiYop/mh5y82J7Y9wfnB81WE/Z8787eil
28qyAhY7qGzd94StIxHVv8gaZVcSwb8ZdCJO5QjIIHA90OV3HZ9cvEm/M5Mkg3f4
rIia0fN38BfLosvFD6W/DXCd97yvShXxYgwRzbBqg2ZHaITiP1F0HdxQWueV6KLI
zjml/jgvHyvwpyR5ry+1hMqlSGwijQqe6nHLYqWuZbNjWG4J1gulOepqufTAN3yE
UcSoLLb94l4ByOpuvASRazaERMpPwmI2hP7VAAcr/j6guDjv4KPr8D8teaL/6qeF
`protect END_PROTECTED
