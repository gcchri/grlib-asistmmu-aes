`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7OWqd5i+xrm2a2nPvj0N2jvm6Y+KVwvyCdWyZMQan3dShITV2/wZiaOy3Y3y2an0
G7Di8elsrkEVUMtkELcnCGxnIgmMNqX0aChdrmXRNYyg2sF13XlOS41hneZ5QO7U
jAIgSI5wrW7z2uJ0Vc49+trpB+1GPuj0sixLtjeeSCNxoV0JBvxud0Df1Si33JTc
9ZsQrhFWS32yLfL+aPfBlMuDjbZMGAk31KGRMWt0l5VN+OxOcY85+wMdq2We+0D8
q/e4o7i0JzxfCI2u3ZBqSTfUanSvI1hazg+/nKDTQNCf3JyUSGSzNq8RtM3iGBNx
yzCo+HA5X7k7BJ4AkJER5TQFooDcnkSMRJQuC3uHdfVGBFx2D8iCRj6sx03xOaaW
h/EJx81mygyJ2ssjsXh9Sk5/UY7CrSTyUW7ZPBYOFmQefQtphmi6QAQHgPXp3JVa
eUBMSwilxaniRRgwBDRLVg==
`protect END_PROTECTED
