`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1sjPueZCjKBuVaUITzlt1Txo27KwPAH1VMS6ioVMEhQeEhd492hJ4PAqhN4Sea5s
Z4nXnJxusNuB4SHNHP5G/MVCmSxmucciK6a5cdL1OXrEW2HTiep4RdHMviVpK+/c
pOo8WDsPv8tPIhMLDcNmg/q94sHoKUOhogzhz3xKS1EM+H14ehIPtPZoQxXEdwk2
XDIC5x8EliVyWgz7+vZIiMCDyDnZ4JAJWj+58zEVMl+gmZHo3YPvv0yYBHxm+DWH
Ge+re2/V2n3hVQ5w76H9TyYZtbIfpjFwDf2PzddvYniwr+C3kS1gbUPdc0MLRZ90
Auo/054FUgfC9Nvkf/Uk2KBw1B/vkJEif3HoHNEG1W4xvW2t1rMMPVUOl8rAeaQ8
4PpiQivfbXCoN81j/EfVbDUyQE8b9CzYNnfwW6Vllsc22VnFQC+b5UpqsrX/ziIm
0JBMlhcW6EVPqpQwZP1asXB/FpavAH1FwbUSeUkFfFw1MdsIa6hNUp2snMnC6kJ8
uLruzisujcRm66x41gAJ+RFWJligZcv5iA7d0jxa/rpC85yTMIwdXfYu5xYfUYzJ
/wqctnYKo9xy+ho2LYIws/TBohN7K3jt30vQzoXJqAXDQ5mTmiLhZ35O0fOpnLE9
FsoixdaEA+QhavxCnqmln4iaXH+Ts+51hs8LJpbJD0OXfAmC4zFCw3/9N2Jdl6/T
G9e2VVA9LQF9QBVfOxn1lVyXeI7u3dAQQdQnZ90KJcL5156Ojt6Cj9ucHvHY/OQx
YV9dFDPw6ksvjnWam5+OY0tnM0xoUwK+xdeGl3YhLHQ2rZkgD6sOVYOF6cniC8gj
4qvg+NyzS+JMwnXFCWijzBaPFCiz4vWt/PucvDPT7I6bP53MTGpm2Vk2wZtl2ffi
dB2JW/daJtAsxZZIMVCpuez73HLSsWqqv7MF+4PLtG9vD+9TWlHCxBJ4opZP7BJc
UfwjGuBBSJD8VtkoEIGWdmKUaVg4tDu2uk2kCphAJ3nbqt/Vj/zcJxbm7zqoTQbv
JgbGknFbQX+mC4Ety/y7Z0aiww9qmieMbi1Ko7GVHy6QLLVmiBb88JSSgR3csbUt
XwivQdJxA3JyoY79AZQUC7KTzC/EYqETzZmo/XO4gNq5asprUT3yF2coHcyrMPeV
oNJqQAEXuTbYgG8p7aJU0iX+29zEnPI0OCZL3V3AuVmJexmN2eWZ5hbmpUNBODyB
RJgySXO5ar6ydNSpE/4d5ExPIptPZweOpXSAo6yVEg7Ba7URWGSBf+ktsl7O+CKR
JHqfjwQY025ze6k/7LQi2h3D9qkfeqoNUTruV3G6aHuf1FddIvJHwmtWLZmhsgWx
iy+GMsopop5voUn83+HhPcO8nhynd+405WElTmzF3J47AGuc7K79PjIjCb7rolh1
1P01NxDxYmKsipumjABpMU1m1c7RdAadu1AF7DK7o6BXS2yQ3JsWs2fOwrp3X0/W
ggp6ScWQEJzTt+DM46Bj2IKyfh1t9ysunCCzA/Gi1dHwrjbEZlCM2ISawAEFmVNC
fyLQldPZo1/wEKSonPPvpyx4Gk468Pk9yhMDRG96l2HX1mW9kmSivp6BpLtsUStB
nu5M304OCwcIE1K+9C72CenTrrYZwcXiAakfaFszVYNOReOslz9zsxO/lNxin5v3
JrQUGOrFjy6YBRdDtimId13PPutE102sK6la7fi3YboBM/el/T97Ig1vKuYgShFX
HkA6DJHpAZyinHP9nOcXXLXR/8QxMP50BfyKGj+CBsyNjUbqwLaFAVjPRpRJWv3/
6sJsVKRodDfxx0oJ9ASglL3/OLyGVJtcAVODMgoDLI3FhX6vDH5RRgi0BNuyRugs
E4/JnXUsTrymRHrq9GQByQLbhnrT6szmkljKI3bAxbQorKpN7qOjwzj6b/+r8QVj
5nVR/nwnbGFTRlG84/1IF/DxXWnL5NuDB/Xx6faw2OIquXVp52vpArQ4WaslWggc
sBzI7is96Xk5ODsuvp97ZiFxTLjKj2baoynG+wzzoohYtRnO0H4mHsb5ZJDe5cRr
lvHo8/UhknoiOMbGQlKskaJ1MyfsWuHXMeQkpf5lBLS3/Apg3RCUVnR0u9GnKmag
efXQBDKEU1xxNoD9HIKIgWLtgH9jz5mksseOHzl6HSV0EiNZELbVUpB5YUyw+bj4
m5WTg/B4iXVUIuk0nP5Pu11t+3q05kXts7dh3YIsJxRAc/2AHVsGVxMvmu4PBEJh
86X0R/sob42t4ox/mP9TJFvWbSKaSI07maF0vRCY22Ba+3ktGkjtX05zpbkjMKkD
AUFVZswljRz85nFgjjowJb4H9ogiW5wDzyH1Zf2u3cStHoiyi0pYYQ9IitxkGgD7
Jz6lr+yQDvX8pLlMlTqvqYn5/VDm89xOAJ+NaqcGYX5n32q3SstFUYnrhB/15bfJ
BdVNo6yg6lwrSMzwcS1sfHEwi4pcLBSzfVEJvywdtF+K6TZKTONDAd/u+rnvA+If
W5COXPgX8AVpFPzH3p41SC3FI/IYdmdEWND1CxVWPaCZ7eGaYoqQMb6X0p2K+c1Y
DvH6aLmBlgIjqHjLS/GvtPcDCEzHN10LBYOEVVG96ypgmDLbyBeBqwrvvAWXxbD3
A8PvqGdU3ihETcTN0bmtJgbc/LgifeTkOOjiLa1kWtcTKyI3DVSdSukZtygmedLE
nGrfmhBUt1bFFGzyLwfuzO2Dew4VEW2kp39zw+IpfyTxNweMlQ9GaIVg0YlSVfKo
zfwwVTE/NjTgXbJxl50rBkiDoG7gsWbvpCucnm8R7M8aIU1gYeKtwWCZRgjXyLtd
UFYi1ExvBOCxOVBq98cTSRE7nx8O5i1/dyVJFY1TfYPJO7vE7hoaxdWpIlLJgH1g
LjI/c21d1+bQO7pDluoylkEAF6364C9W6CdLHJEpTJUuhKoIioV1ZGNXk168eW2h
pbsWwK8zBj7VhTfyJYi0slvZ+WP6vyjjTivQA5+ndvVF8CubQ17q+c4bb1VMdYFl
pM1p98VS/DiTSuyY8iuzel/7nNtrTKImt+y1I3hXamVD1Dy4wlqgk7v7SQh7pGCd
wYfGzIw9ncRtukhOyTTNAQaMOoSRjTN2hZTfyQlayNRypFEg3sveZmdLeF/iLfZt
zdUl2Q5lmUfFtcM3yH8fRCvo3hcwom+6N95WrIjjIVtihothrOWz+gdjMu0AHNpn
wcLodEPHp/dLziU9wa9g5AOQNa3+szYuNdkphdHyPi42EhXbNaMvmvg7e6Lf8Wq/
1kyvRCbW4u5y9T0hGk2xvJhcEWjZaiqxfWfSyTwaa0lJJnX7WRtV62ch1epX3mL3
b0ENenWDq7yuzgtGtPy2W0OODOeG4I1q16oIPslqRpS2NYAbFvSXFh6kAImJtk5e
Fj1tulxYNe3fAit8qWmlzwKW1C1O1SE++ImoHAqkZ0m2m+/rwA2Mwrc39M9RBa0t
FyjOFwfg9vdEs7AOUedfh4jODsRIULv1k9m0S46qvgKn+/4DWpRa/65gAa75ipBX
utl7EcJ+cJ470FYzKWifMtZKTXwDcEqEJpyC+4vGKbH4cRHUQMe2GHYJn2W9WQL+
2UAImILim3HVSzN5h9do8pClxB0+1MovD/kisaTrACKUgCJFdgOWA0VJUvFLC7F6
oMYRae+L20OCn3nfyTZtwMhv69lm3tV7AtOSP2J0Ct73n2DVfMsGNkhP6sufmMqD
RUxYDTI9uMrYXBsUdxqnXIvwLIkWM37Ib84d61IDhgrO3hoHSeCKT3GikEKD16X6
UPpVOqwBV0WcpP0T5UEuHchH9Ybo4uAs5idksWXzHqzYwEq2ua6Qx6IC4QErSSFA
lH3XOlFbk7UzDaBFu5YsugzThuFUl8kuju6kOaG7L1OqvhtvZjKKU2NdmwmaXJr8
mEBDnst+QdL88Z+HWjtWfHKqKTChr5Lszk8D69BSy2hokd12zGsYh5KykX+0phEA
VQUTQ/8ISNoRhy82O7wqnG9ZBh+Hj3mCyl33IRmh2C55pSqorVF+Ly8qQvzux+Y3
PJ2a1zHTPtYwf6tzozy6gZTdB1QmFdrhgDnL/WTSwqq0QhRjJqMDhc2jzsnSsJCK
3hkJi4t2beImTiMyT2Px4xo7WFSs9T5BGTV4+89zQCQOXLUHUHobyQD3WMAcSJ1M
8JzTFcNc06aYXD7DK7ACDIAIbXnxX079epGczyxvLqLcWWLlFpcuagwkSnHBQiVl
M62jdrM+ouEyVm2sHQfVK/IX9y3q+mSTUnzOoHgcw+JipDckjFvUdvKG5IvF6ghS
JccQKQ66VzMvAGoFAcnwBU+tSXLc5l8iOcK4yutfp9G2UcaWNFe2kEIheou/lQ1F
Do/qLX7SIouKANOj5Aeg/J/NcfbjnFN9sgw4f9e7bikp1ZODA50AFYHStnRT4H5X
wwJbfnB6kRFk+fjg3VSt3dqTNxO2M/sshlE2z4E26IZBFwhSl0eTWYhK5v5p5Yba
L4q/JXElCPkLxztB3n6Oy+b6Qe3Z/nvwY6uf8QTcFolVHFFEx9QHAKPG2l0Ttpxt
KhdZQGaL1TaoaHAIjLcfrd+nFbOcdP6tijIxMmXoLsCzlV7aQEh/+uVXs91Z2Q52
Jhvvmvgdgbu1Bjhb/xpqhow7cRoZavvM9jqNKvlj61cviV7L5kBzWFN0+mG7PYzu
U6Xj8pOUKxbrmHXDe+wi2SmIDtXXSaNbmzBmTynzlGC15Xyltey5/EEOKweIuowv
E6ZNz4oL3YVHhirr9pYV+XdWyVvzOz2aqXNgSF7+yr04YWc+OrcmP+rRa7O38kOD
ibENVD6oJk0KiVC0dA2okUPcFovro/QwBkutFpi7QWsHDxrsJWQJqmeEyuDmkqhs
1ShZ+2DyDsIiA2xNlqwhOolRrszPSmuc6hM4RXwTEN5bhvN49+4CBdsHuTBU6DC5
kzHUEHOVO+XDec1FikRIdpX72Na0CtzKytxheB7Le4v4cyPFpX5ru9yabnTJp0BM
LKtF+na0kDje1DRb5QY2TsKbgCTqaDntnXHWCpnLaHwXTVdL35cAGQFRUizD11/1
5tilRKNhnyasshwN4u3n1m4gcJsvg1sqL7NZ6vFFQ9iXpPWWu3M4StS66ogfmhM9
yglMCsIt4NW9KauEc/4PR7KP0EDW4VMLxGBTA0QSXe8yYALE2vSv3KP7lOxGn7HK
BCZ2Fgrv5ICOMFGVfquL1u8GAUlowsXKZSndbzboUtRzz/N1m6Yi7iZEjd3c1QF+
Xge72UquXuo45HwSfnHbNCtP2YlTDWehrr87DhDRRB0rJHN8b37dQ82lc2Recr6G
fWMCA57wHmpLUnIMAUsApLDtxSzKdyC0LUc9WrcB+NbBojGbAl5LcnmGGpbXXeqy
Fwt1mubWYmBbQGf8csTaD9S8L7uEAWJDBvFZo3D0iaHaTBQmz/+MGOy07ARSM7b/
Shs/+rX/k8oOtL8iUVehr6NP1JyPic5B78qxTXCJwP+HRY2UICW4i/xMUjAR62mZ
wi5GXl4tgNuYVXTGD7v/4QHHzK/SLgmhc4iIKowEd0m7ohRBSzAemz4z6MdO2dpS
IHgeengP1tj+B4ZY2rHaQvBg/DxpjNkBpzpdVhunqWW+939bi/MH0x+YXoRTQs4f
JaOM75lUrQ7pEI+yLj80hA96o4TKfAZ9tPIJtJVXkd0ZI4nC+X3duaUj0MJgHYQO
MiJTyH8vHWD7IIcekHeG69P0mSgt8BOyq+7hCT4G54uKhg3YcSbiWBL7VvjqQwQl
Y684utV9KqMSwV4Pa27gYrbhQZ9k1zT1bpnniuc838crT77+AxeblP9RwGgrwcuW
olzXNnkh6AiK8w08ItagR1jxgHkflNOz4HwtEB6u2c3QuoZZKUU/L+RMmIkLEq0J
GUD5JXvm2DpiTjPwjO8YzNtjfBht/F1dA9gRidvx3K0NRI2Gxv7n8J+0rkf8+RiB
H00ph3nDhOYrtD9c9UKoFL1ov5D8N1lGCHRFU07jShXDMlWwL+8VJRm5CJay4f1Y
BBGm6iexdSGVRlWiookSCyniaL0PEEcCiqpItlzhreWsILNIn3VUn1ojbwOsBAi/
KveJ6JbSXPLNoJtN4XRrzwMXLHk18a1Dy6q8mJ103N+Zzokom/verYV09VQwY9fQ
2TdTtIY4sCa/S/nN0z6oWmPVTyl3+W6Yr+C1BGEgkLuRtg1/YxRxhCMlLm+bJUeZ
uYgKUImEkFT2JmxMm2Im+vH+ZISR1W44fQkCJmOvQsBlDXSB29JbgKkYSVr36ngs
vzB+MX9PrifaWEXt17s1MI0fBwMImqalbllNaE0Oj1q+OM6KekMPcJ+hH/0PxVvT
CEScgLzAxF6S7/7cyJrH1RcHhBDhZIQbuey0dsiA79tD+QnlKzmXfhiaHImv2LN7
pgOPxe97ppg2i23MG8pbsP5AB4hhYDzep87vPTbdixDTN66TyM3puJgy7wTnqrLB
hNQmbpzH/UmUTyEgIB3jvisGcrkOIrD6K6w20djdlIin8TMAQTCQ6poHqaml1yRM
C5yX8Iu3pVt6oQu9dh7lBm2Y9UKW0dghPliYhnsUfMfBre+bhxMfSmGubGa+EWZf
XCyj9zVZtL4t8JKNz4UTgQd63IQSH3ZHRXNDQ73mqhXDwXCfIKjxqVk+ZpyYVVGH
Dfjv+mGCX55fUGGbHiktzR0hMsZxbodnFW+s0nK1VjAhg4hCSOY86im0r8+yT4Tc
wzu+qdVq3vaX6ywGRf57OSpTvrTSh+O+t07n6joMUXIcSFekKUPMhWgcuvkkQqYo
/T/6gRxbW/sBZxGlW3vYG2l/uokD9fzYs36YWxIIfVZZYNbpc+tdrzqO4W6ZfXZp
XTu3dofHABNQiF9GPsiARGknH+SyZt5vfZEwBb5PskC8EErnQeqZDgK4QMmFStEZ
/uO0aBkUoFskrFaqKsGuQPE6FAQFf49jnm0vf/Oe9jx1DKPsejkTv/a30866xlsB
8TBa1NbEBT+yTGdt3EeoeRdYQeYbUwDsLKMJm43cxUlIFVys289HyqAnaMBPb4L+
0fzocyW1hHCJRWfNC5t7G3SVMbBC+nPrQvGaKALBy8lU9lqoWvpVuXgSrfjA+rKL
m98O5DAiZ92fANZ1DuqoTrjdnqG5Vc34f1ZQZgkGffp9v0cZi1U2s1qgawV4FEQF
pyVc4fhdvisYz1IMum/N4eZsISwacVS0hnbKja0AcOg0sQ3qpwwsJxo++4sFbE/G
v/a2Qg6AwF3TvjBuPtkjG/2e6mK2rFoK3LLWz9+NZDqWdta/8uMDTWgcly/bOH5S
5qsW3QnrI1lXXxrJD8dA58Kz42w0nbqYh0nCheJjKGZzhicWuLl0JvoXGp6/v3Uk
pKAUAdsA7zznRhxUVc6y96jdgp+hdpBRHRZDjkwxfuYC0INX+ScEp2UXgtC1NQiY
W6wZfsEEg8yaNzcISVFx6xDR+NDlr1p+bhqzBB5gze1c80G6OONNFctOMW7PdO3Z
0G/FrtEe0uIpEbDmG4WIv5If2pntae6KnGSsLpW5vUXoDogOqGyqbpByJ3GSZ0kU
Cv8IBA3DWYHlP2hoJoDiz/jecDuBB9OsPVN8w/LntfqhIh/fupYQN1UiCjQRzTck
nwaIxPZ//crRSwKLUcgj15A0ILvqaTPimRI9L/X1yH75Fm5NH3+RbEco2ts0yqrE
Y3W9AX0w4qhJIOuX/wBUsbvn74JjAUzXRNJxAPoFCW88whZelOh1otXPsbQOrB9Z
HK0KkdqfVc3qyV8iXRZ9DJI6e37mXBNSNgPxMpVeH87elNOZuBPpvoD/+iGRHk4t
MCis1lIsgbXVTNZ4UrspLpiJ9gTi9ibb+RYJOAtuJLZbXMK2jyUXtlt9HeqhloaD
xhED7b8cbn9fmmPqCch1D6e4OnulRO74/QuGuBcFlNVL7ndTIa0q9WsAhmPVTMln
T6T4zvncoR2Gz7tRBAOz+xtaKAq0ekWSdh73eNJ/bazF36BQvMZbpmicNNpkAlnT
dln3qCg1sJcxS+kdhHqacC8GqOYECNTikyZt+zgFoTC3BJ0HH5axP6F12oicTnl5
cME1QcmJpIlRkNhVZJ8tE9AonCJT0C3a0ckZFgQRLV3PCibP2x8VEYjEXaVBZJ+W
WISUA5V0965hHQOKbM9j82X2aBfafNcdKdShFZs/OSCAZsvvT+8uBedUyfKmCQOG
rFSm862g1eVEsnJlRQ6MpV+YiTTLHfM0wDPd+ythuw5eqE3Bfjrx0MsN5XYPameS
poJgOezFT7Y7VmlpjC3GGRSBh4GogHtbr6mhri1FgFFTAQUOMr+LuvQh/SGltsmJ
Jc7SbqLSmuXX5vZl1SufewUjhTkBW+z1/lkLRUmweIlvPNJ+Vj6ZH7AoMOiqrruD
ShZ6atEUNhdBnoszLLCb2ROK/Js8CoOdhd2dkOo9frKHwZQWH3ZyMoOApzZeZWwe
utoT7dEL/syStaO1geJbOUxys8bTW5wxRVq5noLvWfzvp8ZZBU/VYjQ21D8LWwvi
VxKlKUsY+Ucgx+gjmMXUXfD+5a3vO2kp/PtDtR/884zzJU/BKzLeVpInO5cTiJWW
H4zFL9+aga2sPwI4EWj9E+t9xXVGgVLkJ+PevskxFL3CvsyZcko5w+EuluRjXESN
rZ0mslTtmyENPoqRizAsTzezw6hTz7RDQeLYAkS66VVtSliaho/lUSg9QNMafcnb
MSyta8u6MsWT4RxgVoghzGfJuDXqc0EV1Ok+KLCOjxQolC+OIxWStw/Slh4WhbMs
onFvWj31JnYkvQhyoW4m5pIGh1LSWDOapVQCuqcf0k9PFTVCeQ8B12mkTTgdtgJw
5Rd0+eKfevFquNsJyktaJ+BD7oVnD7Xr32Hqzfk9duY1wkr+fQqvN7PpPrzExE6b
mvx0vnfjQMIto/x7fva3S5Nbjthpqk7LT0+PKqbnpNqnq+k1eQr8XI2xrPjdi5TP
YVM47O+4eY5xWFMNJ6WImHHnHz3SBkgQZLubmMbl1DwSmLzQH+AF+iHUm1oMRZmP
kLceyyhRHWqkHjq+r6nOlB3EM16LNmxs96x5ser9wi7ok004PeD0ZWrFYi5XaizX
YilisSe7zT8DQGZrxBecZkD7ZRnKnLJQ8pzL0GJ/zaCVq7QDJQOAmta5nQQfvXbV
DTFQ14lsZzD+I45eMKW8iiJAb/NTBRWqRrQxEDynw3GqgtuxFWs5XDOykdRxpXAx
d3ZC8/5j2aYFrlKBjFI+rnANKtv2+3E2/Mmg1rmv9LgQWRYe6AXt7YaOIeOuahCK
FDs9xmvsM1XK6G4oud5FV30Y618RvCanu4vy8K8iK/id0nI7xKDK1/drtPit0y0v
se5kgzRZmubx6G1y+dEDZPxcWikLGyPoHIGBxeY7sAFrB6XskoBHdC/4XhrNmy+K
uTxVQptbb4XgRF7db0Guty7Mz3Sd0O/GtCrcOnolNuw7uaAjtUmZR6YXrZceBo3D
ULbpqkY/vbB8KgoihXRABt7GGgDilllaGMY1Ya2HcG+1P9DeHeV2k2NYt2IRiE24
8E3NMh7BziIKb73CiOMLvyMzrhgwu0rfuK4BgLwp0RadqxLeZ6XaT/GkSwSsb4RZ
mD6pvUAg8AFdtHcwRExAFTTXNBh55R9S6911ZK0g5AEPLY5WP0yoMfdM/OSCPbbu
qddw5Jgbnx6oGMV0tO6BxpxDTpB6HlHNY2nNwt6Hp4kLpOrBq7hqt3lroQTK8IS0
lrSRY5bf8XBK0uBdoo7ZTn915xgjA/ArVmtp7qW4kXxP7ZcqefSAtVVtWNWSBruS
pVj2koP+Pozhr3SNxsyQk1KaPB50SlpnEdOHAu6yKwaOmKiaJzpwWdDT0CXo4vao
XKj6E3R18LyZozMBvSdPB7O1CgsYKipKr/NKmO1yOy5NsL/EmYOcze7TG9f20kwc
RgNb9+T2bkgweL+846FyLk3GlsMjXdV7yra6fcHDsExI3u6fDe0kdGDsgM1BlSlW
DhoRLFMKwNjak9f6pj8koo3asSyG/9teyTE3Z/uhgjWrtNx/4OD/J7uGW+Q7pOg3
5PvAYTp4IZLQI6I035Agd0NeEjiUnUHd8s+Ou8T4S9EZDSIZFfyRYquffkTIMFDY
PPVwfAbOIv+QVUCTOeOxhaf25iWhbKd8OJ3LGOV3p84Ksd1JWg5FDInR1gmB29af
vw3Bp006ceyQDQOHc+T8PixjZ63RZW/6OkjCJEd9NNB6hcRGSBHz0TFkGXPdQ/JD
cRLW3e0q+nyCenGiEPitZt8JdFQNBcEYxqk5H9Ex8n7UtfpTJa+Y6yu5KOnxU18j
tv7V8h6Sd437kVVTWxu/VXlMnR6M5OCNLt599tfhqDdUGQXgLmEzvvZT8V2oHmgN
fF7uYwRlBbyObaTMBM5TjDqNVzVc/EsMrWWbm+90xVV59wJlMX414Sw4W70ZbF8Y
EoIueGcffPceoO1S8/OtE3diTScES22UUYJn9NFGjHVJwc8QuL82CyiUpkr/ZKRP
1nFEL88A4oc72VnqsNWDI3etBZUr1D+VbGuUslDwlj6T7MBivu+hAtBRe8AORJio
6Q88KUCD4gXmo59bKWpfz1+FragYBw9BLa+RnPirwGEUEbDShiYcdcGIVoYHSjMw
By7Aecs19tEod8+eqKQTBzRieNbotPUi63ZQZX2bvzYFgeoUXZ6ySWWOL0QrYcZF
aX3mJJiZLooMqIqWV4cs7Xji/AQcMjvkz1N4MhLMPQ67skoKYucES4asYkRky9zN
V+gMZlzzpLaN+YyvZW0FtO5fCbCML8C1Ir8VaLUk7IEzdaKbfSE9Ysi1QMm9chMs
1YJh2BqgLWlsa4x2/5ZSfFS6tm54UtS4bjBNUhJ4VTP9LVpapQLfoV/reuI4EqE5
8huiLyaKCZDMawUEzgT1z0gNdegbORQJ4czWar5j3YsvYn9MiM8O2Q7R1EVmvY3s
/W5LuVRzBucJWTmdjSkAfn8rRvUssS+uHfcoD1dZgZaA8eViulJekarnLM9aHl01
Q+RSDrL4ZJXaU0rzAjvKjOkhdY98xZbDjt1eouX0nEFNarRC1ckRGqT/B9d0J/5j
LAd3buIp+EBQ0PEnAZY0Gh8vD5zvbOIr9FSFmNz5BrNkCt0rgIZRkd0bG3uanZbs
8JcXf0eZOy1zaYoDjiiE0EJfUUFXxBdipuTVaBjECwjIf5OaG4tUfO+7hEKbd7xf
ehxDY3q+w18YQAG6yv/0ylBm67d3cnaMlKiXdRc7n9VLLPOpK1MxPsoAv1lP1z6u
j5eXOlAAMV2irk+DagTTyMvx3h6xBmCF65iNmDXlNogw/Xjkt2HMa12GzJ0nlNKn
4R/jJFWYBwk3zUxTv1be8IDRO4N9Ud8iXYpoG0roWY0joXGPG7C2bCZyQxltOWx6
euqmU8mQV+yix2/Omb1DAtx3R9ODStPCnMkaPvKLRSP5YRy4QY1wWM7G6YTjg4cP
iPDoVQpYa270E9kaX3TH6bA5Lcqs6ozVSGAxDsNeUP4EDpHsU4nCe+XPSjYZ0HG2
vkQ1/x+eGaY571yLeFNObtXLPfRcbOwT1/FixtAlTSkO/wqEJl0W6+T4i4f4WBpJ
ALaud5Ed1AYHWxTER1+8c56JJVC5bVoPr9iezfgULR8kqiPZdzP6JDRWedR3+thQ
dGS+9doTJUKRydDT8MBjcpSG4c/vHJDoQsJ7DCb3XPy8ZwGbbIlRJENIV7emurpn
1QQoiiHUzWO4l55vmIq0roX58Zn8lLvHRVTcjKrSWnigUpH4hlnVqRfrJ0rYrn9I
yzE/7yZgDSbrSf+WPf8+t2iZ++YlPCissIb1d0Y0S5qofIO4BApweTEGfWdHKAnM
Aa/cqtTsaXp+JiTKBafi+QYd/aWHUvObLk/P1PG7hjKRfACPDzY/MB3Xr8zsW3Ri
Lw8zXY+pibsJkCATV9LlBabWcMDYMWD8Xg4+kpQQs23c62vFdAnr71ERJ9bTSHMB
KWPxUfdxXsu+Zq78YJ71rgiEMS3oESDG9XhuGVpyWvS/95rcFgQR2bhhnNFDr/HB
l0Gry7Pfx5i1HCw/of2ImezK7pU4YD0uzLRX///E/8dcOdsYfKmsBoowrCc7Qqlq
Q0leAqAe0wWdINqyb/3lOBjaCwmJuUWrRaoUmkTCeQqEUw4nTkOnrFu6CAtBxWna
X+jkG+JTllf+8FTyRED55btayY8TZj7TjtWYYEbGqOxEGOazZaaJy2Sn1OVl4uoy
/f3DmFMLgfkldsSs4Ry+eOwTjKcCQjXmeKMUeXrPmT75MUWllm5buXlQTPNrNJwj
BwsUN1GsfxRV9Y35AlUBwXI40N1FQhCaphGdfMU1fIQLAOVeyIlOOiHO+8T+9Hx+
9ipQBNY1drWX/HbQJf0fYZGPO0Jy2713Gr7iIyx2ZlaH4b53r1Q8XSCG9ExXPqju
7sBaJLqcVEf1OwEYyCjjJG6RwNaXyz7xYsVD0R9YUcITkNF3Ca0NHKobMHWgFVQU
eVK70vvKbaOCuXcZGGiV2vD3rR7BiZ9BM1HaJkAAb3HcM8gJPozcGqrIn1cuW5Rd
E4GIpCuSQ1qee2ELE29fODddIenwZkD57kUR7Qfxjdq3mSg/awuPH6Y8YBddtErS
HJ4kc9KHM+zYQm3EgcWFNlzqwUFNMlXArt4hq+r9pWYaxr90tzMZHfpUMRh8uE2E
jo1OdK/6i/smf8MjjKuCh3LN0q9dyNTiFG3A+0087Royx1vOdsr7UD3oEGCBjg2H
TCyJvH8pGqjClG6a6OrBJKv+PRPfnIFU4+ogl/ZsPj5oBZ3x34F5Z//M7mJ8nJWs
+RlZAeqQGrLQPblIhVneoApgXhhtGXjowCJ8PrDVKkm3by7vI24m1bdfSyUn4yDc
nBF8rbqzItCjOehsRU9bcCR5URcwjs+DkQT60l4J2MDn6tpwLUs0lxBS0u2HWbG4
jjhC2bbwd41pn4fLidatczega3kv8BOPLgDTE4Hq4goZ3nfp0wlksR6w7oJDvhq5
zxfQTasBG0Ci/QGOUkMfD9ege9s6BN8BRSxEe1yq0Z6LRE+lV8APD4MXVDGXdq/W
F06ATEMXJz5PczbAF1P6Tv1VDg4lDLibexE0WoC3qG5tUawsAxUwYbq5Bdt3fER9
vXNPvMUN9Y+JTNI0jVXfaLhb+/LiC6PG9+SWURUf2Qpb0dQFSJAgIQVEPmhBh52j
Zpw7NUkjI3gnFhVfCTWyHCEHv5LwxXlv0k5KO8Iz75bzDc7LWlsfqsH3oFSOZBYe
haKYeMXu8w0tAZskXEriPLc5f37y3JEP5WZhaJTPRk2o9aMH5hUFige6uXU6sBUr
O/n58dddHkdmtrWtqAfvEZ6cWkn56p61AVT9FNDnomZVG6Ww/+mQuSUMcETXCRH9
8S0BrJ3LgKjiuI4Ajdu0mEphb9hD0BXY1/nLH/YdPcDSY8HMtVdTypJFqfQ23jos
INIFTjCyggB2IOHVe/43Z/PsfFA1DRujva8e7/R6y2XxykJhwuXQ1h6P7z2UKfBl
Hp6nVHqrLo+/3myIhidHq9EJa4MYs3H3TMbntHFoARiH1WgjdpmxpU6zrC/iz6Gu
0OSXzIQHDro/1jG9M/vvaSbsWZeFc1zXvPT1PmMCsoM+bC6ZYJdBadYgZRL0n4Ad
bvFsr21l46YtuXZRmcDGDKBdTCUwJYOfAQ7Gsv1HL1ghiSwzUu+uWacNcnV0fm3W
GWX2JyBDjIR2C6VMnJ3kUO2sIcuqlSSJftLXJUIUDK9FEVAfjewHgiPExiUDochN
Dqw0Wn219JjimTyjUGR8E7XLQeifgenrvlS0ce/bPNEIcNxOvLdpBUsmT9Mbh2eE
RlhkSkTarJGMlLUfcrUM5/B49MYOWLnbLPAPgyj49S0DN8kylfB05mps0N1q0xkf
x7rszGEnv9nerI8FGL5CMTvu71ngptovSYn5KGlDZPVLP/BCtRoDolNdrlyobHBV
n/hPKtoYVLZg9OKBTW1WUPF51J8aUb/jqAvG5CNHi6dfL9QVzNNEqDR/F2E3nvtb
vFR1G6/J84Ki/SB2J754vI7s9SFwpEWclGu5dSr68OsjsUfbisKdlr8qbN2cMS/z
AUDoiDilv8jrrZW3RrYDgpf6ijIEU+H+91ZAc2lcKp2fJ5mxV5b/2s73F4Yfz0nu
1Rvs3yVJuGfwd7li0eNAgfFe9li73ODGjyrp3qoXXzS8GVOKob9yKkfaKTGhwlpN
rNWUpmK5RCN1i56P9SdOpuPlB65VaauDT4cloFJZm+jzPzb7SQ3QDQFe1KxZliHr
L/XQHJuAOThI+AjIi/gVzJFr8Pa2zB1+BOY2AX4WG6RLOSxFYQH+PS/FKvpJ3DJQ
WdUOIWl1LuFo/jjQklMQvvHeqQZ1700iIf34OlN31xYL38GBEMj8WrP7ZAnkhMyI
rxEMrKnBiaejtbMyyoHtAo0w7qOKtEEYiIbnd15IKImbd06sIfArcvZPSVR5IowI
gWk/i/LMYhImXxVRX9stHA==
`protect END_PROTECTED
