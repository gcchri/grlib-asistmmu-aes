`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3tPd02C6t+5XzkuBkj+blADVkjR/qHz9CVo7TOEVkbFmLX4K1Cgp0/a9w/cD2qhL
16zqRWPal0Gh0xgIOqcoWiQ6X4YqIaVFGtq8FIG/gBszq2zZyq6cqTowN6iI5YwP
6O6w7tElLZ86dyKmcG8eOkhKH9LY7Jn26Cey3NpDJ4X79tStLKRSPv1eS7jkZ0+3
x87JhvAWO0TOx6yBrJQFFRFZ5bavVATfjRMxCNTc0JvQ+JcrsiBz37dS1OincL7e
ifTzqBUcyM3OAnEdmR0EFdBf7D0Ux9ywpg/kG+5RvE/bHgj03TSqUIme7qbXV0MU
28+KTc2glQdp3gbJf98Yf4vXNCk/dYZJ9pXNSuf3tbjm6mkcsQAXy7DJMfmA1hbh
z9088PNAk+uXnXPiUNQ+ca8CC5EQt3gqvqZ8A3r0/Hr9jL8+UGaiBjzRloW3RsRT
g3AJlRQy1hR0hB+x3NlbM6xmhARm7kL6C79DdK3e/qwWNmUtal1em+jrrqRhFa3l
WKad+qNW3NJwgqv1Fs1qy57tK7O1p6l7/qCePXT5C/zbSnzdUHBTnA2KU/T+0ELD
sZ/oGVgpdRfB70dd1R17H6ln2Qbj0bab9wpEv0+hmY3UNzswNYxs0w3a1BhE1EZO
i0QMBbn9yWWejrnB4btC+ow6KQqk+i4hXmG97hcH2d+PR0GCnoylCsxo4rBK53kh
p1wE+A/8b40C/mokInqqtD2O/3gdoJ2IGtXAUtNCrP7WaTolefXx85Vm2KRv8HA3
RQrO5mVZaQlvUFvFk+wEZgzj/bRnX2gwdSz/c2uUWchwKgcRfFxvdb7u15m+1aWM
Fe5Zyyeh2ya72EzI7ljOuZ96/qAYEgcVGFbAUggm/1srwY/6nImpJ5gIvzNue3oi
dy5DP9nG4Ry2PX+cAddHI9Q5pMZHvuDaDd5igN0X8YXh40pPwGmTrEHn/+Rit+nB
JwIC7B/ieba1HJUSxUo3xLi+AVAJ+dTA+PPKSkut3/WYvkpCrwYPCZvwwqrvvj6r
waeZtp7Zls6QCizBMvoAzfnKcAyG2v/n7qxme2WS8ns5W5XQ+s/FKJorkvuqzHHK
B3uyoXe5kK7eRiw2hrldQ5TiGAwEnluWaRvwHSSWJSsqeYUhxtHHuHsaLwiX2ZoO
qxKuctv8RIadGHRWglmj1QcqUOtOmCIzaDvHceN+YC3dkMNA+WspQ9sG9v9w/QMg
IR+ENk3gPRaAeJ+7WFoDB543Qz6mxv3TLl5DrD+zCRSVH8g572qiIPzRo54MeU3V
RUePQuUEEUs7CQEjNhShexuDhJxCULvjHWYLnSUbGIVdFA47bwL2T1RZcEifqXBu
miTbDq3eDtkJDYnNWLoFArXTK7uCxrYsgxS2LZF6sd134EVU3joxO8L+0vBX1kqV
WGt77TZwAvkn8Yqxs6lOB0mKyO4QR1ZAKMO6AXpHBbNYoiXK3KYPJ9UJ63vYOcI/
xA12gzKJl/iTEVGS5OK4U4lTA7Ube2JmN8dw04Rq/NMKS5WIgMEB6StPHok/yBvL
KJA0rc+yahuzvbQd4aW9LwWc0ZilOWoZCznxqnV293C8ugBw+ouyBkBNOuGk8d9Y
67fdLHUfOpWpaL6J1kwmuOD5fWAW+CJo5PmJuOXMPnM6c9LXayTjriy82k51k7nC
dfeOxnpIP28R4XAwIUbC4wQ8dIugrZz5748QWYSlBF+yGTWxe+ace/26UxWqDW5A
ZsGDVVXYS5NwLsElbTOuPz16XSHkcJUtWJH2o4n8DtdGhbDSMa6ktdTgVpyU5eHX
AUOxxZYnWmNNgX47ufD3HFGpXRsegDMUMPl/mie2sY1g/KU5T578oYn2TKoc1XrR
CxPpoFFpyWIxROFJ4VZHP+HS/90L7rVpEyDxNLZsA43TMkIx0Rqh2bXS+MF9zUPo
gFS/YVr+8nfYG4iVq41eU3VM54wHtnB2LkpQRScEAd7s+7WgGvd5DY3ns/rIPJQd
yJp8mf8/FI4t9+4p2xQTJN0OQQStSm5O9xosX6Tp9vp74x5BVVtjgl6ZAA77f5K5
UKBNQz58ZeaAW6xosyGwcgiXuUv9xN/mJmwsgAcvl6b2+twT1owqXNzhdgE2t4Ag
TrZlGq37Zhbu775yyVdpvfjKVfLbluFVBtF7EPb60kcvdbSkwBckjgZTeYsZZsGs
NfD58aZtiF5bbvPavxvVDvucSyHmZy7RfpgclLts2JRUazx6EJDjFEnLYuSFrAyb
UEIXdc0/QIeFra+E0k6ApSQVmRjOqkHDIb4jK0dKLpHAwCV1srqudCCLo/ySPfLF
bXnPnZJiPZBiwPhNAqnxgVHag1CpqzicJe6URloLIg+b/uoAQ2uKhnSsiUF+9oi8
BfzVeng4Imm3wWAx/4XxFWJWO6lMz6lie7JHs/ct6Su4sa1Q6gsUC8BOqKpJtYZ7
oYFz0Fav9M3/fsMRzei8hcqnJtJpDn7jqNsxoZ/8jHzr4fdXXAj2Ns3G5dq+N9Pd
CUmII7AauGUFDqenG9M9sSKdTDBeR+8nBn8pSE3POVg=
`protect END_PROTECTED
