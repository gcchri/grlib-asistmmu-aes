`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iDYwB4Gc6/lJturqk0uhjZYBxMWumjw1yRLk0ARcmzHxtgshov6YrHaSetqdqqI0
Fsv7AZOw/s2dccscMNVpRXMuc0/0B70axM0EcaN0udY+DtAU8CyJJtcwgkWXjPP8
f6d0+mr79nXlM0XnZ5Wuqj3UxkDCCp8sSWqPUOwMFfcbvq7MNJkGG/UYhqqOzLEL
YnYVUFRbui8hjZ632fbdKRgh+jzZbkAN4Pm3bV/w7ymhlnX0TxnCveDhUWzaKVzS
CfCiNEZ/MWdNJz6PYr5b624ktm/dsmYJUbQlgJC3x20l/5yPDEHBDXKANZarBm7Y
4FeIJVosEnEROz+oMulUUDwu2glLBRyobZ0WIqiExzEDOWBc9ZeHRjVDxLgkpEyK
sLwX0U3rNqU9wu461NX9xcAmLXSPrqsT6E4GG9rlza+eMQi2uNl1547Nq4NbO1ws
a99G11u1FyoRXN5Gkj9zDf7QzIFMtMYF/IfcMsrdJRnEiFHAY2s4olb2LexMu75v
1N+CFugKNzLOTq8PmUI6eXuBg5GpF7cxZR+ZrDKxVUfWqbGLOsHdXgP06ysSHaTm
6oTkkUyK3STzf52FnAa1Z5TCWRV97S/qLX+Hj4Peurk=
`protect END_PROTECTED
