`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y88MUxKvEhrAkx8CNDL7DN+AxTw3bo4DN/77J6Xd345MDbPM8Nqht66KsyK7KW0f
9DFwHPjSnnxUry8V88AvZ5tzKC2zlOwvxxR7YRd0evRe+4IxR2tvT0wzoLbkZ/xr
eDRAYElXechXgn0OzoHI0oPzdSWdjv9KN/ErvJtQxX8bbpsA54GNtrAwhAcOb3Vm
aFANtekw73PyRgGRqGkxccCE5uGPp8dHbxS/4KzBj/AMP35aEQpUi6Q3CgknJA8j
oUXdOqbDdfe7P7tcb6PPHkD3DAMFXIYzs0sW7jrFo2vzHFnqyGxYcEHp5kf9hMbI
SCWWzhEzYkseI28uOWx1ByFFvaHrbZsopsJ42YD3nJ4B8r23ZZWFh7qOxvCW6k81
`protect END_PROTECTED
