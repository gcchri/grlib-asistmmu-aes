`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b7Ih6hvKuZuXaWEFAW63nB2ik+zcdnBj7oFiOVBnFPVKUbfyGBKAwkB+egHjma99
OKsl6uLbTHoyOv82k89+mBxipAaBzER3BHqJjBmdk3PBwfg1d/cJpxlS24Zi+lay
V57AtEPWI8Bx8qA5drnF7R5Rohrf5gE/0KdvQk0hn++PxzUDCuTxUHFhdBEEGkOx
36dq3281pOfWdIOF86KIqN2qGAVrvPMpWBK5HkkxsM1Q9YqwL/mDzkZQRuVa5cb0
KAXKFwseUpwevjaHMZsrBL8sErhNhJqgJ4AG09f16U4pVXWe/wRIumMu9zsxWIcI
Vhc5v2CsOs6iKQH4jtiw8kiOsu3e5o6YDpuZ0Z01umiLK7n5wOKxEM3K/cgi6PSq
/JbjuQL5ghmNGaI9caZmvsK+R39l/WEpsFf4JpRDWJQiB70PANqKgoz/ZrMbmgSS
dVTS042gpfszjVc0m84OpLN6qbbrsoCjQH+Zt3cFhnlI1PavCSaqIlRuMVSbQlpA
K3u0NNrF4FgJHIqJJnfJdMWWE2cyKlDGL9jyror29pm2uV2WJEpv1ZKVFeeuXCYk
gp1mV+1MVR5bzMtK6MhaY+FUnNygpps9Ds2wrJx5bch1uSCP9BLnzIPI6Ja2LDmP
qFhJTGEoEOOl7ePcw+qafxnORxX94t3srnudM+xSEr4USHNRqVpl69Ni4Sorw0gT
OJTuyyXviCZy/IPgnKMgdGiRWB4jgnPBl6O4l7aUC8/kS2IecClEA/QI3gH9LECI
2VUKcm7W4Rfheow5gYnN+PltCsoNlUtUJZZMs8MaCh3jR9mNwDW6lPGiW2cd4QPC
6/PBRnnKwiFC0We567/nnqEUtVNbXCh8Q5WNqRn8lWU=
`protect END_PROTECTED
