`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UWJuoACfxBuoa4Yt5WVdTP3kgjzIjz/5n9ysuoXxV9xG4zR6T/x3QfccoTY3HlzG
5QYLhHBjpjCqe6Merhz5hrPSH6iseyfBBqw86gKGBrqj9tZ8XJjIEksmyJXe9TyB
+KsFiakdp+JTl72IVLIqivl+wV+PwK2ep8mVVdcfKpI2iOSHji46BsVnRNrtQJeM
lVxVXVng4GyRrDm2qywpVlt/19RZrig/qh8KwT5lyY4ETjbHy49/IPbaVXqg5/OF
3L0JRj5Il/BVxJ+Re6jsdnsSVI4PwhCLc0NW0sa1sFK+pvd7cCT9FZhUB3fBW1/l
GKIp9aSGIbc56dAzfvLQmCXwbYj7QSCfdefnb4mxno4=
`protect END_PROTECTED
