`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1S8PBABPT3qSqLwjha6yKyJ0NMrv2tSNCIZmn29J6hgRvImaEAqwMzD4UFfsBdgG
dDbST7GKmBB8H4lC60j8neSyCR4BFScFYe3WYfmpleb/la4oYTdjFCKYXPNWdJeg
L7+XOgTCdEeu0AihPxPabIwzymdklRDwKfyT+x4TCauXUnXpwk8c67fqtgjGLpXy
Aw1yZOWvGgE5vvJqaXup3NMp4wN6VGuCFRqCkMUEshrDVAzH8iMq6VWG61atftiI
elVEOJ9nvbQsbIVUhC+47/oi3ainjn4rxQT2NaA+znt5AcTdo+rEyAcK91Ll1bYM
O9yw9WfEx9szYAjAnpEA5laI7/6JMnFrF3jzOlRHyGGSeQtGS0i9utbU/rVHFTdI
0u3+lSbOZfoRakpuC2X20iiNBaAkBtrSJVEb/bVtfCFEu72euv3el0EAx04i2aTN
d/Cj35nOqigmwSeHtSzA6ZU/z3s1i5aXWRfaFqW3yLI+7IBfQuUTHDllag6soEoS
TKYokkn7EZcKoOhBYvNRTE0RnDU8F28zNFhBLR7ExWNZVbVGRzCVq6zs7RlpUdmQ
`protect END_PROTECTED
