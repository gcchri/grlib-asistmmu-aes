`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0uqPeKz8K876zFFleGIn6ldHNFpoLJRls3s7k+rAdUkRw2Ae74ocj/ZeyOjgCXG9
uGHjCX2cBhj5bcEeqrhzrzKClEP2KE+NcRj/73PqIGRu8v40/xhMh651GZbyAbuK
lcykcFBdu7Y6NnVCMZ6BMNImlpp2JfgLuybG73is44rEFbMgdOoN4FiWapT/gtCz
6MSXjaiZPhf0YN8vp4yRliIYxXJFYjClMffypI64hIihBNBJMqdTZeZoKLxfT/dY
19KLEFkR6Tr4kosanYVi/3CNc+vXc6UK5hc4R0UX15t/0+8ETYlInjJFPn6IPB2N
+2+yIhuRIrEX8nXEXZ/jRI0tQR4H5LxVBJ+tzyqLanhnNQp2/AiQYRR49d6k1uxA
7ozLoaRYJr4dZJ7g3aLG668rj/Y+7/rHQaIoAQUYeNm3e7cl3tB7SBFWn2EkZ65k
5rVYJXQrQ/GLb3mJNTlWZfcaADXAKlhebOuR0g2ZNe7wDjTHzHbOzaMRTmj3c0jY
`protect END_PROTECTED
