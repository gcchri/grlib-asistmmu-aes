`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N4FzgHWyY6vCUPCgsj5i9H2SGnxqoyGFExCuIzOa2DfhmyNr5t+UvJMNSS4ZiQNJ
XlToLciTOtGm2eKc86ttCunGV8Cpnv2iLXXvG6cq+dT62h5lZJIapwzc1pL4s1MT
uAbPGKt3e17fNLbYwa5q2JSP6dBEojivlLtKGQfFk+z4Iioyujo84GuoZgctMCuE
n1oduIuLwXpR7fow/azOvubXVbq2bfz942PjAyT/Mphyy6EtLsh7q/gA2vJwX+pC
YTFb2Mey81nEP010jUVGYrV0I4kXP4VehdbJiuMWkODWwW1cMsjyv7WRRLjZQ/y6
XcPdGLDF7dyoQNGkx1YKV+06pO4AxaspudMO2G5Z7H+boKdwdy9xJGNGAliPylej
JhnbvQCxWnZJT1jyl4l9d7gWWLnq0sMAxQ91SUUABHTaway0ghhR5PtQdTWXl0W4
uDhEE/nPILxGc9obS7k2l1fyNQj15mZxrrc1WVflRgKI5sEpp/SiKNIuICnyvkBL
l/kyThAfTPrQKnExX9sOpta0IHCaHNvIBBKtxN1zoHyBPhj0TpIgdbGrWjw+bpnb
ubm62VsNiXIDHFhfMnVX96y+nzYfaF3hHphu1c3sgphecdExmHi+pQHHxg4Dtvuo
JJloL1z50zPVi7+1pbtxSHCpkSVfBTkV2y/ko0LOaj4=
`protect END_PROTECTED
