`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FHLtDIh4vxuv7PuxpAKNi1jWqMeIDxhGC9LBwLD1J4+1+3HJRmnN14gbYksLZfzZ
6j48soQ3xsCzTSD4jI2IeGVGscNnXuYWSQYp3MeAfWKYDwYQgJTBWHf88HVBHxCh
Xw18/Ze9f3lYf1hiDw1b30E22xmkChVm0XUA2gx2i2GKnwO1o5W6SPx3StVqHpYp
e6cDnTX9Ego9dQG9Vnd5CYGM2iItK1kJbS+9d3A0ZNsSL3JKbBTf5QyM58czXTNw
7pLwi7BUoUrLAObD1yFSnd2x4r+rGOZpZ/dJx7crpxBwOkYw1R0EXDh5UQJ4XpbG
u1uZ8eb8RsLwdf+SzyfJ36HK8QTsH0qCA4GWHDoyKMGPR6PWOB4zvQsD1rAb+jtZ
Fg3N1LgXRQRyszOt85/cbyFNPTugzo0BCKn/tF7AcW9ZP2WBBmrZJHC8tcKPKcjk
shRU13OCZnPsbavZRErftO3PUvgOeV7dzpt6dTDlbW/nS2hmFP5T9PRZVFWH7d37
sImsxrBnpVWx2w7fVkrUDdJ8n9KGjmFhLeoepIs/C04SvrXac8S/J5R+eLlLLkzw
`protect END_PROTECTED
