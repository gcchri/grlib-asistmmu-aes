`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H6ilHCam8/lYh5AARFd85xb/AzZAdV/xMcgH/4XWPVSFsseFn33xI9rFOqIh25MB
YLy43aybY8uaEj1casAjs63cCavV0Ic0rLdf/Zd5ZI69itd34FyIdfUBsHh61lWw
4wPwBLVHwIfUmJNnuU5UnNUI1WcSJPDKl/8wy++SACvn/Zo6rw3YyZ48gAEskLoO
C2Y9e+vdNdurMhP0gFC893gwDFQF2scLNugcGFF+CRzUJxBDOadUNX8XNHDRkaVQ
EAIJSxFGneHwMZNTXxtQPAQwYSCv7K/5xYXHmsbfxyBgFpoNpHbnCJnRAUdjSWz6
q+HCtiXAt90jllX+wGoSAZ3udTyZsh0mDS40lVR22oCjLfWQzT5Zd6YmIKvyTGUW
16F6Ya/Qy/9n2mt9ZdCiMOUIz5AQGxEWsacXGMYAc9LF6glzyJJaEU9XLYdR/qCQ
f/0M0CGZp/jLvLKlsf3JvsSJj5JopkcwgWMdG7+Ts1eRx8ap3gkYvYpSj0kXep3Y
T8+R4dl2kjWrOLrbTvokqqpxw45vMg6OQYAmsftp9Vt8DsNkPrI3vWQljILUgqrG
y69Xm+tqGQyD7k4MZdhnv8K/BcngKbb1m2DyG4EaMDVzCPisDiBNj+geABmp2mD7
FV4FBZ9gonaO/ZjwlAyHAw==
`protect END_PROTECTED
