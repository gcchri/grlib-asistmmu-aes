`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UDb41VasYqaLxI2Xt3xq3vr54bdgzYaf9pIzHbzkYOWmYlGmanvGAoOvan7RlElg
GBoGCK2d7t4pV/g2g0PZTSW9v+JD+ACXtDuWMvWLSj4Btl/gOYak+bnxeX5OUzyl
AoBmh2YP3FMMtbth4dNFijPbI378WA5gPfkqitO5ckfWnu4d2ghjKiH+ncaMPokB
sM6+RZ6gQXYWV8IDmEUeaS7k43Ku6l5P1gSF8+3AGS6H6ZFdUgY972amjPaQuLiT
EkH9puovL3fo7E2bNDWMYmWCE1KjtfKKTjZ6WT/p5oBO15Uk8wnDRJ7rR53kUjNO
ht63BcuGw3N0VSLBu6iT5mgJqVRaeYtXbyO3E3s6j59R8wliqpGLnBPmbuP4t+Ns
jARznNeOvxj6RKfUGjPAb2d+Ju0vSyzDSqay0tnPE4rLO7KGZ0UQh0EbGiifoKzL
bG5BOrH6eWF4t1C7x94eVainVcMzIlYLf4478hx4GCDxQuIQVHz2VrK1WTdRwB8K
DESV7Md1mqtC9A9QT8t0gbrNcQb8K74YrHiv8RDXMAcnZatDteIxJ9jxiQD2WaRJ
u8NE5M6VaASYemFVq0xgvPHKm/B8JOXgmGMmathsXSjFqcNTSCWuBISb1cpPD2P5
xg1pZdfIZ5b0kpEBlk5XmBYozcsz15xdpQYJ7ZpYezIzrt9jOUYcg5kFD6LykPEW
HqUXDORsdXnSiLFsgWnDditItCXs5Hheos/XW1zJTfSFqvkAFe/1/R6pu9Jk2tNm
NkGYu0Y7UcDg6NQQco6JuDsZTCEX31uOi5wLYJrZClGbuYvr6D6TfvDIc2rWzOZR
UFQ9w+eSXux86a5JlVcvxm0whzEb8KWUyGJJoDU1zWVIEUEa8x+IKbRFKZ14+Oo1
oxiNxCZx2KjZ1xqQ6+D92AgaeXTnTMZN6qKOxiaGW0PZtZkh4QenrFU9jNG9YZ7r
D5CgC4UQB6PhFtfHb8RFE/tOHitMmW0eG51+UDklJocf+w3cwn9kzN7DDApWGoti
hznhBVdj6/Y5v6FJchXZQa1OCQEHQ1dWCSRr9JxBQJAI5xapOu9VkNqONq7IiziS
6DZPYYpljnQ16TdhK87t2WRlkgff3UOQbOMNHEkGaaZqWoGm1uTGVJWfEutoZJA8
VfmAV0/4gx5s1VkabYLOpzSgR7MdOZKGxnMZ1nw4FBSEc9H/GX1OOVDzhK/46lUi
jJP1OOdUx8r3qsxQrZU+/pVC+XIFuI2XLgcIM+gA3NypEAWeVy/6Blq+LxEoGBmg
DIWIpqj4oJxgaOnRhGMuUyzBjIwei0xC+DQ2iNkKFU1YfI9ZgMLVgR8LR++Vactd
7w+Zy/WcwZAv1rCNPz7BtapmFMeehvRGOeuw1dZ90tqL3NDe56eGoHH2N1AXOdB0
rJR/6V7tzFpdnmUtTg34KgwR8t9NorsgZpzoQlkd3v6R2u5bxXls+J1FtJi+mOhu
cnpBbrKRDwyTxm9Jt9bXCMAkeJwksUHVm5Em6bHuY25E7gaXzyKMHZx3F0mKhV6h
6NO5p8tHqJeTa4OTzhXpfhvlr0G6G8+0Ivua5T/BJH+eheoBesKNFOB0upGZX0Al
vuWoD4s8RRNvg710+8lQKLdEGDFRuBHiqMKzTo71r/Nk4Fr/TItZg4ruNeEMgHiy
3qI0huYz3vz5TeMvNuBZHnFNgL7CKaqmkjaqSghH0U95sGCogl/HtgJfja2iDPyT
mMPwE6NzeKtq4Vp/zgagXa3MCZC6y0lfSXoal/CKCoQdgdR29ACWXTdP9z0ZuayQ
/J6cImMcyG2aZ1yQMzbk3PZKMTTgJw+/rmjAK19z4dmRbq0tttO/SWTs8qHs7UOo
V2Xng93lZrUZDWaZhpm1sWktItOoKjsZwXIS0sYGI2zCewqP8WxQXZ0rZX7qAksC
zSKWD+DEy3n7x2WI6ccej4RHQ67HGJnwc55+nurSZZDU+4YUjzg6hCgFjGo8kJdv
y6aP7x+jWUlZl3r0O4ERjdRcgjfsFlEpsfz7JM0jspNd8WWHEnLKWQElSXLgNGjk
yj9iH/KD84v5eRL+ZwDqOU8fK+h3q8MUz8wIfXbuktpuFRrvo160ScyckH66sXvg
nkHsIgKOUbH7astTGeH0Ji0I0NkPrS7xREi2vEXQpw9vj7RDIMKo3opDlqph+zG4
mUY4031eq2IafG/bJGJel72BPKxaEI6N4E1AnmAmo/37LJKA7pkriI4IZSFK7Nb0
83pi9cz9+JBl3Kq2x5094o/paXwFuwIGU8nF+Wx+N4HGHZ92GclZoX8iEZPMdl8U
MraKhgM4JdbZGdoPkoSAW7FnmJ99/ifD+uhqfxwz07Do/OEbj94I846uuyZvsc1S
38ZUBhMZleQtgKWkOzk4M2A8VDWz75wqoEtJEpoGo1ygz67VCtU5YegSVwBe6H2f
Lu/+fY5HlvqMFaEy6MBTcL4Ke8OGAU7gA+1mOqo+spow8o7pFyZv9K4eCgvEuEC4
/P+xk6eYh8WoaO+O9A0+YuveCpVR9f6HQAgbXNOVp9uImwhiP3xW/qTx4Fy1zta3
JKXKooJX+Xa61s04mRXQ6H5LvNZy9PZsrmGUWpB78UUrzviqt3TDS9WqaPCo8oys
llrMdhCS8cwANvSRP8UYFtAYavK/Z+m9NyV8MF03UFBR1K/v0k5stx9+tRgR4xSN
zS9el1ji1weeaVh//t0YLkBE4cpI80FwwgkAVScv9ZJzjlqGAHOZjjj/G5cDKqkO
0Lu0KKaTtsQe37GxUHnxj8os9iSoyiVNqQEnDEXuNTmm7ebxitkj1cIR5sUakMaT
riIUR9EjKW4vdylo5ubzc6wvrc/05wB8GYpzxyK2Oczmnz35nu1+4bfPvDXQgp2m
SU6EkKLnUvlgNWepCLowFTtopGgzYVkxWe6Ne6JxQzfuXmL3ryRCNXTG0BR0WAdY
S6t0ApzCDD3k/awpqR5ET+VAuwUC5Cc1ejJ+WCF0WTcDoWIbA4EK8OiLWjWedYy4
+Xv7Ue5KLs2Lvj2ZqgoLHIJ4/AErKKOqGqos3ggBMsl0ozqVJdm/eDQxjl8m/qwo
uTnnHbsfogeXjbuf5WS4zHZSzONR2zeIo+tZbSaZ3d6HE6kUEDoBpneEZ3rVdN9z
laOPB4nGybR9AMgqCIGueM3RXizKOF7eusQwyTBcomPBorNBVIOQLQpJ+wrezDVt
L5xJb9YuFumDkhsuewztfirjMvwkILW5De54wUnQicOaD8maJNOzjhywkONLCZGC
0LBtkPuQbgmOeh5jwsxvma4v7NaGEWZhk5g/ANffCdycT6TFwq1gS0usjvgfrDeh
sv4n9hYTk9rRR/+A2S9JVid7+4F28ktMWTMcV36e2POk4Q13PM5MaqcBdeD5fC9D
deeK7GtF7tQUt11GNLehm6NLVMadmVjDWQa42MtaC8pP1K/7A7oz+w2TUp5M1gpM
hRDGumpTAk0NZ/lQMl/qVXdWl4V6tXdREhGJHCupDpq1QZkrmQiLI9K5PfLsctiJ
Kx/CnYHR3DKlgadWoN6hIo0uZhwbGH/iFYZCsUisZf1b8cbG527xlFacX8RyvvfI
vLUWggm133IMzQEApvxz61OOnwgk7v8q087p5st73+j54AW8ZwT3/ouv7y9CZcZM
q5am6C9tbbxOH+LmXPEs8PiXk9x0DoqgG+YMY34bz1Ww6Ne54umztvjlxcQIwjIp
OGNc1gNsetp8Ba157jpo/VzI6AOLJ8QxAC7T4v+6gW5Mhd3C6GwbNTPW2m+HAeaY
CTtuKEB1T/Hj7TGUOAJKhsOaLJ0CoG8HgsLktYxGcPc=
`protect END_PROTECTED
