`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4gQJGWtzZq24RX2xaNsKinoZVQbI831ldJuiTmVcMwRBGN5WqsxEzFoleXKAgJG5
nYDGMclqClbskL8/7emw2dZmNgFIoEddmI4onAbTwOj0+IzzI3YCxUyJlGID4sVA
HDumV3+c6UsXVHAEtWVW8JeBMhdgcrYh18/6G6XLh5GVK94qu30RTK7XPPNJQQad
SlWC0Dl4ei+lAwOoTZT6H8gBKOD0aIT4QtEqe3bYfMWJg2U/VLypZckWeX56T/Op
TWGx1h3qO+GBvMzgy3dnzQ==
`protect END_PROTECTED
