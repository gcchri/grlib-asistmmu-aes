`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cwoMpnGa8kMwI9jTgLwrqbKvK8rYDVLsN37HDE1q6ISXwhE81caNrDpLoK13Qyaf
IlZ7+JImyqdTSJTyzl9/dUbjHTjdQyubu8p6ywz69rwGXjqrE6Kaz9zgahMpPrH5
sShn2tLPWYjfL1unV1Yr5x2uQpTtgOjKlc0RQagZkyUntCibJfuRFTwI+C2BShX+
CmNXBK8FsuAf3pjJpxUBABC+ZEw32BKEYVZQRt9eDN86E6w+VgOLkP1pGEe1m0dq
eJOomPwqtNL5LLBn9NpcSUC7nnatxaSSRW/nNIGsfOYcgL35Vbn0vEZIPH9vhVXN
`protect END_PROTECTED
