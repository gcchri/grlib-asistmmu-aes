`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UkoGfvu3qNrKMriXJW0uWg20ORrvsL4TRplgcuNBOGDojZI5PJHODhDuIJYuQlaC
amNXuaGI8FoG826YI1X7gXJXSD26xQpQiEsWBIGanGbWT4qaM9pI1e/Ey8cbCAuK
dwIN7oK3lQJGABjdx42ZtvXscXRx29lryep+gRcEisrChT4BueZB2cw8Cp6wJs6e
Z0fgUGBFtg1it5l7gQryCQiCXt098aOqxvwa/pUpifAvBH0rN6RWIMCzO71cUroc
+rXmiWpk18mqLdGqO+i32Gqqy7MA31dBwzCWmfesS4DhgaiTEMrTPwkqhB5YVIeK
VGXG6lkGD9OI60sQMQ51mPd+6VRGrcjrJIPcnqTw0k9oEm+Kkj/MA2bFmNnj7Kfe
/H5pyRy3U/TeAR0NzuxFtathuM4skzBBmqRZkSzXWJfWwriSIB+xInP+A5qAS6Hw
/4Q43epMnbnNh27t7K5HIMPfY7jT+4pdUqmhiLbc2RC4HnIX3skzPaLkHXvYZj5P
IkdLzc9WNVdtpJluVbdR7mhaifagoPrvFG+JhqiKuszDsEYFqnggHEQRZoABL8Xw
`protect END_PROTECTED
