`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lUthElBKvhqvApbLr3ThUA2KXiBbsMPEMKj8+bTXfrQYdcuafjkCZDK1juuk9oNq
s9fFgTT4eWllgZ7wcI00NIePcEtwol+7OT1Ae+VdH+kjcxnf0fz7ZZ2yjSZw3voy
CKsuzfQIhDmJt8GwoucrJn2e1ZBNOj6Fh3PhSRKfaX7d0uO8WepHM/x70RjmheD2
ZjK1PdISEO0viZeAM8YXKz7xwnpIwqnV94lHnskdtxvDhjngo7+YUvN6n855ushD
KGa7Iwb2TZ0c0yBAUXabM0SafjCf6LKyMM0xoe6nNczW8S8N0gWVfFOeQVb9Is6K
oh7u8rGrDciWXThYAzbdz2apg47mQ6wvDoPDsI26KZ5ANxLwUYXzTqDXitiLZ7Fx
iAJbdYgvh+llyCRJqGeAD/KG+ubUVfUYi5Y8YHP+QHw64kEwOv1Xg/Prhg0ZzPtw
`protect END_PROTECTED
