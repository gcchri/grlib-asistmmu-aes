`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f3V3+oVBGteTAqN3cS/8eO8daZStKsc1PMVSGnbWDS8FHS1U6alXZr43bYyW4+fl
296xjyQAXYtBAspEJOsbpfhUk8jXpfPTXYTQkLJUUZXLmmqAU+nmVyYhgmGAgYSb
J+VjTs7Kx0UQBDToUvZ7ENQI2276oPuaDZLvClOpPqJZocQHYUPDjRWG+TA/S52B
bkU3KW+0qJNBUVRwVOHtfjd26AaCiTWGXuphZfYmTUbVBLKRbAOeXO0LKO3KXJro
8YHQx/yLsP56OIfGfC6ix2A5qRdwSdLqG1lk+sXUXil8Y+Jtqg/CLWfiOOWO4TRe
VH33mo/UpEpcJIQ/nr1h57oUnFEOuMGGQeD0k9+IU5ynSLwz4TIdUQRahOHu2I/b
wGkd5X1tyI+2/iqx0OvNmrBlOI6aq3HKBcHZU38f5fmk7oGZ3qlK9zRyXhJ9YLMD
HNznN94n9f5TaPp0QXsFGULtUhMrajzcEJt1kQOKmyKZssImL4kY8xfZm7MhWn1n
H2FMoLjY9EgoiMrWvZrzmbbPHAF2rp/65gSBAtOt3uQdO7Tw6Fsc+XIHdvHAuGVF
kHoV/r2IM9m5JETfxpw7fR9NTqhq5k2jf4UxICeXlLuf6xwRwyMACSkOTq1o0Jr6
gxJjdnXw7E2pu4wplU8Kk02yst5lFQtTJaJlzRPgvmPbIWn69Big14lqQNAPzw6U
wlsOJ8CmHNN9tprfv0t07ZxpkDZxoQb0K+rG3Qv8Bj2p6SyMipi/vrSe3gasfAd9
CRcuqftF7osxWPJbUpqHYA==
`protect END_PROTECTED
