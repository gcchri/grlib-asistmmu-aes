`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OWCxS2d20hd+lPdwkmo8+0Mr9NpJ60RblVmATYP6bpQh7PbrOdm6mhNTE/1x9vP2
ECaL0YmQW1x4EeTUim6470yIcOQw8g4UqBLz9IfwUEGp2NLvE7DPSAE2RmCvSkjX
vuMM+MBKmIpXI3XFajwNJD5AdVUbMkC5A6I7whIKy6TWoQk9vc6WH8od7+0bEXOz
2er94Hln8OPwHa30dq3qfznMLmaIRTGxdsKMwwO92ggwMRGaiXQ/2nXLI7gfGlJw
o+AGIxhl9R5kHd8UZzJ3WUttfmG0tjVqw6D97qGjCa4FCe6QmK+ggrg2cankCwt/
i2I8rMOyCPADCtiXHgh0F6b4hpf9kMnD2D5lVb2LrV/7U6SVBhIilziMV6Iz9kfo
PYNIR5Vh6DbpUVl+Z3zWjWNpfZLoNM9U5/2Ct7FBYk1Zef5y8KrTiw3iffMtlvT0
f/NzOY1ss+VhYZna2ATCitr502Z+Gp5kybQDQZqMEqPmruBwSOl6+b9+F8G+AztL
9gmeAJo7MNIDnBIhArdk3niv4UnFYwC4b0KQPYlv2YowaUpSpjJtE7qcoOsFcfGK
F1bxLi6IJTRwiyqrNu35tk/OXYPtP8THVu29Dz/nxMikUrc9iI+O3OlMTKrmT7Gt
5zpV2q4TTLJeKGnPDn2qMCCfMPfkAnYr/zYj8ksm5mEhkBKXbISRkqtyi4BZbcTe
Mhdg67hBX/tr6E1DXI8VtEYBl8MsDbIIFhMImmDxLTRp/7/FIOqrtUW2AqsgLzEk
E3afq164jV+goF4lRwZty9X+tYYm2/7GELu4Dj/IHnALCc2vT7LLaoyZ8GkVEerz
zq9w10QLTuJp3kacxhADeEf50ywP/zdVJLbdkyIkxM8=
`protect END_PROTECTED
