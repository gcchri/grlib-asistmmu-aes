`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y/1wLg2OMb42+eELbkKcpdNEQSB0D2ZhsVW3JDp7XttrQ14bT4C184EcpsNyUFDH
9PNZmDqCOebeg9gERZWsKexdPT3CoSpF4V9pBiO4iy9cnWDvk2/uNbHezjMZ5pXB
cmdM6ck/WotUPUBduKpuX7VM83JuSNH7wLq62b08OxXFzQAGIq/Jr0PGKQctbmVC
JoRikDlnQP0063HKTxbHkHZ2AnZ69P+oWk5oSyW6dj9rNXONnEbjjcyymL/5qJf1
O3noS7pg5Zm5qX+hRu/5EO2mikyGHZFreFI0Cpxe2ooZwscY/oJ51OozcODzGp4c
jjH6PPpDGcbbY7LrizzO1R7FyVA8vszE/z5nos4lPHPVM/il9BcNknNcEMJcU2ZP
5/9KGor6RuJx5ooeB43DfUysNp4OTHKh+gBjvWNR03aNyCwPnD5yuevfljxcSPA7
2ysaWo32M+/O/2uBRBwKajq6E6x6uAU216Z2nhIqD7ie7GluJSMZAUhN5JIndNAi
dZd2TeFuY40BYZc5Hiw2AOOQHRUH8F2cn7mC0DMRb39BTWmM8G4c1OAIz/Zdlnwc
0Lb6abmToUHcmlz2jEga4E/knY/ivBMW8oIyRQox/BdYj1L6JJtLByR0D3NsDwTY
v2GZNqD/pW5LtJlQl2rbiNOe00gdg5VCwxW+uwvne9zBx2QyY0Wb5NX/9hPkxKBQ
QrRLw9DElT8cwEa3Ka0oGT/9veiky6UaB0h9UB0mTSW5rX8QpConmp+6Crzixnio
i9TcwZHaQ9GUcxGbedC9XatS/1A0RcHH153lQKmMMtHDf+h7bXqztKTw8hRJ1zdP
C6ZHJwIGU0AKhh30J6PpqVvpLih9s2BOrimbD2T/7sR4t65qk9ThyQ9uHA6xoapn
yiaf2Pgz+rCVZ9MXuZenjw/vfs9zfJJfLqsZyS3Yb4FEXnw70C6F9hFMDe/lSmWj
oH2qfH8AREnQRoYt4OtU/xYhPHs3zrxIVw3QsgL05u4E60nLtPZ0hVIAXNebwj2O
gt6TCF6p7QUaMZIr8+ZfecWtDOYqhB738VVQIpbv3QM3dwIbbeww2U2/AAPEGGTg
WVtoOon+IvueWZIGXsKuQZV/dDBRXmQXqSxsxurzVZS3h3WmqrIsAbhAaCJ15Let
3jIJtTAvYYE6efDhj2Q5un2X+i3xXGSOzixgwOQDA1ASpFhHhbuRZ+Pv4M73VOeA
EMlDXzTJQkE7fbFbECNzDcV1XAqsB2+/og16slBifdctDwn2NrRWN6Elwamn5Apj
2eCOxAhKRvXH6mCPr3+IweMsWAOHVnYmMvCuxQ4AfrhwObHEZkvoHLMP/1H3c16s
XWzHfqB/IrhxErsMEQsiYUuOF+/4aQ1nHM0zU/VfVE4RcXzzlY4oITj4OAvtz74A
ejMpOovMCCIriNy8+NGyltFPJAf7FZAg/krZVr6esRYtG5rNzKRGmqrZ20+JYPtK
/Kf9euj9nwkaMibS5PFmSt+lD8YMVR1eFwf2ChybdE3Txms3Z7FVbtTYAarad3GP
hVtCwEo+T5/iU9OG7kw+JuAGwjwlQWgz6c/kSnWLPHT513gfMLQbvTZb9RVXdPsj
0Iu4rAh4sJ+h/EHnF7ob0DodV5+hlGFxs/SAFfQWp0kdzz9yjVBSrpDEgTG2LuTw
ms+mGyzkSL5XbKPT4PQniydwglF1w0Xc5unWmmqySDFjCBlh+bNYNg4TLKmBI3xq
Ye+QJooUlYfXopaF4KIHQUxyTJ3bpFCdzZ4fCIRojexn1L+nEW7R9hglEoIAcJvp
K1YxM/FAbpVsv7DaBCjmbypRIlmQha40c/cMRDIb+ghgR9HzJm3gFexNWwJbezGg
SWf/8+o29rpmEkjoV8GT1A1s96QPNVzzamP2bwbAxjbMb0d9qgdRD7hvdS9vSXya
ympADMrMfwsxzErOLT9/7OzWtPPmXBg5HBUiW4OXDb94g7+2wGKVNNhaM98U5pMF
yerN9nVrE/HquC7817OGPgyOvLIB0fbZuJc7QPEz3P9+Ox4YbzutTBJJq01zAs83
FcKlHdSrK/N1hfYaTK4eW5SyfAT6bC48uSPfz4HJM3u3mFqVGEEP6OVa5YAri52s
lsN47AwcvHJu1jbcBuhdpVSSuA7H+N/zgSkEcVv39fzO4OyLtBeKA7+3r9oCszrY
YbKaYx+0x7Jn5+MwoyDKExC/PWDgrwHrGRlmMzK5WNV6LrRgX6uVajINqC9u99k+
i8j9m9edX2G0p+BZgppXvmHLkaz2/1wUmJqEYopvz0VMr7N7EZgv91FqkIPCVPwg
G+A7BX4cwrIYgtq+IrMGBBQMpLd6+6LFxdpO7Tg6QgwwyaNQkDawuYoaNrgH9SFx
rayQTtiyWWCfYEVMq7vOkHezoEODRYkfbYSMAjad3wH2cOgc07PwYwYViJs+hEIy
mn6AZaB/vIGQQuwaIVMAG0hMVw9LZ13At3bHYInzQVkL8wzl8CCrV38yHamjgm2r
9WVBUFt50g8/fWXdIdVt+ZfpDn3SLvmnRit71vW8xo6l+n8q7Ms3+PP6DDX+8vmi
ARB8MPZf4CDD7/0gPvZTVCYY38qkGJ29+omGQJkc6lVlZRyWlTQARk50yUZnyEI8
EeE+Ik/i8C0y+M7bNItfMDPYbdCWbMn3rk2DTwLE909mvpnOkvBI3wtcCNswCtNW
I9ClmmQuEeLm6hgxtfW7GZMx0Pj+L0iJ5uaqUsQNfUI=
`protect END_PROTECTED
