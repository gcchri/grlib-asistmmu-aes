`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aoA8NBUvyooYnUD5RbR5nNf5ohUnakKT5EIdQmrJOBuQvcSjPygQJcjRC58GtTvM
iWNokL6z11SJhririMyImiP/uD7Gt3ao4zpiQ8FTMuf+LDkR4PaBBOChPWTbTWAf
ZXwLaqP7OtdODAQnEORSc3n407j7IRoAhHfnkImVu+voDBvFir3Ot7fCR2cWmkzx
cN+gkQQa7hgKvKKEiuWfmoElv+wF8NaoK9/keGHgNFnarP/79pDrg4hAiVBaUDNf
KR80fV/2lJzEjSrhjRVqOKnXuCq5xYx8LhE/JegIR+8cdHzc6Tb9NgnOEBjAQxWe
rgA6KDJy2xonQS4EyAtYY2gCI/z6hsQPQSPGpAhpkUnd6bvGJx8/md8nSQ2MQVeG
ONmDFFJeI92RKQW5+K6zhe7XpDfKBT9ngYHf8CTEp3tCvOa/687YCo7lesK4VPfh
L3k7DPUNbaPpKozatmrfXUcZnfEBt+AmT2wz7vvSw2+LNAJcgtebFjk0RQQkeTCQ
QLvbzVkPBC/H4vmwPqOAWFEO2EPJbNN17DRzxkreEg6xBJepqPp/8ZFfv6CrPF3B
K3n6IsfaZrT/IsSFqJWScZQDDwGtt1/4Rxu2OZQulY00GijKGgK1tmMN14JW/Cz3
89CnhlS6FG71arlL3LNz1Q==
`protect END_PROTECTED
