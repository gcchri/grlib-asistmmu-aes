`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KJWdwH4yaYk5co1PHZTXn2io24dBgEwSAAGUhER5ShCLWGiZ6L/F6G8VqAFxIZmo
Nskx6vAzKK05wUX4eTTZmL10IyHjWt6Cp2OtLHoD4D5o8JbiRXq6k3xmq392iuNJ
hzw8qA1IKobtc2Im3YhGDiJewox7lW1snHltCCWzYfZqzTTOI3KG7mr8yKTgWZVK
9vEEG25e2fmCeUpFDcQNgLsOpp0JM4sG/Q2lKmkTFX3oO3y+QOUkZuZCNVe67A8E
ThJRMpGaCWJKU9i+7XRcWPXVPhSqhYr2hTZSQRzyoa9twARD60vvMZLeXMAh7xma
85X2Xx3ZvX0LS2wVvCf1s4BpFGcsrnVouwiIvGbAsCVOz/sMXUAWwb5ntzEBLg5T
in2o+JKh6YIEJXAVcIYRtG5IllTwRUh0oR/QNSWWxXlcgPpxHuFrm+SUdP/fKNkP
KYpjBInCUGSKTWBGvauscEoW9hlVBu8F9/2O79vIK5r4AfIJpVvcUNul3hCqNNBe
9+HqmVOCF/yoI8fC1f7H5BAXMmc86jHS6j0YmXbudpgkgtPnHgKBo552T9+8Ykz+
sDsHpAoR8r7dLp2EWYcDYB/7VogJt7cQHuuYmtTpn6rV2oWwatVFXKjD2Bng9T8+
NemUvyEa8SelkVzXW176FEbU4swFeJsghk/qrQbDyp4/YFIyghP8Jzh4QQMX8AUa
tt14PQDgeoLBxJGf01tZB3ljP/KqOlXyOKexcTmUEswtE8zbqklqBV9LzdzQ3ekc
LYgyBuT0+SWZfpKGZ4FmdiOahYXjSYY6t0rNbfg/ZgQ=
`protect END_PROTECTED
