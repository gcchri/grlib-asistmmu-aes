`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CI8xIKiokhxAs96tsVKDmw78nQEfr7a1UrEWMolcbZQIKKGgpVWWtWGXvNxHv/c+
eqaXHsrJyGpigsrJ4vza3F3M+wHj7af9Lz25uKzqpzmtevGx0a7UNS5wjsvX3taO
K/JowYHqbpwhfd1YBNDQwAm8K5SQ3NCuqAfWCB+2czTcyJl8vAmSOlvVvDcx6jbj
Jg9Wjr8ljtt0fUSpwo+uw6g1Nd5pY2Q6b6e3HCwQBdtA3VhNC1nTXBiWUeyxJ4tP
FOzDoovdQvVOh5hUbPKK0X/AkAV1VsQz7lCUrfcA8jyPHB1Cyxtp4iEldYpYdZHq
rRgRTOJzszCPKazI3Gtyv8m22FVQiW4hnLmaGPgwAKV5FWsXmBUVtd238MeCNPZ3
GFkZ/edbVms4zLPl0hh8RcPd7epEi81uPa2gpsQj+WjetOJVfwnpYXwPvt/JYiwJ
MB3d1IdMq8F2jQgibjPlgRj9LL09ARWObVRte0yov8fQrdA0Uhfa5yNEpLCCrEnJ
`protect END_PROTECTED
