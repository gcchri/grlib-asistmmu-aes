`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3hkqgrOkmu4QEaEuv+BzTWd/g2i0rtqdrAWpBi2FajjRQo35z1Szi9/t0/mJkAEC
NfQhLVusu16q/wT50xqVbsl7agJZTZ8hswjwFcxMiSCdH1FYhhyQ0S9ZWXfpD3Y8
Pf+cRah71QLBrvUwIw28yy/eybhrALb5Rjox+ENSvvpumLSw5r+22V6xPNouoV58
M5VDvG8Rb0i8O2Waxyhj8MsbTRqdPA45lR2tJ9+9Ea5dKlM1m6ss/LPGztiVwyto
bf9FufX+pLhktA6eaC+v3qAwNh+ko8msDC+dSMRmCtc58csujzbhT7NW7d6ISta5
6k/dybYKHSx0KsYvAzbg/qXVs4TG2m0knLZj1l0MuAivaEin56HcBaAFfs5z+QpE
Kuay9Cn3pu86M/+yh5TlP8ggnCVpTzyFYfSI/qehO34Rp+4y7KIRCFcr9WCznXNB
l6u7UviC72db2z8bUqVsWwv/SNW0YL2584Sc/h60vh94Es29ILRg29UX7NO/9l2Y
cSFhuM5CFPXUwap/ND6doJQQdCrDy4S+cwXVBEMtHwRhD2JpUzu7gnMmnt6bby9w
bIMAejLJM6SY52/H61oJ90P3xrmgCnGgVidWbX61K+/tXVlr6MePAXd07oN5/OSz
QBMykM9zpdwqjPQba/LwHZIe1OPqkbTcKE7UvfHj4BIv+gJmOo3Ln8p/jQ4/cSH7
Pnr5yZO6Tu3wpE5gnkkFrPglsJwEOKilk07M0gMnye+eHUWZJim/Zvdy5Y2zL1sA
jJ/j37P9Tblxlrbds/CRbzu/+iodv9veF7y7Op3+PE0gYSIx831m9hehx/PDCwT6
JDPmdfbY5nJmxY0oi36lFjsDHTThzOO42Bo82PM4az0K2hsI6FKt0F7vZ7Eh2dST
8gb/jpJhfPlxNSkKzoojwyGgLZmROBEfunHvh8/XLgzhiCK15MRFv40d5awQRDvD
rxsZFGAJ4XHMfWFtHxcn0V2HxvJV+hzlRIJoX9c7Xk3CWi+a78Vh6r33uY1niWoY
u8zKNO/p5HZZrvCnmiVKhm/2YNUss2KPx8RBDHPLvCfNXr4/VrTHBYeDSuw2RuuA
1PPqZS7+ZLleV9RqLSRgxurfRvxtTFehgewG5etb0hZHPMylxJaHUQnRGIPc3tFB
4NRgVrFnzPySNbe855OLGfUrh29mNKUTUScHopQ/de/s30gqPo4RqX/kl8+cQ2g8
duoDnjvD+I8KaBwBKllNCgzWD547TTi3a7c5YpdxlxJ0GJZ3oKPICzMOgTZ4nGIa
WgCLYJ7G4WDvo4w3olrb9omDoDZ4j8WR7uFrkHh1vpuLVxbjXKkcFhOFT6hR+ydZ
a1F+xhKmxHce0dF44jJWP5ZGwsySYKcoQE18uu23koKixX8g9b8xB01H3lSK0zNr
KjyBqmI2LtoZDc0snwWKlsdhpYvl89WX9M6p8zO3MPrJUYF1GznIBbV/VGrC4e9B
jFkhJbLKyaxje/82AhE2Buc6g/S+RUSdnEzux+2RlQbz4PS1w/8dhzNHsyCSWL3x
DbRpnXMhv3S5r/PUaYTjSSzZ9mONKaJWZcE8pKpTThIWPhmWTHaMye0Xc0CZvt+6
fdBjGXKEpLlSqLWpzsNVfNAo5tOaNxXYemPpZg8Wvxg4usPVKVpgLAIvQMEXAgSZ
zwBb1Oyv7YzrTuZIFtM5oRHtHBmxYtvswkBuH4R6SQ0LENYBtfVg6Ftgr/rwNWMY
Q13dfdRqNKvuxLvLKE4EZK3JMYz+inL7MdCngISq5PPyrFLlm6uf2i8avYcoub7d
MxYsC4559poR8LSASRbqo3sxtqmY2PVb1UAeyrZ6GqKXEYar9wEaHbUxTwJOycku
zZtThk3egUO+GsBO2kiReKFny/t+jg5aiI7PTbzHfViAUcnc4NX4USrWR7jpB9KY
XJShKHpu7L0N6+/+W0cZj3/Df4Mhbd43nuG00UVEAPV4axwL7eAPXGi1ztL3P103
ViOU3Ix4S5RTp7hDJK1uGI1NXvlLogZzfMWHN6PcSGpVX68cDjEN5mCDQMJ7TfTj
ALYq9GuoJI2w3n05wynfT+fKm6XbhX1F+4PHzMis4me1NGXnQkzYjWPfO4HAYwye
t2cGL1EjT+NUAbP2Hn7ap2dcy/rjUyfuLbTKbMA+WFqPn90Heh13SK03lJvw7FGR
RGGAMiAV3v6sM6Ov/zeofy4QS7azS87FcXMbVtfNajqmwCyWpWc7Scub01qfpWto
qY3vOUZWTiR4xnFCpo2nxur3N8P427P1TmxdD1Ynofem3B9ZDgkYSfEmzzzK8ZU+
VYXbaieA5dhZvimRrCmBEagpHFh7Es/qV2xrnfGaQGwbaIpthp8O1dvvVPGPZR3I
tBTHY9VM139TvywpoFNP98Bjf9OFZ1WPtc4B2dnLDBShXTBgRWrtkPeZpj5LzUpH
fgLZoRn620npsOfLChnhBptwDb4F3GQ+D3gP9CdMNDtVoxBMj5vEdFNWCbqsctzq
PAnjLOlk+jzmDdK4KEaW8mAI8sfWthaqqEGmRQYPdB/Nro3Z4+xpZlaMdEXbG5FD
bvKjtdUA+gCgazJyJMndvlB+ULRPzsebsTUo7pDbmkHt2rZ+OscOfW93O7+gQXps
tSrJYDulueprOmRNeTZCV8ohB/qIZbEaq/DIMbpNTrw0TzzCcf3RBMFidv0NOrHr
4/nBTyFzQGdbU2/k4WKAzSUVM9RPx4CAV4HDTNhoAQI3o6BftDwGDYUYNUcLldR3
rEn/DXiM7DTnEV07HW+LCPPxjhRnJthE0gaApqIGKRYnXtD4bDPoURqMRMuTVv/U
e+x1bGBRNtyA6RjgEZ8kYPGBH9AUD2siOQBU0nQuWDXjTkPeG1K6IKUrpSDR30mC
1CL4CkMBAvz0cUqF6BPjVOmkYIxWW5JRjXYxoMxY5qyfsvcqRTPoZssb4dBvwGRJ
o/ho6MheyjDK5zrBd/wULlDDoROJaXzInP94fhSWMw7RLSY3lQtMvg47D2NQcffa
8htb7q3V2tSEqjB5t4pTUGfW0uQsGrocfrUNFhseSW8KfgWPnH898weNhWc9O+uH
E6EBLF9wTWv8OZ5YGfy81N1rPJXSUS9OlsWB+bD6lgMPf4UEduWhyoOAkhlDXSNj
w8+Il5pBbXSnNl3LxYvI3ejXUwLPCid6XRZbgX46vSP9BIutd96zy3sB2IPfqkah
HOubwyGV4wcyzjjxdCNbxXJ4VHFzowNJhx0rNgmZ/StfGiOSR9TwQ+09P5auf5UZ
QWN2TldecQXwK36JDBG2u7bt8XsNkXAdI4an4caETPzEo9Wd+FK6bA9prpJA2Voq
kVYFUV5DzAMw1m8dA9DPW9D11iEqKHskHAMqFQPzDkuir+9IvxoaLKKRf/LDJhPZ
Rnbn8hFNOtRhUCo1cpz27k2QxIIhyd6UwiwKYvKhbDBfulTUAKcohiupCgO5O5YV
h3gGeXCSjuCesVwvzFJBrLH14AhFftH5PhS3DHkwFv5SSHG8VOlAsLm2pw5SUAzj
AXzBpctfyHy7PMMaDFIjFdUG6M/jG3Vg288LiYCsq44nu/FDbi6A2pfnIm9xA0Ol
sCrRM9PkQGsdoMVU6xnEjdh/X85uhp5vJoc4GNoCxY3+WSDGdB4poM8UwvBJgOP7
u1Wk4fDZLvinBSyJ+iQ9Zgh+B7yx7iW/L4yYMSECBjM/0i4QMFkJBmqGGrQjd3tP
U76yOdF1JMLKeA7C2NWE/K1CKp4CnjvCDMZnzbreHyEoSz+pP7GVcvhKdR+q0MQq
pMBD9uH75QX8cPn75lZRZxZuvLpNGExlWbkPjv3s5aal5qrVyKojVtncbEiivyAL
eWCIfbMyOAgXSMvHkJL87aG3FETcK6rUz6D38aJgGUYUGpnuk43IJKWcFgCTN5p4
ClzAV72jCTSYp2dGtoSK9CFi0GOArwNZB5BCMRSKgb3YoylWUadjD5SZUhdo28SJ
NA/q4igYtMprKiWWxYmSSJPDhbzDUp4ZfOfmPWD+9Q9rg6krShNOKqp3AjTPUGr3
gVEkDgm8gPZfP7hsW7MFnvJ0axYja61o2UoPiyYysTudTLRk4bwcynRmj3UT+X3n
yETNHPA0yQVgPZE0eRoRyLyVhGuqVYsEkjZvO6A1YPBLtuhq21rR74fDhm6IY7Vs
n9bg86Wov22FsRfhJQ1UQbo/cCbcE8FGHBcDxtFG1Fj8aYnshIna2xs6gI9d40m/
WbuHBbToSOfXMAQhYXVPNg3jmBttx6EX1+yFG6kPL0tg2lWa1Og3bEp3vyq8sPVu
5MQGvbA5A1iYIUQhnI+d5iOlA1UDZKAwxh1XRVL8XP+/WA17bkoX3asX8P7aQfPp
GG22hyyZINBbZf/edv9gS49K/zhsvK7+3hLOBR5uKWw=
`protect END_PROTECTED
