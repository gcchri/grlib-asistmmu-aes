`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ir9UL4MyeX1fCSee//u5uM9kX4x5Gl/3B/BUY/hIGWJ3/2FLPb4BjihXjDl1+vig
2rklIOH1a45KKS8+IW59ZryXVIaOP1gnSz3am0GxjJ/vTZL6rUSQOk/fRVl/tud6
kzLdiVnjHFSv9IBozcZ9YBnaVLR7PkAcuKsi5qCz8WoxwpF897JCUZRqzY2AquzY
3ZIIyKHPwZEf1EY6TEiqJWbdWukxuU749CdkYJikzDbpmjqjS9nYUn869oFAos9k
2ib4Jnp0BrkBI8AMmyJKUsTGR6+ovT98L7KEv+HfG92ugv2ezKRWOqqsryTqswZH
DNqo4/v9jVFuZ6AhO6Qxd1flwMEEtrA5WrD4TjHu092zppnI9eWGbhbuHDxg1oRl
jhPYE+mCXDMnjsLI4et+ztaMOmAFAUx2TqGsFLZx1zw=
`protect END_PROTECTED
