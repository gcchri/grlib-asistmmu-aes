`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QOO838AdObB5W/l6HmBR4VGISk+TG1mi+fgBv93C7ePTjwR4l32VESut7/SvnzBw
5aeOTrvMQfIQS0xkc48mxOLQzVnzDVUtL/PnqK60rWQ8mG+pb96oA9sClKDeIyyI
otr7cryG0Fo2EH+kh+kx0XTfMv8XaVSdaYHvmh8cLNxCLswQmAeLs8WajBurTkru
X8oPhdf/+/8JGXjY69q6ruiD84/RidGvhHVW96X/OtxKsED2VO8SQ+0TggT53bAb
bAxTjK3up0PHsJ2lRGez7fLXOrHvoGZTRHLCnok75DNeKTbJLNPOEXKjq/YcGBEk
RksEYRJBO6V+tseAcleZxlCefu1yUrwr9UJoOB0b0YTD9aZxDL8qqixpBzWlfu2X
Olrw1SainpnsVXmraTHCOZnh4iCFZTyAqb6fL13QGHO3YULGs9VYTACaFcLK7dzY
bRxZSaObSkNUpW6P+0sUtfNGC81IlSgP/86uLZGQ3sX7dxWcskvP6LGYE2jNG/YD
w/IspaQd1GxWYNEhcvbx1E4oazeR38hTOg7LOOKYgl5OORYdXd+CcqHuLZmml6Wi
ws1CQAHXp3YMByZHaZK3qZbgXfp84XJFmweYODacbOXWd+87FfDBF6aLxYWfzYuy
ts6jRWoT1BEVAKEbUKINvu7/khDd5bmFEqsQg6FePAR8+67ZG3UqjhwIUQ4TPpJN
ZqasEhNvz54rA1CCzPJhWGqWJf6L2AiU/494goc3OBC+JYYQ5SpRtfbfzpEvloov
ji9Q9ND6XL8CgDATFpGA0droRsB73Khlhh41IeQUyiBkrWtvYRTrVn9+49Uso/YD
byWedDb7UTDfQH5LSwQwO1/oQ/jA4RWmDTZocZt4kWrTzUkuSDHWvuLk2fHKd19h
YArM5U2uw8c3kjg3AMvVOB5CMxjn5gx5oWIClS91R+c6Irx3hKGUk3l9Bisaxee9
mI8vbmJx52vYrPMwymgM3lzSU9LYkmw8vimKwpLJ+1sm8cUpSn2kUBy4Zf5wQy7c
SOk/B1T66stGnj2eEWs6B7qRM0DaDQCHvlmvdSecUEM4IDigIUg5ABhk4AqZgQNC
ZXYvY33WXZfeQSBwUVW0SPNukDXhHe+KujxDnzgHQxOoOIcd7mklUMkcaJygo4bZ
VmLVGg277Jh3BYfgbSvpwGpnosWC37TVqprf1Upz5LrjCoDVg1Bze7WMnS5EkG41
yKYPFXLr3suvh+aZ8yU2U53oi8vMq7odVunzWg8j21bzD9hHC3xZKiR4agKuWsDu
ki2z/FGZCv/8Z03TqvXdu78WliWiVidhmoKxbkVvDca4nfHYGbKgCtwW4MrPW2h6
3aXgJme1CG6A/acWfymuDLeLHhKZZpSpsw1lWoUN/cFj9jiMQTxQytLlXKawFaXJ
5vCcLHJpRkV0KG5R1IAYb8Ygzl2QwlvUuUIBq/omAAB+qQfhbDMYGpQGlCAiIyay
aL1Yij9UBZ17IjhgpD98uzUiasSOxD1u4m0cUUjfbZwMIc35zjrLU4PodESbI2rq
HiQV0PWe7CiDTM8fAIZqZIt5HY/dJKCWia8KW6cuN5mUN2+ahqJRMrhzyRuaJqZa
`protect END_PROTECTED
