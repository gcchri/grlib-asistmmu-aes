`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N7uY+bBpb8JnOjE2zyFaGbdxjMe7j9Gq893JUa7QgPqdhnFfkkYCtq8j5KMvFECC
O+v2FFvftNkDL0Frle2A5GVFq8PfiiLi6bSMUoSrIpkuVCto5ZlIcIOwGkdbs4bc
ng940/rh2RszeL9Ohl46/+a8cmYYq8HEjNu6s7gheQcxK9YrKfZEojrldipqFMpJ
3kZsF247l9zUKZzdQeee7fzznZYcWi/JMZxWNoLWWZXcr7h10W3woVLCSNCoEzoB
94qM9ne8J9UBuG4jJEhUMc64uu4+8pAwtDHpjJz4a8hDt2swJeiuMWkA0O5J5+RJ
Y1VnOW3Ja33OwO2TQajtf4CfNzoC/sltpt3e5873lJzm8W/miMGlkZyaE54AhnsY
lwbW9hn6omNR+GsnApVOzV6YUm9s5L9qn7KNyFnpqemiwDi8nH5P8rT2y3wPMolr
tq1TY9hpE1UnINeGl/BKC6EfY/aGfXCICcPZ1W/ftXWVQcGNrZ9Dn4RY1vakyYL+
fuKU4shTyQYHw403DLF2wOfIPNM1gStjr1dNs/YkNwA=
`protect END_PROTECTED
