`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dClRfCysoD2xac1eCReStBMPWq2WjNmzd51xRDohe/C2aHjutkqEQQNeHyGm4nWz
Dc54Vx37eXOF00Xzhm2kWMjPL51EyQHLdQv/BDp9fsSn9cfdiKAec6kIfF46R1E6
56vlTO+JeYD2ftG9B+kmrcQdwZ0NyThtOatExZ4fYWrarPrtB1NtqbB7Pe/Pqqbq
rv1tasL/vgje+xB1ikqNaN0CdN1E493FWlVo8Lx69ImUMsNu+HbgwuFzJQP6wrHm
mWYo/ySM8BB47v1ygbHOFMyCrnZ1XcU+qxmmPF6/tLgnd0SOpdEIX2HKvmZBnh5V
C/slrCBrWLGZ9tuzwwhWWCgUJdda0/9/VHtGtRpyR0Ac7kuV7wEZHQeRZdl+qmgV
RwBxZLDalgPE4/RhCK4/hEOoNODgocdANVf5qFrYNsqV4z8iAPjYMKFp7Ji4voBu
KX0GFMK+QAqXXhUv3BL+4dYkafPeMbjgdsJO12sCBNuzcagCB0Kcio2BfRycpw5q
DHb6oa4XAMk/kRdgZ2UHdsu1j3VtxPQDcr17pA6OABllRXmnr5vaSZuHmCy6bKVr
eKl3wT+wSsZseKtkES7iD4LBUxAsR6TmHM14K4VwoAM=
`protect END_PROTECTED
