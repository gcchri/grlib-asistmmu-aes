`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
czAbyxZb7cO2SrMRmVvZjWjAvtjtrlpK7OMBVcd+m5RhqFCTZOJpqtxNONjayHqy
FwEbA0ywzA4FmCHZ8TXDAr6z0Q88HOVuuNb5xBuuQNhgNRdLhnPeCH0VI709MBjU
X/rjFEZqyo3E4XFfBm8jZooBOvs7iG7kA2e7ICx5fg4C8HikHfVpEaJGdGsI/Ke6
ut/plN1BF3tO1Mrwk38kDxWdS7Wg2Ud324NQcHtWGMIMt5YThuF0hINPRykvAncQ
lupLntRyTELiAC0XgZCstTvWaDpXUx6J8RArjFvusEPfV32w2ZK3gNg6tvDYpiZy
rPd3S7gktmbWTAdDrVQoEVsUFR1b4Pi627aQZ6fccFOUTXQNXtBwIML8CxmTcroD
1YrDYW2trmFDyepuelQCEHqvtVV5avNZVQYShTwMANsaaEGqZQ2D5O4pstH12lBL
nsBNZ9NSFyCIbU1m1aeimqGRD6V9edg9aGVU6Q78FHGvUi1tDNK3zLMCNRx3tr/Y
`protect END_PROTECTED
