`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g6AdiqnrB+uYPRgfRkoUjbvClMpCB9u0tLz+o1aZmBUtOQyWsXbspCa4IYClMlfB
lg5kh+zTu1IRUvBgAU1+9LF2zyXziJEcpDDHEJWeDGFJw2sMC3V4fBrFfjjm1vCK
mXzOwXwIaiAnScZA3MoYVZfu3dO8Kmr+pB+LfXolLMBNdv3EztNdqUwc1MaIylrR
1FGvaYX1Uny/1a1SsQ00RtBOUlDfh2rdJngKGosL8NIKgvxuiIJ5nJt3/s+dwovi
V9BrwS/EET3XlKuMEhWrcv4DEDwiL+R/tT7O8bC8Fus35Nk5zrYFXs9r8SKwx24p
tmira5YdBpf45OiawAD7bwSNwIR5/nLCicAVlOHs0xq2Hnl/5HYbjkEVNq1L1cKs
lkOiNtDnaRdLYaMts0SHJsAIdBAqfst94O6RiA9EW38=
`protect END_PROTECTED
