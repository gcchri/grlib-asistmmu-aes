`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
in7a6ul6jZZhIZ6w7zLt3Xw4XFEVsows6Qe3NUWGSwRUZAbKPnjAK8yEpSx6gCKM
KZozCji3R6Aw14FOFB68qjTDux+KyJDdfQk15CZPfijH+eUSBL5L07f5qEkFZEYL
/B3Mh5rGlIUszuEsOOheYTry6kMqqLjDx4izeCoWIzn78GdQnH5eOiKFu+FtsNsi
XGAlfrqjtnmmkjhK39312GrMx22XhfbQ/dORK03KE2VKhnhjJBbew4gAgOe4v3xp
7CVXVWmgeaF7Y3hXMaFlgSn4Iy+8glbSUoTGFRxzybOIa+LaNauxEwbmPQHTZupS
/D8a/jq+XMas/iuLgebwugzMbghmL0WnvAAXsYYOWJjHmTBNdwkc/g1kF1JXWA0l
UFv9Jc0+CzXbCiTgpMqGFumoFqVQypXger7OqBM5Vw9IVvy2gDCB24yJJ5Zk5zzI
RVBsLOFVjHgHlj7I0z3z2/nvEIPOFU61EP6yP0U+9PvgVMnzHUKcsjDDv+DeC6Uk
YNaf+xGEjZuBOhkTNIUjYHBa4lHIOlGcNysEEeAmwILYTIsvVJ3NzUh3C1fnxakc
E4iarY0DyTO8CLh/mIYL9+k+Rr6PC1PS5/mRnk9SK8jH+ZMO6ieWVF2pas0h6cCd
1nFgJw09gfUSUCL/smN+5OXUH5ik/y/sxkk41rZg/+LHNUjQtV1L6FrxWuQvDG7k
RNlIiV94oiSArTfGI85+TGW/JFS2zXBScU3CSS9Wm/vbWItWKCiH5yYf6DB1frXz
0d+UdUvzUfMeDH+7qUtrbfR3LIeaIwYOKkA3b7hHvozbpVmCZu2rkuTd2ppchzzP
OAygKTRxRxu3fsf4Rom85Q37RLB1qU41Itf0TnhkJuIaBGdSsxt8o1qpZbXHFxaL
8mQWR4gH9Wmc3vtvikLNL0rEqZcywIUSsh0LsUP8PgIUsf7xqaaCJ6s1Czo83yJl
V86vRDdDAptjqL3nyFQNLJQTA7icmu5R6awSMJRdBADK4ARxUVaB+GCmWIKw98zA
NSXgrxvBKvaU+RjxMuf+yEGKKrNELLkfKbEw/kxFnQqTOJ0qh6w4guMl2i6UJoBI
bixUl+GGoR5bq2Kbbn9doSqXPcXTUZtTQYUsTbPhBt9JXK6BBb/pLgaVNb+WAn1h
Tx0Hou3fvM+pzvADcZcN8Aarg6xDyx5vhJxUTesQ0jH0pY6H46ke67HG6FN6UbIF
OUgTydj5v0vQ9Hhg7ois5qE+U1tx3pw56u8dlGAPIePH+xXVVEKvAEVsql4SPofi
07i2d7vASN+L6+09LwYLq6blLTz081+L2SjW3Uo5WRPLqjz4u0JQQfH+v5QTQbCo
lsYt35ou34VPcCjQeq2wsGVmT3C76fVDWS8QudC1xcebsl9UxC9gI3SH2wVC2X1+
avnSXnfs/go1Hcs/gHxi6CO/sXVNwdl3de+0ppMFuyz/SkSjWtmiM8uRSoL6HOWq
ufqAY16z31QEe4mZoWbL6vq+zEHAg1q2x+NQ8J7pe8f4jpIfS3f3DOcWGGN3hn8E
ZuEL9ZVO0W12xSttZEJLa/KkdxuTx0qL4/UI/sBuX/qMh+RMr3YHFNizjLtWnZTx
vEUW0NPabTVzwf7Go2B/bNotHR4WyqxMtAjtmEsEnFh9abyV/IhGJYXzDtuKebx0
gtUtO+ixiaCSAcYn/SV7fAbvf2REaNnYgqunAWRW+vsI7rN85kktVwpjXw9Q1yW0
`protect END_PROTECTED
