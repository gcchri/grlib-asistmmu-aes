`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lm66a4QRH8eTYsKPUn9wPpvIzRb2zPfk+2T7AOdP1oKGJZe7JHOPifS2MOW0W4JL
rpjrZgAORQqVfVCCr7SUVYgUPrZqYSuJRxOtz0oDTGwcmgNkSUn1es9lTn1MLGcQ
5/2WPfZDkA0A5cqZD64UxJJCEs34PdsXIZPSWhPftuVUYUKuIc+bHlvrv01YKvoR
ekQ8Vg4zsNrMf0oIfKl4xOw1wKv9EoMYSnWFyPV7xfuDYhJA05vCKIFla5nqsFPx
NDgFatq/7XxOLqy2IEdjDthRjhgxnejWhTBcZgZJxpz2LOZDM6XXOQitNfM+Ehxu
uruahgqgRaMqw9RaxatA9j6Zv1pMRa4IqscRN/a3YOplHHJxbBBUPn9AbIjv23dS
rB5F1EWLhGNtbmJ1ge98ufOpkB2LAtxSe1bGgNj8U8s/gsUnf58BRFqMAQZDCPnE
1zsk/xa6YDDZJxPThptuTa9dkJJ3FySXC8PY2cM7fzrVpvGXVp3WN5KH6OEC+GdE
FYv1sNYmMS3/glY96/0nk0vZIm51paa7tB8h+fpJj4CdlzfMLwBMyZncOcpV9WA9
zc/dc5Z7t/IG39xAiTL5xFaeDUeJFnmd2/tH8bJ/IqdQN5Kn2L5UpeK8P1t3BQeg
7GuFhQnLipcDQXE/NULUnsX+C4wv3enaxzbryHF9MKLqqlw9AxJMoIB4TMhyi+or
Jr5NvzduAyiB8IsCBnjDxXRiWihqMP20kox5XcVJ5WwpBlbse2gAX3ZK+ISi828H
Ilwjfg2p8W8dFJ2UeQBq3AgW/luEagD1dqAXxArS+/iaarX9Z/HUIFXX8edwqRbM
+hnY8UHQynui/zk2n2JirOrHLT5cFFsQeDWctf+8uctRrZQUIjF2hl43Uey8UQWZ
u8IrN/Wb1Bh8RMh6CriMH1nnzhGwrC0Mq/jwtnBt+Dd0gqvm/c6hVVqf6JRavpTH
q9Gk5PmuEHHiMsNfDbOIfKLq9y+ZOxm5rNtmjj1ZElAk3kAPzQhW6ySO6kbz8DYh
DyeL7afd6600mS5RU8Zuj0pDOaJJgqlEfV1MO1Q3ZH8X75EjGHtYFtoaYJUet45O
jmwIqQW36+l4vMQOfHstqBhoaoCm8ZgMy/Ul1zo4X1tHRCMtQBYPYpt5pCethOm3
`protect END_PROTECTED
