`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ICZ7jozgbNk7t1zDML5zrKrXMSFRLS3I0uy05b/IhxgWPSB22nWELcsh70PxTAMx
T7PhTY1bOVFkY0IY717grK0y/3mN/0DHZSY5e7dUGcgvxFNGyumE7IGc2DDs+1ct
C1BU9HLhIhwnJ0vyTIE1vcWUR+bqAbTFGvWGwltJCPYLx8ZaIgMjcJEE1SkSUBfh
1r9TMxdHKLWmc9EjOBLruNbVSZNi+juzPbicwJ0pJt2JbS41+03Dlxfit0AnWdmC
yuZr34Xm/6E89YlAo5uIn2CQcAS/zZcloSt6oZsyj/6v/CfDENdXpffoWwtgAh0u
pcVEdAydYBUv7LSL+0A/sgNCMpHHB2zSO2UOHabfYS2mR6ja/4mFgxVc9H0gQWz2
z4K+eCGSei0bSaMb5KNcu8iBbUAhTGx2lAGHQuVJpa2OglnUKbhNv5fPTXdY4MrB
`protect END_PROTECTED
