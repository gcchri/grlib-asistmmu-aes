`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YfPd9jxpawwpkFP/Tcv9tTWgox42SWllOAsf3USUlYlZURJZJe32eVmFaQl7BLtl
jJ+qAoQLGvXkmNX9Lqy7ft5xBXKzzn4lkqkPi35l9tr3FH2QpOqSC+kuZURegL1T
1oP9A+YkvBllS4NFJAFMb+CZlAIVlwx8THA/X1j9MA2qDfU0wWUSxcLnUpGoLYiw
flynr3eRjqry8aidXqlN6GfLm0XM3/LwhnlBCcefmfYWvg98/dfEVfx4bGxsaYq0
gWE+pi85O4lVs8G852ejY4/6BmbWNhWFQsEPHgUXW2aM9WCN4j1APBirRN88toi3
KDpRjSjC+rpW/F/HWRAjxG1gS49A22MyvMdIt+ByncvlEfFevNHbKKgXZ+pZJ+n3
6vKHbsXLi1TacYLDhw160ecAcFqlFKJXrF9lzLgq47OOR64W8OcCXJI1uT+dfINl
LVhrpYiWQ+u4SOdp+wq2sf3FzWBCmuyv2JXLtLJtOtjQm7023iJa4xROpIzWCX2T
HlS3rGqgjnMCzCFmqHShV/Zp9TKUU6pVCxxGZYKf1p4I0VbuHMMrZXFFJc5rAB8J
JFVZ9NXF8QLq14Q+8ADQ8E0DuHz8+c0/4/i2+8AiTz/8fnElSBrXvIqAIB1I6WO3
9bkldUXMOItB6QQFzy7mHe0BYaQKeK/PXN5PxBOOj9nWDaiuhSjmvv5S1wiOhCtZ
kad566KusS5fupXBWAhhbep+9R35nruj9RK752rbqgZKZyXWRCD2GMJOUVrs39bT
M+SaOpZqj5OlxYuI9OCEg6o8CDrn1QCdtgAtrlR0zADlx16KuL7qf/ZJuitU9fu5
xtb8phFlbBas9Al1Y8Y9Fg==
`protect END_PROTECTED
