`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VOTo/t/FqJmJQf7BbbOWlcWKtrdX/sT57Nt3RO0R/Fq1An0mosAZGXE89xltPxQz
7lWrCqeLnA+AVJL2iDFV1vg3FYvjqHD5CgDGZekt2GVoyhXvxvtfZmY5jriKb3Z3
1e7YhmcwfPh4rbsFU31KYxBKYPpzYTzJ24O6jcWbCDJqrAZY2+DP6PTjfTbjEQ/I
J0kHMZn8BTMIoqfwbM57qdO3Zhf3/Ai5/aWG+1RJZKeKN/jJpIfd/bWZfAkhMblG
iUVQ9bhNi3sXhR+4M1pMnOYFh1NXqF8S9zL7rtcpMA8uxtpG6GY1eCOoIhSxYtcZ
i2oFijbNbbnw6TnRrNkVY7vxsRL8HSebr9x82ezr5v1sya6+tJ0aZUL1SyjJ7xT7
arnyguobi20wbCIEVze3CuI6WKfdFhwyYevuRW2ss482rG4k7/slH9pj1hDY1HLm
h7tCIuR4JSOsaPbdJkZFs7UtRW8Q9GdPUDholn8kDAtDZIn2seQ/C8bWwzmmkCTY
pst6LhqGzDC5tGl6ApgZfbZSTYIVXhpKoxdBnNS/rfTxUfXA3+SKzBurb3PZnWEI
HPCeSES8mV78pQO6zFGLGf2Vq+8NjkYd3S0os1/hMdlDfcq7mtiaAeAY1NHSUzFd
LEFXoVBenF6Mkqzu/AQ3Y+Tqbjo5UG8zq1o3wbeOrSghsGLP8rsSBiSognXwQiXX
g3EUGT6Vf7oMD5GMzJzrnsFgI/LgCA+cx9GfP4Huqdn/7jfnzyg9G8U7XawnCwXk
Fqk53UY66k/nncgA5JaX15v7poiQq0XraZQVs3Do8bouceqBZUCW3BmKKSRmIYSR
ZeG5co3tDR6gfo+Olv7AwJraoVlkf25ii8dyFZFWINBX9Lc/RwR0rtZnezlmAYqk
062L31gVwmxcUH2eO2jGdaj1S7S+qTImIHnCxINPuZvHHE3Dtne8m74I8UpRDKwn
C4Yizv50WLux2R5CDq25KUYfg0WIKKIfbDGQtXxRM7I7COmbokzR7yUnavfirJkT
gSIrudYZpKbm/jozn/FO2nKUNRaPrQH8vNBI/eglfy3Dypln9H/ETv9/IkmWw0Xp
9khHeB2c0d6kA+JirLtw0v5sMe/y0avp11lJX+DZXdav9fKA5gT9YOl9Pw20E8Tj
`protect END_PROTECTED
