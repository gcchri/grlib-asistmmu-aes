`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K/T80omDhN+IvT072RB+cQuo+hrqOW8vN+dhInvz8TReVBj+9pB/BANRhg9Iuf4p
AqK+ApliGY+PVPw1sYJLWFWvJXQFtETsr+9xADtZ3baB4M9Nly4dVs6fTInaLt1y
nLL3hnEw8p9Lem/3OidLCPQmlXhrg/2tErXMJaTizRWMLPqB/BOBRR0w48RUvgK+
q1pOQXdvmylr57lNpMGQvnAex9tl9+9gmr1gR28spQM1EBeImBIZIJDqgRP8h1Rq
Ss8DDv/Mq45QETZNcvXCLZzP1SHIXKBYAahIaSXej1Z2o+IxYDeMN3RHmShW2W9q
41lzChLsafmL4msR7UGZCaTLpVWem6nGIf4hnC169G8BbTQ/n5BbSulaWzvGed3Y
Wb9ckp7xg3T7bkK+X3U99qOs8e7s7y2XtI2mo1DTwpQlnUpQkS/NE45K75qcriOp
2tmgM6BuxD8czC7hB8Vyqse71plwplcJ55dR96Hca7SCrOSAR6UKodGk6S3negY/
+ENdAYytNEUwjPcaXHlXUBXIHXF8oaD0JyFHWF8SKfuylsX1mzIC5eRrG5LVuB2g
nI1KX73X+43M7oRnOyaRm5R+h8hBXgd0UTJODGvLiTiKKx2euOY8h4N/59zzkIOQ
jKgDCHUIjL+tkWTD1uNd8w==
`protect END_PROTECTED
