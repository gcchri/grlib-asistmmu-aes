`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jVyI3Xa9MRU02Yb8LKijE4ATXj3Y8CXBdcsZvkVBuLU5PPHOcNSygNGumjclOE8X
40qt1UR56rUMUkPPPl+7yF9xDarpDpEix+fllMkFsYnj/I0PCeKZG+Vn2ApCP4V0
BM8534mx400GtNXVCOSwccOt2vEIZNQy87txTvHqvt11X23tvfWuXLeRL8qnSNjI
WXDGY+Yyg/5DBG40l/TaQ3t7uIg4DjwfpX+lPMK6rMT7PYpNXYNo8BmT0BgYsyqb
wb3DyuKaE6p4YiaKb9AhR3uv8sjRZqGBPro8LrN4TsZXCZGxTBC3DLVwtam9e7Fv
QJZ9Ghkw85jgv00rqxwxoYPq86rY2tb8pkUCim7F0wLiNqwKjnd21YFhLZbTTU1N
JU9eEOC3wbV9ICfbQhAzLEIU2weFaY/0sue2ulj9pMqs1LjzVqVnigFrXcBO0fgv
Ja/cDtWxIzdnJj96zRcfuuv+7JylvRjVzCoi1e3H1pyxscDPE+nN/SF6+szPRkL9
rkhq9zr3HLzcr4nXyJNPSFAPZai2V9b74FcVkKV+PPXHU1KaWfP14PyDqUAQB3R+
qW7nI6fydf/mQhv2X07xC35GrlW88yAM4Qip3e8Iq2oF/BiZ6TGQM2JI3ubMUmpL
G4kIYuS6/Km37Snig6gHWti45nbDdBGrJtqzagXBw/YUJT/r1EVSHAwGN/ZVTWFP
zJ/aUdenF5HKncHbc3OHepRehEZgo1xDRoHVHH4sIS+njb8firqLgjDT3ICGNo3P
8PhCWLvZ4pVSNN8iCbiDpXSW1tuQxlcGH41HBGyyuHzcz2uTdKlyFsmDuqB/1V6E
Q1F7F46NBdVLq8co2pvZ+jk4gFChlDOe7A3tWYGy2K75ZPMfzbdAVkKfiPsZ2zKF
87Ff/HDNql7k9hlNK01U89wGas0WLtfbsdQOjmTlemYXZdncq6gxWOT1VVqsL7kD
/dJ5ofrN5IvLmmkpYsnvL5syBjJtM3oxZX4RF6+NylkzxE+7YHmL9JK8gxpno2kb
k5GuWIFIqwmf2BMw3HlxXA==
`protect END_PROTECTED
