`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s69WOMORvTlUcRKKeP4EVTJw8YnzETiOd9vb0w3QUbGrwnyHwNvvmzxq3qKqwm8O
IdZo4qBZohC1Sk3IfZnH9S8+OA8ysmA0Z9x4uHnJwMOoyI9GFEESBLEvssSTHCgl
S1ak+XkW1mU6y5qF8BBcH2p+IpLzdSkY4t0PB7blFtbWf7QY6/UW4mbAPoo6fgq/
SFHPcSrl3TY4RacjKU4PgdL9p7jc/Psahf3FUb/ZtUw2h4oRbiJ/bUjA6aT2fSY0
wJB59SyoauXtELK0s/Ct3GUHXPcIUe9toiJDHGS5S27dpji1vAeT+8CEcdZ4XfN9
enkLlddvhvIGzU13ZDc7TxVu15TUUWzOEGki46vWL5/DqS5mu7UeWwCQTFffkpWh
ZD1JSiXPqxAkXUhlH2Bo3DPGcsGULS22WG2c4n0EZUwRXe7/fXhOxnljb+CtTvoE
G59KE6knA9foN5jslOM6D5rZQfJIFkCuk+DZ+IIsDUf4WfVTEGRtaetGzyqRxovz
ZEWCMbfaHb3OJV84KfyPu4lh2WcJXZsg92I84vsdH5vD6whHa5t60m2X/Mb4EXo4
BY7U7wE2o96QX4OJ5BSnkDf5zfbEMnVrw73J2zhOm3/wKhgPdtCML0HkHQ5ILzN8
cdD29muRzPWnnq8XAwb8O9atFnHw69CTz9qsFPCGcW/FX9tWtA4/CqQdO46mKzeD
rkYJlT0mq/f8LCbADGJF8QfFxtZ0W7JOzzqeTVnFZ4qR88E2fmUpOsr1qHMYYaHe
QEgEoMagKkND224iwmrN00X09EIIP0aEf8DYveHIrNywO/NAjep6Uj0S/23n6uS1
beruzUXYGLyqprJKhcCWgyiVwi6s1i/w6ECx04RGiTFqQjPjHChKznftYrR2iQ/v
FKpl1+Tk73h0u5GVdCdTFh+lrYhXvCr4yEPZAYaN1ScsczhplsnnINkJqQ57pZco
i/Mu6EVgO1p+tCNKdqQflLGOmstTgTBeNR3xqvS0rx97UNOD0lm1eplVfFHVsApq
seZKVgkNPbKqrIAwTxwl7brg97T2mYOtU1iFRMMSNwK6lI9fnrw2Qp+d5q5+kMeI
Oua7ulQZInR4uRw+D4sHUZjszd745O1DK/PRM8sDiF/oUkFbdDjYmBSTXCdecHFD
v55EMv0os+dBDM3/9FWpwcLyj5xvKz7FPYpAAenjs/ljxd5nUuwBXbswJPS5eXDv
/qUxxXHZeSGrYCOSIOlw1jAvVIDIaucV4NGm4AcX7B+dPdbtG/So4LH0ldtnfg3k
0mWfcvuf/cYAEqneBqvTd6PuEfYnRs5niwomKe8ySOUtI56E0zAgS96C3r4ad8Ar
5u3y4pCf1mzfRkNCz+atO7cK/loG7nD+th+3sIzuf8y8B6FPaNsDwWDrJavTNt2n
dxK1dr0crcuZJ+4m7uWk5d/R9mk8hANwRPvhNSHFjNNVduemwhpyidT45FJDcPv7
XdcHLHI5PAC+Al0gb5l9gjjPNqVFUr75a8flvmdsZlaSu8fzVu6BJijTDp5PR9q9
va/VCrx9yTSHJKeBVSyBcB6qF514/5/nBzWV6nZvoGzVnRdwIwPYLzXXRaUMxnD9
5Fl1Y2rKVf/9LS3aHsepE8uZehKsaq73NwfvpCByI13UBmxIcms2R5/QQTOt3uhv
g4D9B7WqXABXR8JaKWySfDyJqSGnqRgBXE3pKv3VmJI=
`protect END_PROTECTED
