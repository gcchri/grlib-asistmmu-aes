`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
upiZ4ybQYdwJXKNTKKBxndwTzQm1qArT1kFcBrp1m07ScmaGmgp89qUbeNxUG1DH
0oedTKRan3oFVoXrQhVkLonPgzYZg0Umyg/BBspPYdL+DMyWrBP8YcDnG1RitBN4
ItXxVteqVEt0elfLIKlCCtyE+SbEGpu7V0QLaSoUXDLF7AtUAx2f1YAaEVNsf2wP
XXVBArJeg5J3cvqei21YrYRovODl0slIubv3K8gBt7b/2m4/Z7R/RHqNyyeCAN6X
nxr/y0ygPaSnbvGcavcOTgSHNKbZBr9ecombYAGFB2RZuDxYulyFAFpuETcweWqk
DqeuI7Vi2tdPcxawBgJbnpQiaf6GAwxBfy+YVtBmokRpHbUdBDvn0seRIqvF1pIY
Sw/yQQzropjfB6BYdrS/zQllfQQub/kQhOAzCR272mEBfd17eLdb+bxQ8kSkw2wj
EQomixkte9DXja0H4u4gokLFfDRlJfjGHzGbPIoTi94g3XUJPxNRrvHpDQ9H+8Pw
6/gD6IZJtNMEbsa8NSBa0EwbHA+YakmQdyhyAgCYqzv4Q7m4qjT0wHIAbdTBmjcT
ujoEfMGHwFNDJuFB3PhU26/z6uxpI3wkdr48u13Ra1vrXUjni5RCkK7HMqkNtjY7
wNftDztfxZGxV+B2r4IilxWGcGcyMTuYUQBYGwjWe05LB5TY0EH89Ycdt/b4xpdt
fsSMTVr3rOaw4DKBO31fGCcfyyoTDZf9QWUcJ1DSA1rWtWnw8DOBSlxydAJJu/L9
kj29jH5Knpgu46bIwL3DgOUUeVpfUa/PwU4cqrcZ4lqSJl8wbfgwYgNN22ICw6CF
7f6zF85lmrYsM1uUMCZJAEMnJDKRsicxkPJzXGwBkNU=
`protect END_PROTECTED
