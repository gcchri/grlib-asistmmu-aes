`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K0kbeXgD2M9V4slkVTxwhGgTEW/2h2fjMBwAp3dMYAf24K0EWgKZbpsbqX1W4Lj4
fWikaWAnk0NXpyf6CF6qqfu7Ax+Jql9Zu/IMmg9XoYGbW5DnzRmd7gzkvqzeBkPv
mcKHRwLVhFimc1c/Tj0rWy3j8F3xIhAUAPn6W558UPW8KZrDD7ZF+U9ElBcCK/9q
DzlbqkjThN118/790VT8ECMAaK+6El5k7zlGbrITImoVfgUkDaeR3aehW9pkIXcD
gu6+UVpjHh9iTqjiuOBTEgqCWUvjEs6uE+dSHz4M/knAwMryUhKFzX/xLoXxtghc
ToqHknsHdM0ne40a3o+OicKywO7IZvYlw82PZ7cpa/McopZqFL8Toh+dETfLJ8+y
cNvXICm+T9VvXTtjLZ/NFan2BhhnwvW/+lZNS4+m0F/DoASn//SxVAZzFFuqlJNc
5Uwway8hvQhaB4LNrSqTYVknO0Wtu93lYVCoL0mRBm9NWCU4MJDrUkBMa4R1aj2o
AqVPuoigDCsEWdp9DJ2O2f5rqAAVMGv1HkI+n3sBk3YGbZA0tgnxq4+y49X2oxGh
T9P717WRGJjEhuxUN07Bp+obG8HYhuazSE31lyalt65B8+V7fqzeMHw/jJmTPDWg
6m0K2Nq90HpTBxCqMFOWbmJTqc+GGzLK4+2z7vUCQymP9GBykG42zOvTD9nd5AOz
m2MZJFvDxYOlRIqVFhOPJVefYne5QS86bJseMyE69qYnVQzLLw3Q13WVXiHtH4Af
rWDwfc6qalDAWScUOGBcAXC6WTA/BShzkogXF2VNZgPKDDwek/NKgkNInnJY1Iz9
PPgu/kyymoISeN/MDhy2Eq6DEmmJi5gtstldWOtA04ILfgDr17M5LuyChVAN3ouo
ZoAxurAVYiSsvzJT161jZ/3FZg/TkkVUw7ftTbdvy5MrSndFfSxoSQPkDHjzC2LU
+HKN+og2z+e/dHkHsjYYGedPWvx/PMU4Wl8vHuuqrezmtqMdt7+SS6Cozo7fV8Eb
jBxIBRSAQVcKz2l2MZpGRzhAqLahhjx1+zaIY69k/cmHhDvYsQdn79pSQrRjnL2R
BhS+NAAWBmYz4KDPUzZiWJdMlq6zScpj5OXjDtqgnn4xi9dQS111zj1Mcc52kXp2
+eYibGDd9QURZIpu7g/WToqtqJmE14Pq5hwIUrlIanZL673GfH3RBZkcab1ZxvKl
SQSuI/J9gm5SijzXi3f5FNXLNdV5JGZuRNCZvLyRSzpqlFkqFJXV+m/A1sKlsroW
bzJ3739oZsCcyPpjwaNx/OqUoZ3DRtoL7FQBoBNbUAfajTooSQnNOo4PPKXv1JKL
dr5/8IlvFj5+F/os5VFKkvIQqusJEzucsjBqS5VOtORVMbl1DEpydbkawsu4VUi3
+m5L3c16xg/OY84gLsbE/5GA+tsFUgHetY7sa+eSl7gWfIa3vFDoSGuOCs/YGsz9
MQHUxGXcZ+/8PyoNQ+pwug==
`protect END_PROTECTED
