`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D+Ph6SklG28nls9zWvH3+IhS9HulFJGlaQWqOLGu1Co3D4k4fiMvmya+11WGBeu+
0or1Vj/z81o9JdkA1IsXNWfPMfid5NvSpfrE/9A/1CStAK0jVon/10Kz9h47fdt8
8GQ+z5pkPjbeHYjTgTPbWeoStzRyRTsM9+tdVWbGNke7R4Iz8YrwYVUrbecchMTy
rtdESKFm7cfvF3XgbytI+gMpbmICYhcwzqXzYQiD8Vrqdg+GL2splUPcSf/b3Dt2
jeR8oFh7JEDJTvBDycEqCSA4RNGL/YZIOlXw8maoI6rpt25nX+rHWnp7WrVM2zEM
rk+3ylmpPw7N6l3FICyFvD4CY0jy2DSmUD3v5HmD/aY9OiU9ZB8g094HmmXs44+g
aKMCBpw6NlrUddUXmS7NWe59XP/oZ16o5MrMxYDCSHFAsrg+TTDEkYskZRHmL+OG
ktitsj0OnqkSdyoZp3P4mbNHKsGV+DKxurkUjnuCopMmPVghYWpEvvfyZ9/YHsE2
`protect END_PROTECTED
