`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ztsE/T1jNPewxAwz4rXnFmsSUEbtQYlhJxkHyk8MqSXDMBcYpT973xebtHvp48A
xIKlFcvTBDjAGXB1Nt4Uhlv0hKBf0+nwkg0O0cm5QevYwJxBnUOR6NDKLaNFPtle
8f1PDQrnIGDxW1z6f6LN0TaVm1ZywBdoprKiUySBCD7OlEebjq6rlzSiIv2F+39A
2byAC7lOD5liPNTGcwPc8B7HwrUcch84cQ+rDWrn+D8UjoUciljqVUwZyNgHTGVT
3GxFSniNKmksjBebdXF3Y5Ou+6a4qtkF8XHI468oxGoy8rIipEzgYb9XZTI0ibi+
l92PhzqDVfl6P17fR9Ci8o4NgzukQUTc1OsfJSTAW/olhHgkVLwM5YhQEPwAA85I
m5N0Xj/a6pOcVJWbhqqoUjFIb/z+LXyp+W5B7xVQPUmrC82mn10auivjy7BFHZmi
xj3WGwWvE9npYFbcxssm8lfm5eVpxiz7YMGfFmxt8aiaBZixo7CHQD0z1W6jncRG
BMjYRhxGKTHQkYxG71L1YSDolXH+Moo+vqk+9QdbuSStiWAmIOJFMXeIbQPv5Sr6
`protect END_PROTECTED
