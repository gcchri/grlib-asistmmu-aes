`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rFlcGaB7Wmg/6dTJKL1rt0IsID7lStgwEpLEW08sYELf5MmkIRHh17mUTUxlqUun
t0jel1zqVeepJfS0wfhaPWdBSadU4qn5sJL38snZC5MMTzu2eM7iTitTvQyS5dMS
uAcNymQPz+OUnoqbyRTLvCM3V54lpA04hyPpK9ZKK/tDlokxueYJFF9zQl4gtTI1
187CQSJtzorEGumYpbytPQTaNR+d/A3UWWkJtKzPjv2mQ23BiylSqySaorz4gMhQ
4/aiH/24khgECGCo1rXJM/3X7esvGYtU42SDpQSfrnRj5pW9lYl441MpDnOLdcjM
UYsIGkXK19b2DqmhdD/hkQ==
`protect END_PROTECTED
