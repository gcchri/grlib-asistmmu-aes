`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ocJl9qrVONl5oeV3SQdLg+iamS0lfN8yCM1UM1oMTu1FW81HPXxc7CJ/n8O6t42
Lkb+1uLPvjVTiT2NDSe/PXtS1YAuZn6UQce45yvLd3dDgD6KHSNEm/8S1E1fC530
QKPtISFca3rRwROdd0ExoCTkKtoSjRyrOBnG+t+SLxcWtxNonTr0TJK1Ojei6lQZ
a4hSB3Vbdnz8KXXqMX5RYCMVZ13JaK7WyQhHUmcZObBBWIRtwOTHyrBcU49WRxgl
uGT/KxC3ms9wxErC92EHl1XU86N18CvYchS7YATSXl84TtWPmzR7g86VnPAowTmw
tS8c8WTgA9psNqqo9SmVi8i5Q/zi+qzRasefOj2a4dIIARnNRzxaWg6RY2zHp4Us
q1q//n75GBHU3xAGTUczTwIBVPpB5XbiqH18JrZdLEvuTmenSAy8n4ov93rOfJHK
qeyHuF+OMNrQ71vYMxVyKEtXrjgX0Idfm9spG/SOghgWHwa9VcbUyjJHNhXwhb34
`protect END_PROTECTED
