`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MuRtVn8boiFbNdz2AZCylFhl0Zd/4OZ8JCl8xLrd8TGkh3M+48S5RedVr+F5jv5W
8McU7gdoAQR3w/S6ftt5hKpamWLA2UjJtuxxL1ocFQlDN0J+sSvlSjDQBPPHlpsp
fbkpPKCu4FUfF3QIBh3WzfWafbPQVy4G1XBrptbUsHFUdRf6yGBiio1g5LeY2T5/
lA4fiA/BHpbIBHK02SVKvsza+v7PFosXJ8tSBJBnnWTqwZS3/MttcFLJnUSePep6
nFyeoa9Rm1mIfqQf9nnO2fSfgAEjCY0w72KzZGBBjxC7St/+5j7pEyFZlenDTkd+
mT+T8KBs7vlpuPJMV2Fq7l6WsV4OaddXddhQZtbyOndG+aqVh4+yGH6U+GPvr2pE
XEMOszWCxhqOIUMXQe1Oc/QPgkLjUp13vP4wMEEaQYH3auI8J8Ez/WTRhMf89Evh
clhuPnh+SiFkX8s+fdlp6DGjoGIBzJGuFMHaN+erhldrXuqSnfpAnYrBSu/2y+YP
DpYpinmosRno2RfG1FsdyrKFTiGrSZWUDg5Ny9hScLnY9d8wuSvWklZR+ZtPk/Cw
3CJz62autZ3z8pNwNfNe2yb0/8i+6hVSuucBpDU1+CD+Bll6q6TidnAse8fybspR
4KSoaxIEdRaWEpvv4LApiw==
`protect END_PROTECTED
