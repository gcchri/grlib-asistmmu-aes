`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L/0lgBLIBkZpn+E39z7bAapaAVMPc3gsucm71SOgcVXz+Zb+0IoShPzbYoxXrqdt
MRdkg/uiAOSn64y9JnR9dJSQLTR/22O+sk6EZCRV+fHC80CBUZ3880CKyGAzbS5d
CSWNvCkPLvSIIQRfhXwv60kCRZ5j7mRDhn09FeV//EAygHrXhl4WZC3X79/aQNQw
2YjSYfV7G+szO3NZw2c859N4ojRqDRtK/7pycQZtDgY7MZ7XiuyunXAhpOJLhqdY
FV4Gfvi2RJi0xO/VrOGxCijf6r513T/SYU3hehAFFcxtTdEGmZt5+W6ZC8XYiG2E
Sdk0j2SXmOarkkLPvilnhw==
`protect END_PROTECTED
