`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eh0eKH6T1BC7CMgSu6h2sxDAxpmQadQqpmmcMB3hGyS0NxE0JwLCCUCT3TcEI3lP
HJHY8TvycRIitaghQ58gKIOROKRK5Fs8R5Wzgabw1wfdt8KyWySu2CybwSJhiNeo
QtAAchnTdyztUH0fLuxBv8/p6TCEnAtI6e0Gsj27TmZmf7+T1ED6+DdtUpDGPcSj
owofw+Eto47qUU/vRGC2ZwiShvvutXxte4Y68rX28U2mB1Nw0iy29szC1y4qr2Tv
0XI7RgYJ2SM2T6fq3c/nss7sdP00AN/15XvvUpjKTuV3aqHvv/ZCFoTYzx3N4f+U
riuWg17w9psMfSfWlri4o8yA7f1BMCZxC5dglmTJWviQgxaTLlRIaz9aopz9obWl
kWcph6wR1AU3Sx6yzIiphjMIyioIKhO+lMTHzRF2DqqSJn5lw+loGbG6n4+NUVXa
ubR2fPLQ8x/ZxgnZ3/2LbW5b+nSkJoBNiAvBHcB75tvoeyy2WzOJJgpxOgY0lDtM
/INIHhSHB5SCzXwp3BAU5P4gwAzikZduTHmqyMahTg8Jlge3KJcYP+agG5CJT96e
07RGEBSMXaHCX1oJ8r0rf+AkjrrSCKCbfmDxZJI1GAvvyfNgUnhRaAaEzKo3kolD
kUjMFlVomh3WbPPXcVPUemG/wWV1eReQdx4lRgzIaM8dFGdfkzo70ixZrw1FhLaA
NjmFkBzYGPLPq5PxBEzpO7V6OD5rn5ICwj3tknSATO85W5D23mIpiWPZNx/mYAV8
J6TgVfcd6wJZVMEKcav/s7A6Km2cAmZVVxNK8668bF/sHOFKdLK2gnd9mOZXLvji
8W495S6O9fCEd39iwgcrcINyPUaRBjjDE1xI6AtTxBqLTS1Ag3NNY4n8oy4GnnR7
yIv0LhOCyxIIqDAzS/RLhYBWe5qBf/o4cwtetp+eSv0HLMIoikael7gk3v9/FnU2
1VPk//mt6l3N/W8R/qj7tnua3qmlpYB/KGIm7xX7eT3f5gIlbapIWqOb6k+fHsI9
`protect END_PROTECTED
