`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BVO5xnHqW5a0FJkZYhAso6IWrzwEijaloGE1Ag5MRv8ql0DomlX4v/Nos730hJll
M//5SFDYLgoWGUOoqC+dg4jXl9BFyGyfJC85Glt6lOibdyO5XYCbI4/BzrQT1cPz
dTrF65yFD8ldW1MoHxlMoJPpxxWhXMcAA+6WHIQEcdLgfXQ2rQgy4w+vleW0qpNv
DKVdGjL8fWMDY/qUD2BkjzWM+dUys0DrKP82as3EB9KkevyyiiXrkIWErmvgustm
1XlbZzZNjvDNl2pSS1PyEILcAp7K3rPz4dfRFQ8RbMi+SsP4XqyECUvI4W64iVHB
PrVujiqW3KB+csiapIgxCQJYeKIv6I2m05zr0pr04ucBgKh4vITElaip1yJopgqT
4YcZB8wrRbqscYOF5IZKh3GufEV2hzgkVM8q2jyViY28xwmGpO4hjZzqWWZhFEMC
sKblmf2LyE75iiDw7Povip+m9qSlN4h9q63oTGhs7FMSxa7DXHmWbHEz3oj/wko6
4UZ3H113yE1+KaB+NZQrzA==
`protect END_PROTECTED
