`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3K5uEX9McdJwl4EUzQjrxQB94tSXihEID3wYfAZt3BV35Ib6fcE6Bz9nOZoGG0XR
klB5T2njv6vHKyHgDYuFyo7rbriaJM6S2dCHV3tHkE5WICfTY+f0m5/rdQvklaTK
a5cXz8EfODBQIbWayOIH3AmIkPGUgOVuyFLDp36dqqqjvNB/aVM8nWh6o/NPVkyD
Da0lY2FELsbzOKUj0YC5J0Gqx2cT+mC8O81YmwvOgfbGK3H3oSSrEPZK4CmWsZO1
VHZ9z765ao+cP7BFdCgce4Oqi1BwttfqNNJXYDPmuEqndGN9UC76UpEQZboPeSz7
2/cOPJsWWHL9jGRgGXaaOBZYZZjk30mNcj3KEcWXtBc=
`protect END_PROTECTED
