`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TfgI/S6han7bLKuI2Ct7f7wdBRTD1ZTIKiZGUqC5+uziYJhJXoWH5d/EuYfIzq8l
vOReSZqmgxr2wFAGT5deghAWfW6vGl6fWFiOFpIwxcoNrR+eoJt2GW7h53VPdWSb
lXBMFOVHXhVnjMhx2OPBgQNzSelWASA3TwozcTwmfRkyAOzkDCpBPa77lAy7/mIB
6zvo8GaVKV58NYeQq3rwoVSB6O9oDOhiXj7pwBXbvHwVRlyoKByinhLEZQKzGPSJ
MayXy0N/WMMUwndM6q2VfsfSRO9BSWxDPW7I4E/Rms4zsixh7heB8EugDTg5DSjZ
TC8qWiNc8oiN4ubNeywAdbRGK4i0LxdMvB/X8vR9+5OFK5lHDm1b0QJBharaoLBN
ENrS6RrZBF0bQWKPidsDiMWWE/jplASEOn5hO+TwAmNJhwPBroiJYrZLX4DkNJqU
`protect END_PROTECTED
