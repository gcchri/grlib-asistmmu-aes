`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tJNEooRClL/Ng49kiQuQkUfZzwFUG50cXfeOtjV3Hk1DjQIe+dmtTw2Oo0YBRWCL
J5c60wmvVEKi9oi+v7xgJIPO227uYo7LEDZ4xl93wUWlTSt10L1lGwhMVxooBfAW
3XwdpP5Tgo1a4S4NbPfwHqMEgiRn/KFgFBlHCNnqFuOht3OqhKR0pOxE8Csd1dfe
KS1GTOba01s7snKTzeMx+h4hxe6bWTKZlFPqnb7FydtZe3BPbS5mIf/RayBQgj2R
ohTPvB24MliQNb9jLtgM3zlyUJ1xDWtnXaLEXUoYpyYJzesxIaa12HcyuHr64z0o
0+EvMuC+8A9PnvNd/FD9Q/XpZnHbolKyujiLXPmMknzGsLQLA/oQVdqi6PtfoMtX
thTUja+Q5Z4Tddq6uLydog1yzk4cGoTpZiF9d7emqrm450cLzFg6rb5vb9//yXOZ
`protect END_PROTECTED
