`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BEOjo4xHL47TXxX+XimMkcaxlquAgzji4IaeS7T2tcxfXZxXXe1bFKKRGjrGpfbb
tXwx1Ck8JPm+/yPQb3vJqJRmifmShReIE0vlnkaiICbk/tBGILLJh98/m6LgxgyD
1pGXDVpHVAQB81mT5ZXctNexBUQLugnlcO4mq+cEAis3fnKwmVVDsmBE/xd9H3Qj
7pL3QR9oMuWOpnrBqHBVTt1ZsI3cD1VU0sM9VUyvNCCS7GXeBFsm4QASEqzySuOo
apNW+nD/RlY5+X5ONoYFySxakd0oyDCs9cMsg4O8QmUWzBEQYJK6r59ncRe1MSgf
mQQVGPZYJOpctoc610Fk7HUk+mdC3PGSkocxPKgRZOx/yI/RqoRcirOyp6mKAqn3
rMxDTsNWD/e2Jvs2gcYSpnKkJP7Ow3x36mgYK+fkbY5AynBfbp6VTVJJW/KttmkO
hmzsopSBB9nrjQitEwNTog46VH/34xcbuhKlzXkKTqU5zQwocJFHUBPiMEgGnk8e
`protect END_PROTECTED
