`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gOwcxZibovQv73gu15Q8TzAkm+m1nJswDJQl82VBBF9YCe4RzoZoAkKi4AFc+mWu
8FuQnWhfDF8JNp3rK13a6sf+IOGiYleXPH0A+fkRwloGNyYEEm/rZ08WSamwIUfu
PFQ7DicKrRfPqmDqag9xG4H0jKGFRLpQwGBvEbN+NUrt+/j9CP/l5tJIObaj8esq
Qr1iQkEpur8kf1p0+E0mnfqdo7Vscag1hnlwWGHREmKsacEhEOarK9wRQBwaUVoT
23BTa9aVt0B6SX+BEZmiy4R7qtErkv0VE68L1v7FQGkG1bWUgDhFOHClkk+zbKxV
MmrZa3cTzQim/rkTuSbcbbGTox6Nhp7w3EQZ5EUDT1bNigtKTqH9QVqiB+Ga4OXj
mM+QvjDYL4Q1fmZV1p94WjioEvQw8TY071Ew2BH6EOjBdvBnA+23/LM7b9n8R4zn
nZetN7vIb7aMbCKcgsmZVZTdfcGRPPBNe0EJF4waY+1h+qVv1rwBG9gHXI1pbd1A
AZGli+WHk/V6I72dYv69KdNzuFwqg/yBIt/VrenrW1OnNv86SxXULxT3cfVDX2XN
epEcfsHOOEs8Dl59lJsO1Hyy/KcKSUiNo18DP/shAArblUqem31/KxDc1rmodNyD
owZp92z7WGRSWgRnZy9Nsl48ew6RnBkm0UFo7Ty+JiLzEi3JMEmxzjR+OEzB44iP
RXwJOgp8Li428bpIM9sTFfAlxJB3cvIuQdYCMWLyA5d73+2KDcylM22551lMPdl4
lCD656c7KfYPvyLaQ3PE5x60D3vFfv2FcPY4oFByaAtBjkkivMLVKiGZsXCPaxIE
sIgs20Zl12X+KnkSUQa92QZN3LFybzC5eORIzfPeg6wIG34Aa+XG1Cy8SaaOE4YB
wyDdHHgRPlekP9vsNypMcQ==
`protect END_PROTECTED
