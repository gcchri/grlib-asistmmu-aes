`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6RmF5Lt/huTTPgqLrOdnK/b1zpbS/JqqB+iNR2+yI4M2A1qrZUpMldQnkZsNJ98+
KM+cadRkFqtnwEQQags/xYiK/PyHotql49B+2TwxzZovvQBlIZ3KJHMpuI3FK+Db
UCJMAJzHWduh2JAv9wphU6ikLt8A6yoUNhlbsuUvHdAwzGEpQS224PJkz3CPJr07
lLesgGdAX2am4tm6OiaG/GrcuVuo+SWb9pOyDMmOEbNjpha32eF/cM18uu6N3Hjy
n+7k/mmCOgCYnnmYX9H31j+brCHeOO7FG8h92U9NJCx6LWGUlDUKztsrU+jS4Has
CzzE2UA236nOd/UYc6zKF15S2JyemyuaJ7+xZImZAIxCzQaJmXDdzlRAmz4xR7ai
6qS+cKmiZt2fUebz3OEDmh2yeaRJRd6UTHhUUIsPG5VeHC8qC23HWOARZ5jOGkR8
xpQ6w8ac8s4wEjY0EaTRrOfBSYhHTdu9HNEhzYhiSd1qzJWW+FA138mKUtS3ROcb
d0Y2UcyjjsHnWvrLGhZ7hqkV4co+PuxC7SiXn+MUN+qNwPp+ctCO3XwlQWxheuLG
uTm/bcVnYplnfbLnanmwQcpCYfGKYuEReoG/4Wz3lKmWeUjAX5zMgF9q/DtdQUHL
WBfezYPo4nHZKk2ob9Ot2epyDtmi6xORZFxeVaj5YCET9AQGux5kmCIV1PuayvgX
BifmhzG+5gVbpo+BjWae7sB6jLRUiQVpYHBEdwqPKU+Dp2rgxJQqdmM1SrOU0UNF
v0on3UfyoLikq6ewsYiMFngtkeuo/RtuVO1SgB7gBQoMqrpI9aeDHzaU1FevUNFk
GO+Pl/xoYIBj0jr/BnvZSpify2KIPv5b1jHpZQAiFlZ6dGMxRcB7WmtxDqDXoTfc
YnqXQOMqmO8iTdiWaK+jMTpegPPtl9TPcvJzIp3JGqMMf+ghzNF5+5PNiAhdnTRY
+0boY7QTJ18coC+KuJaC9n0Be7LmnSf9H2FYDXPe477/nCynDxDSOgTYnGd4/uNR
MhK1ehbxvl5Gq6+WhVRc/3tMPdaqzfJpj4zmDhuent8=
`protect END_PROTECTED
