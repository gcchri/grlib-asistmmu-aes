`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QvmRJ8sTbKIoeqtgNOJotBuZup84ltjExeGvm3EU2rCSsdve+v8tmQ1lpyc5RRXi
LSA0FUxE9ucfqx0R2p/GdIJan3EChCIaxlLCNRHtB6cyTcLPxUCGcbkl3LrsXu1o
9rZ5rsR7Vdz/bw+OugsbtygSMBpjf2CJHcQkHQCSEWCz9LbywVgTyHcw0r6Wyayx
NLDfBxZw51s0B1o9kf6UpYYrq5ECmvCiD2hTQOW18HoeWf1da63HLj1SLJG5xdET
gyRLtQZ9YNq1dTxaNuV3v9e3dMkYTFomlOiFrY0TKF82sRU9T0sCyrHtrE2ifOqL
I0kLrcci9QaIDt6Mx7fFjA==
`protect END_PROTECTED
