`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n1+WzpTgjs22xqVv9dtk3NVqQDjeVayvUeAygGemsWRWT7jovnEP4Te7PVtYvh+z
Dm8p3Y+z8ETSO/oFrW2KsfgWbUPrlMcCBI5aTUMxDkJ/dAreYwMZzDyOj5Dcmn7v
M3emqJjZJAiUJMieTnJQ/AVG+QR9yCix/GPFqJ/ocQ6IJn0wyZI2QqfIj+pgQiyS
KQ7lQIoPiZO+VZdYwGWaECEcevKF6nFXy2HtAxd12Xax1GiR993MZp/oWsYVfhif
DRckBP+tA/OFfZ0bjtWxaBHGgunKkl6exYRdzOkVVhAtZ9sjv0/PlYBcyV5bjf+r
TPQrnqf321FKqNqlLFG62DF9o3YuIamHjINyqdTGpF9rzzM0tMRj+yXNEFLTz7dp
lYqcNS+MPTAxU54DHRmhZYzHmSfMiR3/wutLNymH/j6e8MQOJtcLsRVLE2dktqPj
F8Xifr7yCuSf5S1iEUBrkrOyVx9enN172HArFxTQqz1Lt/HphilAvc+rImU4i+DK
QpZjToemEif8I+yaF41o7Kj6wqahJOnoZwUW4TsgYgCqjSD9Eixg01s5/OHJA4NH
iToJU8t+2I6X4cqG9l9ZsmiJnbzf4ZKONhGIdTIpU2vQCRQKtlriFB+mr/5AuuWW
aB+PJW6Rz/XBsERpKeXJ4B84vKzhaFC1v4of2AsMu+KG9wsxuIffo8m5Zo6izHW4
V7v/xBv02zlC1obFhG6zQ1aINjkb/8iAZpfyEQHkbcbFl9EyvXXXvzI6Wf03Wmc0
H2TVxZIseWRdMquapxXS+w==
`protect END_PROTECTED
