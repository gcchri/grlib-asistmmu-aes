`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hF5hJlJZy60zE5sLMxHGZ0dgEKjMGwLGJHBTUF0if2/l8AmnGALeUgNkGu/aGFUs
I/BdRhSuK/te6jWw3zlg3jUeFVRSq8n7fVN0A7ia9mOkF9M/eJHmtexjUweiXPNV
x7gPuuMXrt5KDfSECJmNu8MmaZUhpv+MzsAgMFgQYIzaYTz1IfP0HK5P/Q9SImtu
qhJd6XUmR669cvBxf4mHwpLKFbyAq4O2cODok7PjI2cdcIBshzkXuFoxpOv8Dk9X
KBVFq6SnlRjm5v6192te3A==
`protect END_PROTECTED
