`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tu116z8DfOQ0DGJfzXb7bP/Ic/DiNYgmje/pWYTeoHZzhNDshdoa0I/TlSKBdjE5
JFuwPdNmsO/SP/h5RgbndIynytAHysSd6A6bvayYVv+Mm3dOIiZI/23o4nrjln1w
VxBFX5FFsbzN6/uwvwh+o52cJLnV8regwPScYeHxSyB6edEw8eiCn+GAYj2t6x2i
h8GjQJya2ZNQACT28QE5Q11xTWJgGZ/zqASEdyhNoU4ZUxua/PjdLJ2oRi3sntm6
42E8WnzrKSnBMent9wXONxUDjYpxil9Av9L+vpSgpSjSiWbEPxFxinAXvgXPd20R
py7TU3yeA+1AbED/ji/Gh504tFMpuNpcBVZa38naxCT7J5lZfH1uj/A2RQcXwWbi
zVvRtma1eDtNy59UFn7fXJbD0fVCHcaHa8FL2Klkmks0QRk3TVpOj/Bpa9C0iMMd
lO8j1hZ0Z4deIdb+BeejC19UqUf2CIHRM8UqzoFxlnJNMklXJh+8U50t9BFkZXIs
vj7YMA1PLkzqraN4CSwhKfPatWbpXLJXfpkrdppnPzhVWvWWXV+e+c1HpLm/OfSN
FntuOeXWphEnk3HduJVucoAPd1HGm04t6a68s8M1i5ydx8w4kwoc6zUqcmJzD4lA
kmILjb9SmB3ACbuRsPs1O+xDMvpwhRtR/z9JXXXEyrHPqSwh9xs1XoGem/Y7Jseh
75gsbve2RCBf7PO091LGVgKIwBo6k9uS8v5nvVviXarjUUpGdHZsEehDHdWr7hVs
NL/rLG6Rlx/2tOrNnjhFlg==
`protect END_PROTECTED
