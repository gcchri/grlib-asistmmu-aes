`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7aP6E6TY2glX3MQc/woK78Wge4oiKof8iBPwAyZ8i5MTEWbNx4bEdWtcylUMo34H
n59Zo/GDVICj8nDgDQqqUEZ/i3chPmrnnE2NxQfkCbgiKk+mRJSpdkF3CPB2bHrr
TXoKNAlqoHXXgHajq+Nd4TzUpOBlid1gMzROOLZJctd0vbGAfzp+Rmfief9lc+Pc
E84Uduv5ZmaiKAP931WChoreyrm/JrfO3o6fAHULCrbqlzCEL0K7TJQFM7D58e0O
TJmGrDHEQKo5GooGYPc75xJ2Qs3caGm6PEQf3ueIdfUu2ZgIb3RweVwNAncZZrrd
bjF8HnUdm3U5g05qnbuOLOuunNnmc1kcpSTKYmwRSVtTz92SqnSQUhHQ0G3wRAQh
njNqkJoxp5So10n0M6enJc/XcXxlka4Ko5gvo7CayoPTRbcbebWlbBtS2P0tYLB9
hUAImUtqQcdyI3Z0nf1ewJ9KiYTkjIY58XyBWw11m34=
`protect END_PROTECTED
