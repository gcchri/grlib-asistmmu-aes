`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0m7HUijejSDWuXGhShu0iHxFq0yPsiiEeQqVO0mT8Xc1+I98+q+BJvVC19/hrxgQ
njn9EEQO+p4DqXwgXyhcmqxKK3LgirWGjByOxWU6gJOXnCpZD8TtjMe3hO8XZzaG
uhmTOOvuMhPU+CyJ/qEgyDZB4jZitOA63NFbhiupX6kEQi8LO5o1+XIaIPiV06MS
VA+8A9Su5SI0F8Q1Nz6/8kuk9qjlH9M0zOlj6NvjQxUJ892YIsIRhNsFYYQh8ote
C9w6TFwQnLL9UXq63Z6RFqCOtjlJNS9W9ELmPH09RMSeUQzyasAuQsdZ22IzJu2p
jAfC1jepDFwIt6c9AKxaR5cEIFiy9mxExQl013ZCKJU=
`protect END_PROTECTED
