`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CbzIoPK5Gvw+ceqEctIJXkgkTuct3uXlYAYlH4Ng58z1Iy7V9mohpYCPLc9LD4IH
peik0mKeqGFbVVuDUSNMKG68THaI2altO4yfWuC3nJtDy86Hcx77QhwW3IUQ4sxe
sIM5UYv2vkR7+hZuztSh62keDEt/AdMf9atMBhgxHolBMcvhJ3KuYbXxAsNibs9Q
nG+BSeQ3XCoW6sXxRgX0ZQwktH1k7wYFPjPXn6iLeAv6zI81g+rGKSGJv6ZpKQfc
lNSkaNSgLdsdW+QoOop6LF9lOCM3fYFsZ28Xfq++3uJSTx+B4Z1StYrY+BZGKuMQ
XOPNMT/Bgb0qGousSVK5/9P3J4sj0fV3v8jPvOKZVsUNOs0TuCUEJPIUTQKmCAGd
G2azXQClFouA6HmUEnAXRyYuPzz3g+45JcDdH9f+sKfCNxGlWOmozvJlhfOTgD32
6ucrggAJZxW5/hnkMsQ01s2ofvzOIPnjGyQjXcR6MP+wq+xunNSIONsrlsjl7DAG
`protect END_PROTECTED
