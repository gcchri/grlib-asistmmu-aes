`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KIjoREwT531yhoTJz3/dc8qYs6C001SaW1KyMQ7d2MAhijvnQgbp9w1gYW+5++oH
b8xCGZzrDEaBuZORDnDrtJDp4fm19e0VSkU1Mp8E3SbrDsb+m6kg309QYrmYTEuv
LDLdHVDFqkuSjUz82AstQrptlDFE6DfwuV6dicLV40tEKJ1uCYHVFt6rqJEm6Sns
HS1rs6twtAZgVF8uzhIpI3AwbYldwEdpulykrySCFQFzA5fvHx+dTJYCepSDPE/w
OXpwc9sc7HKRTTlRcB9znY9ahUniS3nw7/MPOpewD1RzL568eDCvAu3T3e5HMUsY
Cr+tSUOKAxnnSU1iJAkS+sg4+gMz6+x0dgUveJ6FG0SbQfgVRYSR2Hzqzamxvfpn
3a2caA2Zpc/S2ZNlmui4Ml41R/tduafZJMxXCttvNaAUtl+UI0827YQih0BPz7Nm
tTW67AsnZKc8BY8zypw1T+L5RTj4Kpmdtw0W51rHgH5m/GUp7g/43gyZiGarNavx
`protect END_PROTECTED
