`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
absveGRx9fr815vE33NNDIF9KwUGOJSNrHILUVeutCTRqz9ppDxYxyvS4lhuqOzp
Dq/4WyYZBT6xfG7hogf8dWaZI2wE5QPlhLQCFzlhSy4kC9/yb9Wq3NdqloF1Amwg
xUMUpN8R9tbXX+vuNl8wE9qSHYvnnZCPukzxFApC/Ty/DFRNrLIwByPWgGlO+3lZ
CpfqLL5WTlq/HwtZlJrrANo6ZEqfDpmau+nKE2hKGkJA7Rslt69UwLIuYlvZ3ZX5
Rm8NyKnpZUBeOT2QU5jaFPoybMKXH7tUR0s1NokHhsGoFG/uMNoSnMipqWedmqDv
X1wg5NcVNwq860MIcAl9wNvdrPp29BUf97ys2BCYu9F9W9ZU5uAga44I+qOr6Sal
9y7NZrLX+1xgILR10pvlwFepZQnXYVWEFGQXfZ/vVenmJ1dC2LvH6qRBIpekNg4p
DWBD4KVAQrWh8FnP6+z7zZ0lf7SPLjHjMtHWye8ZuFDqbhtKH4WJFin8PFIUw9ge
L06ujWf6dVZ0GwCFd5l63SoDf4JF41FbcSfkjX9sxJ1xe/kFSIkKRnsQkgN5SzRx
GfL41y9DkWHLfr4rlLH7wkKas7cybR9SR5d2zrzj2U57OGDLx26xOjHcjUjop0hM
TfikvAq7GCQrT7xYfZEAeRWfrSrzwhlE247jtdhcm+Gx+YO5XzgnpYUaSvBFK+hm
vJJTfOhbOnthdokjEsSN1SyZpKXpVcwFy5bFcuiQ0rxDbwsDpDrviPho9Red89n5
B7L0X10Hyc19CT1IdJS2yswBS8mgqvr/Lc9gn/AylYXW0Dj9IkdMOwJga1qPh5Gz
VbUNWJbS4hnKf3NGXhvJFLxZJBIcwm27tO6UjdBAJODoeB+d6brd/r5qIcWBRDrC
GDSN0Gelt9bRqQDJakiF7tmltQbxcDq1ITBbuSp+eBdBs1Ua+Gkbp5KNu/yyCoLb
IQACmF6nC4noczU/yjmLsUF3pzumyAn3DFRi+ccru8xrHSGitRs/KDmEWEKTejoc
XkAJTenxQCw5zY8o/gsxA/E2KYb+Rse+qS4Sis/KneA13m6xmywlpQRVLKDa+UZo
I/GiWItotxxT6HKwQrqK95BRjaerd78hXGEmSwx/LPqUPeKESJWUExeb5Oklb9HO
F2n2134U/kCVPlgqNWGXcQtEkIHb2Pe4DMpT66JDpqq6wEAv+v1lsDv41zUpu1tf
5Uy3uxCNBNYQFWGmt//Zu0FI0Jx62QUO5Yt++J69YOXts27EU6PSqFqAfPZ0lVWJ
S6BuKLI/lOgjUHuOn44vKOwqiyHyq5JtfHSMVSTYFvRctPH97rwqa0WKDnQOBbMm
THKTufrhH0KD6YGFyegWi2ZYPbtgIV4X/bzoElQDYZXjHdANOhtpuga7Sr2GYd+r
0LSsSGhPxFBxaM5jSnE4TYBx678GRYhPbB4un0z6hMMh8nn5llyCEds0rfltizDi
oJ3B0w2X08e0Ihn1n60ZvuZqKOkgiIOFz6SRyqNVwjTqFFJ2p6SX4PdNDjc35Own
/G0SrMiTN5nbVsPBg6Rh+eR5qr9dYgy5pvbLDxzryoba2UyJ91hKx7avRz6J6AlW
8ZQDnmLmHdYQT3MWnDQRIS7opOxP1xSAnPjxZ9YgK2J/9rADPFFZ31D+T/1qxX/U
ZTmonq8AHPaZwgaTtLFCXnoF/WkaSHX9X1f6RMpOHu0z/t2ZH5G1hkeQHV04uukm
xgdMDPJoUzmm45IE5FIgycxTzNyinhTidJfR7PFb+Faefq7g18sJ66bYXT6Ubg1N
w1evTdLgNmJ0q3NrV86IoQDq3wYJpvGCEgMtjlJmTJ3x4zUih7nB1FI/n2laKTUH
jR4RKExtv5G0guTbyOQkuzlWNLIgy7pav7Adus5dOurhtKfDlk/VD4bm1AxrGZda
`protect END_PROTECTED
