`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8IJLl/pxuzvGwanEy6vuTvFz3voqu91WvqnZmcD3Vfa7Hl0p3JCxljSrPiGAnMbl
CZFKQzFk/FRrkC1QMTVOZCmvux6y6JrHmYP8aigY72gNI3JW9FJ5fMkx6z3pWPWm
CiiWfifw9stHZnSX/DjcwUn8rR43O/0C9I/izGc3mr9ekpPoh//MBToHl3irLVz4
4YZ452IyvnyexzNP7d7pWGqXpmRKG5AGUo1HkaWL1ZMzL67pgprf79tvVrXN2y1g
TcefwMiFcyuIH4LXYQ4FIgYVHPb7WzL6KewPIWAYP4MdZZ/UVbF8r2CayBcUaAh1
3tjGNOxBHFDKRyS74BmH3w==
`protect END_PROTECTED
