`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kYCf9BNMV/dXW9k9sPmBA++MvkHzTGzmlVYd5rNoa8+Kd6JXDMWGLY+CXWGqTw0j
CTrPzesiAtEHwGYddI7zdjLq6ABd6WvfyBBoRvP7eH+eSCA9mZz8/28aXegjbl9n
uNlu4/0V/xUIGuSXGpUIDWkZ82X86VxFDK16wLp/kyxiMlXQ95w7WZvJONL3EvvG
bMegCq+YBoWsZuTTSQkvSThfIB0wfv70An8MHz63h+IQBSdlefrdpgWDuq+AdbUr
MSU2dC6k9ZfmrF0mLDY9B5u5oi6AU/7TwV24BQUZdgA276P4Ent56UQncKqYgzKa
JUc56GQe/r+198RwHiFljXjyTyHbcKAarrDMxrZrKM7BSjM1IamhUdEZR+rnc71i
RJpFeDuP5bKLlN1k35b+Ell5mLQ0OXjh0AgbgFIIHfBbVYG40PUf4PK0HhqFtqMG
VOPCd/NhTByQx7mSkXVxWvw/GTTE/4+ehVUJ3vmOJQvKYXmAA6Jc748ONzidIAmk
d4eoF+v9lVmPRZD8WYuwSPn8Vfbx1A1zaLxvea2QC03TmvE2IFN3lr1yjMwZ8fNU
4FJSN7cgp9XPXn54Na+SQVuulW+QjPF0jU3Qbn91Q6j29GzpNDpJm9/uh9fm32KR
D4tja55RZ5Cv5PZROKKsApdmW3lbi/iGrJlnIZ/vrIk/7McqEcQLZ3BZeWPeNWSK
Qv1tL3QluWHvgR7d1wRVV8+Aq6XP0TWkVVuVXs57BUvLBNqiMxiiptDAWuSMALaS
+TzdBmlc6VwQQX2I4CeqzQhdXbgIf7vEVYF6LodusXW3O/J0g0sGoMjFXC05xQnS
kLD6YfA2hB2wAiFdpfra9/D6J7Sf85lRZoGWdTPOwAvCw1rtfFNTUTnCKI6ZwSBi
nz7JAAXuwk1ykvVlSHFNPsufQmU1tT5ekmri0Ua6Mqvnr6GnnGBcZwjjtTWR4Oh0
TTHaeZpZXSQyoaHMvZbADU/N1wb8oo9zh3AJFXsEh47NOXQaqitj8B5sKLKgnQLn
lLKXEMNgqJeKi7NttikpH3PA/J+rmVFme4m78aDXRnlzgTGpY/84efuh04CxMhkb
LOTawdkRIJCd0YTICrxRS3TgcP1Jy+2ZfDVSj2fbxtDMpzjlsOaeDyXRzl3IEGsU
Hx1InjTKAbVKIBJ5r27DjPZ/jjubJGMVw2QqavuObnshKgc2YKFGqDkx9zn0W8x7
lE45BL4bhDqF38gEbMcBJuUp1sb+W26AvmnrZGqK7tOlJFwJEj3KvrQsJ/PxERj6
BoMiIiW7DQ3oeSvWZPo1RP9QmYN9TGK6nomppQIurG27OFGHpiQF/WkkqrWiM2P8
ZViiAnQs+3ti675mmpzbAVjmro3CtYgsJrqCV0kjUEGVbZQ1xY/6W45QOk+2T3Nn
8R9Hixcw6bD+8G6LaFiHl3Rfsiqh2mxZ/2I6vXZiaqL12l3SBzszw8O7GCPn8iYH
Ho/lNiLiSRue1xjDpWg7f40X0Hb6Q++VaTDkepXBC/ph0Vbf78EBDUsgOntMwT4M
dLkoNOubJ/bnor9AfKxTv/Dso84Gf020a06nAayfRmsdFEg0ExvKtnEqqaSFINUp
dNjdlqk+uVDJDw2tYf5+BDv77BbMgEP3clcmzvRgTDyslII0kg4PDNJPMBOBeeyo
1y6xpNFyvTKnIPOZ9HuJKkJUPbAd6nEwxUxl/G2UK6hLRTWUmY5WKkx6KHp6Ctp6
c8FDwIvCZD/jXm7UnvB/GBnYMJ+otDdeRhyvk63JyecA8WTMvEuLN2jzQa/w4a7s
RUmYu0QPeJfa531yduItg4wSd+KBKMWa8qKXk6v+B1i5jTBOEh1dGppuzVQdmU5j
lwNqoyc1O+uTSFtxQMQU1S/REnbJyZ8uf9hjLot1OBT5EjG+EEjaT8JFFzwUrJ7o
a99mHrV2j6Xx3ybiRa04Pjonf+nDS62Xjjl5NP1rgxCYaAcCOMybnHw+yVzOl0RS
eM0CZ8Zoh04cXEoVZKkXWulZE/SLEDTlaCGdWZT5ugAbfkH0aQNxT+pToB2YgyzM
reqDOfPlQGGekSnnh1/iVQCOIKqgm2q4u847fc4foaZ2RkhaU9H5K+Or9WlxJuB7
SnkJ+NrKmmIqRia4iGC9X8c45c+MG9YXktjO6i0zkj6QWeBRkoHm+R7K5i5uPwFt
uNj0HOL78OpdvFbkZVIjTHLQWlkJAGgQc4I9+wICi/dwYU4pQEiKMcf+joCQSxj6
giHZiku6pinTqqw4Nn+1+tnhAyDKT7qnF7a/cp6P7FGbovHFZ0rIYcDUMbqdvE2T
eprRTtp0OLhEVFnS0faKpcLvdFwwGX8dss+e7Y//AcIIafl4E4kylsjdDIVmAXNt
GvzxBqQtaprgBNlARdsvvdW1iEW9lRwLDow9WHlFxkRlYz97Knn9ZbqeZ5A5pdIm
fxPU4gS8ggfUw+1hTsDOSXKRBFi7b0/s4t+IeLJKgHcoYa4bN3ugoKfGG0t7mNAT
MfIzknqLIoVBgYkaUgTtLz9LPAxELTHQtLNKiQYYh8qTY2jchqd+gb+FZULMHwpW
3YysbO9S9s8gRbc4X0HBSUY7eXKhUfZoDxPkSHgZEtO1ScK6vmpKTga6iyTDhmec
xFqtR92jw8fh9JKqsj58C88t3vA+qbSkrrhnJTeFobfofcGn3lwNdlMub3b6o5VW
XQllXNzOnJugSg/tOMaYF/G3Ia7XXhYyXkkK92acIg5FRF04DLyMFCRImaEXnOWY
HA2RVDPx2H+qMswVjruVSDZp1DlGNjOyzs6AsHybGWvBLlxkSUDoz0pNV3zPODOj
LpHtJf+ViYQQh152IkCgHB29ed8cgZkHB3fB4nQvon8OjnECbeMyafvyIACR30Tj
sZ13IheZArk2iM/TBPFIG//mqczWXZTIFnCVWhmYpi9kmRXrGK8iFTFHuP0E/K4r
B0sjgjpihRe1ylJ9HeTuxNQQh7l3OtTFPSkDrywMvZQrncNIOKR9MW2/ZsppM2BM
c1py/WxCHNCLUS4jvrrgHYutONaW6xWYcmCVUchn6Fry2OZS1yR3RChNl5X0Hguk
SMfrbgGPUgE28ImNnRSYGCI2vNJiW/+oQuSwWCbmMaAigZatmQdk0gjfeNW9H3Zg
jCBw1WgyPLvzBzMBYgIVmRVDetsIElCKXYyes/5TjEBmHWWLyDag4NUa7VzBKu0b
rs0eWZqw+1uKLSLmvLwJH4PZi32Ph/I90PG5tBidEVQHo5/BRGNNHfUOS6iKhPyx
zJeQ+jyRaBK1mSh8/nURXQH5omPLG98XQ5iUeHmi67UjMDZzhjUJE7mEc+s9/qmp
HhkYSG9xsB+OW9Rl2FZa3M4bVFMgoNS+3WAivMQKeL88MOEaqZeBqAVaPmrp48oB
oXjmvlR3bzXUWBQqsPOaFVcoiGAjzLYJGgGmXuPHBDYUza5gMBtX/P0rK+HNIOuB
0eEtGYwA7tv8ECLrc+vChn6RsnUaDGSMgz06R2ZmUZOHMWaGLyjxD4xgUD7LhENS
q/ewwElcbo3xWVk7fpqXU8o92hyb98HhsTUR9bsXaDnl/Y+7vIKl/seRn3iMH+qF
JTIeCot5KQwTLGTQU/WmdX9NZovbPTFJQKJ/BXiMgExCT++WJXpaVa3YJ8ZffRdV
lmKlKL5i09dIimtUSpAg3+opgpJiJOKgWLyzHCvNwr3GvXYAI5rUvpxrpgiVUiv0
KscuFyGZMA452O21hSE50BC1vngZzHnk1Cj/NCHDPZiuA1V9bmMyUUh2hbann9dG
9YEO6leGQW3K97w1/qTAiENbKU8Juj34tDy860DxCuz4ZBDPVfOrMDZ89Eh5uIap
fXmYIOwsofBGilyWXYA2Ollv9urCEeCD1cDURD95Zr+hEa9LEREJvsPOd/vCY7st
xTvNxWVRB7nI3kbRFyxh+HSknTMJuYAaQUMpsN8o0hAXsPZUGNSmo1aa+RbYcRaz
GsHpLGpzNcgfwFdVCOtHDf5u6JpnilmcFH9Fnos4xdzOUuVuHI27vlYlKSKyQxMu
tQceVAovdxr2wyoaAvO+KxJXJLGElcmxAPaU4VDsaQHQewjRB2YK73IpwvTuw35A
NzigHNSIAuAJffg8lJzxxRT71wg5K8DFlrvKBLATaTv3b04eY6TToxyJSDZVmqoW
6VdSsxye0IBJ6huODF9Vddzqm1T7eGHU0wAI9VSGNtJQzyPgY1fGIgcwC+CD6I57
TtqeBUyBGc668isMiynPRzqMFmiPcQVVVyyxgXBvdqIDgNb1NhyHUzijHppxupzY
Cj2KNFwkniudmceS+NZ267anp9+zczSQv/tJzIq6/t8xVTkHfBMSf5xaruRahCn+
F7OhEPKChqgfwwW5GrDXyQfHzO8YoHwpSv72TO90/cdkt6a+KEnqgF0qvRS2qlX6
oQcKZ358yVkj/5dKZS6fR0QIUah8WtLQXri99GveYtwtnjq+uy7lz1ZM+PuDbA8B
lQ4FY8I6l9BufKQkT7lNrM/FrlscPVYs6Ttq6rnn3e6VvxfL94b1lDZPArwgRwqT
20WLrk+UVP3llITPOdc/DceEfn9lBaOMpp72gr5mSL6X9JZRi292Bk07Q21v6hwH
JU7tGKmVlijFZ6j0L8XNLf9XB7ynM3KtBsu2hbh40xW+yi7OUetCVAOvfTg+sp/9
KaC5yJk7JKgP9Bq5G58hS1vUznq5NQHKiVliMRGulVsv8OAge9nRzeVay0yeO5Os
3pEB2PmJ3kz/dL/TnTibMK16/H5uk18cbZmCHhvCyxOO8rQAckvd687zDah/iuOn
OMP+NHASMOB5bd6M+tXuw0NTtGXzYCzALx0TNm7Ul0bNTrlR3abF3DWrxLsvjpeh
CjIyEaF7vwzO0NBaPOeQGrYZQO+zSGLtplIp5ueEiXPNDpKVnqaKZ7IZmaSgBEQ4
FPseE7AzDtz6tGBhZ6Ogydc84eZ0yMHxjxMe/rm6c+6ssycrptYKrescZWGKRPcz
nLcptD7qivoGa8gJ8IQyl7zdoE0BjnYe07mlNEprPowGn4h0Mk7I1yphNeAeIyZI
Yg6d3/Ok8XfhiSdPQpZ1MNRigRMnk9U8hmWAiYtwZ0CWI7nMnf+CgfyC2aLf2Mky
n6Z6s+p8kDghT7lq8ChbnUzRL+9BP/dwSvNP2A6UOObVHYUoKjK4R9iZzpvuwr9S
NQ4gwtlSWtJOm5otIamy864N9443rq/oBfpHH8rPbQEBsjRZMN7DvoRExOrcESOn
d77oH582vZZ0qRx3urzIywQ+moQC4CdA+8YCpjSxBvFQVycn6GQcWXG4YNzz4LFH
1TTu1+P+SvwiFi+FPLp8IqK5DOJUWWLQ/qF2u/+XWaEtJCUvkxOm2O2lEf3FcfN2
EYqrBLKyn+9ltJVy8f/xSKkwO7E2AwlR8f3HKtwGQ0jDIFd83dzwCg96lwxGbW4S
Cvgo0qxcM1sGx9+MARanWsRwGOWagHoi+/CDpl7kre94rL7xoB5risl9+9Pd8/jz
O/Z+wkEQHU8RPbE410LQUL1mm3fchBXGpzsWlxUfinMyTiR8JLX3nRqX5dCIdEgs
nIBpQXE34M75jXrcIJBxrQvzJLNWRZSZINdcqXDGoacefIi/iaaIYkGrh6slBHXm
J9cvKc79l66OZrc/GGh6/insyAeg0WvqShTKIFqyELjtLdoCa7Nbms9Rnj6OgcTw
VPC9kdjrGMC5UdgQTxIHh6iH7OGq4Sb+uy8MKjJ8VnbLNrEm7KDCwO4STancc9Km
QaetTCVu6tA2xUZjsvW6Wytpx5cBcNyL+0ZzEAH9aUWoZaInwJKVfm9UJiF+Fjf8
kZDfcq84uyi8hk0RV2MM31lwXOKUViJ7GoL3tuibhKNaczXlU0t66/O43yPXYjzD
j4yM50NPLE5fznljco6aOvqFDDWVTJIzWnLtZTPs4MvAEw3LVzoI+AUG3ERLvOyz
qeZGG1Y1sSiL8M+Kpccv2z1S/PLaMBPEeV9uXomPHxvtWVvg7LV8PpjX0BXTWFko
Unq30sVipAocDZXAAgx58xW1m4dO078rUktEHsKNCfq9yv73jtIQ2Mv0+mLarnxJ
2VpqH/1s2/5yQpPlBUNLBV5qPehllreIPgXa5zTkby6ccCR8s4jiXkfQ4d9buUzT
Bl5YNEf4vp8ObDvXUg5DiSDiluxXELIUCbkWFuZKMgX4MwHN2r5DrgA5uxNZRHz5
ls/gqg873IUUinmMxgotgQXufVocITKHcgFuhfSZKwqWJAJ2LblpUxXNlTXDlpwF
hxtWtK1EF2k44PwgaMqbBIyp3OyCh9MW845AHvhf+LwSw98wGECnqEdrmetmRC7p
buyuIGBVGr5s1USCQoD1BmvUDNI0eDkDu6Dyr+37relQGpPEgpQocjiNp3BLWR+v
Mxa3pREltwWlw/XhdnR4vXml+n+BfTFBYFABDdg1sd7wNVD028+bLD8sjLX1W12W
ZoqJvLPIwJcjoD3s/huw2oAG1q6YbrW5enKBOtlV+Zp47o/GqRPMkog0qdyWQTNP
8kf9puh2gUup0Ho8cBvmm7p26Hc0zlaZPNxTGcP1F0sSEA7MYNan9XW7LVBj+wty
LiEN5vmRq4d0l2HqJy8s88YNZ9b7jLURN7hliY35sgjXqxKDKeOHN8z89PgV4ol8
sIs04OoRqo8G8WzLPIw+qIF4CHkxrKLkY/ypBtTVsJ6Dl9WzGzUU7XI++s5Y8k7V
3GrwrGgsDT8UmJ5i/ST8xOItMXBaVEaZJ7upUyGLFaFjL5ZYw6WdTZWNvpytuu/C
RoU0KX8J5jQ+JA6uq/GKQDJSHiyleJu1TDGCfEdZJhg1lGJkVfPm7c032NLYHlV4
gtra4i4j7Miza7X/jf5sw81DeogLrWVyNKbB+RUMXz1/2JsYfBM8iDIOTRzZLZ9U
qKEgi+LeEDrDWlnnrCbR3mKVGvtn1+flLbM49UWU/kxj1SLbRve+EfHVXCIHsKxQ
YqJtuJ7BO3QfLlSSGWjwhKfTSRmeLMhRp40i/Wrfy/WsekdKcguqBL1qROLQMWeT
xaS+Z6jHWeGKtJZbnTimsHFhMGIVmybHT8ZgDlS0k44jQDAGWWUewN0vOdPRJWcJ
QEDpMDGsqO4sDljRawDvjOOuvyCnpImPun8LCSJ7I0pbom9q1xU/+a6j795Tl5tg
wZ5SsvYYjJ4KHywTuIs9jvKsDJcb5ca1uyvmN6Q3S51Od085BwtNBCQqUTtDJGUb
sBDBKOypzWjRzldaghn68UZxLfOLFRyx5Cv5SF5GAYXbSvta/gsKABYReqlYkTJj
Rr82lXNw8pnXWoLoXu/GSA8aQEmAkdFsSvZK+D7+HMafLMKF5KX7MKo9TWwLKc9d
pxsyfZYU06BxbIpTM+9jo+Zoj6UsiSDJdDNQ5MOlq4LfK0hQNx4u0tcGKDyg8ENY
JpMUeZi6nPXJPDLhcMPY2ehQfg1U6Mirx3wAGUADy2TyD77gt2ICWeyyt9hjj3UU
q4tKdzDHc/qJpUFEQVPI74U8qoSUnIYj+NODTmNNKfDXGUwDZTjtg1e+cMhrcGXd
6DXmGVizF5wZWxEhc7gzJZ5Su2drPA/FcQdbF/E+vQDCYIlO17HocPjSeKV3fWO2
eWSeVcqhjko7RaATPkm+smioWNqkg1aiBT+/Lvt7Ek9c1v6a+E2mYlINrEtYYPjb
vumR9GXQrJCOOwWvr5tFPKB3DOR18aqAB2yMeHgSZsbupBCS7eoypKQzR3KfM0Ft
v0XawUj8gSwrCCPmrYXcPgn0IhTcnHS+OIIpi9TPN9+Bwg0jgRIXHcgS3wV9mZSB
o96UbOYXPFXP/i4BcbBhdx3uhwusydp1msCtFCZbaQvmGFoh+zDR8GeRCQk8Td5N
9TdIdl0m3s4e9Q/IsOYOdHIkA6Z6XvDGR0DcWqPiWTudcspIqeAcO+4qnvsaBFrV
wuGvPslNRFprmNeBYisvPGld+zIty45x/gR1Z1eEepJf6A5PVmLczmSYvstx0QiU
/O750yUZaGym7N4E46rlJsr1QDIL69Xb55ROlEFZqCmwvVhVFbWrWcj2V4+PBtj0
7XJYmDIy8FMNwHlKmX9X5PA/uBapQ3nbfvCc+vArrtMJEz0MXCRIlOITJ1fRjiQU
UeAok7OJxJ4bhtwdQ3CAE/vCNBmDJ69PClhLD7uHKj3hjmX/vlb4FrykaVC+g3+C
jwkD705/jgR0ve0viiTLq0kXD3K+/qrCCVKPdShf4xakZR0+BJCh1FJefyDDqoRZ
HsUr8sng2XR+6Ujcak5MPAFsFHorCk6wghboX1JPALyC6Fn1uB+rw8WGg7cV6PJs
L+tze/zqOnuyTSPIW/w1Rjx4YSvjtZgS080FWhx0hYPmKF93nI5meldP9HrwHz+z
vfcRvQFx2Imk6wG65+hFa9XGQuVf6lZIJeiQM86DkYw9OBdkKbEgBbA+tqZZqOF+
IgNqtbvDcEbh0D97ld5AGXv/PlfPuE7lafjHFdSu7kiEIFoaZzLe7/sHjcjqwFyA
FqNGoVobXQlxt4c3Q4GqC2/btzgz08XUtmOUXxVH1WjG+8duRg6XJOZhrypM8buv
WqazMa9uOLTikb5hd3XQhb7mS/4/iX4o+rcTSltqj0OtdQe78a7PXNHazjpQBn3S
BWiuyEk5ikrv4sXwDo37/u/9My5mBhKvlzVd5NMLdRYOA+FHm8lGCjQUHp2Zf+Ac
NUsLQHt24nzoQ3BYzp9TlYWj/3Gfs+IboyziWhn+dTZ6+fY5hCYyMmww9PKbkBOB
5vfW3psrp15MqBIbtydZ00x1U10bO46uygJhPcsRLPWOpx5wLlLX/f/dADe4ERKF
21BMLQCzwlvnXWN5/E6SYIfcJ7sDEi3FtMryOdqWVOza9JuglKQMAbInThWYKzuo
XzmWZOxh/4Fbxk9SiwuwoAuEbJdFUrWQoa8w3uJKrrWhp8Lmd0fqn5npP+OE4p78
S06GwW9KclF6Nh2qZdMuM/cLKAADHG+rwii2wPNLTzp1xw0w1Jas3b6ZOwjNzzC9
kU5ETnOgibTSvWNA+yfAwv4wHd2ghxdCvgeEBvWHj6dX+puV3jXDnA3vpnAL/NLW
Xk58Rouo7qbARytvYSi2+TQyiBJR667mBjWZ6Z5bPUK9L5K+ygqEvxssdQ20VtTZ
mqHZwgZZVxt+DIIc9otwgTi282BRaa7FX8GuVdlAXj5KqvO/FbZ40flm6Me7ZOKF
zR0dFKwEpOz2OqJAHq9bmbFz8CkSyqLFuBsaBtd3GQfzHzaFjzBwAMwYcAdofQbl
ay1dLmG6nSsH78OqGjFCUgvrieH14eWd8RAQboTLaTiK5MMNzjVFCrP1g/IDnWGz
/rJjbpA3/iq2ijtxFw0AZgp2O3UqPslej2reCOrEq3Dr47/m54McyfPqpG5X4ZOP
SH2ds8P6CLbd+QMAqdWrQmoIkG3ZYXga5YrxhrL9b8Q0LL7f9U5POHdXRXUhxs+p
WFxI/h8zruWS/Z0AbpXajOh/aiSSY+8IQhp94KhHGNx4HEU7axgX8gOszkx8KOdx
JEGXbo5C8IIkvchThJ6JhU9Vull3v6wrygab6IqeleJVRIwtTRSHAiDMlL6mRODe
7ppvOvBhxl9VlZsMHREGHBD5BEocgZsqb5JqoVlyQvxfh336C/i9akw4aNM4IYOt
u6/qW7z2iRkwpsDRpWdTw9SZaPPK90j74+Z+5zUqJQZ3FW0s6bnxVzb3sdMHAhrt
eVVlCX//3FmrqYHtjk5ZuWIRUZDYdLCCmfFqzTQ0AMNLLq0z8tLao6/QcmAftkHy
V8YCKL6pUFzqVunLR2hpyX8545/35TNbSq5tzHiXKvOozSEVANkuw26BDCTq3uH/
Voq4TYB5LAL4aYzVbVuH1mO3iGKbU+28nAjgZhvE2vHrwgx1mYCH2UQAC0JDnH9l
TElkTrmfh+Zc5bdE/01MiE5p+Hem6tD43JJBNFmRpCoCMP1x9aG5TxLODtoPOXOX
lvHmeHWtno6a25/FjGW5+rrdFElyjFIe7zyNSvGh1VZEPAGlNFiJIzjawB+9lRYc
RoDN6mLyJsf68/8TSFDX37VifN1zA7SpE4+/bvEn+g4T8hqBNRspNVzvvqxmv0T2
+62c2SQInoc+jpWwZFqXxOvEJuc3SvmQhUVxlT4zQMEirBPDBHXcH9m26UgiPNI9
rSut1IHRUBjQ2wmEH5PGr7kKBPVtW073iHPUV++KIS2cJx19mTJ7R9U1UaNVLurk
kfYqJtTGUnfNfNtiBEz+AT1qkg5UIDHjmaJFQ2k6wwwQ8owg1i35+Yl8LfFwNiVJ
Uos3+bMPpR0hUOXNr+94QSqNZO1snues+4uHs/LABx53RyOZvCMuYxWfj5O9ImQg
W/7ZJEs4vGYwaIWfOaArGvRB4q7KikpNNzSxOtIK4oHsucgrmPOWaL2balIs/1PE
kSdOlusbNlm3hW7Kav30J6kngz1F5hC1k8h53nAfZv8AFzLV5IwnxXTq3AH+/H/O
DwNzKpgN7kghgyybWuA+HmdxsEdIvJG2i3CA5lIRCFuEHbqcSzimGNeuRHWS6jaZ
MPRQpdV/QESn1NUZxvzMaCo1wUtJJlsVaOe/Vnt1pN8+Uo4H25CJ8NvFmC0KCJ8p
6dTWsNQSvnYAc228s+xi1ihWalhGwBpaEeGJS3thL3tFcFWatnFo5VZlfdwnnRoi
XiJBUjliIzcogEG0Ucv3gMQZe1I8HzPsZqYtPlQHO4sUqaBCIWj8ldFXsv5Hz72G
WxfC33qgpIYawg63spzflE+I2FtuHlqQXsFQ46p8l2/17H3ostrx1aen7vUp8TKS
stJ+1NORPj2snildHFFT2tkBmfHXCdRZ+gMoro6q4eaLA3ctGIrhrfNYT14NJPBE
zwTnd52SAODxOX38WAug9VAmT3kqwmni1ezVjR0vom3dLzpZV22yWDognxEtnDQl
WiB97w3d2RUh1nRCQH0nNk8u/a4i2PaLFfG35OvTlNHRj6s8chRZsAcGgYeUZKNm
zAzydc1x660g1kISAizZ1JE3i7y7qjzwNqZtzwIsX/3f5bfq+StC/geng8kCRWLr
zCkm8uF59K2dzh9o6RVazeIgndRUNIrjqTuN0KK74u5ExwsWu+tNL8z+IkUuzTAQ
ZVoWqTKhcB/mj8zFhhiAO/BlvqQ+lDCjdTrAEoA3+SWTtl6/jytZWj+0OLKFvIzI
irCS/zOek/sQCUMfjuTvxmLGnViuvNzvpWRbvUyqIJiQHltk94but9IwrSqiD0JA
GRejvC5jUT4v/lzswGR8Ftir2SLE9HCXRCvM66P0yfuPyT8WCaxfAYGJrCeAiVpr
wMYiyxYV/VDceArJyBhKK+NeC/BI2Yx8lu6rbUCK12XgSd9mVXlmtzLo6EsDW3a6
cqfEBYib1IOKzdq8CMD4xrK1YWx4Ddzp352nDjo00AoahGBGnK0lSDGrV9jPU6+h
+eXWEbo2xzA8OVI9MCDUdAtR+XFbUxzGbGwgD3B40LrVVy100vazSdOsY7aFCodo
fNTt5JJuj/m2XTpYAO8g9QbTVwOn9uH9viDYejHF26Wbl5l9zhQpwUtdhAyix48R
vBapQ8B3TPQNrAWY9TQjj2zZO2hZ8QuoVmaCg/mN82HWt6mr9dQwa+iqwBKDrBhF
U+khFIwedTE5vI1MsRcIcuEPz+ISgJqD4Whgla6jwfamWKSTUs8kpZYCxj2zMeyr
0d7/89MuZwbOXq6CIGk8DJD8U0+y9rPOgLFZhfMOQRInqqHYX3aTb5PFJ9IgVJ79
3Ro1XqkeN2rilNRYWuYrbh69JahvrlMfueNnCvPEEP/fiorypP1bHx60hwqaP7K0
LSwgZGlie3ZMa8PB5s0IZQLEwj8ynQs9xMCyrAbrEeSZNRCz3Y+8SwLr9vXfVJlT
oGx3HpucqeATvwK4gTdtlHO9rmOs8PQAGz4v3yi7v7xlseU4uuZFD7jooJl+7Oun
o/KGs8LEIb4U2Cy+ksv7etE7ZEjMdWe0YeaUrPTg8ZBJmButGeh8WNf4yxLcQZ8U
5r/dH7XyrK9MJtDIwAzCtIFFOCdOf6H+TX6VSBAqhPs33Tc13wix6ZeHpNWd9qCs
GoGuni7OZ1vKosYYmVqK6F0TXv3j1TzM4Xlq+pYN0IrMM7WTtbVRi+MC3oS3AMud
JBbcCnJvWmaQjAboS4m0EHGYtzWaeceZHO2a4iP2XqSup7w5EhlxVEHkWjtWGwin
vwWacMKzP8IFUcT3pP2Y9TkU7jZnPtrmdXmIDyHVvqWo3W+TdgBBWNmRE5sGbxP+
BKNOgyz5UMvJlmYlzPAhnymqTeFOs5m3mvvw+i7uSHzihIu8ccZEK4t8eBJ90gU3
+Mdv7eMHTpmnrREPgdGJu+n3MhbZruJ1yDzwHfwxNS8yqYWGOj4UYUX5B8S04TVS
rmszUqXYOEMlrrqSmezFpdyg9PejbeR9aVBjZOfso+QR3hPasA/h9yoqiuawPjm9
X94y+vEG++BFEFtZm+Z3sN1GBYAKWvto0omf9Nsmp0oxBTENiBJQPUekpKUy11PD
BSHtcwUzl3lSBBLH5R5ZnrTsH9usHp8GA3YLFGfWYRebGzmmFORKl2bOkriMAA5s
aXb83eE3v9NL78I+JxBaZs2g0HUD1GCEHuZyqgp5zm+uqaGxqu6NL3OZwqWEQRgC
jZSq556m3SF7gSVx9Y0FOkIws8JXK0esU/0JCw2glwSvPDpwGhSboVSFB+7cAW5T
angcNvBwBed/Wj8oe2dTv30vSUh+Cm+VhdPb6AXLtTUA+J6emvpfuKhu6I6fypGz
j4p37+ad357BfmZVq+MYUcej5TyeVFQ/mK4juBTMz4EyiQtRc3T9937Cjwndtgu3
A+4PcIvemxsTQXj3k8A/BHojWFWB+rvMglQLWh001Kf+ENsVxt5Q77WQKlVeuHCi
1MJXrtQV6vN+i4+hiFlGV/JuFGmMXt1tS6Nr5Q7Il4cPzZ/KsU4UAYfcAb7Qa+Gv
QToD/gtv+zsdFLTvMGZwBsXsGj+85f6iU2IPJn2pat+BmrY4AfHvsZVhvANn3W1K
qJkyfj9o13JhlOXIAg3tmtKk+ua1qzt7lhuCi0yaJEecl9ceh3lkFkqGPmQFk7nS
yVQqBANvs5+uKNjIZaptldfj9z7khfNp6GQ7jKUEiiYP8HaWziW69jyGect8FB8m
z1YKglP7JZLgwkdQQyQiLbTQOjW4I9DZsBXkg1JvIz+QdDDXD3s/QxFmgWJONUd4
8WKmBN1Zqp4YsV5/W1BecqgwY8i8NMGGDMOA/3M3EHdSK9CIBCF2+kI6NjDa7nVu
rXHexTQgGcbvgDdXcENSNPByApr5iu0lOw3ZvbvYYONl2Re7hdyVQh6XicV9BvXQ
Q3Yt5NqCyZ3nrUpXdh1AQVVPzpuwDED9xp3W4HwCTEi1osx9ndyuM/rxz2JL2hjX
W6fLKQI6UVhWa4UKT0KMpegU1VYkJgEd4ZfFBJUMGV2vMS/2tEOQA4dF6LJ7LATc
BJQ4m2xDEIJeGzfbIwyZLZuzJ0rFvhn0JX0Fw5gR/LOIeI6D0BU/wXtur0vmQ65I
Rdp1p68PdqyydNJYlboX356nqt8QQu7VxAmjFe17JyGshne4q/0oBc2A5sFyhsuw
EbyLxqElXzip0jgGS+tzm3XpseyKRgZkCz/cZDNR8nnd9K8qKh4fU44RVObk2eEx
NiOkfeZWqEJ2bxNT6/rdUPGei/JJpb1arlaatm3+xlevkHuUvB0sGupyeH7fJnPp
4RnCnirdINujVGLlXE3Pp0gX3+mAXvJGezGYCRNYfHHSyM1z9jqc5k1vCwQtFENs
dvczN+mqVwgpnhvsN13R6HG9egU+C2I+T40rqiBL0AjeA4lNYFDLkVjhbw3fyF90
3voO23D0xl7O1Wp8ZnwiqpxV2FUJuEaj8nWe/EItaACg+gCewUtkZp1fWBZfgq2E
nz8PmnScN/73/gIn5hRtMGDLLKtI3f+WeoPhbXGO770q6jj6AWmRAHFe/tWmMh4a
yNjso9rlVunU+qsepu8zrHUE0dzgRqGm9ZAHR97SjTbtkWrj8i5qrR33miApvrKo
oQq4evYhTT+303qjfB2qRN3BR7VyxthJtMIYWNqCOnAnOZQB6FMRBZdbFFjIir0w
YlniOwRWuirV+r5lz2ZU8dOTkPT4/ouLsvY/cnEPWfv0gPXFOGwMHSHL7D4DFcgW
0ffkHBiYPwhzcNCweH8+61w1n2LeTrA9fXpDUU8zvAKSp6STujPYGJ0wSNF7CwR5
nWWbXx0GkPO24osDrySHI/m7h1FzGdHZb1a5C6UYNwJMIjhWlHoFGd+YasV/dl9X
vKthsGw7RE0T0L+a/yo2INdyI/RofSJ3PAstGGmhCTxB3GtSQZT3QPU9AniCNyjS
ybBfjI2dV432ejVORry1FBtBJwDa+ceUVDoecEKPKasyDz9FJOmsaSVNTbRrGZEj
rpXh1P7rUenCSE/OupLr5HJ6yQlWELFePn8+jeLOj3TpKJc7/blmmbANJHwY18dR
ssgpxCoYnQd8rfbCR4yQ+iRLln9PxL6PxqUjeM8Cl4CG8DUuPzYdrADhQkeRCikh
wOA0EhgaGNNRzzveiDb+wQLdOSYJlivNPMW/o+DcavzCDmRv95hDVF/PXXCRFW9K
UpR5RLE8Qh1ikidnSZ20DTQ+08j7DpO3ceFzXJ+0lLSYglzb2gqlgkd19IegoLpZ
htmwdeSqnShvSybb4KoNPvZraSNtnqYYImA5Qt1eYssbnnNck9sDH0NvziLsiIiN
qSx8vTzfJC8OK1tKgUelR+DwvVkkvC9owJ0s/Hs//ZLB+CRnB73hZOaQCrQQ7IMv
5iudZDXmScrVAwWzY2gF7YrDPkMdlOJwnLlPgj4B5pX6DSGVSG3V95ZLkiQ/U/07
rbQbs/romsWaRp3TxYT+Rr9SyTFTFSMjNunY165K2Z8i46PR3JqfKaXYU/qMUseC
pN2CnAR4vO9OMFER4pXRj65Nuk2ZuobD0c02jUDglX3BBfWNFa0KfFHwdKmaRGUc
QS93w3Me+b7zi/Flb+sMW8S3RZQnaUkaaQ1113Q9NdJSUbN8Ku2SMkibJ2AWgpvH
LUacqIBGjsgmi9XCQWo9UGhYuqHKV28tv8ZV0XpM71sJ0TzdHXXdJY7N9mWfBFsg
5pjFmyGDFQ/8jhdW2N6kpAMbJpqh20Z+8AwfcReiahvWuAFnNth/XmmtKaHgb8DK
Y9iDAwLbm2Cq5f1wsx1UXsnwhScXpdXSuSsu50DWIWvqSyqFJUJSA+/WJEqEdjV5
wetoT/Si75tqU17GFFL73Pzlw5sh7VqFN8uISuDduAV2+/GLLJ7hDLUihqJv6jGC
BF45+bxApvmFiqNhV+d5kI6QX0P+Ptpx3Cu59eb+PXkB1+B0witmZ8c/AGRcl6+5
EdwbntCLSdsJNnykNZ6V//wS9lgfyEXddwfvYZK2gNQMbqhilh5Fri2ScaJS136A
le/iX18kEU9VkSfebS6UUn3B/pqievh4JPIBuiD9JAtCSXxipFKh14JtsqntPiCG
Y6DUa5tpBZNLBECvLatA0fYHnF3YoTWqWLWrJ/PqSIizLoHuhVeg9iFsVT/4DKiv
rAe2JdTiDXEEw+Iuhj2TRMONXInE5HH2nBRKDjfB6b4hnGHnyB2v4WopGFXfObPN
9k6lX6rHJ/nxDX3VH3oxj6iPDekPfGGE5QF0iASUFWQuUO0M0sZI774tD6PeBGwB
7LAaCgDY10/DFRxLfVfvxWhR+y966rQ3hnvwt3Oo6biWD6mReh30p/jRWy+PTLnC
75kj5y6Uyz6m4rlf2Ad1khazPXSC0eEJcrqNbHkc2tE2QOMLoO/wXlcYw5wCJNoR
EQWTXx7iECpsvuqQS7qs00ExOiNkBg5Eg4qrOaGhZ0GMm0EBhIrylwhwdhLmivfw
hhN/1SXO0q2/7h255GXP35S1vOS5PklF4yrdR67O0emHwp2CcymLNt1k1SF/wJMZ
4aigtiiCblHPRSK6tmF/S1MexYFWZk4B7i4DV9ggDx8ZADEHrQGkcH7eIKRgxc63
WyglTUnAwBZhwoHl13uzciYiF6E+SxcXbFYhVmeKYHqIt2UK4pX8OOZ6f3kgHw+4
1Y+UO4aEuc4VIrGkjL37BBdYaJfSx6QvEtdv8ZHeeW8HEXQwjCfsskyyknzefFl6
E3lSiLT8EvII1PUe3x4JF5nuYFRcpJSgd4can9QIeGqqqS+A8HzF1gX0b3t0IXGe
v8FCj9G0/63vWUVRgL+JYL0/Hve7SPEK8tVLRcVIqywtlGmNLeOA32zKQzOS7OGl
OxofMYxqekBY7iVL/NBmPkd5wfOVxKBtWQzjRFt8Lwl/57plVCUgh7BY5HntcXhy
VMialoh3BRv6ax2Mfk4+MfHFZVmBL5rQRCOyifsgI02xCQMvrqISMiW3lnWU41SV
VvaHR24getXIh/QTIKxNG2rJeVt4pnz1f9mvsnXR3relVya5UMUvoU/Rjho76MUt
xbvCo5TAPQHGshPghNAPpvFnp80Vtew37k7ev+Qc7MOaKlQsW7CbLqREoT6Y3F/L
YWat05MvcacrZ+WrOWwnN1knU/wz4D6sFDHcytIYs4oRS3Fd7RrbxIKnm1ERjXlB
jNGxLcho3Ioy175S9TAuO5xxIQdQ+TXe0Gfj8E8VRDOoVY+/0hHGXE+y5dMb9RjV
a6z/Ut4XqHg7D2iEIEkChKz/ZdT/sxuDxYNxyA00HxG+StRzGlOMuvM5J4PA6yhv
xxEPEpDy2zgz67L1I0lar8ylE7PsItnUPLp8Y6CsDouTW0UzKrE77/WSCKWoLxd7
GzczrqrbLW6crzJDOtFRzVSHEadpqWmFwVewuPX6eT4g2M0vJEdQGrf7bGih0iJ7
GPzBgeNru2OKq967iR6R4e4m+4Ug2D1Gufx9QaNaGfd1/BEmvtDzWEAEvULVYm24
/kjoBdFVpNTepCLJwGFBMWPXQBEijCGHJ4qDcUADV1vWsj2xj3L2Ywqj9b1EdpX8
16aPW3aTURi5H8lLr0vuJJ42vNR7pQTYcTFDmbbZE5C47pl21al/+HY2vQ7/YwyT
vziiMsPF85gPd5W7Gzztaohmk8A/OSdlEit1SwgWnUbkjHThx8J6fYFoUBL66LlB
BcqdKxGDkDOCZdbSeTBMSJiwkiFEJN9NZlBb9THBJ+624WrTajvlOg6HXRvx9rub
3pGGTkEoe9/Ca+kjJTqjDl7Vyk8bv5mpHpWPMeSeYc0P7AMKa7azRJ/4QRnN/pcj
IcsHCZjlmLHi9gw263uXHx77d3NHoxUKwjspNLvsz+v9H6ohstashFd35wYuQqBC
mHSgsA+AhuOTi86K6CqzyImayGh3D7k2QKcAejfc4R+k4DTEaTEmN/G6mS5kP4Z0
lorXZn1AGbMMe8mTT/e+KfzMUWssa04vOoW/023Dsp8Y6gg3zJmWtE+fZJYMZn/5
qhLotd/ychG/Z6hiBLllmePviIGZhLQU56FoYjqa/kk4zhj0jMo0wffcSOJQhWaG
ZW8O76tntt/o0fFYVHbILGb6YfUgYWdTPCT+CADrfnBlnDbuGH+GyJagci6XXy/F
dwq/DoGqNL/20MpmgQKzqneOjn1qhkZSUcBybXWSibj05rIRyEwLcECAgmScdeir
DrmrzjgV4oZIqV3A0tUuiKZTkcF/QjX/UTw4RHKhk9AXA2yBGWo8m5iEO5rW2yOT
iaduuFZH95uRLb49EvdRYhHovA00EBsdB4/EsnnnU11PHybcUHwUxtnIGnw8KyVe
21X1rZwAySogBqX0O0Wa7Ccc+EFD+5JyRXCDr9sp2+MEBbKJEq90AVED8MxBmcOj
TvP9yQ+nT8AsbMRn6gy5yW9uwEsVmD9refu585HqAfbiUo7v75HKh1za6nOSBLhP
awHplcwZExsAoUs1LRnKmCEbTsan4kZRpPbM6jUd9oYetWda8DLADJUP5dilOYZs
E0hTcVwXgrsohmgGqakglNL6HvS6xVFgIP1F4Cr20SKEP2v7J/aNqRSnNMlve1u4
dv4LaKNxQ0fLb6DBUS93ehrcaYwiDdn5ojHsmufOYfAwkM3nhEgFMbYosBIzrGw9
AOxtjRr5N+XhtJDql2KcxuXEe3ZOdPT7mLkudykcXRJFHimX5FyCnDhxqQKaHb1c
Z8P6efOyGeeaZzI/JzzWgIZQKcvBrgQrIsdu4k8SI7ToTqDnanOFJblKilAuw5IZ
Xpq/DStdoBlFdObGOv1UgBJjoWGVJng1qTh9afLzz83boAWj7LzhmRMLzJyeARY2
SNiy+kZbNtbjsyNPtn8cQbE+Hrn+sSxIV7LSvlnQ4F/326L44PXPfrmXEpvm5G0U
ZwozJr8RiQ0P89eZlExXqSy7GHlFDyGWubBGCeAy9ad1iTfd5We0V4zAI76nezJp
YKMEXQ4u220HyB1Ap4zY8UeLkTtLVUyfg77IluS+SLRkfvg9622P2RvglP2k1hq4
w0yKkGbMtk5dx8WDYLvMl8r027nkxGvtiN0nZUeM+yf+umXN89ZEYHg27G5+hkcG
yPKKDw0ddKwbgC9Ma2cKjXgYRXz1a6k50XHOgfKckDP8QF0oEZ7CC7P8trOPuMV0
T24f7+xxDoJ94VPl2l4tgGESsxRnvsX20W3RMWyTaFpPCuj0EoIzrjK1inBFEG/j
1IdGY2lGd89cXu1p9Mp8Yfb6e6ORrL5FTzaQn9ZWMBSMx0BZZZyxgUedhF5JfyFh
6ABullBdq9DED/FF91aLYeakrp3CBroFT/wCmDMNvB67TyFAXT5SsuxljvjH3Whx
EjtgjgvW0fS/XyBtqwHl4CV7IbI0BbKlVj6QaIIrUOEl0Y6YynfhkBWL56hQMeKO
bAYQaL4Ctj5spXCb1e1m/+dVanY7/a8Ps0wQmtzhFLxUgeL21QIRAYRGN5sW4HAH
IK+SlDyzZ+6fzSc6fJKTvZhNPH+iN72HwoS5cFapWSBPQpRTd18H2MTPkFEpCTB9
3qB1utJlc6CgPQ9lEkrL9O9T6p6pyIYgiM8osAFXoiQPD8TkI9H4rTNitcvn7sQ4
EZS5jROIGihWeDltgdrCCt7nsIu9VECnrvVGJFFV7bFhaLeuzDUOwM/dtXRS58Uf
r2vbBgM3Mn2SOK5m27IkxQH74n6yoaqWZjL99q9jaF3Sd8zUPpyYJhcUfuPi9Ec4
93Ab4g42SlJyraIZ7ppNocOBPR2vHFbsp3EXcEHQjIBZPnPb2wrPFiYk4AJUHYHQ
8Sj/lT241H5teYFNJECri0zuz8hzVwD0d/ZFX93Hc9Zt6exgACMGQglkM5FSl6AZ
TTPxYfCBv/Pb0BGYCeuE4LvVwXXzdXtD339T4KeWJZ72zceGbinmr41RkI9Xw4x5
tLXRYOHqStdesAyFSD9bFarddy7wU3se6uylpJBnjiHV/cbx/amNCY/MSxPKHU+F
CMQm359OnjD6OOJu97vdM60ihnYBc2VWhuU2bTn/6mYzyg/+zk8mLQZm/gaMwNx0
rA0SnKs+wbHiS55hffYU3CcMYWZD65aO11dJB4SydTexg6Q/sNCJm0OGFkt0qkEE
/PvxXtDPTjPaUe5gd09E/aBzo420PC3V9245llLdA9MhmIf8gReR7zdkG2qYcbcR
2IyEcZl7FUpa0NQj0RiS3kkM1R1s5GW0lcUGOnRIn9yJUJGvPUk7wK7smzuWXg+Z
wVv2joJNb7McaMLVDa8L1Ragz8StRWA37BHEgOfGMiLmg4Ru8Ac5bJB/S3ntSPhQ
OEVN9W+3hYrZuPA+gTRwQcXyEFKpc7N3/ji99RM30V5OU0hqU2dIpNaw0P+DlQAp
NK2JzYxsBdl/GeN6Ypih/RYayqpCFfQRjUqoPlCcDHr7+wQNRAapSXac8mO6235I
wHnLIEeI33xwOCVIUDP4rK5EHP7sY/TwZ/ncXeZPjBxLOF3UYZfQmJgvqrKuoCZV
jAoz1M6tmDaUETVna6fIC09F1/ojtRZ436WgJEu7l8FsOBpJYCqzn+D1WovVYwAg
gskgj0fzgZp4sIqmRN0ECALe7xMka1JvoSDtY8wDOMnPUQd2zLkM0hPmqg1kPkGt
zw85IRIm+D9HWZqyZDIbiLwJ+dplH+mLu66flWITN6/K5dQNzFyVUMQBH9wXYg8b
hV0VXowGsYyrvk8NNmaihlniJQfBkIglnXXra6k9j6NWBCl8UUOlNsWILkR1B2tl
aaRm8CnNzWjALNPzpw1CWqQMUHKgWBcUNOXLvzCGPxZLUca6PvVwZCsdPQWomyr+
4OtzhG7Egsv8+A1qG1oAJtzIoRr+5pYLCihdDSIIxt1RE+/p0BsxQfNyrLhacTDy
RE49ZA8ipdl2n/jd5LEYvzol20b5d3xy/L2aiPOKM/u6zM0E/NYagSVgAas2n0En
ganq3NZ1JnEavEL8fpVg1M8c8eqA8hZTb2EfvW+LhKY2XwA5H26PEjRwPIkgQRN6
msRpYvTDLMFUzPx2GlsVlwv+i256HRAZb+5HBI4anFlxnix1xyLJt7KEHYohvUW5
dzvB/y3BQDQey1fBKT4UGHfbUa9ZgYjZoZhMfTnwi0kFHawMMvmINxVv0rX/mIsH
LfZOkxpi02Q3JtWCyhSzow3oUWw4mVA5Vni8KR5UvfsfakQcfNZNlED0lEMc2Q82
IbdXat7rwjee9wqLyr6Rb43mbIxjnexJGwAiwqMOYXRAc62SVNYOjs/Vy8HsgY52
hOASuBS6tTOf80tAcjTmWv7GYbxfRz8MD1Up6zkDk4OIMiYiJ8Ui7LJPVTmFNhc+
LxlFwa0CNTN/0EmMtsnxTsocpiPzdvnsI24mpo7UYJQdsJtcyCwleyO84Z+FDner
QCBdpAxxctdzHQHqI7Y4kwbDSP8Jea246zPvouuXlaNfxKH8Fv/eRfAVW+uv2Atw
WFuHZ6VvnEmgfoRSK+7QWiPBP1WuRENyZcDaIIKRJU8Nlnpm/oszOw++BDi3qB5u
wa7D6jnOexhEsD1+9j9ufSpHj+lIhIPLLQOXF8PVlG/Pa8XwJzIlXoWOEamDrE1f
9lMKxdbgg/Dassoe70euSgKQPyoti5tfN6T+quxXNHS/Hm9/c4OwqAVxrHNEkzRx
fRI4c90jyzrzC5gpucq5bHLre1RiOzOUcKV622TIarMLk0vyBnRfjbMLgG0eF4Hu
WhAVaAi3b1+niOfPNt0xyshj4MAX5BcHT6+nADcrpz9V/n5uUkoIFCOEGUd66gFc
xf6cPAYn/cSgpFgAb2Ce3xy/RkgHJnXMV/Kmsuz0gGgYZQE98Jb7wgngVxe+tSjd
aFe7me7AzRXEcXWL1skQFmMJol42FwF4EGVro91sWb4r+FzlWB0o7obmcLWcP5Ts
D7uBf+WYnjMws2g0upSpWn3NM5HwhllnV5lu7CozCNF+Sk8HEDVboHMgREMv9v03
4DXWDMaInbyH/X66W8RyneDaBkpSj9VqajRhvsN2ohRMnR2zsjTnr4CbJ1JileAD
5JhpHhFKww8WzUDhmNfHsMJcbOpSdElb5t0r3NhuJ9GN4X57+WUl84vhmcOCbfqt
WOX6qZvBkzry+7PbC+GzQoZIfQxUB1TBuAvz6UxkvaYq2dVTSUp813USbGyf65cy
VkVs1RuzBQvdg6j1/jwAeawrl0u5dFk2qRBFkO/jb4VZI+YFOUh6Wn+MJFKn8h8I
v+3m36CnMJkOLqocam2sf0Dpf2tRXD6f70PIKwkCqv876fSY16dW/ll2pGLfcBVv
WEiS8QXL1cfXGtzU7pXwr9MQgjrM7crmXYXc9ZPJgWQnNx16aKGjvnCI5BblXKzt
rLLJEC3zdsQ0HLcSdZb72ErJD3aIydauQDSLFDqShTHey/PaoSoyUEIyEtwv76J+
Bgsi4lxKYA7CT4WaCn/BEFxo6IXQpvbDSpEiXVFEWqpTxjPIF98k1GHVsj/ErFH4
dOflbSHcJB3XbZ2B50xEC2DvouEssiuADcwO7HCCeSSUq3oae77rLEEcaLoSYuqN
xADSHetdocOkPqkMoNRSrTvF28JPJauJvSLuvR6aTHmS0YAbesVRRrjcyTXmUy1v
4ImYLyyS/dimGJHkQtQ6urqOjFyOmToQPBu7ONwfGdParu8i70AmzPkkW2qRUaIS
fPmenFzlJFc0tBU6mUAbu1muHpGjfqwiJh2I/LBFWO4IDkMdfljkeTzPZnKw/uAv
Q3CEL6v1c13jTk9D80aXEaUWZBtNxF+aBAYjPCPXT19yNjCuWQHCLSufyB/z02WF
yZ75WhniMBffSQmsXdyRSFaUd3Km8XiICzCathP/OK0rtsHTbzk4JMLJvkmorZqK
YBZlUke203VY+ZUWmRvmW3DoOb4gw/OqBZM8EeASD7CBfjicbnj0DSr4+8CiLSmM
HrfMKDdbraAVqGP1BMC13EgrTdVWghx/ekmB25cWiGAnIMeDa5JmBSX1fmltK1rv
Khlwkv4rmE23sPk+BJkHuO224ZUrHKJbGl9xED2ZLMSNqw3yJO/4rhQuEP1AIVeh
Spg+DqTg51FQvmO96Oe6a3CjpFxV3QvRy0nEyJByWV4SNGCP3yJT8SeYE/BTMtYI
rd8CY+G9UKijUlk573O4jrfEYY9vLQle+XCh1gpM9OujBXh0Rh5B7/9dQBXaP97c
E9QS2lCOWRPaGFUMofe1IQK8DHNnYVSMot2Ctp/FvHL9DNOGhlGQ9wopeXZenR8G
3gbI3DieCRO3EKr/enVYs1knRukBDyt55JtcSd+NhafkLytAh7seuqdpL3hmZhyn
wud24Al5RtKgHtJ1UcWQ+Fl9cXwjOftCKI56O4uVUAvWR7oIu1SepHeEGFkreoeH
2EtOpQF8NFYaaShkee5/NFpwU13Nf3Wtq1aFMcUfR0QrdbMdyo8jgYfrZN2u39DL
ITV8k4P9Ex8ORbL5oAuuCah1GDstFawtMLFwJX7Cg2EDM6UWfkX8fcTQ2FExb+AF
xANRyNsUpKppN/eePNJyeozypNUlRIDrsgmsQJhk9rfUMGq2+f9mMCvCE3srJ9jS
5nAAx7PXVwkpCKkB+UCV+6WKnae73TqFNvYD44GxP0xNe33kvPjcpxB0/W+NFqI4
HHeUFEwhmI2twTG00sUwJ9ygmvLWosPxCvGwgCeqgynKyFNPiKlUho+w0tpEGXps
ovp2GJkDTfc80m4r4F00AZhdNG2TuQGiEjIJ1w4pED9k5Na9Y9Y4Erlhxruks3Wf
vrOh3IflPlxRnjc/fNoDiYqdlm2kR2m0zwWnGo+rrSJAIDl72hx15iWlACz4P6Vh
TaNfoUaufbARqtepOENLApjy8rXc1NBN5dM4gX9eXjo62UtxkriqD3MQm/YVIMvL
AMQ3u6q7qs/miYlfyxxHkt5kLdgLRO0ShxutX0PlgwQJ/oaiDBOklInkeAD+AxQS
ggqq09WK6j9cbHHmyjFNPHzc/QnchYflVDvFEpNGPtgtpON/zopGNbAGkL4w6JJb
bx1Qa4zjV+0ZEz02a9PZbJe+EyRHsfWxWtXLP61GQLfRqNba9Ml9kiiEUsfoZYK8
RgYIR1HEcrXX1xd6pOAw/LcMwCtHqF5lAOhiiFSmmzXp5154UiBWK1CdZyWOno1B
BPxm1HaUPBVACWrQpGsOUaKdtB5n1DNny2hONT0RFegn7ThUodmcFinRkQAMvoZZ
GC7DQe+O2Ppz7zYQIl+0l/ZxxLAf4TTuwS+Om8S0c6NyEEyyWXbfrnigpKNi7IHY
xxGwa6cjlKkaLxZ/vOkfrrAd2nnNXCh7ARzisG5hw3CNJ8K97RFWHrNh/mkIAoMq
BGKfX0Aksz9+MC1T2jGxphlevOe48ILO4zM6mEp3XDjTHT5ZggLfWtDh7402/jan
L1FSbJSohvFrQRtm6WKPm8n3JA/Pmmh7AtvXRgF26ohJ77m+GkDn3qOtHLjOusY8
jDDzQjilKc4B7lEwNNoLToLcpqy4ZMrlGHPrO54QXwVRek+KhByvuBqofztWPPne
6evx4sV9ETeQNCUbti/V/AIcZhm+baHZoGpceKbv89dYIuJtKnBYGcrlQGT32tJY
LNv3XkJgecO0sMQ3pAZgAcUFD5PWZ9vEr4iORsIJWyJEXFbZWVqJbnXWAmQMnDd5
C/UZ8DPj6xWnri2MZwUg16axF4Ra5j9LHmjalp1U6GbOI3d0FoafMM4W+G9LjZJi
J11QRGFjf/iRgy4svOf3ZvXaJaaxljY79bET6h4OmsZhvg9zXHGasqzAoHuCQXEd
iWPVgem6OT0ePl7PSv72wURi7OBPg5SWXEkcp+P7uDsizXQ7HYnL8jt33u+yN2zd
fzgOYGBjTiTyEl5hf1O7Tv0/6/HSwzjeum7dGdekGmL5mE86L6EHaaP0bW0Zh3VJ
FxGG9ggWyeogxLgCaexXh4ZhJo9lvdGJdlCKvksPc3KdE7DjGAiNtBW61YRn5dYK
yKFKyepSUAZTLXUbLdaWwGzfTXDbxOKtyGn05ZtzigIuoG3pDMEJVoq5y+1yvLTd
QVweYsckcyMtDQQJl6Uuo7vEUj3rr9s4nksBEEaLna/RKar5RfYR6RK0+oPFOr/v
OMQEXv0k1YgWbvfLpH4e0uW73rB9UEzc/eb3vwGXEK700TtJMwUSz1Tuqh9byTzk
pEd2grlsMmvQtz8JL3Sb1+PO+ydmvPC8FAOf+AlYmTrQFOkM91eK6h5i9PqyUnDy
rxEA6FyQ7yIn/FWjWdUuNm1NzL9jAWeLo/qjAGeEvpgOsCmVm1y7D0YRDDnB9Iy7
8DfWss2xAPla9UUjOEHnICj2zCVQO9TVRWgjEwSj7ayt5JySm92TJU4IqhT7U4NQ
e8xIKdcUXpoFPSq5Yw+9tum9UkaQ28QxRR76mLIoupEPE8DxRKAD8V+4Xvci+eyi
UZ7SxQPp90br5kHfY+jStCdcHeaneL6izgHgEMVcG8fZ8r1mgtOzU3w4O0ff+6kY
p1o7Q2NkEqexQidNzlaIfhvKsDDlLdaNJ3FyJ+1YyRVm6E6i9VEtTyGx+p5bQKGD
/Uyp3BTeLEOQGK2KGAfChBHnhf5ReHLUyytOXZ8ve49Ism57SOIrZ2MSfwsuM+SL
wYu0ZqiwufhNfo73drvd/5u4hffFEdQX544/Kae/WZUNB+R9kuo2WdzbDvxALBaE
W5/mVWrtHAinNhMCD0xcXzZV8XS85v6eUqFjYFXvqr+4rYW/hAsX4iU/nUy2PEcz
Dy+8FBS8YPW65i2yjwpTUz8QXzn3kNxtux58GyipcVbctsd2fUug5k5D1eClU9Kz
Lflg07U8mvGgefyqz/AQ3alTIgTN5/dk3oLozyn/BqErk+fwcYm+EjAaQv9rJvoH
hGMYGKM+qLtuEbat3j07fgog5bglbO33k1or54ehXFbqpIfOye0gbcnoONpq/heS
9BdIaDpVN5iYvT1j2q7SXp0WpBdFJS32srZsCob8ZJXrdYxkHP/NAxBxkusVGx+4
CgLUw4WPMB2pBNTfpj33pCxH7NBFrX2hZ8vg3wN08VRwVz4ZYUypKo+HIp4QDra/
oAztGHi0BVFnicSxvIYi5EjkwCxVMr0jAQZqlPYlY30CmUJVGinJEHQhrAieq4VW
tClqc3mfzOWedqfZzcBhdyx7UFLcj5qff2if94YTL0WAFq8s4eqz6DusPcma27YJ
3T/o90pGk/BunBpbgbsHpyH+Cmroa39RzILRPkDhiqNH4fXMEUgHKpmzA0aMuLkX
kGFssk6Z27UVL0gXbvz/qWDuCKN7R3db38nW9/j1/INtZ9GPzZlwd2sSIwZcGraw
xLxuWvatYx0qWEbDzNdMg0P70BEZHZRyVFZVEmAzvqKrt2mHb4E+gCA+QFn89YLI
AZaVBTgKUqBRLVGsqKLcRZVllX4MOHbwpxlxzAKlDoUoTPqESGOcK0eyTyHOqdVl
1KH4mcXbrEKUT/WAZ2en8M8t8jWwZOL8J+34oz43xYANjSStPcGrXuCSvLdh/6BI
9vKjxDFPRNaCmK7hIrW1zOrgIXr7aU+tzGt1Bj3VYvV9SqIBZBlAx8ocF9zH9Dvg
RmL/LAzQedChbm/1aL6AMzn+yoVLKtyI2lkBGU6xJ4uP4JUDAIbAKW/JNriAVGFc
yRRpGYJ+dWFZIlTd0g6DZTZDoTRVz6Imv8t5O6ZA05l6yUfPwS2w6kKn+cy/Wnya
hwM5Ol80ILZgl+RLrXiNBbvGHysKzTEn7ovaSqnDsmQZvFkcn4Tt0NycoQpBIddA
nK9q+SwVLyqB8yEJwtoEkXCTzypYX1XstpXi3vjeBQ0N6go+EAASoDhgzvmTNPxV
T0UZkPrp1nzcLeRTgvIrfMtDT6/SRnofhzFfidaT5+CFORBODrChXbo5RfkDWlIL
xNAGiC1eKwqXG3vVTE3UBOk9bUJCetLt+xRuA4X0AIJ/42TsTK0ssFEwcx3fJPPC
yZSou7wqMO6mMKccHpPr85gfW+nRY9A27JzCDAYRoSs8lhDGjLYsT4Pc+0vZ1ieR
Cg4LnT7gCEL5m81Zhi0D9ds13ozbRgXM1l84zh8GBMuL1v3R6SlZ5Awfk9dL5PfE
ysF/SEHdEmV8cSwJBnrj6oVNdVRMqwiXQyHZKCezwUhEJup/bGrB1ds79DoKgbLI
33giVwajJ9PwuGiDY9w/poKtGDBoUyziu2eIrQ6A6UxtCikVc6Aw05GREsmPl3xa
Q8LBvB7Qx1Jj/1oebCZw0wz9OlBe6zrs+Bcgr5GN1ro1uQ34TqTTyufq62Lo/bPv
fMb6O23V+HuhM2Z+K3UzFOEOs1Fm7ndgXvHecni6HuAIEDqdfYbiFBTU2x9O2f/9
pCf9TLamlOIxMeuSir4Z9aj5tBI262ofqOqAYgQNZQmBYr0h8Zb8EpqZJbwzIYxE
IGqF2eDi2YExTMqDeTrSxbRS0xIy30Je5FzgOV7khFqNw5BCd3x82Xk5QcgcHfLC
pm8Zmyxn04hneSFwgE2bxUdtZtm7eN9HoFlnEDcJzGHEcY0TS7eSGFG1Nv5DJ2vl
nKZ8JFdQsW8j/sNPLfBjJpgijS7ZyB3cGSg8ylWSa3Qjey29Rx7LKQqw2GrAt5Aa
zaqAKSylRcY4QR1tdbfIC3HS2+WdR1midiSpgkEcamhPRzkAj0Z4wDC6qiTRu6hf
o764qMy5hTDnxNbP8BwdMBFIsx2M5AXDLRu4MiJW7/TVNiwtRt1ep0J69b/1H/rv
nbb6+6lFFDnHs854g/t/6Y0gxC+Yqfb8osekl6WbG+kpUGgYeOTlrcNYPdqPs142
rJEmn5TF2WjQwaTVxzdChmRGc4mvxHUOvrlPEWoPvUl88NgnBPyJ4NU9oa7u+9V/
7z8Nzz8qRq92ouVi7XjT9abLFSlKrlgfKgm5S5E0aPLZeUjSaej8RZtyYsB/J2Yj
EgoLCA1yXy5hFZGvJ6+L8YLsEtGyu6uPEn1M2WWyt5Iq6dX5dGoldc0+7+nLe5ru
1zODeHvIX8VVCjMzvqboI6dzEa/3dpjkZzeHVpQdiwJ89m24OO0TBFjZrT9VN34Y
PQaeE8lSeOaAcMPwurWuw5qzY2N+cMkbPD1vrkHXSe97nxviQNoyjJ8SqB3Z48WP
u0VgRDzKmgpmJJOSbGdflDAYFww0+A4YT3BhMjmPUHH5uQ0K+fK66N0naEEqof0z
+vNXqDzSHd0mRVdHRs1vY5aDIezw+Xqvrd7CJ6sVisNSaqP9uKYAT3TlExww9DD5
IETK/3suUtg40/U+7hVH6zumoXRA5+goE5YNwsQGYOzLnj7Vf6DXnfS2i7FKSJ+y
TZCPsTE7/V6Qnc9ghmPyL2WTNT7ob2dtVvZW3ltiOT/NCUWU4eLQ4sls5MsdACyk
DykfCRg1yDnYLh4b1xL1xUcsXVQLJXJatB9QJhq0g5cyF79AuAfI32TRit4WzQxN
9p9ePHzSP7bvAjtj2TLSZDhnaQ0AMvNanpyNmSqIL26C0yBcwnC135EGnMZ4q1FN
qzA6X4SY1YZ4jRWVRsBTSsmkY2zrmXm2uQbjexHRKkIiLZVnofEGK/yG2ES2V7+J
VNCjwz1jZkJT8J8LnMjjC66t444PcfpBhXhQzm175UyymkTsytexe9WFSfenGVeD
WrfQcO4ZmKJng573WrqfRe1rKrKAp7aqRVaPkqfsnoPfbfz6O8x1W05pUcqgwSEe
tJCca4keYlIaVf7bj3+If5XxhDM1rzh/G3A6mSWpaFejTO+jY3wH+xbFFOdWLXcW
FVGwinqPMDVsvRB8shutKBGcXiWwKfON1i0lYgBoqof0A6t+rQzbqzStzgDKaI0X
+UakYCESw7OACwpOvq2i1TdvXEGm1baDBoPyqxEPcKQm50tao9W7xU/3NzMxKC6C
KytenEtAHp34fd7/+OxA24qYIITD2I6mgiEBOBwasoOEbPIRcNWJi9iPj5N0cy66
MRR6s/igqaaKq/pc6oUF5qjeOotAEJf+2qnqr9uW2bqw0gx9v/yJCy+y0L+V1Dt1
YXMhNQUBp23u2qo4ujYPY3LcL2FzME30L2BjmL1Fk3ij2MxoLvdBmOotTZYjZnvZ
C6KXps1gQ31R//+6LIM/gLsA4ggC0IdeCyA/3McAQOPm1QW5O8qmF6ZAmCBGmF3u
/WPTpIe4Mz66X518iiKWLaETJpYz5Sz+XVoBGPWjDzr4QlQGXputIlgdemzl5xBP
XNHrEKAsT5NcTqrqu+DXsPFIdgcVxeRIxFtRueE83NJA5bHgaZYCtZQqZPGKwwWq
rHx1j6Tqa2Ll9oov5nAh7+mj2J7OhqgkQIcQzZ4E3nwd9KmwWmxKU8/ebFQgJnXh
kl4+zh68N+BTm/BwHNOCb2ANwMVbZ91yNdgdN187f3EVjlCs5BiO2nDqgsVwOwrC
EovRg/tLIWYNVq+HDoS0/0u6blK3uyiLDEAjTFGHWhaha1fw9Rseu8tMy8VS2JYR
FglQ2DJZNnbbS+oG0k+3UzDAH8pj9i2sPoojD5x1O3BrcjedkG1AObNyJJfKt1xD
9W5h7y5u2MJtiIaN6VHb2l9Ld5fa+ixxOPf1UsgpqoQf7zyQX7DCjtWuOwgRA1SI
+A6ZQksuOYMEwkc+bZlpQmnkxVRwKSYJnULDrVTrBTW3IwenpJklEKtPGv23fato
3+Km93lQB3rQFS1swYeFCl2L1Fl8d76d4Js/ndgcT06K20mldn5ydAghRP7CaYKY
huFd8RXq7jfDIAZXt60AeuFDfGs8+eCgVjfPGjXFRkWOMf6nd/C6rc4NbWXXHzSP
B8K+joBNbmUzNt75cjOIrQsbUhGKUEcTmOpVZbA5Cr3KcmGxoU1bcbQ2lEOtd8aq
2Z9EtLyb6bnNsIG6L95Hko7pnS70v6KbcrJplN4sZq+wI+jnqOOR5TOktQNc5NjW
duWBEzVSsO7iUkBXg3XC+8vt3kX3NCqDTy6eBHsx5L7zDpBlJj8xx3j3Bl41j8fB
E1uTrJ8oX/XD7e7GCxIYmN6o11hcof6KQHnd+udmdzVb7tOML8px4byDhwSvXpIR
Pw6SKK6dMoQ3Ce027q0OsTo3q4YSd5bZiQquMr0v41BO2cOwpiz9U8A+sjZW7Fsd
B88pPcGHJ+omp9PVaeZ4YsncPjQSEwH4ECiRbGMJyA2Hs550/A3AtDGAMB5dff8Z
DygB+iQAOCk4WTc1gtrgSsDA2Aj8Ye2BHhoZDFgi5WCW27EKyV7nFkTgj9FERyrQ
YWz6fY3GQig6k1L6WlTCZ+Io5gL851rMXZH+6ePQaHhqm148T90nEtBr82RwnE7m
9oQEdKOQNPRUrDNyaiqS2ZoJaQrZOlDTugh/SX5tnlGT4AQlhDJCAprB5/4oSTpv
fj2El9mAPJ90HDiD+44VfRucmwemSEV+mcON9nVamnM=
`protect END_PROTECTED
