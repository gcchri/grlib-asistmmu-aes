`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V1h2AOrlWcnQ3IGDkawO0w/2kmdlAeHT072LI9VgIg4Pg1SCo99UDg9azy/JXs5j
10b+yz3mcsa9UcHAYwfzKphyLECIWBIYNHcLsfvXcxpcUVrERiLqE5N766P+AaZ4
/R91ET+IUbp3jgolySVcYhOF72ghIF5USbkB2hpn4r8zBx3UG+FW84aAXZFANUTU
WoEFOIhrZqEnFO5nSBixmBGwn+CP1bdiZEpCX4XIQaVZr/4wkOpK9xs1kh6AqI8K
sW2TNYvSC5BOOJmPYuyZZO6SztmrJgCJQkBUnx1//h8EVecDb+x/BBvKu8pawwpE
vAEFK2CWLPM7tZcRujd68A==
`protect END_PROTECTED
