`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FG0Pwl4Ijh4far7ZvrFQTki3kY+MSgJ9NQehPYM2TC59uTIuvamoOM4gr29wggSD
tik3M5dZZBh4ln2N3axXjW7ruTi3tYVthP8RMAIxPiI0zcu+Ua3GhtMYjgLYQVlz
xSC0rW27+zKxazLaaADfA4AN70tQeAjpJ+KKwicu4Aom/864uri/ancmDv6ImgBQ
Ke5JUepLZ070Pz1wzdrkEWWdrEnMjIdJDShPXq5fBzTgahUCCJgnF6uyNGNAEJrH
kYqVclFwLEHxuRoDnV0FfLDFkbFTqpXXJzlWjWphmlqMGd3l1sTeksLfwAbRrX9c
TW3HYo87+QefCjod7nqFByhI5cVWL5ZzvPnYQ1fdozdUz5FOZCV2ycemzaVnvZMg
3rbrCJYSj6Q8mA1frbyNkz/F4PzhlsOGJcDcn69hQRA=
`protect END_PROTECTED
