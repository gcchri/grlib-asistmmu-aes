`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jlQSw8nUfrFi8jQayq0wH5Y1U9HnbUfQ5dx+lL0AZxTeJdvB0dNXVIypuUexEhk+
CUzdXLmT1dpiKi/Yj60CPT9/SeSAWdknnyTxGZC5AmAh2f8k9RDuKhL9oZLAOwLN
FE8LTW8sg3hdaSUdVOZt4VAwwS1aIMCdNDoyldtln53KIv/8WWC9QhEDLW/3wNBh
NBpj/WO6wcMboT5Kn0PsPCA4QYiyb6/ctwVdZp5B9gbmGR8voEWU3JPB+ayzPwm9
ik9o143cuGJOuCuRmMoSbcEoeZPwjsUfMDjIRejdSVeBEylOBwf2kyncfrdz/15Q
TtewhdEwOo2cFDoLjxf4/A==
`protect END_PROTECTED
