`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NkNS8bU5trpf+UlHp+G995B1AS5oRYNCMDhJLfPl0dAQi0JKek55RlxQuNeEG8aR
EtSBk9+CMNpN/Bopj56bpd6H/SYw7Qn2SrRS1XsqCPxtIZwxGPIQvr6EH45WVowc
kA/u/5i4/zyASdbb7sW788XvCHRjvLKucZ4UxoDnXtPN2sHneQAdC+B812AJ9DlI
NdLgTbTGvmjYPW4+R7ox1HGuS1dcVnsUKOoEd5c25rl20fBfi2AWnpP5jbBoHmBt
+U7WDEt4Z4ZqGJs0pFXIKpHdWRO9/8kQams9/PZY86hGuEM8QfTXLKcV53W2oLdb
OpAaznMacm5D/RbzN/bKFIWnYi9Sx3v55KNSO+IF/RnquQ63Triuh++A61ytIRkK
npjKI7uT2Y6GGl3vv//aE8Tgyvmx/MxzOkIz+aCFb6M=
`protect END_PROTECTED
