`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3jvJueIbS9BUDOEEOofSl4/5rkheQYX4N219TkCYXU/zJA+4uu1FZ19pGqHMxenT
0inkHOP741fnK82XP8u40yDcJ1C2z/1uvB6192Q3aBHqW4QoKuM+34v/tnzenh7h
OSkFFTuqgJ24aUTULYHp45suPUaY492mCTZKJSWiZOQjV+/DXruD4xzYZUfHveXd
+A4Llm4xp2NThbJzmuQnZT7exCOh5elYgDznm+U1+KV499T8AKTApgldd5zaP3EC
bJMYLOILi0KkAGYXAZlU9uq0r0eoP5B/m73jmgZFPW7fS9HnZ/d4YRpsyjvJcFte
U1mYUtsI5T57wG7nyiTWg7mmw6j9izmxoa55Gj60sHa6pRJJ/n77nv1ubUDPDMAY
JLvoHvAntNg6SSJL8lQSDNKxAgm5gzsc2fBWRs+0cbapgPwJ311HvcpIxUCPZ75n
eeH2XpGk+Qj/2nCdN87lGBczjVWOTp7c4+B7upP6CWIj3FcuTKyk+FsyQhSoZ3q2
HGJhBlaZi7lNRi5LL9hMk9L4FFgUhkF3Fs9C8p4286uROBHGARprF1Y6S4LxpMf3
5P7G+32+MmFJEU+Ctu+E+D4BNfbHSdlRfySAiup3hFcYb2dq23NyC/ePsiAemkCA
6NBaMGrVC61HTTCvORlUc2E9ABigwHHtBE4ynFQ9lY2jP9AkZ1yHKYGXoHS6kYFE
P1JtWDsetwD5gZCh9x+WGDKDjauMM0AG9Z12y8b5Bk+3K9ytwLiaoexy8RrYxuPF
oIq6x68TRuMkRanhuPhhljOks9TZ/JPuqWzoXG6j4s8HlYTjhFWnzOGqH7/prOHX
1lsLNnFa7sIxxt6x9zyG0rLQI95aVAeEBkppxZb3iCItHGM/dUqgDj4i/b3ZwpmG
EvZ+Ik0sOYPLZhZGvbpMVcGt9uN3WZrF30lcWTrQbVw7r64BR3VdrGdIkDd1nnq6
ay+cnI10fecaIiEs3w/Gc0ktjKs4En0JdJBcA4E2z63PAES47yBJWtDFwE2Xol7d
i8PUCx6mjO6ng6wNg7mJvD1pECEP4xSQwIUStkMbB50h90IYDlylxCU0CZOkEHoD
Ccb9BNG3c79SDvIB5tuV795edAUFTQl6cjqEMsWbV20+hpPn322yzTZLPv8DhVF9
4ib2NeS1oTYprkgIBmCwfmeFqk5lESkNcDImzeEdmNsvPDy0VogGjn7d5tDtAdtB
r1+CbGJ2wzXimXtKC8qLyXrtMDwNolyyQwRGmixxhKMNq3um6OT3C+Ww8QQF5qkd
FQ0qLDFEqwynIbby7NSPDmUivhn1Ns852E2KbV2jq7ty1LpxWqX7oI3sMUxbcH5t
`protect END_PROTECTED
