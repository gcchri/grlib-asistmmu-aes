`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v7MncmIte0RXtS22uLu3SNwQeOVp20i7yMCUfQscJ8G4FLQ+g2K253+JsZN3xCRm
6ctJ5aagBF2RtmbiNwRa5XUmFSM+Z49+/COtTGSTI4EEm5V5rB/G1HlWlSFWBMFX
7/ej6AlxuO6QU+OVCF8y+UNauqeLVIEqed7YHZkLenu5RZAVheIwiWlRGvmQTrBC
PAR9xEKSyzmguuDZzk0tQnFef5we/wMUPWtl5lfdgE7YIpgwdAGtOPzajb88aCy9
dqIrhXpIjK0YYKCUSnRJG+mbz4oXpwHl6459fm0H6V7QrM8ojPbwK4Cqu/2Cv43R
pjBSjXpZxZeRNcmKPTyAm6zaXhcclc+eefAQi3AYAraeEuL4nhaCAwBOKR9weKzg
a2ejNDEoThZ5CeoMDNShg6Tti0tJRei5BQrlXcg2aRWHsrVdmVlz3Fpeo8piWZ0M
FhxoquBSsMfC8S1timcFfMcQArE215cbxMF4BO9LHcvoqP7q/p2pXFQSTRGKrF0N
`protect END_PROTECTED
