`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MLVoTSx+nBEppAnHL1AvXrA5TqcFtAwW3S9QpdtWPCnuaFhYmePfs5dHvcgHYTw6
OrBtxd/RULpnxl5+xqPj1F2P7YVmojb9t4Ur5WkARBNt1K9Fxpq/oGP99tTWarB2
5ThokeAddzpOXIUtioG1+6QRcGNhS6Yzohfcm2KrInIEcy4pfHpufUrSeYqzFGcB
UF4rLIqcHm5GhQeFShvAasGYwUBRtqGf5XfdN1Gp3CJtaFPUjrQEc8dq3tGi3gjz
TU8puX49Zh1OeWApdHeIFLjmGqYB449smt5hRk7u+b/tbBpUyV3ok7iokIpcYxUH
OAT7wT5hH4yU9KbYQ7hIHQ==
`protect END_PROTECTED
