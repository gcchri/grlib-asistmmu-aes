`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t5zOiLirldsMpKd1CacYWLvTOFj6QS/8VNZvfgxqewZ6wjvzFsbYjbqRZ5+8QqWn
3Ny92KkSQ1w7LhPh6m/RfrkHPM4G2BP3LQsmJvLoH78evgh2UtLAZnK6OoudeFUj
zfX6PjEz6CPw8M6xiooYN8mVRka17IeFO3p+wqX1N01fGd08PXeO8d7cU71h3V7D
kuSKHlhaZ082d0fYlW/n29MhFjjIEuU7H3fxrS0ZZPZ5F2BlRVQJ55LrIkYbkRjS
OD1t1RmdH02/vnQ8MUogB9NyfQekUHSJMRIE1y5SozaQ+zVD5PFXAjPpmHroP83l
gB0xg97/ZvlG669HOIIZisP1mpVTtDa5aK0xSjDlI1f5l0BiNrlx2po6EeS1ECO5
ZDp96gJ0HiUXlNd0S0kMG2d+HaTHB2cna5cIKMkUB7qs9hSTyzhe1LXBVovGyfAS
rpjeofXAfItnbgfsMorPbU5kF7R2YCQZYrbF4cOPLGM9XQPr5C9JVrrai9cnvVnS
gXNCp5PHQ5p8usLm954X6lcj73pLv3nrXZye158RvZE3hgDZqWnPRGs312h5wMjq
wX7rmdvzXjJGxXrYE28xD4pA0TN8439IIUnfHfTy27mX2StL7rBFCk+40rWSdI7g
ycmQln4LaWDUCdPPcLNjHKtT1J9HhMCIEkESUTzU/R4DtKUERYqfHFfJmHP3kZfv
NbL/7cro/AmUv5c5qBvYi8djcvscvItQ/yWPYcVeKwxEN7KdECEffq44Kwo1p9Ve
aHe3oym/d30Hzu3H1vqjRJ8Uschx3x1t438NJxPtM19ldgHdY/O1afaycLFvpz5r
YgmerZyXW7URsL9MJVpO8g==
`protect END_PROTECTED
