`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S4nv8ZTuDx9EvZ63z0JP/BCVD+1zCtV4qnU57KEBesvTeqXwT1kbmTAEJPbeG9Ww
fDpb9ifC8sVitnchOr42MZxEtFmOO3vRXkoFFoIjIye/Ek2Q63m4sMUQtcM59zLN
Gcxbws/LJ4yJ+7ncIQ/yVX5rTGUmEyj1OJh2Y0ypDf+JpcQsMNOlz4kNpwHg07ie
YX1LD4W9fvjLcOaaLxpS/bp+79xFiB6Z3oVNc3Rpz8X2/yF8uZyDwhdR8GiYHCIt
4zTv96ySNpH5vSNENaguM41g1EPI17YSrzPofU9EYOQ5y9T8HE9sQqu/qQLATIOG
9L0isNGGV3nmo7vnKUAo+60sNTG3oi465gsSQmJSdxQ=
`protect END_PROTECTED
