`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZTqNrctAMpnsxZry1Yw5Cbx69z4s7+v7lv2Ny3LP7688UlbKXTgGfN1JaLmmvbkA
xuXLhcyGYgmdtXaIcMrX0D0svRf1dIEs45vVqeT/3w41Ni0adraq/To2B5kLrkk7
A2uRWiA4N3tibOzy/P+a0f6ycGCDnBtJQByEou2+k/jzTTpeSOVQ+JPIJpHnRDTA
lgH25AWKpOMpunS/s+JT+SQIJD8z+aPIAN0iz9VoyhJV4wL9bhOoYCYnipSNUWSW
Slk4d3wQnMQYPVDFVBankJrBAkDFsMKqoMZRmUqQ+6bgcr6GIx4Iwp8C7rVBkpjJ
AUWIFcGHtD87bu5JxYwV0q+QkYrBFlhThl98bAF4gma/IblW/sEvaovV1YYp5EIJ
e5WWA8E78aLvuj+nQMM6eyVBXNg467oDZqEugLyxh4IV8yTi+834mo4kLOhZ7E9+
Drc6KhRzF1V0M0psZIiUkZE0Y3StAMasBzeDj3TEZNGnJ6Uc+wDM2EVGzP+aSKM3
Io9usxZKb+sbqbsE55MtDJvuH7Na0J1zewOP/rNjRuA97+a/+QWD/VZqV/BL14OG
niN9wzuCUUq426IkrTzPaKKtNWxl1vI3l/RdM9gOJrSCXrLbRBH913G5tdxNQCc9
6KgMvhzkjOzsBfaJdXPQqAzPBKb2VWrp2+EOjy7NqQ6md+ZI4L4DKElkdxMc6iy8
Bj3y/JDKWl5hQkY7ckhi9PLtq5+EfO1TxCJyiIz7xS12Ww7S+Ag8T9VXiwpRhuu7
iL6tDN2y+78orSPGTpUO1XmTQT+quv+lKNdfSwx3Nnz5yeVN77HcUyl9IcTh+E6Y
WKHp+2P/3LIzA7x+tj/6jItlJvePq3NwUtS3O1yJyt9w0P8ocPo1iF+phDrxsD3p
hByklTH6Adzx+HQW1n32Y1U+bVcfAUZ+qCjzghq7oQxJmFraujc3UV4H1IartB6t
KId/BtyzULOlIFVVfiXhc02Vb7Oi8JSBiA9gKHob5lP/2VY68vpODgBoKlUBqJBv
94/pedEg7+/HbeG/kH9LQoRo6Hyb8izFe1r1z9ECoi68dOPc494AwwhbJH8AMdCc
OJLl1RZDceRZbOK7jg+PCfDYoTg+zPriWbvxQ4O9w2YuXJ2sBor1uUF4LNczTnyW
BtfNWdbmwkJbPXbrGLRJN+DwNpGvy6OROwL3JnAZQUrTFPMdpAJogpu3I9WUD+RY
qmnmg0S7GAzPdwS2fbwEHtv3tifapir8qXmhaDXDRPxHef4Ku9aySimqL7HtB4ae
aDWCsOlDwA70MlNP4SMPYIMQUscvnad3xkw28SKqd2fe5sg30zfxY16FhMr8tqcb
Z4dBRzt98S2/xGrW7mgI7kYdJb4rRI/wDOrkwJ0/JbMcMRqU3RZlb9qosbR94Duo
GsaDq702B87w8/QVlGJHEPny+4r4xj72KimQ50GTJ/Kr1OdflBKXWM/gldIm1kkV
vB1l8M4mMmCJ3W4W9phcvmS8iUEYHk4LTXG59KAEp3R5Xb0/jog1AfueydOK0064
QfiRQaVSZpPmjWXzEHKyA++jByD/rjTM01QUuW4JeeHOKj724plQHGrIILcY9Wj2
2cC7VwjaXPQhdwD58AA/EzNvFt1BLWGudwJiEwr077YuiMF9rsMBfWm3EUGUQ5nr
6rroD4I53Ic2fQOze6gNYlQPTqjjWLlsQVkxvQjXuUSkKZwaxrT6tfoxc0wDuEbR
2kCxabD9+P5pT34XSys1QTcd9zQMnXiZIe/HUwzX+ECvWE8BX3G3YfrdzkFy5BbA
MfvPUDDnRJcSRYOgF1aUHgfBzubcp5jVw7uVcvcLSqmao1IwLHwbtXq2ZZ79XJf2
A/fBQlkQz4ldUS1AziIlXA7a9uoPxVhnjxM2rbfzJVFOc39qAl/Kwl6OS5lkAIAz
20ql09ABiYcAPWu+d5DqPPU0n9jVgOqUVZXVchL2Kg6RH97k500RMZRVjhzn2UBK
Y9ClyPjZIgmIGobstHhMoWE3ITDaZAhKO2PHppjVnzgJx/PucaXQaAzIYFC67EVC
ld2tjayBQGEo8O+oUTixggiUglcmiiHg42ZpgPU1fxjsH3s88PrBx2/qLjukLKcs
f5V8flDInMKx+UFnLse2XGBK6uKYXs9YTZRl5I3h/CRfYqJcBskCfHKarQgfXmiK
Sylg9WlRkERDH0jDGoXiNrm6cWaCTF8JQBsYBOlk7UrqTSYMBH5UEu5ZqIg2e5b5
lqLKyRTb7ffxadZSoQqTuwCBZJIduMZ7YChghzlkGarJV3nmCCMCZC1QcgOEI9Sb
+hySuP5Rcuui7jMvJBvgvDaViol8qtUatMjuAd5puQs89raXvVnbyUkWAeRDPrRK
pcjXHI0OZvnE+oiKbhxW2oSfvc95UdCfodKTcGEHTYs46v2UxPUpVs12Uxrn0x+3
uY3tCJLGtuLNDPzQR8lJaks5buW4kdcYB+Denwg+ZvMgZrqlVg6CdZoMmHeK8ZRT
XYP6QC3LSdniTDQpcgxoG33r+btSMnX3oSUnH1s7iSnYUqyq247wy53M9LWyctwI
kafsvbY1PoqGdb6YKfXFrqe5z4EiL8opD/fSlhCau8mUF3cBsPxwv0+/C7NFhD3p
8Swfuxvn4HwTfXTDTXL3Ok8COXm56bjxl9sAnq9zgkp4EbmSayhzimBR68lRNnBB
DuOKyUseh4OUOLUAijfdrCWhogFJ3OSAwL/+Qey89vI8IA7OGm9CBJUbfTr8MM8v
/SC7maOvgks7ZnHhkvqowXC/PbkXO6nz0KiaYzJr2s/Srw/M9kPdILjazas2tWCh
ZX3xTrHN3r2pkjjtPe1diCuKVhhWUlsB+2mmoEo6nyHlRYoLnakqG8O3EMRYGdbf
LukQ3ONwMulcoVQzN9+GjuKrAdy3VXGKf0nuCGUYKRbgO3Q3PD2zJLjJhxwa4iwu
7JXtdR7ZA6IQlesXQh+6cKbK8CWEr86njR5MbocR3Fr7bOGRbjnCV8dyJN3T0Hnx
Qq5rNSbqqiRJYpeiHFAbUCirfluwiKLMnyJqn0oUbyw1HsaY8/e0V54Ux9ydQhCD
aaZW6abIxTakxwoIyF6QF+lgGWeAhco1k5/1TBeog/6zXn0rbKn8ESubfzsowaC1
f0J0JdCGbHEr6kxaqjlBDsWocxqJVp8GepbSkTqs7eUJG5t8HqUU/0irNpMlUraV
J2Pf7t++xI4ibG1aospoz+pPB2WGv3Cope6CmNgvwhvaSInEi8nlfxGAXCERgfpE
fLWqI/UYYc2CdkXOlt5dt6TkiZJV3g6jjRyqM/O7jigQMEbWYY1bFO2APZegCUAD
pi/m/gaFK9GOYP6/Kt4POhH02NXrCLIBMNCrrbrIZoGlh3pMOvIsuH6sVMOWbAwI
QnTQZe67ISGTo/Yxo4OArVxTYph/14vFW7L3CWqzuzVhlSldQmGYJpAZubDw2Qkx
dzov+EaW0zahSNej9pSHArWnz1btv6fvkdrGizJ4oFFPeu8cAAgym9bTWD+3/Cki
Gd0l8OWorRZ/fI3LdDEJkfeXnmIOn8q4aVVkwt7V63sx9ONOO9zjAR+9NnYPbNmI
JEXhL8EhsoKG67YGj/cHds3zq+35IIifA4Q6jz2Bzh3+zTm10YL2/M1bk/KiFKx+
e9M0NFggw4q0Xk+V8BFb6eaSigXwB/chSvVsGxgRgJRT8DwJDNduz/jsUEnWF9Ym
gij27OMUAwD7VYNg9FRf9H5BBZVwX9le8vwatiDN6/tHzECO+EbfrqCcxdIgJ3YA
5uTsoavikLfQEFF8pjaRKPBVzSQtEN0WnikTz6bl4lbUBcdcuo959R/q1wVRWvVm
BxinRDC+aBCyyONkK/On8a7xp802STT9NfDLhf5SXZZ7mhWnh4ZCnRm4M8p2ylFt
0/l9vYZM3g+s0FhRvZ17+a3pVxtKfZ5uJp8BEEUXK/jM2SJi3eOEt0GCcjyw9LTr
XQscktECuWslWOQmOhtiXVM4tkzz72yR6PJySnYWG0TXkpiF4i1SJrP7Mw1vhy2M
fzZ+Q6Ad0qvzHxfbH+Ex9fQvCrD1dQLfa+NWeipy23GBjpAHEs+u7U4jwQUhce0E
fVHThI23kLIafJveYY0q6+Tq2YwGLmjwOr+s2AB0ItqiNR+GnHuvbBR14vWURFR+
9y/s1EkCv16x9/lwcHikKU4AjTuaiV4WPFeUCFDUzdhZmI8lfIb87XORJCLQqJht
1O/hmhV2X3x/8xZgNNhlXeOpyvm+g2CXHafGCWMfqhFC8a62fC1sUQ1r1ivYgi6U
jOCaHNHz6x7xSbodQcyBMaFgE9bO7QNfGYlU5b3LazbMUrbWRW/akLZq/OMgLBiQ
VX2R5PR3HSgfQzD8H3RQ1f6KE8jg2VlnDk5R5QX+TBlpEqjptvp/tHORZZLCARXw
TfSghKrGPP6ilKMhqSKsHHlfTwsRBMfc8vkngquaXOPYK6p7QvDJWa69NZ1tk1xP
+xwpw37NKdX1FMd/JtzYxorOCIvUL5tjjqV+WfEkPeZEqrlJzuBFOHGo2StIThB/
JHbkQWbxaMRuTSXU3DbrvzrlzDu6gd7ybTIZ3ho1uz/QBraRg8dK4ercNI3LN04j
UcfZAAUxd8yPIUWPOkvX7PFN0Iyl4aIWrL+gYdR3QDc4n8dT2M/1FgcogVwN4zDJ
agFS7Q29koTAqLLMBm/PIfTCzHNix4MRo9V69f69L5qvOTRONojJ0xHpDsiHBnFl
vxNHbMe90iC2y8lNcJXcvLFb+AVeecGDk9y9kQE/KaD7zHlnXzegYBNGJDPd/i/r
SpnxpN41BUbC1IsksvgUO2MuQUBjXzeHhgCZDZMShAqGiRfLv0uuXPLb+aW7qkwl
tbABqqNhCXvdTSEgYDBBeb12BLdsVvuDr/1K86sAo7l7IjTQSb5nqqduGpWB5Qq+
8oSXY9g85Pob3yXMpRVLZds1Bo/f7LGqi1tmp3InJ8htLS1KkZiQPRiJUC9Br6O2
KGNRQb6xmq9Lvy5hFp/ISCa2DOPE8BN1ZQCWN4gSl7iHg/mNubRV8QevLPgscy0J
Ln+enrel8rwRknVprwxoVfifrHe+ZrkN7x54PuqXFadbJK3N9i202eLlmUa0JGlh
HKGHVD9kdgPuzXW74WcfS1PaPeYMqCrRIrrnSrFwewfl5VUucgVodCYupStVEZ+e
vTamzpBL/MLm7JdSzfg5Eixu1sio0+pGrYi0ztGTv8g01TTfvTB+7I1r37/UZXR5
xK1OwX1rkgiB2VfowHI/hoQZmX2QsGV4TGnn+MCG/hCkaCMqU0s5otzc1z35pLYI
6rj7mRi7thUvduGhf0CnYzwFR1fsxTsHtF6YapaUZ8xDC2hQ564OkAJe3Zqx4IES
tDVevZqeYcMIx2uK1YMfTOqe0fGJm9RufU+68NTs7UFgI2l+vB3mV8MEZ8Tx78Q+
TcSwYkzNKzBY3NXCIjdldulg5l7C14bZZer49W3bfzAXr/qut4M7o4KmxcYNUndO
JY4XNwRrDPm1r/YuFeJWkK07E5gklX74Uzac/8HIZuI1+RHJn0suzaX8RfKDuETl
MhiNYx+T/Xi0zozfKfNXf1RdsWZSQA0Q0CkMAn9GgaBiIhLfuGDx9WOItS/Qi1vV
LqrOddgsZOZ1a2tKBHkMjft+gWyLEyHU8WJKpxjXiL2olo78E/gEQP9GNcL+1NkP
5f1yLvRo04ezq5E8NbyJDyWoJU96ykiwfYcWcMmuPGG/ErClauPLBVFuvMmMaCLV
4347WaJEjnpzOaqXwX+3nYiExSKTSiAyNwiaDuH7z4vM7lhqY6uztVnQRSYYU0Q7
b0DyWS4JTYVJiav7SCnhvpM7PlTGTTQT583pgSy5fWUe/AlgN/as2mDDCMP+tErx
6mVP1sj6dpc9Dtc+buyBU8k3BLYA67hJ9qTPqwRXoWqIVGZ6ReUadhLaVtvgXBRh
sQce0vIoC6HNEQxzt0XgU5EApk8QDZxXs2vCZXFcdLEIed+F60DF5rQH9geJUb6B
FV2vKtTyBemZST4QvNBwCt9U1eEj1/YCGCUbBMVOTROzbzopX0k38vY8pe/myJ/H
oce6pPcNTBXbbTlFRaJqUky7Ee/sY4u9oiYLG8hBO2DMUa1bLfdItdImV9aBsPbZ
dhl8tcDi9n5H3m0UDWfMTs+kKmc97TRZ1mKWGp7Bohw8EyjuMeUnAqf9XKA/jIo7
X26sfQAsr0VvyVKvkwc1Est/5X2zkl6SKJUc/9lvlOE02vp6jyXljo6wAyYINjw7
Bo/gbpi4krP33lO3eA1WWPDFQ5oOVreWUczFx+2NMNRMv0HcL/ESQwejQEqrXX34
+J2P4nUOFmmt98xiDKbGMuLwG0WVSuoeB+Txj2cILADPCy/aoXRhSuzmHD+iXgzS
+StHvdZrGtx/gl4oTap6EqR5vJQBtxX8lD+OwsksgUl2Hg9QkcOILvyPaPPXbUIW
9+biHfRikrZ462QvgQESmqgoCIwdOYkVSykef3JS9XnwWr/Ij2i0GqyvzbEA6MEQ
tnNVhiuw4BJ8MbE2g96rElZCxLKLiJ57X6LhZworLUxFpH9vLphj5yYv0E19XQIA
AsjePF1Gh8dQIK4KX+zdFNbplim/clD7JdSHtQ2kQ3L8a069rcsOVK1W0lT9U6Tr
kctYKSKs0G1saF3PWyCNLtvVnSfGeIK/7Wcs0jtzJgoFTjvRzn4nHxtNjAluob3U
xu9Hwxr/I3yAtH2eQQ7Hcm9Oomju4goyccI6TbXGOsfBIEANvqbvVKZq+dxG+Wgt
cZhArbfeX5hj0LEp0Oj4l8VihfDPPszV/lEnvL5mCmqFYe63cBFugAikaUkbMJzl
i6iGELlscKY9D2Jv0VaxqRDqJPH66nl7ooPY3/+ISCpTXaYd3f8ymQXJqJ99YCdF
3/8Z5SKqX/mcrNFVra7LkHk1Armsocw9X5xzBXLNo7BscciN5NJH1BTOdM73d1tH
6k8SJs4Om90WqZNtjGsINQoaFKufFU1pevyitha1GxwjOrCWJz2cuGGoiIPN03ar
C15lGlomfxXNTyjIbA3ACFalXpJTqlknn2FNvZ96kruKoEcBJNCGUa4lltMOBR5y
L5WQE8dMNMYcT9LfLFwD5UnaNt78jBgtcVmuznCpf7ZfLeV4xLRs9+fqTTmzin26
cCpWO390yMjhSQ6xUqd/s9RiMMYr+fPUAznVo6aXKJAqrke/ttAkwEj/y0d78Sph
uT8cJsi5M3t132cZLgV+88uSrccz86mIrb39SYHaNNSmjyG2aegyIBCdhXd6JNH/
Gp/kxbKazouVPppOa/aeohKA1UKy/Z1HV/S4FNJAz/vXXOJXe5CxZtYfK8A2Vf78
uEtzEY/990m8HkUBLyDZ9tNFEBPAaiOtlSeQh9/OBFvKhw9HAP2XE1ypTlx3+t+Z
GUM5b2Dyqp2PSRVKPn2KGI9JEAuZvxia8nNbnL6V5smhyyvUcH/V1i5eiiLtIvDX
vQ205j9HXxOSCGwhp90EDWTHYx1o3IPqVoJkvqq83UY6RUMTmud43e8ll3qhodMM
ZNOmVQlpVAiNUoanSrGKT8dQcfLbqq9JMpARA2nSWd2+WkTK8fsd4IIvZqXWu58a
siVAGhyBgaS1ddunFy4FSVaQYTgcYL6hYzKSncGer+wxOzss/k1bpC4H0VTboElZ
XI4OI11qKRZYuoXWVHT85FgHjzu4WkPM2y7ZVeIJeikBhEfbruSL0Dc9VFbHikd+
8h6pOdFjeZkyPQJG25A/qDhi/M2rrdRW5zDjPQX9/6ZokP+sLVRlsFdrgVh4rO+n
yVUimaPzmUQE/P4sv/dPe4mpn5c5lgYJ4SS4F/qCl/kGw4nYrF9R/sLf9wjWZuFu
p7tfQ/FGcIJCQjs+Wy3u7CHpiLccx51KxSw1y+nAWG8s9Vm/UjK80/ybMqo6z/aw
433ebcxpZ0fNLtOeAWVVAk7X04f2pJ1m2YEuaJwzvnPIbZjBQ0mVwcrmJRR37Tyt
27TPlS8TW/utg+H6zhkACYaPOTpJr2X1JGCHnaoWdIVlh1LCYySeMF03glGt21kx
GH4wji3V+eo14P1vlIJLcr9HWaZ60zn5oKiwdMq1SM4BLxE1gP8IQjaUdZEiGIU8
+cnqwUkL3pCVOqUyTw0A++n2h0JrH9Z9S/zJYy0Z3Agtm5IG5U1oDmRW3kGi/1Op
cv/yjVd3kpZejab79u/Kxa3rKvBQFNJ6U9qZhKIS1ZLiXTgt9C0/T/1kmnp3Rcw8
stUVcwyklrfe9q0BQs0xUSCQWZDfXwLuXOMkMLDPu9SOlXcPU4MrU8zANo3mUao9
usfG6yJZLSmTbUiBdxXf0ydhy3DeCvHp+IrDTpCGmgD3oLyajaP3Y1q+5I2SyMOS
WBz57ml+NyjBF0Hb4jovvnOzPQDJZaBdCcbxgsUGWrWhEbOy2uC9fnKml8BVtUo4
AZJsxV/BYCpbWoz/Jx4rneggai71uLWF2VYxt+yXRT1oEQ3YfUPe9HihKAqU6tZC
3aKkqys26BxU6DGE0CQW+dJ4AA8kZcdqYuIq61duGGxpW7Dwk4kEXLVwXRM0PkzI
RM+4zTw11Z3ctJ4vISrjFJ7Qctv3PqkiThqSIInD6oCtbp4Y6IVLSr85SL3Lw95r
eVhQ5Fob4dRNMRaQSkZqBwCAZLeqGgj2jhu8u3jq9SYIglwQoS0W1UnQb5LOZ7FS
pfh4DIpHA5FqlkAeAQjydj4S+S+v5evkk2PJ1C42vFPaR9qRJCWYARtj/ctTBnw0
fNBBE6INrxj5sSCGbPtVO8gWFOX4pZiCal0eRnrjp+nZ3OGHOLJKk/+ZM61GDmX8
Db1IjzGt4re1WYY45p+xd52lPFmLeedyIG7mr37CvC+jinO6qSy5uLj4sl9NoHRG
wFtB4/aIVuocDCIBX21Y0Vgseysk1yCRHcTxcxL7suulq/AXPabKc2tGu3ZzE+67
DtYafs0Qqt16alDeUFDMqqbMX3kHoC5YWt+LNkluVJqaMjA3BAXToJVLZIUV2Cj0
Zq0AEV6IDRbodGb1cTmMh7eJIajHxbGTek4+l2NnXrYGlg3DK0do3IU+2VrBovtl
ZkrxyYqlNNAAAbHq4FoBbtPk5zuMPbCNzkxD0MKgVCKJ2icDNDWMw1lysHi847XV
3dfEkJQg7hdO03L4HEIOXVDtBiaNDkMkNt4+X+jV51A8UssZXOL2AInpV60FmK8l
Gcm3G/EBDCBTDoZ8xwLSIa9p/CJCVgweWszGqzHZEp8fHcEZq8R/XlCFD+tcbG2B
Cytqek3xLCyagaDj6HCzLuNkxzaNUcfgxw17HyzKZkmJl7HoJNCcwVk9BczA32mn
nNHwrK+ImO7HW9xSo8koBwbA4PCwKS+wLJcz9rUeSHvtS95psGYLF9sUo+MKVvIS
drQP+NKUH2uQ3nw9dOU88uyRK7JmZfpdtczIguXuDTfwWeHbVN9c2Hwyz3AmSnOe
Xx/lYew3HUtayxGwbk1rzgXT4o+GfTdg+EA6ZZXBOrBLrNG88QRTacnLy03jNMmm
TslvmP8pkFj/ZMtzkawDGNbmDWIrYUyg3fXPjH5jjJ9qPTRtXcJDalwbGKrB8B7w
8UvBrtjXyMP/ppfSzuhyG0Gk3s8HUd6y4EUC3maO2bcCdmmns9SAxgJAJcf7j61i
pptP4nibSpTr4mIVxewnnGw8pD6h/gV2HpNNxDw/IR92DaqLzRVCOvpK1qYbd203
bHHMubb56ybVyWY0NNyJkrUu9xy1fvQvw2wG+c6irCqWicEV/TCYwIgLnODYw5ov
LV3rxjW9CAgCc3eWbI7SdarGKeQ73aOnARonwfLgqETNQ+DPWgh+FTO8EN2lzBhR
BHvVh9Ql7dOynq31XAR9TfdCdAt1SXggBH4NS0M5c6fg7IPIREoxH8R4ZgfINpvY
ARKAcXTS+B/+zU/Y1K0xxzJQNMcqvRdBP95St84i1BD5pUU04iOPAoO0srrsVawh
NKYDr8DuVt8fv7EMoU6i/AoITKHoOgDl5bQzcZ2ZKSCFHsg/2XnH0HGNJ+vxJZg7
Hnl9ilEdfSTRHF5/kONw16mZYlxZzwYa1afJ4kPR5ZCp9iqIuVwravX8W9fWJXSa
n1G7M9a0UsiF6/UfvlMwBNU+B4DP3IG8MMEiGOLZaZQttTwjMcGJDmiVixWQXWNb
iDqLqO5vHq1WXZt9BzzMStreP916RRChCFK2ZYGJAEoBAXZAwFQ5QErxTuKAMSOi
pYrpapmwPTLUB3Z4vySarP0xB2uH4FIy240U7L7tURpkVRlo7r4QtRAZF8LJQoQZ
sygTAG6QGmoFiAbxum3RLxteSf5kXehe1QHDFMGd5uxeGeqa5khpriNCBz1g5+/8
K3USKKMIOVWpSXEkricsHOpnURMNukrW402MtF2uD8X7SF+7q1PLTP2VLvOnTSco
+as9W48LXvIgVc+CHzWsU9LWBhzTWAeRmSCPeoQZFQ8SbPA0HwWh0JZv8gjOFg9u
Dvw7JVX+dVfzIowsGE6GpY75EjIoPW2wO+AQlqiL/RRSW2tjaV0XcjJgObay6JMx
QW+nJB3S3cLTnmwSXb4nkegU1rYd1gR3qjlNv5U4zrh8zfCmORjmOYKY+/mYk4yb
qJe8mXZDyWVevID6tQQeiCWJkIj1n4QIogPiW77Snn8XlYvrwuAojoZLc4OdM7zY
pxI8uE6B1KjP8KX0udjArBjIQoScTm97gZ1iZg8O/0ABz1/p3M/vDnUOMfHmWebJ
bZ4ITRRWF8+RVzNn3zUTm3gqpEJZgIliczokMTBhX0MaB00kCzt8QushimQS6A9L
ZUWock/79PDYdl6QK4k3KpeXjWGTQu3ZGMgmW/l8og8cgLB/D0LVDjadhyFqlhFO
uTjHnuiHepnVjq9rmf3bPRtfhb0Ceel6YUQpYQeWxaL0RXJgdqukuWYj/3/1t7ka
j4kl0bN+3xiuKjhJNzYNAMn+U3pj1Y2gxL97yi0bFs80luCG/WCv7E0hsLPZCvJ0
aXBuX6CfnfnBxg6v0S5C5uhMssggrcIriKiL6IjTaHql6T91H4FKxn676cMv73V8
1fPRIPLbYfkdj/G3L9RfQcZKGObSW9KEfZ7wlCSZJ8MPQ4glQs8zeiv7ghebX86A
fFwZq97YbphJZ4oEpAkO3kMsVzRQjc450PRfPjzTnfyJfVXctXpTbHYt3V+myRzq
Kb9fnIyl5wzRz7FRjZIdq7EWhr/AQbCbBwDkexXo+pyW9bIO7Yz6KSTS02SWXUhI
N9vMJ40aG7Suu+HaT6+0mMbIng/qUxrbpXP7oOIlzkO//F/Snrq91gBSAtVDpNhQ
gDdLMh5aUl+NxCWGHe0v8j0eKAKif2/UZykkQ0lAgGW25vX1e2AbvNwBHVfPQJj3
6/Wtvhb6H7myf8FXrShWC9kOlK1kvJjL1V0tgJHQX8erTO3flZ87TikRnrksE0WF
DiXPTYgE2bCsvVD/9XPij8Wwoqi8Y2eG6fEIS58dsiRuULMlD+jC66l7XnLr3GKQ
KrBHJf/qYKAr5uGMmoivdQ1LKKsnRoKaL+ryVYAgD9HpA0AmaMjbUGmsCoKHASTj
Xqi7iKePJDUac/zrSddNVGq9ePihA88NUJG8wkaWBwnd+a0Dkmyu+HL/KFPgaw+b
AhH4hiCgwmFt1tl2QBVf3+HCCiFglzvhkuPlXijlyCeY+Tv7UWX/oc301Le2xFc+
Aa3n4n2MYEWXWbRC8J4a9ecfeK34shr6PbsCzI0oSXUD/S3gP7sgbrZ855KXINNm
uDyV5BbHyBDfWeg2ToT4aHQ7H61es3KWpjgQ0ypqhPt8efDMpzKLrqmkZkyDAkgE
W3oxuu59G+EDcSkp1cWRFFRav1igWWRdrs92TMrrQqbDKnxMZ3kR1dU1kS7j+CjH
KSsRkEuwr3OShbIb3CO40Vf5pDEqzBI5Fv07U6DncePYxPQJcHKk3XSb2pLfPBHM
JzaDzmg81Vd9LQ/02exdqr6YQs5vCtui95RrbYkEq/pjM1SDUBGAK/Dc9DS5bFSe
/76/oT4tjtPTHj5u+7cVvodS7wgD7e83xjI+FDlgVmL+p9xQzflAIMyJEceiUv68
5nHVvXdDuvV6hHBD02ktOO9T2UoY9A8UsyneyR7K+4eAknY47R/wH+0gERq0Iudo
zRy3tysuehYRWddHZX6sotq2TyChN93jT+XYmV8nxpLtAC9PA8kCRjJ7TPwapL2A
vLPPdBrJyVTu3XyTMN0j36nKd6nRFnBjo/XBSZXggVAJn6tjltenEWjL7Dgy/cWo
h5cht0pOyri7MeHoOBMNzAXbfN2c637eLSQX6a2DtgIqbtm1nXgCl5iTURr+kSK5
7BZseOtFeiuedrDNR7LYCVuShJ54yzkaCDRaBzz551Rf32GXoFsvcQvpxtWCOoT2
ZktExo8xcWtFBzuZIS1Su1D0Sv3cp+WCcuKHEBidQhOseGG86N6v70cnO+S3VjQA
RFgmX44DoJDAmLBwofT60Uj0HY4aVLeO+P5nrPQ9LjEliNHPwfzsGpYEOiz67wnw
0lH3iUPTAaBQA/vK81ZHNSh0Fd05Tula4FxeJTWXp2UYffqM2o0QuM9+AyknDwXe
T5lx8Tv/IqVN8v0w0DjWddQaPvbp076wt9IkSKjBafy2A8Yd8qDlM2KsCUKqCCEF
wWDmAMQ4cUAKfo01IgXwZSo2JY+Ai9NkkCkU0qc8JAroWOawOd7OtP0TnDvtSuP6
U3xJ993c1w65sowmrl6pGXH5pTXzPZx3mkS9YsXE3VDORoQRbmU3XpNeQ++97iCV
pMcK3qhJiOHCKgFQBqw+nAIOQwgVl5eUu0XLFrm9cFfJEejkEKOmMBpeufuWJCk6
t35HoYl8RqdVMNEQwUOH57hnVZyx9EZ/z/RHYu1jAPnKx1Pvd7w5kKOscSG8utCT
pvTMp8znoGpHsaH+xJNqrKm4ch7sEyChoiJUiiFk4cqYy5c7vLXt8QD3zWLXMuE/
EsyYCdqBZgAXnFQ0DtjbkOHaf/L6Bw6XJtuxCcyPkqCcR/iqDgGwWM9/h1zkvNfS
afCfXjWwmYaLgD1AjOqmFdUuFr3RfKj5vDwgjVgQgKqSJagih2YhAcnts6QiWSaS
E+dFOeVUZa+j+6UeMXQsCx4DvFW9jXk0PXoHbTLNbhgOcsFoMy1ChlFwSad5UHxi
J8swPPPy/IhbQxBA8+85Ptqc2aSx2ZrjArqBmc4kCqz9Dbi4t2gSvDbg2OeQ4S7C
PTiHZSZnpXmphNqY44mX2ks/fgODJ7EYPM7hvICj1zYeVwSPe0bT9qKwMTZwDWFE
btARmma+N7+OWygAbvF3uqDKM/oA1HcOLUsRgFpA8WvRJYug/k6+3UnIk3InlpER
cukK8MDi67jmFOaCMnYNAHZdqkZ7XYHlG3W4VXYUqC9z+AH/fU0UQOTUhSy4znlG
ZVulHeELhV22yyV95Jccj/GKkVzQOC7gnUiH1KEFM0HDN3r8MFAyJEi+ff5TbVNx
E2SrQ7hAO5Md5F+7u0IpooAAsZaF+aWpZ9Lez+bYTvJSQXk5G+WxpZH2l+00sZeu
2utjGyOlZKA2dRJasBPUIfvUSuyQHWp5rniAfyUCiNdgHcVOSNgKTKg7kuyYMi2o
8RnuBgo4qr7AIb9/moooXVmhmJLEGGJm53VZ14QVqk+RPpak4hVZCEO/mjCk8U7d
QDrvU6MsK8RtXG3XdUxXby/kQEU2vd8z3Cr42UvM8WmZNfukSBgP7k1L3Nb+PLS6
JIKxFezIevBpsdS/hSuAE/l5gH1EOrPBTbTuw8qyRzRD3AWdUlPZ4yxt4JPu/FpG
cEIbsBfSMS5+DqO5b6qIE2ylkQXxMjvpnvHRsrzZJbYd8CrQWOmC8ESpsWF54BdQ
1ouG5wVuEhNArtzu6n3Z2hFUdu6tWT4LNmc+4ff46w5WEtu9ZLHc1o2dZBa0SEA+
wnrgsHeDccPQTK0YdBeehTCe0Hosgn0RWjGUDH1lbVGhm3hoik/8AtKKZ386hSMz
9T1ok5Y3g0Cac+nKJ3vuJcooW8/aBB0fL6Sd5oVPgG4SLxXkb0e4PnPqTgd7s2m2
DzTUqgLCJyvtkqAFPign+Unx2Drn3+MuNVdvCPYh04yNcwrfDPAPzbBqMXQs+aE6
TeGsZ6qqy6xI1ZpKdE74jrdWXJdk4mJk5idpHsF4QJWJ7aiolorbS/pcSZhCQ7c/
XdGP8c6Xnw/SbgOC0eF1Du9yFev9FNwSraDlcVT+rjYGqm+/tRTtvvJ4GDPyikxa
jLNrfxCRkL4hHuazE40l0pmDauJdAmQiZSSjFmo/EAXPImb+nnbW6oap4oNl2bYW
MUGwaOfbfDAAKZRM87z3GLjavtVnH3jEWbc5SR9slNBAftseA0MLnWO+Mr3EQTe9
vMSaZKX79KFsfmL1vYGUZCyhKy8K5kNkpvSauEHgm/8EldsrCNFDAmxpVADojWQL
CwHPlI1cNM5HjH/n55y7NNRx0cpWNOeQO8vv1np5YhvOWFwaNz4gXcsgIj1BjTAr
umUr1Z+hRrCJcwvHMaPpE1d4kYLflWXOv4Q5ytZklWQinyZwd/whRC7hFHt2ho1y
IJ5zDhAjj+fyltUcpTZQxmWyV3q+971yfzlJeBzfZKAXE6/l5YfJPslDyvF8wYGG
2BxVxx5N/sM48TkJQ9Au9ZlkS0NlYKrN0mmST8l3RdP/ByS8TiCJuOZm6nLg2WgF
VtlJlftJSzsxatgp7XmrWq75dlld4x+HEo/7x9t9TiJM2xqRR61JBneq+eAnp2Nw
F5AObdDffcBELKeOmJNcd7rpTOTAwUs6WUMOz2V5pp/xji1yjJLPMCuh5lMoTsN6
ThFFGTMJ1W4nxxiH7w0hjuJeNpU629/98CI26iYKfElTq4M9Ajm/h6rnNz+/bOeh
4AAuMoIZQahnz9oV38qFPuqJBu+wbpIKbr0HFD4Jr0mumsRZ96uFqaLFSm5NpE4c
xdM/QTKlNk8XCM4a29aR7pe6SxMe90rRNZxEl0Fv1riHRrGyYAIalLOSm4cUS71b
JcF2yB9QU8w1fn3jeVquCWleoMMxtRcWXFC5quPsxf32Bs8kJ0loFxIUbo83xRh+
KgZhkIlBZp3yCLDKkl9fykEOHc80y2rORhlFctDQnHqIawLyI0DQZMN0ew39/9oB
0qCSRDee/fms1V5c/mKkEnkN5zBG0SWDDCDy54+N0ljFEsNiMPIkFuhr9rSwMZG/
LIT9wMbN7wwcVXjpZdvdA/OnuvtvhYBav1n4J8pHxDuel2WL2PRmUOHS+X0oKnXg
bCCt7ZTgvOITvAiTqQirzonhjJU3d04eSbyg43PHX4Flz4gmVrHz7NARZ6RgweyX
rULcqmUj4U79MpeMedAwie/r+dHd+jv9EeVu4XkLPtG/tOpGrElKAK/YnBCuU9ve
nwFz4runCHaZ/ZhEqY0Wx4cxrbl56sRcM95C28Uq4LuhOxfwKb7S3nT0iSRw68AB
tTLhbL8L8/VI3fWEp9TWkUuAyetum6sA8V/kIpahoBPT1xGnkpim/9tUKrTDSXtX
Ijq0V1Lrf36KQgQ1/FqZ7Ib0hR1Fi+Vp4/gZ4nOI39scGOsQ5X7eRRWfL4hjwbtx
XBjDk88Rrq+ZO+j6FSCU0LnQZ8BYPrS5cOiuk7R7ib6IomBmDKNgktXV4IGWTV/U
prqS0DupSxUNjZeo9asUtXjBU0hyaQkLJx1pAAW/l2xn4CBjEN1vgsseyUxir4xI
Xy8nn8Ho7PCPKMRdW5nUSBN1Dj0NfbXTiaHztIlU+oRXrksOWHvULaNtIETrSSJW
KVo3+h3aGMAfEAcfjojluvauGo5rB+77mk5NKoRdt72cqxHGEvP12Wzo2DG8QB9P
8Lp/OuvbknYK1r+Sq4QV5zVq5vKWhUrFGIJF3xTtM+MBJjnvWrB89vlVc6yvAbcU
Nl+rbIZx41Ayf6jQ4F2k4F6wgxmr9Kr0eZMLYfW8deEl2RTWVbdnXOkQ2u7SANz+
iOHjbapz3Byi6BT242Qaz7kdzPbPklKYlUl5Z4HB//HEP4avElz+R1QTAyIVJIGT
uELS6DXpF9uukxvmbPyMXOljUZtWp9yseurEDZbH5U1ZsTDtekUsKhQykPwPr6Dm
2NMOvKShNtICLqwSiP7s25h1LXTKiUPGiZF7itiiJU8uBXlKnnedEH9n81O9ReSe
28spLZicRX+LGH6reY5hD60WcMZWHmxs41fdNGfWAVA+FwmJ06miKKCu9ozQkUnS
cKt156ELu2qxGmEs4grYDoLZ1hL9nTHVAY726CynFAD5rDzTCioru432PbVzM9sE
ZMDXyPG2XlJlocNfUoDoJMuUQnzzbZKg8J8vfRGmAL0hhvh98Oc6FyUdU+ow34Sh
9Z4pFc+1LMKzqKyFX+pSFVt4NoNTSu1ZnDuOZWZ8AWkT4McRNWrWcJVildTL88ax
+IJrOatt/GnUm9oXaTqTIyrtdLuKRx5IkhMLSOeXmGedZIovmsiqQ/85YKZ1uOVI
74zAJgBLTUhDuqC24pPqxgncDpWhyDE/BfrZ/PifGLfKB3lWrwMFRD0zYQxObjbx
HU7FFYjBeMzFe7H5ZGu57B+pe4JQHv1aj3uU1YkXYuzzXQEHMwYpNqpkm7zsgwE9
61F/AT4DGCeRcpJcwxRPnqfhjt24IgSA22/405VjCoNCN8zMF/VM63Z9VRvHXOJj
y790o7hdcxOpTVU2jQ1O7PL1rmyeAMwob+/uwyaVyAKso4yfMxcqLFscw/wD8nTn
zRrVsDaGeXkWwvTtvX8QWPm30knstAS7dSYaWmTxQPj9InlMDjvIdE+RGClntEda
ICioLpkAb6J/UKHJV0TovLAHCEnb5gST8l8GMMFBYxpEe9QoO0HSithwufXsoZOr
E+fQD8J1C+a6b8TbF6xOOgTekmZ5n3F72efrDQ0maO97ctgf9vLZKEdQXryXQcpY
PukP/bFqWcXKcdRpjKzk3J9H3F4xFqo3COQvXkZZD4x6Jag46czev0hcKIRRRMb5
1C61+k0PwpD7CCR9izi8fqrf2BgldlTxmhbOVZzu++IeeSspGyXMBK2ZsFzAyDRu
nKreeBAM6+McsSSxoDnZZ9q5JmSP02+UetpfRCUgaJVSnGfVHlfeOM6/Q07unIDm
mzHDo9NSiANyMZe6oRjixw5bG2hYw5sPXRrtL6mnDqLg0pFFwQb6abGLTTHpDDQX
pkKufFxQit4rwd/is83rpHqwnrE2HrTatH5X32un8yjw0UuY439nhwUaOYoxoWZl
EpB7sUwHwtdKRo56R5cUTaGpnZIL8OUpRMIJC7gObGZ0uxANFIkdY0VFn7wSO1qG
tUT1iTlvjBRzNgNZfQLXMArbTc+6wf7FIu3cCxO4VGP06r+oTnNa245sEHTU9qmL
v/Gbt/bU7VJz84nja36yXWzOmPH4bvcsRayUKOqkEuaKsSF3oWpdmKZtNkiCMqB0
56L+rxNuDF/wdZXUX8vXSph1as6fexnPCJ63hf/wch4D4yCquWLJaBEhcxTsQKfB
XGOiXGu9FbBhAXsn6KjmBoJSUkrxH75ARd+BkeWaTadBMo/Of4oXnbUn6ZWpvriL
KdZF3E+cPCABBJV2EwQQ0ay5oLuC/xm2bvski2pcsRFMbRFZVeLm8vKgm9SrnJuP
Ru+g/sydscf0Ks1a97Jv3FHkzdoCotz4yY5mkEvshM29vz1tlhJVniOCqYuPjq/5
yy8GtI9kA23OepEsa7z+GfVy9vSeTuV7+A83bOCAnAzMnHDVdkRHItvxTf+41GgM
pRnUmrmsY83dFb2eTC9cpiugQfMZ5i6TnX0UsYBTx9Bjc8wTh9r2w02iGJ4JI2So
ilGKS/LZJnHMy/CfOg2haOuaS91ZTG0E3QVVQKsk8d3uX+MYPtRtf4mDwlTj+ksN
17my8CYGYJNVuwqo0Z0V3IvWnRBAABxOZosAf7l0yvvT6BIzZXeNB5zEwum65wlL
dKyAOVZLvxY9CgcnXhs8ALpzSZZu8Nu1QFxgewMzEzS/hgC+Nh2bv1NzlmzooXzQ
IUTjGAZeyoq3U8KgcwpRcS3cNX1iE3iM18iHLaJ4DGjvy/SH8TyM4ZzpbtOGx038
jxTU3P1d24QxHq3Qy2f1hq4A/CtgElwIFRrhh7esGoRy1fbPZ0T6stz3Gm376bkX
rHk6RKPMuH5eat9tdSY0ngKmUykEYGYEAOp5rrYw+ozcDtDHRYewrVM/jIyKnu4O
zSYRLmsDu2MOgjTKB78xYFc+WJKElSKbC2EfYBkdksOhb2r5WRkSwaUDcTuMSv2T
avIjqsElDGuUDy6KCgK8VKpU6kkfkcP2GP94BDnjLQZ3E0NPb7OVT3ydDxG9RJmW
lFjsZSXpkC4HkR45jehSnpbytHOdZCEGrl9mXKY77VpcBXdXgjTW8woHhl3gkm+P
MQqXgjunAPayp4pYBQZvGLEfiFaSsoFRPSsSNSW3TL/JIxQ9SFhMKAogA8HE4Ter
AIfl6ZLl3miNEl0I0y7fzA1OY2ve5XmeQlYXrGYOStTDU9ZrvY5s92GZCFuu/KU7
3JIv6R9P6YYjxIIZYp1gzSrncy8j+3yKxbl1jGTKH8ahwZ13uBXUXyENDTxt8hU6
c3bluLRq7eM/FAmr5pZ4bS+YUAL2WjO3qH0w9xhD42LDsDjvhQo9dPaqqjVG5ePF
oBUMkCaleVosquNjlLbR+g==
`protect END_PROTECTED
