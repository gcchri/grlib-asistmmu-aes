`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rTbD0iqnfPDF0GOzlKsuYsDZhc09AooXqqTf9IVqQLWJfz/OpVSD9mKLYjG5tAnI
/KX4Ecb9IUkQv3j9JwW5hGYgRMUzacrpLV3itazYwxVccEajdO6FOibqFaw/vZp4
wffseLqFk5hVzE/kHWvI7MB2sorh5l7FNDH9JLQFVOEOfPzhutiBI4ZLXKiW/RL2
1kyhR4Jzuxl8oIg9qMjvfFF07qWym1Z/YxVqjfESrrGnuHgq+1zUG77D2dWSxYhw
Wn3uGAE3yq//rBUy+SY5tHRwxx9maQSiwYl7ju90qjVj8gNGDjJfkmt8XHjO3Uii
X1reWfgA+TR3WDJaRIGaJgiT+Ov1yMSsEPKk33itfvBGhZ6TbrRrwFG6V+1Tth7f
D2Cq5ohQst+sk0yeysRIScEjBuBAChymi/6bVS+QA0DsT9fvVGETELFSUsDOYkdb
La0oy3+ad9tnJEmcsinMhKUoXIakOqvGqruoD7lPNRWT5RsjbyKMGCiVK3I8+lcN
o4ilYXjDeV67K6NuQblISGXxO6s4B8bLzvIEqLUvJYIN7UIvTGf3E5UMwVTdewOK
g9/+hRWvE4FhcMctH+f0W8KXsFsDj33UOn6vS3zTh0JT+biCN/otfv3Xhotb/bPC
5ninAW27Oknut+3zQ9w/EA==
`protect END_PROTECTED
