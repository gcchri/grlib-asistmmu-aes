`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wXcfaPRHETnoDksFa1fgCI89fZuCmnCXzLs7SAjr41TBcrrCHWphl5cRh6QYEvAJ
q7WPtdSn8lyzuW1bORTp5ZuCLvSYcxFaGiN4c02Bx1qS2P4rWg57egCLm00RTKvN
jPh0BjBWCrHG5Di+EEDsFPgR3roZwGDE7+9yh/kqu/MZ111u2QlJP1wIjldPJ0Us
6hadNwlXcWufvHJRH7QW3EdX1B5rll3UbNIFHAiPP8alSHFeJZyoQTbpNI9a9tQU
S02/vaK/60vdL0ZEC2SiwQx5zYmsarwDgonKfVx6qVNilw5dbnvW5B1LVRTw7Vg+
V61ObNQ2pXJy5EAOheKJpRQRSp0z58JE0i9deyNK47gVoBAtGfW7hAOA8X8pkaV7
GnFNAdLEAI7t/wmPCuVU0s60m1eYvV7uNW0B3MdXgQ1rnFVPsDwMlkMwYUh2InRy
qsWGM1UjLUkEuCHRBE/abg==
`protect END_PROTECTED
