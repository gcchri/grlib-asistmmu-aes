`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aR8z+fwbaJL4EM+nmE7yQSpaLn+e63wUYmADBwnFbqOj0YTiHdWMbkH7n7wD2kvy
Tbqf+b3/3upUb6doqfVCUSz1N1LXv926brTdlGL9Mt+HKlB0NExUJMMs/fOw85Bp
KZ1k3xaXNmDP5sP3xhjnCUKRt3gJMErBknYIEU4jWPNwTfHhCJboBoROUSZs8ejw
NJLU1356Sxs0KrxmPK3keiHFXKhhHXHSlImvdUd76y4OUTHO3/51WLFG4THtHEh9
4GPlcQSl0DSdj2jio6T9V9DVHieg2z5K6cwuDyt6c3XE5tDtJg4VK4OeRbGy+jr6
7kCCqRyFkfoaQSGdNvQmXDdB4si/kP8iyiR0y7ncVPKlKIDN3odHCQAuuSuwydm+
jezTel8eyZGiyoTu5Gy0gFCZv5+3usH0yHUuL4ZOIZP2auZMcmD64iBHRa07IaRX
pXMRlK6moQdNC0D7dgL3JQ==
`protect END_PROTECTED
