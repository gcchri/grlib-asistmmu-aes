`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6caVs90v6ZZgbppHbDiPHiisswxv/24ktzbtPDkuFFXC8uaV+trrQIafzTElqj7U
fA8MgTZMqrFn/8+oIPAS2TkFpB7iOYZovx+QCavfZsBZaJaYkVEfEIMhy/oAoPSk
1get1rC1em/RhvQQHWqy9KbUXcLFsFuLfeFOT6gF9Bo46MTBGjNvGgjxRCQLYWFm
m3zRQxG73MyhwaqNyTIGoOv0uOFNHxz5v0U5x9y7ZCj0lVwXOCypOf9Mvr8kryrJ
1gM+mkHtyG2oWjdhPyoE8xqcTZffspKSfkvvwRo/sVHw8uCBCjPse3zkEdlpUfLg
DCN+PP6w/Ws+alulYF5x6Y88LFgdjeLTyep2olV7bNqVXhOVVcU57Ly0Z37GoACo
AcZ2ISkwcyzMbg2pkstdNXAI3JS9AQKASqix+UWnBcp4WTBOI9Av8AyPVqvoQeKe
aF4JevJ7BmqVpMjeSP6AX2rTpN2GjGsmR1lB7bmp2/nrXTsb31FQBlP4EylobAp+
ufXGCvJV3eURzAvWlFAauOousxViZ5UF4lNzZYqxbc12hWoUACUql1cvgNxjxHmt
n3yoWlJigX5CrwkK7zejNMR4WQvLrQm3fZ5NBfFgn9dTZXMfl3jZRDFKACuF1R+d
cWH99iwjwiNxksenpn+/Ug==
`protect END_PROTECTED
