`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9vGZfHH3oKZ9l4qihCExpr5UFnKa/7iq11BlbxubdomlOYzRj19VLH7WEc5nE9uI
YM3h15Y4ikLEez9ps+eYxbsVGGNOktrmZ3EV8F3q5vHRTTnBAJHAKniolH1w79C5
6wL1bKuPdU9D14N6qCPa1miL2HMXJHbCEHOqQBZkkxPe1Sk3S/rd/xmkPEDoTAKc
SFC/k9bG9HQImwFKCRFXBA/8sVqfxPnG4kY0+9KUnHKsHkH3LtcOghGBan3gbNK+
ERi4pPMYvBL5Xs4Q8gBUjHZ3ch1EcoF19REQXKOkjTa3yUCqeYoNxU+/kLhoflRz
pjPo45XaCtLPPL49jg/OH5ZFj/YmPbFxcozUfMN/yNxb8IgY2B4ag6+xbo/UHh9Z
snIEi1K+4HUL52dASJ2J2H0zI4Idyfq9S8ybHnUO+lLQXakTfZESvJ8L+jYb4pom
BBpJvESZA/muPSqou9wKyi5Bc8NBU1JWWkAWQ/eNqIDiZxyAPLA23ps0gS14dzyQ
R37bq7gwCWOgxIxLDuuvb08vhoKyR3MdbBvxoebXLCBXT9JqBq7NyxyBSrmDaAnV
`protect END_PROTECTED
