`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iUPBOAwdd22TR1sjC6pkbiDqR9So26VsStLTx658ecl8dCKVbCmZuqHH00gdMT2N
xE4nER3yhc8JH9AwLsIkaoHhnZDdzZYXvrT5WuXrfH4n7c5qBD0rrWC5HNzikiM4
wcPGIclqjZf+2rjuXGxvH3Vv41WQUgZLT9jYyxsxLdGWM73ktI9o/RjJij5S12wA
JrP/6zRm1ZFMUUFFHD4OMRnyA1ghYxeD4UOAqb4FMwoYtFNipPc+CSU7RRqGL+62
4ll8qVA/EkXoQKWHFr3IVYGsea+qkbYuB4vb96BwuvoGBNOPEIUvY33pm5uY6uvY
ek8pA2bVr8yd1bs3kSSKFZFFj8nAgBzRZvSKSSUveezbECZft62BJH9De915hlud
5nYrryeC1oevQKrhluv5duouKgC6tfoKjniYurVE8thpBh7jnwyQDyLYDxtYk9G9
OJ+vhyHZVBDBc/amoYnWE5623exfLksPHc/43nhspBqj6CYj6mJR7bn0Dy0nbInz
vJg3fli9HgwmqgVoxmoQ3pbhaf7ms7QjB7GPhFQCNUSrCxBPq7Rs9DSHl3krNZag
PKyqKa562Varl+VCVT0CIfO2gzG4QSAtpINKvc7edbZANwuFjv0MzVeVHNnNYHMW
MxIOZVbQkoT08L2HEvKKtEK+knC1mn1THvvTHc/owi4aZEbNRUPY+FeghzwWGah6
hz024HBCCRdmicu2BRxHwVFN6l1/8B/L5uuMGpiqKSUlBbGBAuc6mtANtA2WoMSK
+ibTfiakTYxwX/vX9/0qbC/IFXs2mX5zcJC2Hk7jGZil0FchBePW+fbMK6nquh3U
9CzcFDTuLpuGd2tJpzylCGdmqc+En4x2MFufuqCB/j+TpglE/fkTyn7fZfg8qeSl
n/So5URDdLv109KoJ0mq/noio3YgP35UYSBihJ8Vvf1phpZW2gudJ7+hl+hwZCVC
ZsRWBk4DVQ96KZr8wlYIikqRza9rERkZFHQQaqhlQ9Ir6+HrIi/LZ+kttp7ZBCVJ
EvUhIOO9LK+F/AIeeG0J8Xsi7O9UnYMkyeTIaJykzwV3dk0wOw2cFNczaTGJuR29
7009OTTDVcmKOmrkmcwVpU5pMTH2ynkUYq/fqzqOnSlKxmW4ilS6gj5hMXzPxPqU
xWW2CXnaBZwG/nc7z3ILIrbdmT/8uZ+DdNVWFGmj4Fqku8Eu8ZTyFGQFQOyIUyxF
aDxsG8CyFCLRv5KDfP1hS0plM5MDIFNnsje2itu7/9CGXZlvbWw+y9U55GNEdzvO
FlcsF8Kb8zP9JON6VxZm1PwdvhJkt8fSWi/bI81bNebS0pibC4xhqNHHOU5d1SwX
ciRsqD5sn8n6Us2Gq8nny3wqehhEbWZhofu2c/sRnWqLrQQCt/ZzTpDjPUpI3k5j
u4q29oYJXxxNIC3KFh5HpkcSw0s3btH8hiYInbeT/C/aeE6hIzfGk/sA1Yice1Az
OMiOQOSp9E8n1QpwYru4pZ7NugTxG0JrT5xTTxlwLgvJSBcyE4/cwX1AIEVZ88vI
eaPfTlkLpln1evIwiIRcnAVclxvvSeioCxPLBVqsydcBHV0G6P5kqVEhs1QlB6mI
xJ2Tf/ejnZocP7S4l0joLAdiQUSNy6xNH7D/17xvWvZaYMexDBHy2RQXToyEmTe2
pJygYGHLhZZI4nMUxayBTrR4DbtSmJwITsestT6lw5xOnFR/uZLc0X7hU0vDIaFY
TIRxRcoAxrMiE3oWlrx6R/Crzy3RWMScS3FzKmItgdI5vknp1No1Q/m3/LQefen3
LLF9vJtNOIoGv5UiTT74iQn7UWr8FJGroYBJznWwlK2elhHQkvkfS9Nru0HeDefX
y5Oc54CGunJFmRmwAau+Ups+2ZwPaZ3kEbwROl4Mghdcim54TCjc9/HllnRvlCvQ
slgpYf8FqLCMAvUCxq9tSxqGUYCfR6zuTz0jC43PXyOqA38kgvKaTZIq0zgJcMwT
GGWZKq8g5qqDQQMaKTT7gtaOqvP+65O8ScOtHJAdZVDfWbO1UXqP3osEebj0TQeZ
XByRClf1qvX/iV+67jEUn6gY7/qCtouWwViOZJO4LCcJwmY5rkoR/0XmAXIACmvi
d/ISvvmC4k8bPtC0K+FSipyPEvlK/gq1VLVMfuNEQc2lpg1KU68TMEdoT6PlZ/tK
EoFtLJF3Kdf1P2R0n+EM5t36MEpwva7hTWs4WPnnp7UKc9sXiIjEkSxGu1pNZVp8
6kqrIqbofucxu5sbHS2HbLE7gWkUOFZoR4zC5Dd7Uo+cMSFMnc4O0VyrHZQY0g55
cm60O/JCvHBQYkool6dhZPKlJxiEwRgt8iQSoagOCnGMmKXmnLMOa5p2n1hHHKzJ
8QD38XxPKxaDjs+VTmyADAvGFgxSrITVRBEUmEKBrxMAAh2WNHGA4WlAKODo19rU
tSnOg4v8TCsAvyeduR3wypR4v450PbopSAXMRCAJK4ZolOMblFzlinKiiY6OBqUL
P0WaJrOB9ui7/iWz23YPDE9OxzoDq7/RiazIr2cDEZwWvh9mcFEwRr1mPoVXZhcK
X+nP8crgz7K/WkmudZX8dgwEra/ybS75O3eSOjyUeJkgFUQV654vf7zQJ6uW1SrW
o/GKec3d5XZHdtsIQjjp7KSxFzLlT7cIjy1uNzse2mPyNHh9lf7RvPnOvcGciqW5
aDYwrypkj6gbJ9E0EsSlkggokJ44mEQF63AQ7fTEhbe35ANf04ybWknKXTlJBbZn
Rwy7NuupPNeltn8AMjujDqFJX6RSGDDIT3S8MoxuyrvEQtVglD+JiwpaWr49h0OU
vdT7OdTvjlXvUdFn6Vvr7tNKJil6gSqi0ZhFTkQfN+PqWsZY87w3Yt41hMA8Y3LW
Jeo1PzGBdKKUjLbUIG5eKkk8g0YEe6e7tbU8R8Tp4bOq2VhJcBY4bpqGh4RKvyHw
gm9Gr6H8qIROsyicpV4h3sK/OQRQwzbBdChRibyATyBnveHp/pT5ogus6jCXMp6V
HzZyLI6e4ayq1wDaXvPpNqaUfbVgFUNjqGRqBDxuQecr2pzWsZu9TOUUlnrHxR69
G8NQk+N3ZU7H58ELo6ueQsklSnFKvxySqxs9sfZ2keAGQGC0z+vWdYUMOhe6aMNH
q6b6QBB/15Rngyh75d46Lo/L8TG0rw5u0Mt3BdtNV31LMMmFfPpdWJPVmRlRtlRg
xW/sGHEzLO5NwEcmKtOPaX4SxxxkRkhy2EuqHx3jVqrD0KMp30BOiQvCnHZRZ5Hd
IdIF9a0AYBnMvnPq2s/Uv2ky1mgb9NTN8U92XOVpqIepFxAroxnLvZE+IWDlW5qB
IrczO6Qk08Rdnoq06q3234sbU7iYLPPLK3plOzWU7XOaWTx8l3zhzLXc1uc7GTQx
ZrKz9kzUEKw4AMNnHWIdtzMDyOYRNBtw0jelfNKLXsNgibR4V/SL7MkUtaQfV/zH
x666ub1EKFn+QCA1nrbMF6A70h3oVQJLvZpKdYeb9QsQVNCGPFY7lPCMq5M+S0bT
tFkX1cFYARVJiMShlwTjMfYbgoPOoiRCMidTwtp5iStqxN8URBk++NWQAlgmHcew
3nentz2+OIUSKhq2MSYBtn9hC0g+3vj8NUaa8W2s+8taPwfvAA10k2kEn1tMMwky
NWB+csCA+WQ0BDQC5uAV7jq1UR2TGTqpdp2Ax194UzjR5JTcKalqrYljhGOUYu7u
VBqq8Jc14VNc66FQ81hEjT4TGEcehF7SIUYXK3ugM+yvpRe9x7NEdzNlruQ9jb6Z
SseQwSLWaLAwHzk9PVrMy5Pfd0CjyItb4MnJe0oTTYnzYx1dipIj4tHcozSVnNAM
uWt59SYQhnQTUx2k5IDOWWpk2l16divrsiV6VZhR9Y3/yEH7oW8ZkuaxDkpgijmU
zr6MfJEborN/Jaqqav1WAAKJYJpJez9BDpEv794dSaWtlGejdxdbPr/pg5llX5SM
lw2bRI8Gcwm8IexFADxb9Br6VE37Kqr5hJ3ms8XS6SENW0sKDqUoxYCv0FoP5nj2
Jc91FWyJxF84MB/XK8Gk2otg9M65h6Yu+Hpgqw5abhswO7FKdNSFlzJXo2CzZbk7
wgbusYBnVuZReOA2ilMMgNIB8CNZbiwpW7SXFo0oeqjr60L1nUAYfh3cft2JvFuz
1fN5GMGohKYBkkDcCam3/Tx191/v58OWijfcewx0GIJecWdKpZxfdgx4nJ1Ehlzi
6BA5/aJRwV1/lQEKievWhBQD85ZOGWNpPIgpNdrwzzFE35hfCCNq+zpw6eQX0DLc
hkfJHqefl8qCL0OEJzJWHikJmBOeU6didEKEVhz3eAFgJlHJvJ89Vk7lRNfBESkj
/r6wYXLCi43abHdC9oayugoos/yZ8L391F/5CfAJvHDXrV/IDx+xebrKmQJMNXdL
TGp8xLnD+oWKcC4fCKF4vFeKNlt1awaG7zB1eQAuw4+1gCZ7fHiN/bikcSfkl2+L
8sbdgtaO/wUaMHFjVUJ2zXqDyU9sAVNpmCT2kFxSzIUAwAgSpRvDZxsfcWV2l8p1
NvNIXLnUztvUuJR6ji8i4hDUD7DldNG7giUt627C3TsbNGy/aZMsf248y7uEeTKZ
NlOkV4v3P+qdUbvSpUzCM5BdYGL2LI0oPFOtU34ORDPC+3x8ImZNXCbFlLNN8MrQ
U96SzxYyEi8khcJo98SYBNt2U7BME8GLuvwTHwKa+r6ATpx8PjN6cAI3eye/OMA8
DCTKOLNadgEApjuc9xO+kjA4dtq2J8D1ZDDJwe8BBC+HxkQs79zdyp+7yAxMqCov
JAtg+J6RYNHHJZ7lmdQPkLt6j9Ja8IW2kshfh6QG15GxeQcAvq00RV4teyi4WBMB
K5eqPCg7onx0Y30LJutmCsMxSjK7qrJFC0cqh0dhdWaPf5grteer2xRP9H6XelZn
dYpNOwRslf7Y9Jf/wYSAPWfyYHAPANsdEBPQslm0duqkmWJRRA8HNLKYTTi51wXL
08gT8nx/sSv1mwTtG4+d77++8JfgZ//wljocovhSO5q8es666pHFmKu/lxYBLW59
bi+bqtxU3NTzPjj8EBsnATXvAxKoOq4f8IS+JY4lv4dX4CEZ7HaginD5ooKe+oOU
UlbO44iASYLI6GYQOxMzSQibNLW2+C17hP8jYvY94tt08f66EtDifxVBrNsN/tAp
ud931ZGrTTEWkYmqzNpy/pM31pfXp7n0DQaSFd1B+ssMEmIduwAxMUuxYkQv9AGq
HqPqUN132jJCnuMOGD4yOPDViSPXYR+LpcYmA1Q8hTwj1cPEIfNzT/pyhZSBL+5o
P9R/RZOPdAUYRN/AFq8UlKVUP+BvkckpeG4mYWn10Eo5wxHv3vhoNK6iF2q0l696
dBf0+j5NogqsMUvhwipNYFaoaiszOMV7NYAH3GMhxPyUss0jiAJSd+4tdYPu4ClH
SRKob0adQNKfWMZ//SUMX2WD3Q0P40OCFSCUZzDv0ppayCAE4rQwJu++DfMLXoB+
gi86SVnygpsSm4JyAiSEvsB9E4ZdKArb9UkMu9dNNVHsTsuqVPRxfkLmX1bhRADr
WXYcpGQLApJSy+Oy58tixQzz+cnqjvxQnf+IeSXrEkJaCYtcTUpJAiNRvWpAvNch
sdFmi3GUZCJ7UT6rN0KnuvkQhEHr/KYkFQcBka0yFPclE47jbPGMkDY4DluCWYdS
`protect END_PROTECTED
