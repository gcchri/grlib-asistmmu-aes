`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zYm8Oq2VNNatQ09Rnvcq2rBLTApxpN5RhHD9vNCAMTG2cQJXwVn+Eh0DCzYL40e+
3tyAs/MJqc9xpU6WXuF9wuLQs02PRowoVB5zvCgoF6K3S0cQ3p/4IdlmHxGRZAcw
c+OTv/2CoHjB7Xn3NFOft51VWNp5pVcyfp7ExdAqcUhBR9xWNe1qhFFRCNqkmyg+
277Eut1nDm/ffPusT66zYiPAPcZdZuMuAgDN/70+NkR9EHKL4i8mJvmna0yEpCDk
tn/dYFHEi9tWvartqoJqMCmDAgTNrLrGU6j8W/v9LVcgk50qHNlLu4DEQ6hMA4VI
Jrgf+HFr/DBt16xo/g89OhKWj+fmNS+tSLQU4fqLaEHMiuAmUgrGuBxev+ILwy4E
tgwcRds6nqeEQsekP78S6g==
`protect END_PROTECTED
