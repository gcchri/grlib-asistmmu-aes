`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jjp5OJiEJIpqtcIbSH1x2/seXW0LAqQzPEDk0QINm0zimv79CR7oKSRHz5QeVjvL
bF35SGWMxe7619hoTfyKclOvUurXQli9z0Qi8ug4ZnvsR/k0egd3F831wn8A4fSx
R6+jhAuUir3iU0fHSM26ZOaLqeohseIePyS8IpD2l16Ym9coX62BS1fHnLgeFGY3
rHp5rp4esTJjdyy2lVv5ek/wOu4T5oSRLnu8+TPaKpkSf1bNHRVCWCNvkA96zzng
a0zvurm2Dejv+SedCS/yKdoN3aPptuSnidf5HPPLKMrmjI9PDo2DyEqzVTHwdL3G
jv90jWiTb6FYSBVhhh03xO9B+Q/pScUW6RM+/lMV+uDhPzLknk2WG3H/V1Vk8KRF
jN4BNiSEogl+Xit/ew1OOKq2mB3eZn271F4bqHv9pjHUo6tbldBZwdPfXFdimHlu
927Fs6G2CmXmoCddCu2McxA6rXjGgIJTGzxyCigJ+dd9zs1qCC38P1h67SGtc9GP
cc5HOISrqw8Ngco5vtmQeadaJkldAeEc9G0YQp+1RfC3u8vSZFi80QTY8jbYdTPv
epZNLGnJB4otnWZYnT4qNGtbyVBJ5xpzoMgvYRML5xWtLMUblrt29XTmvCaoiyGx
zyVr7wEAo4qBPSZ+H5Y0WmYNVpCjHEAt3zol6QnMFFE+8Uqy8xXvdfQZjQRkuPiy
YcODuNu4gMlPmZyz51YimigwAXN0YAEYE0XdYHgx0ek042ZKiPMtGJ+6bvkKXjNn
dlZRdyV6zwvEh5Ubm8qDmx/9Vl0lLx2o3RrtjuMflZCtjv/XjDwFqWD3/uljXD6o
xbETGdW3EX8VeqsFZUAS8MNZjblIEOLInoYVPwLR6mN/2cdREY4PeH4YBXj0YsWA
F0vMsfj6/X/uDWAhUdj+m0AsZdzJPJsAPgYHAmtldhbN07NEwV5xxdYbXgFduBAY
lUyMjLWBdUZIpkrdfI7l3n4lBUweUFd8+Q2y3S8hamKWfuyavPuPsVo0v1yDbe27
vFlaEs+jm7OspVtGR8IVUai5Yfo3JryXzx8ZglR8hqIi+z4WkYJL5JrRzWJf8otE
c+vzcxScbmLefO9Wdp0Gn+2PIniuwhbZAp3KXrAZFMq8uDo7LqpcAT/8jDlv1pPA
yncrCxXI26zGpfkBacyuBvmcERJvClkf5+ps5G+0GedTVXT5vde3JO0CQioIP3+p
g73sJEBQuHMoE2jIkjZ55Pa+vq1Y/tAHfB1ZTsz1wS2Q22GznhdXU8Y5AIcRiOzz
XuQXSGFjq4xqiy3pYMv1Dy9QU5IP9WE1uDpNt2csbss8QQ6PrJZsIVEQxR5xnCOT
UTaMMMNoygxcm+Wemc2muqFGmXXoPGLeuBXgOMonGnHMgOxU9e6EWnPuAgbRYlt5
67F0Z1oIgoB9cgKUT0+EpDnZkVB7zphFXw/muXxWhmFKMnsnuU8cLQJQuHsJRP/8
Ldg93GUkyOWB9oYr8mi8O4Nec98vVXd4AaD82cjEAtM+TbiHG1MDdfWjKGOe3j4R
eyWj5v4ib2Blq1C45DMEwQcpzBNP87bqydjDChkMo8u+smi+aQAExInXEg1rHJGP
3yIm2pVTk5m8cy1I+x/eEcadsSXBZTolsM4It7HH99kBGSRNP9c0Mm8gkK3XTmvn
bc38OqihNkfxHbH5+Cu8pza58QZT2C0XRWGVTVV6+9W6XfKRXI+9deJSQi3TTXHi
atPrh6TmXBIqR73fBEkasmoTo5TF6pTq6R0sMvgCt69Jvkwlw5KaQNClNN1q46HM
2foUxjkABoatjSBHi4Kwk9VO+UT4byRZM/sZEj0ZN2b7D/2t/yv+swWjCcd5yFhm
la706xK2PJ1tgK4J+sQK4PyCVefEazFq9feSLdU8L2JMJVcTDU1+N2zNvxdu6vU1
LcIpFjUBFi4jdyvBACB7U+YH7cCJZir6P8r5LYHnaYqyhM48ku8HxsXsWGk7UIwk
5j64qZ7gEsOhZtkTHx66JYweFgCqnN2DdfW19qqUzQYoMwb/45D/JhTtKbRD0Pkt
d+lKnO4SB0LafsTu4/fTi94ML05UsZLHepYWHh2e0M9ut4d31cu0aB/Tz8KLTfRR
daQeyMDvbYvhoa1uGYv42FyHOPeBJrqT4eE39JRy65FoSFjPrrVTb8QD/Cv8oz2D
UKm5zyO/CWXJGy2Zl+qCYK18S7DVLiQJGHj6uPwi7RXrQE6PbiuPD9ZRBOYbkIZw
b2fX6vf8YiBU7/KSWfViq5oa/APoyRDAPKWTzob7GhSGW0CzxAPFtdamKoFniMd5
yKjWx3+cQFAa8KwSMepjwwqslJaiCcSe18gQgkRqQmuUj2OP9uXwcFiX2wKk22Ez
6pxxV77e5lYT3y/KkfLV00yFZ60A7E5fYlqZdeB45OE=
`protect END_PROTECTED
