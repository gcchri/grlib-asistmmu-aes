`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bt7350qPJGy44Y3CSx5sbTngzfShXPsPOoAfbvXJNCxAkYoPryRlB1HwKSo1YKA6
eS27H33eWLVzpI6KvTD/zHU5XPxJgyBhQQeGf3AJyEwtZIpmsTd/OUc6+6yYMm8a
eGMpGCHou5PAYHk3zNua6M6tCbw/N5AC4HimvcbOe52sVJAAQL1QYvzaiZna+C1H
MU1UMXvEHSywwfWUA7CDa8+TGCfmljv211pHfW2FTo5aa7uEVMzwbGsauU9e57z6
gepuJplSFsgkz9OatJICQGWipc4TZs5c5H7kRnu5Xf01IeiB1hNxwqwt+0U1lJJD
NPzW7OA/ce/D2PrY4H93GLOFsC8ndsorNUEjsNXKiQpb7sIybj5H23628A4kjDjM
utUqtzLF5NeZJClYSttmgEQ8th/6s9wfcmpYtWp/CxDqwRFI9sPHaMZ6CeesVdNS
YBUVaEhkbVP4GJblfNJMm5gh3vmInDQI7MUAtC7TFHoCTBRSKDmGOG5So64kkq+N
Efwhir3W/BGmcapDpu+SUpYIuT/bIJb8qVIXKbCOVOav+gl0u2WiLP9xRl/5uDK1
p34tDAPQqwnEWeliOKQQNNT8MQSRglT2VgI0T7sVA1BK5JHVbe5vY0bD+Wp6R1wO
IMzMr3lrCMwk2wzjICGdbsESN9bc7EE3wrwV+9qwcp0OWjlApmCqf9lzi/mQNAhB
`protect END_PROTECTED
