`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/R9jz91JsfkEZU4JTjzmaaYn0AQ04auWQVJCwQ8Q8PUrcZ9RwpnsOQUbQdbNN5Y8
E0CGdomBKuGLKbG/IjKqV9KSDM+dfjyCvndumwB2mSOFhKvu0CFyB9bZczPcE8pK
SLmkBezmGSo4/m5PVrf4AUjpV4ysQL/sPeBioYLEEkVlpDrzkaYyrm41smCMIFUG
wjGOdMOqZmrc6JpWIz9omzeOyQqGXcIMjo777mj+3ikSQtJntdR10avPd2g8dkT6
1ZAHe7uxO8J8rAANpLsUdk1Xmp1UbmG4MXBQC3ApisWc87zLMmJ6NpdgKBL36nwl
8euDTKLy7SY/aLdJX3X86HIskmC3Bs+kKMNL67bPJBWbIk04vHsjrIYVFqfyhYFi
Un4AysNpyyPVGskzyBGW+K/1OZjflUYpCuFhLo1CB4UM03Cc1FYxhkq9hEABHGYe
YqHt4B5+xgbHWzPCmwndoe72bvcvL1q2gbMunwXm8wLA4POpbcTOc1gFATpERgMn
X//60l+kDX+MkPo1yWM12Fgf7G7eS1pXTOGOZu3CbDfaDcn5meKPHs0xg77OOb1c
ZRMrJkZloMl8F04wfm4XdPvKI2Et5cMqPZk4UU1liPdDLdHpDgBF4C3OdmPHMPAP
aF0vrq8cUBlbUNHz2Pu1Af9Xg/rmfud4tv7stNEdoyZK9w68GKfyWX+om/CWw3mM
WIsJ19Ql3WpYYEqspqtGht3bKQCydiAIvnm5J0eleuukGs/PAF4az1JFJeAYgobq
gNnp7Gu2HY03I3e2fDGN7BPQlF/f5ptjtHrahV2w1TIN91LWwbCexZq62r86Y+9g
dpju+XHsXVw7WeoDEedLuAsE/VI50Hi6PsX0EwGTMHWINimGxORne6wd96RK2auk
RcDcSeCmUN0X4PHRNCNWG6IbtNAiItiV+wbfQPrQ1Z/QgCLwWDIc9JNYPmYorf/X
wdhCwDOuxQC3c+uKeM7XJKGPJR93+LzkN4epwCx8/j4oys6cAjAFW3ElaG/VpTzn
XpsVsfUWozX7WlTGXopgjqIDood8J2nDngmY/JwWRBs58X9wmqIwDZPIR7WlaTcL
C9Exn1UOzo3TvGYxTMLiagkbDGmv918nIazV6ZG/0lp+HzoPyzo4OiI1bDyzjRCM
xRCZ7L+y0ObbjDpsZS/oZbJ6xYULBiYGfXC2a5XusT5YtENsU8RMDI8NWn3M7JGK
FpupqpViTTa5ojIO+pp4Qe+IXAZ2NktXTxDnMZY/UGFAtvSoQuNIbxFpGIxyu5Vv
me2p/g4fLGH28b7ot8fuiSydsGSoU1LqaAqnSUDF9Qwt5S+6sFcygUtZFbgVATPV
JPtK2jqrTHLdfK8hAX2HveXiXbSt3aKP/Bms9pyalIXr9PDLaFraSvA0o+Bo3Jsi
pf/5AtmhHOwJUfrcziGmOC98V31NjfkaAPK+0pTx5Kx26znw9Uz0pA+tiQLRrKx2
CZHI18DcvaCm/9Fbn2kOMrEFqzz4Tu0RU+UpyJ/blOZRVFfNVQ4vbQ9Eli4wv/4E
EpBwKgklOU/yq840vsHjYXRUcLw6oKvAz81nPRtVjzQOxHhD8JXBIeIwlTSKR6RK
dKOx1jlvk/Hu3eixi7uaM3jTaMhzBNAYU6MJOguJi7O/RPcI7m8MwLEk4hqBUeVJ
/JBuWM6/SDzwxSrQLBZj/33OKeoZAAZ4IvKwyTqDdno6sDsXrJHc/YxNzQOYRSMz
TtYMbnO+TFTW3hl/t8MvGePpvHzIfG1uk5uvpoz9R9VrjolIeV/JtzvmO0zTaV4C
XxAGig4lVD/UvDTEiTNwdyQwdzh/RiQnICgCzDSgWK5ur7ylMWkhDaZUZ0WiNMcT
AW+D4n+udTsGjRonM/Pi/80F/C1XEJqXK9Bb2p+LCO4gQAfC7I9sHnMmSLhxLBTm
dgbQ4hi1mH/k7KYiX4C8pGpRe9yGvR7fshR1Ga9AA+62oaduvhj/7O0/RAMZVf4Y
B3IVJ5BH7a7IrTNN00E4BkXAKcESuoWT0pwJ8GxYsBjcnnLeC93gmYbBqFpbWxfi
kx0XoC/aypSCXL/fPj7g1cOnPMyI6acJSZ7IHmDluLe+4FIvG70Wvjqest4YTk5X
tiMc7+d9RW62cKkxHEixV6dQtGVa542jeZFYuFXOKLYyB4gMUs93CHQkyx+kI1RM
vOmspk/lJAuCcFRu6+/+jwFlOB1NyQQib80Ha4YkMJlOf7k/kVzK5p4JLzOFELy8
FgsLb3ZwxVKWVCJGe8qTee/OZ/DD5TpPUGXfwWAyE/Id6PUn6VkmmBOK0zMkvnUs
tRVxhobaWQPrQh41hsxuyHyT727NZcZJ2CMoXRCF32brq5L+ERhWciSZFOCnRXgZ
3fla5rmB4tsKGGPgHTL1zWFm17T6hLNDSUVe3k2F2do+93/OKjieeH870FXv/Idk
dmV7Lhq9h6p+L4+LTQsVhLq/EnpXq5gJzHuTVKQV3238SsQC+R7AV/t9PQb8cU7v
qCuKgiel/5Xo0+pJW0Zoh+fqfLwmC8CXeq/nS22hX20D+vZxJqqps5OSAkcFQnTK
OUcgHWq9p+0ds78bvrWfQuJNGG5eF3JMMNtJgd9RdJFZ9j2nHw2F+vMbbAZPeUgh
wduiTNauJ4vqKnGlLlxSVHlCSEV8mdUfddDKtJLWFoxt4EO/dHdvaYna+drnp0fE
I9fG2ASmLGC9OxZLOMMrYa2q3/9j9pj8WsHvih3MJ9is92j7hOIq77yLXUlVYqCq
matdGYSS0CkEtZBlHDn+eUm9xas9K65LpvubRqSW7qf4xTDt28ZqM4r8Uo+chuw8
LhM+dv5BNe15h5K8Ns5L57bFGSWpa5+B22UwHzn08Kz0M8fqdnhNG7kM051lwAb5
wGy8dRBJ7HXy0l8XaAiDIui+AKiDgUkoy7/7fJG+SXZHeqv+zDiQWFbWIyWcrwYR
s2U8CEt4a2FpGaMP4/e8vQ62QDRid5mUx29AngEBOG1sRPwnNvPxZdulH5oQNKnQ
iRYCkcRkuUHpFz8D9rOHv7GyuXVCE/gApv0RLgfW2VKw3lL2/ZZMrP30575/Ceqc
Mvy+WK0rnh+YBgSphreYdvJBwYfk4JCi6JbXReSSYPX6FSiEcBUVOGB+jj6/cxOv
uFokiAU2cFZE4tdeNbjaXnBgTGze7fkGAhWLhRF1X3WwSyz2K6O74/UVqOWfU3S6
PbOCBrjbHTT2tL214y3dDQmhcGEBU69fkfekcXRxCbTnKMiRmx16812RCRIoaIPg
nS44Hv7xgQjx4oFn5pWivL8tpF+fBBH1cTk1z32hJBu2NN2qhRB6/4xqp65fQvax
W/fVzepd9aq71Ij6P60dExzeEzf1XuVaZjeHqc9ECnqOf+Cm80pMn4JAmZmh4ci7
8tMavXeVAjWcioU0ONgza9tVmGJOM7S3hrlWgByJ8RV1o6YsXWlUHO/Vxh1EDGMY
n5QLnD3sG+XgkgfUGdfmbSbapY+eKMvzSe94zGjm5QTSO38Q417kTIJvs5cRAWhq
88m0GFXz7GPeR8TgOGVkSfwbtqA674lDRT8+BBaDIrVxSBMVKf3GiwG+prPbIKq4
pA85P+yfeBFnyaNo2K9QzXsOQgPeq6BXOZMBUMxQjonWw3+Hiz+prJMKwFv7j+aY
OY3Q5eiL10sFMGQVBSIL2UoNVYt4DqjNck5ob/hoMMix6WFZDlvXyr4PMmKDqlxJ
HrXg+k/og53qoTnZKmkMBaPdBkoSdDxf8PVYH4JdQYffhD/JgMByFV5zL97XCLdu
0mLGBrYRxU2VQHto4yc8tcjkC+MkAz3mkm9nA7QNQ1CXl8Tv9ghABYkO2+bDNAKc
3dYcahZrVWmDMutxP//Js+QZbiKf6KdM7KIW14W0F2WyeFhM7iMjUxYME+S2XcRu
/PfAbil8oyjDEq7N57Zmchv0wVBwmyJznm9M+UChbu1hHFW2RI+oorq6M9IKzBHX
KtZ18rONdKj8J+zfnuwsVlTvKdkHpHCYdCn0x1r+2P80sdLj5cQ3oxHyLzOAAbIW
Ngd0/lCMupMKE0ERWh3i5Ui8o++LULfun+8n1efBIUWu80f9t0JsbeLMufvjGn9Z
XOH6tl6FrrXb8ftLfGoU12nMwHENxa05+HdNx2/cPOKRq+DvJyWWW0GpLLHdD1vL
R0aXnmfY+AZVqs02wsopQrgNO/vD48Q5PMWSddRV8qXID40FoG1jHidKmtuC3U8o
S1WhgIBDHHEgk0Req0CT94YVTLxt3btY+Sp77ZyOm2vWA8UF4JQZ60dBcnAE3TtR
AJ3HzNgix1vEM3qtj2RWfpBjRLdNyZ18LKeI929dSe87DyEa7CzZkUuDs2Sg6kf7
QWDsYzkRKhF4/AMtrMCmTcxEX1BkJ8dNcDYjVvSDF8kowD7wmyxlCLMgOghxUjdz
/phm9/zD+6gY7sh0tLJkpym+U8ptXE4spPA7i1iPf7BoLvAXaWCacljJaLtojqS7
eJ1bxFuFS16LQY8WN7jIJ36eDMEUTWjeDGVZhyvKsWNjfYy0a1GahrylfjGPdNh5
KfN6Pb/5oYOb0xxVz7EtPEgrZePUFc5E5TejFBwOixVLn6onYjVlG8G65L/RxhNb
OxHy/iOmzhlF018R97TW/xsWWDN2M0gW9LrWIKHOFfWBdmdegMKOq9SDYo2MGI2q
N3ynVnfut2TC2uLSYdMIwCyfEuWXaZ3bPUAdh46zZ7p8xRlp516VPM+4VYT7oWPs
EDi36YINqnLpj/pd01dqIU8p9BuPLqqWIFepnT0Y1Ky+/WjTDpjKqpKJqmvbm4SR
YpK1EnIWHg8/SwSQzru/Ov9b8CvghcTxCaCwu74hfoU+1CdrzaMLIBNNszaUJ5mA
hoiirx9lsWN67GqC1vaIWVpfst+K0w0JgrbHl+M7pxapLd7+/zx1IBJ9bgmac+Hg
+xG4c2h7UbIIKTkXF7oW91TEEjlgrgeOXmIKBukO/GHV0eudLq9GZMvR+cuWwIVy
ZOpUeSms0OpZkEZX93v64fW7vBElR8Mm34tx/cI4cyIOi0wNVGdzE/e4exlgjC9w
HmflH5w/jEVUKn2IjzFO2uf1n0JskXkhuWLRE2ALIFXb6W1KiaN8L3r7lb+nUFQ9
geOPM0/8zi9CKIqfWEAeIedxY7OF06siWEC/6OMNP7JD3JjBvbONm0jwBIQYpuin
8vBUgQsB/axVNlNyzN3jYyh4c50cuGxpkFUwoBNyf5W++Hiqmv7JNy0r918ojyIg
WUBFlmtqf0EMfRZBmABz2YoHEq1645eVHidGm5LofyIHi1MnXEMn/jEoX1iUUJfp
tOoE47w+Ec7I/ZGifmnwdIG2i7Fz6eiZtnY3haBd16wZYImM3H8ZfINNihG3nfV4
l+usk6TNm9JKOhmstGduVvYPo1zvOfTVMO21zx3rkr79dvTRCIZPfCKLgYHUPep8
oH6uovYiimONd64mEK9Q5eAukf6JH84CzF10lsisM9iIFSeqP5Et3v6VNKmdCQlC
PYtecLuslC40hhjMhG0jc9J7ZECNViC5yYJ1eYTXM22l4gsu76NCSdLQG1QjtH3t
rSU2UetfpELo9hZ6/2X2H9F+l++qk3N9/ekVBIhhaejc/2IHwFDzB+AK49mpxsgT
fcQTZbCe/zbkvCJM1orIIbJ5QfS2b06ngEUUwEl1BJYf4ZZpq/qra9MQOAQWQHYv
mq75Dbs48Sw+8Gdo9q8oP1wW2/11w/drIbBc7C5FdmKij8wX1jVgTk3NgP4VMG2O
ui17dCV8b55PRKymHyXXEZwE7z6sRpnjtcNQBCiNO4Klbdsf36O6iSTXH2YH4uKz
ATMl/Kj6YJGRI4YCnorDzPupaTbootqVq79MIkXsyJoVkpRnehCT2cXO4CFIUH5F
eaS3tDnW+SF6qVqKTT/x6ux15gyLenpCAdgD3uIecu7sqF32rhDfOIadZ9ybHgm1
nSfOnEP2PHOvo7tlDmiv1FZdbZKYc3VGb1R0RhXRmMmSf7BblWjAKJehXp7oz7bT
xFzPP1yhhaL1fHkYxkJ99H5+4SRzjEbCwNt8F6MVsmSlk6ycLNxwbKjAN4UkqJyl
Nsuop7mb5MBjdYc3t7dJKP8jpPdc8KsTeX3EOTdYuk4a7ylKrAJeYFZ2nBzMYx4r
CUyM8G3fTDfihS9VxaUVP+QVdrhxzOHSfhyJs7EAbDUkgnJpuV/lEXg/GD8dWcL7
0ac6QGxq+mhOZHl2NijPn0kc4OPrblwEsIpM+kiqk1VKT/t2zX7pKaOjxaG/tR88
FyBYG6r4gCq8EmPy4A44VScE2KjjplYe3EbbD92DUsKxzrI8hlxu6syR02bjWwvy
NoSEXLuBav4ws48tJ53UmAYzAVbVAtjagVq6F3JE6gROJTpMhuikmMZydjKMUX9/
XydX2WNeehrUiuxY5r3gdOm7WtTs7Or//5kvpuFWiTPPm2QnNZ2N6GR/Mq/NG38R
tQubfBWRbjW0bSNyTmsLmk7Mt7rkFKiW4hM3O8kqFbqiLb89h7Sdg/15HhnbsO7C
ZZa1NvplTgD8lsUjO3/W45LLJO3C3O43kqRcotcLnh4YEGzZKBUXAE4szG5NIvSG
UGLetCbj+S9CncJmBjrMH8sxYuUAv/yyDgs8is2E4cxDie0+LWh518TqUv+GBuCF
udK9GRJL7q6jDwCTJsr4unQHdtVWpC5sqTX8+2XAEMuZ0mwze+5fF0tdl6Cf5NOU
k9/HMaZG4ZVxPSt1GJbKuLtDIJvZy0iKP4bDlN5iWMSy+lVVgX13l7jSe3W7mHK7
tOP+wa76yDTix9rM1/ypRuQIstRsXgXr3aNTCuTmQAxABHU1+yyS1VW3ZVW+GS8r
NO1s0Up9zooDcPb6YPpmJQT0Hj1Q6VJWCIeBwJQ7LmxHUZRJXI73SUPNpmkLWNRf
9cnLCyWFwoEXtsKYzMvautXXOu8sYLUmsKoC1nRknRM9pTG/Ss1EGpyHyIEnNpjQ
1KzRgnYtpCX4/McFo7LzK85yKfpyH5hX6TSNicYkvv9wJ8ITD/2GwSWQu6vqJrSC
4UCMuRtyhj+6DYaQuSEnT7OWV1e3GxqoO2IUe2dE7gsKygBFwySm76UTAEYZ0FdS
kuwTOjlMsHHd2Kf+kl7m4FKjjPmrHxnrBL0ZxG/kRwVMzzeJJHAQNTkG2uILuJZA
mFiZvy2Po2NljkFINQXYocfRhasBSZNynQ/JDcgNQ4paDZ62sEXmvk15lbZwyDYx
/GFKnU56samHMjfsL2XsQ2S0b5Qabqq+1mDChUgWmyZFHHJQhNP3c8K0XXTh8CC0
jA865MOkzz02X8WmNOspr0V/FLP+JX5xGoBWIiywPl4hz3eiNKO4UsABOdGgJj8E
jSrfW2DEa3bvx/ex8iaTBaMv4q+mhYR2SFDf60OyI+0F58fjkNY4jAHJ9PxsF0R/
DH+9n+SRvs4xL7gakbP7yAyrdHwPaWVM+ynEZdd9qfkWKxDUgHzwxk+V7HJ9lEuH
51pWwW9XRJvaMhrOX+KD/f605pVKtZsQS6qjRuL/bMxz9wcoQSKXIUc9Q5rYVtRi
31y5vM/8Ue7Z7hNdZ5K/dk79DKNxhq1GHgmCGCTIIuJ4Wk9v2bBXqsMTkIGWTbkv
hg2uiegXFHRBvcwoeOJnb22JIMM+DgmZLK2HQGttquTGh6rR6FYNn2AzPXPujDs/
KR/PTSraoJ4EviucBV5SOFlNGp2JUm0z2Yzz2vOIpRY7oQPDegFrA6ep6t2gdSGh
sLSgjPOtlDfftOeFtzv4ELneeB91V8ub0h0TtR0etZUHROlN4CtwpXRcMHsRXTN8
9BgMYRSyIzvE02M6w6/ZBCs8ew9uS3ReMbQS5vIXsQDqycR51O507EYQFWEbncoj
NVmy8zoqZNp1F/Esh7Tnu0TVnCrS7ZcDMw0Z3AOuQ2vn3u3zipIlaBN/ozFI0dpg
/ZFxXcX2lusj3dCYS6SKIL+6IruDMkf6UUhDSJoZhnsbvos2QImX2zTsNtojiwjC
tV6OeTn8AUiXIxnMlNvkhwe/hiMfF/J4hk4qKMDUemQowGrkPL+hdzOfp7fxs4s1
8HxGnLFXH5VS0CIVrySWNiyPhMJIYUhsiaRyzp8J1+dIokb0HC+tYPxOkXZXrI3h
ySJIZhN8rj18u3LN4H6nsDY36fV8s1XEfYwTlnvW/m9hgVEQ6VZgIRx5irWrnr/q
7FLUiTUtQf+W47LApspKm6/9eGjwNeEZLmHb56UrDyr+ECNI/jqi3F1zOQTmj52z
/T+zTTt8SByPCSB9NCbCeSIM+mmSFvLe6/r0UI2acU8MXEgiY2KHNUpSQL2ygyMS
LhLPM9XDXUUPj3ODwISwJGNBt0RKZfNJHtwi4Y/2R+NsnVvPfJJOUVSVAF6VE83P
Qdn+AniInZmc8wcZjQQ//VnzCRio3aonIbUQyJMv9RqYtmnHuqA4UhqZ+lr/5wrh
FNzBOmDpOIt2ozsVu4oRkXMSWLLQa61g81I1YGlH+Aar5shMjOFX1f+2gazKvEmB
At+omqpoayqjhomhWRAAxD7541wWyQq3kzQL3ZlrQFo7yyzy+JoZ4f9+KoZm+DjX
eEJKYJP4EJwZ1n0YmlH40geqgQ/0VybXKKgIjLjMS77fsl0ZHXrgFLbRAqLgB6u2
RtzvEqdxam04J+jfJgw80GBAAng7FMvR4rhGMmVF9Oi4mCwo9jbEHrz27xrjj1+d
IbLjOcXd/08bYcRNcLENzUGaWreZWdm+6z3ZEdOzdYNh83wOdwwsCE077Gsx4WNX
JDTGU9FracErI0Sxmh04RTiy9JrAvgxF/AtuD7aCEN1CvaI7hxCrOxpl6pB5y9bP
zywo7tMo2ivD8YDr62yUniiAphNIkzAfxbbi8OEVALfRdwCfYNMXaSCoVXlIOoRb
QeFECG/idziTR+XgsgqMZg==
`protect END_PROTECTED
