`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o90lMNneELrazslQMjC1jmm1FNoUa3ux8wUOc7NbF1pq8iRHqYZiZdrv0f9n8K5Z
YNfoeBovC/iMIfJ0EwDdMIIjhFphr1IDHcZ7Az9arR934DqGxKjPicgwdmhzgwAe
b8jTbY3Ew5uiLSNE51LyZuBTvMd0KSeGkwwGhLu6MwDmI6jq1CDZutaLgkjTxAUw
w23/rUtJW8Hhu/iHSl8+6oJ/jFWyCTTFcR1oD5dXIV5hZ1iUi2LwmuyS4+ruApTw
oU1MjI4yJ3JwFf5IcVh7jUL7ryi0rdHx9FzIwL9J9BA=
`protect END_PROTECTED
