`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E1W5ap82KdzUOZWy0nO7ISfK0FmBaWN7PYJS3b7fZmFXIR7cR8MWjt0yXRRMRzXW
9z+ooayVHo1H3G4WcrxpDf2BaWBPi5l14rd/MRuBh//Zjdj+cc1jjdlxrU82z2ld
0JqSO/5lGoSjXIGpUfzsygVw23bod7z8reKNm5Vz0JWaqzIC7izlA3SyfZ0bRJWT
wIL3zQwKqu27eE9qpTRd+DpMGQPo49ts2pMU2HDnZlbt89AdGGI5gV91HqjWboY9
Haz079Yi0c7ydtuu4kPbp9ANVztsR+huzUAiGccM5oOlM0TDRHqI+bKBIAMicOIf
TmZv2XfMBo6SR7t50yjZCU5iMOAtLWWzwD+NflSTYE6h/UkXwmnFfQ/YPwUk8iHe
9dYczUPYxmindkqmquwIrViuqEk1qS8fAZ3jaDb7imSWGekulpNTPJS68U0daahL
H920RQitWZWMx6iCl2Ol3ttkoXy+iZXHrenZdPrGBAzQowyrOLjt8hlrI+ntWhBx
G5qWphNnWitnZes4UnWa6YchkvHOe/j+B4RoTDZm1i32gH0z9uVJh21qLPe0KqOR
ZfHmmrQPuo5e9cT+xaSBDM7iE4Ow+5zZd2mUxh1PeaLz6avcKG29OsdM0JE6NUq3
rgdPkamLeS5PG0urxQsn74u2056OXvtazj5CocAoiGiD4U3+WKm6SV+kRKq+677F
aPlCe5YkT5oqPLT+lsuUsGXZJc/ViRLFbFdkPce5Ga72lVaVrt0rfpOMuB5+k1qy
OwNAQPQ+bWGKe9fiyAXTmRtw9CAKTiKi2nZMup5+OiZ6a5fDmJa7BdIXsn5XOE+L
HdX3+1/Da7M3m7Oe/dJb6KQi4TBUf1hPBsBReL4bwosjN7vmHVUn9N1inVMmI/0o
i4qEd2RlZrw4rOUVXuDGDmAw7m4Dojm5QkM6hi0USJ4Zbd5d6/sQwd3ztuvavoA+
lor34D9hOU93YQ1nUZ9/ZWaqLmMVYzOugpRapZ8CbMwGgWQHyDpeXxS/DcrUwn16
H0bILfc/9E2T2BpSON5kvRqrL5LDEgRSsnV3A62qETrFrpwhrfZVRwZ24Sl82WU7
nnkFkOiu3AGjPw3+j2/epcaNng+79NJHNT15G5H7h5YFG9isVrY04O0NyQ0FB17/
j6IMCmySZHkZYN3mHaZUa7tqX0dE7Sm3INeNQafEtgxxQAhmhr8U4qSP533RKZSS
XCRQ0ksgPKhHoASdl6NK6RUabdEQGqx8kfRabmzLa3/jOLJJFS49GiiIDsDrMszk
hwyHmo62vS7Bk74k/npZhagRshF+wXKhlB0gI/UiLTif1e77pWAb5DGE7B2+xsk3
ocBQubUzuHos7HqBTceZs5aXjlAXwWAazV99bS0y681A2qfwqGiBe47R+WrRjdIq
vjybRQ38tYnA0o8ALJGhyYGhKe5T/fZ/PeDgJqU/5ZJrPosUu+8IcOs687TJWKPv
4ubDbHdp2IEkKyx3aQ6jLUWeNDMLu1EY7DLS+m9H7nyWs5QvaEh/4ZXipHnAQi+F
wXmNvfaUsFjC4y5m+xEcMI7RX2CiXK9DMYPkdxxqW7fW8qmYDu7Gxvvhs3wMBT3Y
RtGa+kBzWHaOumv1DYrJ3FIBWiPiTkA2Pd8ZLRig6W3Zsxe9oamG6Sd9x/NG9lVD
Hms3n0AnINw5AlPwNN4BT6AplFpOtfa1oqFxHyl6YSYtirAyn5yegL0lgY0wn/Os
i1elHJ9gBjA5qZQ0CnsMlC6QtaX+aqdlu3ttVQbhV4hcSJKuOGnUZqkG27m/A7Wb
P2aUbAI/MbnTzXeQ50VYzUh5mQGXLBS19ylf7R5SYIAB6Xo0tZQn6NwtqmKSOWIF
3Sfc5ML4gchtvXNam4BuVtnrxRaHRUrsoapd1ABFddx/JBnTRaYxcmVUYu25tT5a
J+KTpE5iU9xSlJIUA5Mq5OiAl96VwfZBOb5aKCzbLd2l1+pKTsza1sBVJUIyG379
LxDbuCS7ctL52l222KCWEWWhPTMqJ+BZZBBT92UOFMNqy+gnb/QyiHfnbllMszNj
ipwd9J8sP7/ovKa/acI9hvrktQTtkouert6TN33YFLxuGmv/wGz1qmZoExQ8F71m
bfj0o8gaGoA9bWPO1YjzuB+np1EtYRcNtJDgqjT+xifaEWVMq+M21aeoDj9svHad
o7/16KXrJp43wgikOP+GvbtdBiLmGm+0Yj21PH2MtZJowSFn/m9/t/fLPrlQdu+r
ILv5s6VxzVH924dgQUN052gF1FVuemRAXfkRUTB34tGNuHjHXNOT9osznkSbTXeT
8v6ux+RgPav7L+mrKU52MkxPd7PFEcVWvsjVsP8tujOx4xWGA7emFYy66M1dcbzt
IgWS2bIY+sHsI2RIdGfmZLEDC7VOXP6o/ZtKwo/4eR6FbdQVo8X1KYpJQlT7sca2
VX1/1sTEgTOkiyJ1kfc66RxPe/V9Zhp1qU/enTLGxd9eS1XwZPTorYmIQPpD/GeT
Ni7nxxRKtFpLyIQH6JLWGNMtIBcY7GPhIaspnTpqwOY1JjMWEhdVPOkOZXr5beVl
/2HebYBSFDEX8MmPWNy7v4CzOoiRxtOO7WVixRnpe7Lli2cMnqqdJVTtmeDabmZr
Uj1Oetc2DZvFfDwrhTPdmI97kICF6HO38/HuF0uJngf1B3as39qz0ejXif3uPYD8
/YSu9Vdw9DpNHCAdiDY7gzCDbdzHgKamv3njWakFWVQAn1s+cfJTnSbunOk4xuYI
3QWio2e3tzSyqu/Z5VJKEXwwf3jMx21VuyTT8KtnwbDYdBDByl9RWjWxI3doe7QC
DPs3Kkp+/605TMKivvJ9n3Ly1UMMIJy8yfU2/+g46gtz4btJe8Tq+dsr8Pkoq6qF
dBdGZ/oU2DD6WiGSR4cL4zeP9R8O6yJM9vYOfU7bRHweWDvXVVJUSHrDVCsKaoLb
Ubc1MLgNdNuwxH2Kcsu2fW70qc3hXotiqps4/TQ6hqzMqjv63s4/OuTo8PoUJbXp
mvofkue847qPr3TEmfq0eYgyiMqrFoRFuCd24plihjo4D30G+51A6cCo+kG0TXSO
fanyjYkbcbe0RBk61sGRyS56sQbg0sBEsxb1B9G9791Dols1xFo4Fjh4150XsbVE
SCGoLqpuveGhAbQfiwQLcXjXvK3c3XenQpUJEvqcD0t3j6LxSYXXFrvpOqofhg0F
BwbWUgICmIwD1aQacRJNBVuDPpzrvfOM/qWfsmXyYJuVabiWSvjjD+I6eOMfbmp+
PeZ/3FhdzZLPxcwNmkJk7eDnWUGoJ3NRDmYJVOdtbCUmGmUoKvS5XrDoDdzbYgJW
5Jc+NF6ztIEixDfXLZoi2ytBniOwQbzfodx2ONfqSUrguo+yFdtXbzpNTzyMK0pv
MdEU0DICiQEZNUpirCOBKp6hbn7k33vVs3XR1dZBU2a/u5AQP0YNHbnSOhvrTv1M
zv3RpE5JysRGEOiGfsCeS1SJvpbeltiBhxRMS2Kq00RnOxTTFMnj7kj21sL4Qvvq
6TpO0RmRWlvX0bKZ8poPKQ/oB1H2SVovDHPEGdgZLCNNzPZ8BOBhSra9IRIErv8M
/uKGhP0bDNrg5AkKCZY98E+n+4pI0+0LeoFyKHU3z+jI0ZYIgfQEHWKKVnHLuGCj
rDWO4jR+ZoS8kqGibpMS9g==
`protect END_PROTECTED
