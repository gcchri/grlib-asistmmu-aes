`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T+BKHJ81hDvMyvRGvDayq0bwEhdrAn0UNVLedwqmfkTWQMJX+nmwvoaIJHlcHOLi
QK2cUg7sZtIBxTghlK6/V1l9esq39vU5/QihP7xrF3YNpOQO0PZy4VBmpbqNakYP
Kkf4pqaslPBeNB7/a86Kfrdrcivo02a1gKa9UONc1Re0w+sNHhdISqkbLQo8ivOZ
AEaJ0YnRo6dU3U4IHubp9WbvQCk72W9H8HD824qWLy6mzDzJ8ZnAzlMKYj1ePUFq
7dnxOGaSYbvwsqMg260tPQ961GHoRVsN4D4j/0SVIKuIWz010RMpDNUkTWGGgkz1
5h5o7QCde7vbtEwY2C2whOqZtg+ZYalLWnjL1+qU5Lr/+yZkrXGS31eWfJdUIXhx
PSNjMudeuw7c4ebPRWmsbD5Flf0EnGDXTyX3ozCnaKJljmRvFqS0Rhb4WbE3O5dj
B49C9MCKKvvk05X5N8DopdZuuPUxE62E2x47cOuNxLMPqjKPA9qfu6dmyXYoQ6vf
`protect END_PROTECTED
