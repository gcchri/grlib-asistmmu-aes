`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TcS5MM/bd+RPMWUXkKlvEMo8DPjZYtD+nrwoFXC4rkeOorx6GqOhBsaBFcMUqFkM
fYtT+IBHzzaYYImyS18ycb2+D+Hs/JacRpiqv8UpvXf/1PlmpZQFxQwK9Z4AzLQ5
kk/2kYz0xJhT1PZO4w7YjeulsHWcUgRDqhgA4+6ygunpt9aMLM6QNm+t6zwoTQjM
az8zsTIZhzWXfqyF5Z2Gxv6+E7r3dpCS9uzVggy3ixVfGiyYfTzqv3m6n0yS8aBf
WpBPNJfIENmMBV80JhTnsq5l4NoIp+Xbqj/gkEzDKusU9BeIcF2hiouODNYS2XhP
B9NBPje4972wav12ZeIjAzrEjjoVE4M384CIawY/2siXESB7V5znHbtUZK0CLznf
`protect END_PROTECTED
