`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
riWjdzgFMYDszXzlSGCR0LetU/FphOiMNDKJfR+poDrZEG0/8b4rr0YEUiXH7ZJf
KeSSyrYFtOv3mScuMJkYGsuwjyhHpng/3BNB2SzCf/7Dk2wHzNHYUjGK+gJpix9T
x8RSMN5sq5W4XcSTmdXrTrUnKM9DthgJlQcsIMvLbKo46AHWoVbhci22+7hUpIuX
KMIiIHY641ykQsToLtmfdzbTlfrrZtsxJUkLyFmNwCMfnyTHik9OPw3YVcOo3Un6
q9isvYebK2KF2vC8P0Bi1310i2Wku6Jm7dJyMRhplggXA4NDx/FC/2c00vKwwTp/
zp6UK51WsuDzRfT0Y7g8hgIF+VaaL1+Ty774Wx2VKAL1Xkv6Bepq8x4lD/5wyuwg
MZUgaAj1Q1QJVvTveNqUinp8gNpI0/E2je83HsZXlFMHM3KWR3z5jxlhPGoQVbco
DCGzhmz4tre0+JiSZS9xB6OFYM/wwh/XMPhp5H2VRfw=
`protect END_PROTECTED
