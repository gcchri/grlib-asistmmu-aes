`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0j8MQWsavMfURxeTcbQGmty+5mhuG/bPDujN0LglvHWku0Wc8PcAW8H0oxH41QSw
N2Il6nd/p2iFVtnS0CqIie7KvyA8QwEt5XtS1CtmKd1yrxOzf6ppJ0JFj+978yrZ
AkiA3E6H+1Z4UFfik/tOyQTM0Nrg7ou4arTDFgwfNhFLmDJ1ZKrmUtZgLjyEkZOA
qWk6AvROqCnIVhiYIZ/3SsAh0q96keRho6BHGS5ZV7bDL1rhkuuYfLS+EA+EoqUF
jc4W4fWYxBKm8TCa8w/M8Z6XPvtDi1nCRGnPdowdRfPeaLZRb7pTNKvzcKuOryXR
CHPgz0WOfI8mgjJ3g3DlqDf+F5ulouj+jKCGs01fJ5ntN7zSX+VfER/d34m3M5ua
LHgojlUvPQNPVUEiJ5SlqELLmKTWkKP1g6atjbQgVdZgvDCGQ2jF9y3MpVTIFpZ8
uqp2Q3KcHoniyIYQjtQLOWbI4DgVOYZlMt/7s+p2uRSVk4VMSLoUszQvxbRJkedX
bq8qE5THyWQD9HySLg+fOxm6N+HieyI4no9GEyxGccwb0QriPwkOnDXn2RV1FbrA
PelSEye5p68LftbV64sxtJAECENxPQ7g7QKFq3JFO6s=
`protect END_PROTECTED
