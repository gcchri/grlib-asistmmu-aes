`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QHd6gWnL3g3RrIrik7chlGSntd4AUlQmzoqGMuyGtFyiDba0+i01vr8XSaAQg+cP
f0zLwol2V016yXKo8hjxpvz1YHvHgBBRqj5/Mp2Wbb6NLqNVQnzQzOm3DkRg586E
vyNzPFAMIeRJ0LWyA/9RYtVXtQgmPSq/k74ueYHKXRD2cViTOdDexCWDz9wkt6S0
KYe8ZY2SywbwV9djCg9Wt7mJoBAeszXEywgcEQDAMSzvjPFbUN8QuGpb2xmazDOB
7IyPiBWjG59wC+4T5oCB1g2bHoGtW3DUYKatfL37sVh2ZO/RIS3oGbCDui7BBSe2
MSH0Yef8VYa8dhFp0BKtkCp/OQXKudhQThtJ6Ir7ypHSIUNcDTIvHzqvYkalrlzQ
rBy1gUR783cw5Fps2UVU/g==
`protect END_PROTECTED
