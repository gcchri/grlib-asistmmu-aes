`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DJTuVjwXhDpNglh4kT0JJH292c8wQG+mUlZNYsdh3t5WD5kJYT/mkJ2fIJydJlwO
RRUBN2ik8mcwblhZ4w0AfVgVTtQC0ER4t8Xf8X6DTVpZm7IiMrjuglLNqQZQ4RN0
DkWTc0kshJGkP9c1FC7yymKtyt946R2lFtyRaJ2HIF21F25dht4cAvUW+YEEfG0X
HeuHLSSKVXYK+AiHBTEfFTUosc44hdUN3lSmQ92zPM0vM+sJagogaFqkJgctjp3C
+crn1I8vUa95i6gnFZreV9cPJfJFPs0DwKu/+tDLSTMyD1/0KAfubZW4tZ1x9OOx
WfQLjrazrlMsIt36tvopjV6Z5rhX/Sb+tqFEFjXalLolWzJkola5w7u1hfwOcRR9
/hwwMSUUz18kOM99iNHiWo+xblBZGMFveF1veH8BdO2yLjOUiE5wgD+VBVVtQl4u
LO87AejJzmn7md2hPWRTIV8adyZEPrOvg5IhfBfnZQQqTSKKldWyJAhWUO3a5+n1
T5jatfWzalXeao6JCO7f6xtKtOTOitHD0qDNI3kFtuz9U161aCq7ijv6SRDJBceA
YT7rpd5si4rDAoqYy+588hXS6dd4iQZupVLAlhFyV6x4ECK0b110P3A53UQbpwFc
D3BLecYiS7tHS9ob5am7MH0zytEYTR0tle3L0I1aoJNXx73mk0mvFpVGzUbKTZRm
65pB9D3A3ZEu/IJGPABgakYFlq+P8Kd0NiqXmZkb8+awhQXWR6pxHNTTsNvpTezf
LYObKatP2kDZhyloQAHO5w==
`protect END_PROTECTED
