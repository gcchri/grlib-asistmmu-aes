`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PTvWqD2DfC15iW1S9Cvur0/Y9qsGJ/lrIVmyGId/rI1JI7+LMucsfL41htreQrix
cyI1VHqDqpTYLL11RbHjuZEJXgvv2D6CZAWKpU/SD9a/fRR0eDrno01w54V6a1t+
xR2dc2CYe5VOruFNOyVzYUtmyLrlO2UJJE4aVv/xRaBYyrHDgu4nvIWS0vK/lJu2
5rA6vz3QxND23/oXE9XLhM/oSKjss8d8xVeKItaWn8w6AfjHU5wrTf+g9wBDkTzH
jfAuk+H6kNdc6U96/DXFILY7oY4d28sgJWWK9eiS2fWENu+4Z0VHlVIzPMrNuEoQ
QiDRLjc07vYrSejbb8GONFpEkuXIthP96fTcDOGmZT0IHx6kBUtVSDzxNqtS2O/7
skNb4IgQZ9IbvpHdp4PUUlu3YG2TOGhpaWu6+nmT/SLp8mpszRu92OmdBWWAzzDR
j5PBN9QPeAUeJ1UhYt4BswiOGhK6cOD9GLYQ4Sp7F0G1cshqDEMJfphpcqSwUaN+
KAmZsmOAQUjkWGbbl7lBtFtZrIxQnWK+3Xugodr/rjEppQIwOfmJWhxu3t1rJMd1
ShA5nRHIDsPxydkkmjO6ZgjCffw6XMhRtC2c+uVWzI5F7zxGHwMh9caq0lhkHXPh
S9TLwTprMBkLBRy6bsf8jXHoEUJt7oekjrB2Oq3UVIEi1Y1MZtJgfc+7nxFTawnK
byQLX93lsCadUA/cpr69hFnH81xlkZVus86/3qtLJwS4MloKTgZkJM3opG5HaZ0O
Ni3dKBpay+zUXy02vUcqxO/xQx1JN8cKAuQ0N6Dq2FW2/am6MDrZzQN7q76iAmbW
O4dgRJdoUYK2AkOPmmRM+A==
`protect END_PROTECTED
