`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
isGokU8vw+BjCiSHZZ5gdHYi/CEOhlnlzTSZmz8yS/M3k5yIrFUeY0a3MNmerMBq
plliL6i0bL6bklZeszDF4I1ZadXrW9sd2i91THNRLM6NT723TlscxmjrmsVbkcg8
sLHRxw/D6QZAzNsv9G+jmZoSbNLRtmzN8Sqr6DSl5VUEO2ilZ4d1IC4ZZ8DO0mu4
O7eroKjwgsmu3BAwkFhReGfx6vyzY6Aur4Foh42AytTWE9JeSvK2AVOEl4/JgKAh
w3bc8Fw1KC6f97oXl6wwT+DLDa26URRlipVCq4Sf+2Rojlrzz4CaRNoZytUBunF7
1K7arN7ESJt/v8IkbJnW1Ow0fI0LHEbzk8bLZDKUukDodqMDnV9tZxjmFYxWkkHj
z9FOJRaCnokuan62vY0bwlxxFmvRBxgJBrH24UdlmNU=
`protect END_PROTECTED
