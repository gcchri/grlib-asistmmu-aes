`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C6bj7kpgIoX7OFxo5tL13saGBSA4/3PzpTpTlKnTwQTVg9wo0FbCQ9/nrzIeo8OO
Y37DTIuOA1sXuRVRh9ZUroE9vfCp1KBjzBknyB3mM5JdtY1vIKwEmaOAVgUhdRbR
eR8LZyhSkmDfHacGcsk4RkAWnWdVjIRGw8IDXcW/waULasV/ZLFGFw22k50zXqlK
2kPxROk0DOqqf9q4/aq9nsyCil/k+n0waXZ3NoEqeyeaa8kmqznMq8Wci4lII8JL
dsylXPqaB7ANT7dpSpv8pMNEE5J1VUaiCbEZf1710hDLH513642ix7hIpHXUJguf
i/iHqiuMyfCXDdHIglTfqjuBGWplrxJrXMhPKEYVzF/E8cJgD4zXb/JONK1vhqB8
CPXYk6CkduQ9aUyR9imKZLWlOPdzeOWxmWev9EzX0vqpx9UoxSuoFrWq9hx7i8PA
`protect END_PROTECTED
