`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x9GG2lc9lElstUbjbC4QCs9ae5hTwPi6mA4EC3zdo7fcg4C/3zV24+axy8JReSQS
HTZrVrOYlofK2bAd5Te0DHcgf7+bzXK+UNrtNJ+qV6fp2Wn9Sl2ABS7Dh7RbO1eZ
Hl0oxf9l1weu2eFhwcYqWzD5HYgivqYr1xj6tzm0Pme1RBjutUZP5Rbj4RYUcgzI
ICe4fiNjtHyrj4aMYne5V65DBmNuhLdDPREHj58ly6GoQg+vVEPvdW1JCjy+zl23
Lis87SptEAMJbBPc4zYmzhmvACVEyhrYgwIDAnvi4cHYMd79FullPfjbo4VCNf5i
cA+MD1ISy38Ahbnc19JN0dxbgKip5yUuO4eHyS/q17D/+9t5zeHoKkNm3HcKPN33
n8oumg35tSXUgYkDrdi9rIwV86QKiMo7T5x+bgzufSSc7ySegOVCHrYYeqt9aKpB
WdJTaSSGTh52G1UDfUdFdttV3q5kILRZ4AemBuFp8sflPeIJtJT7lNy97a5a1R8j
sv9+CrSpHPveu32bH8ciekdDDcfNag5TdZl5JtXBs0mzZk71HS8DRJdMqxMM2hp1
+NG0KDLsQBPc6WI+FFuZVnSOgbr8G7hBib24+d/8pAIg3VeyB1gLzEQ6mpOqI3dD
jZ8W6l5c3FGflgzQtrq2lefPyL0Xvt/9NVBQAy7h1ean2OG+DyHxsQai3oH5ueGi
`protect END_PROTECTED
