`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/CQwHX+SF4WR//isObTKXSSRAk7a41z5e80uAtAQj3CPxU2dlZCy5p9IRNgCwPJD
m/NPZpxS//gMQRKWVgFOuISew9xUg/Tsgut5iLdiFNdGoF59YlK2OCPn4s9xLmmL
IkXEFWRzB8hscL90C4e0FQTAMa4biLAKq4Myw2A4alCxf4HtE0nMqDWDkVX6SzL2
KJGrI8JKWlTeFEmHkHZg/UocBCMbQy1Jz1fdo2af+GoWCCPzHCNe3ozEXU+4qXa/
ngbWt04yDv5R0W17iOTJ0Q==
`protect END_PROTECTED
