`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jZ/bGQK35D/2V40s1MhhYLh0aGMAxgEDkZ+CIzbAwE5FldAqhojots8zXEjaMhHZ
A6Vn1sl9BlUqQe2JgUxY6jL6KePIW9yzMm9EsNQfsNqmNyjfUrt5ntzp0HkH4OpX
Sifgbrgwi8MuHn9X0ppaQZdNDIMdt+ex3YrtVK9MB0YgiUK3IDHzVJizXWu6Vrwm
wciMUmkcerLa+4p2zcJM1HxsdD4qdYI0CU6oiDc7btsg51oaWQO9OWcp1lI7z2Db
h7VMajSBBsMPvrFhNSYqb6Es+Z3zMY4svg0w6QV8kVm+QEb+otuJ/Yn1KqofbCy+
FGAqJyPOypjenyMVCuoLZ6Pde4lOcclGCOWBoQb0d0rsoyp8p2owNEtEZDsGqB8s
nPUFGCCVuKlMG2Z8466uDyXPj31WHHrSwfPHhXhNPEzA6423UZOkr8POzry9CY6b
/0Ph9vMVZPZ2jI1VXbJ27fkr+MIokk09AuayDf+SD5h32agV5AMvfQ7eIx2YsWMg
w8aYGOcavXmQ4h/fxbbcrOc1UAk0s/FYfwNxgW3gpwOYLpLw4EX0cpsoleV4Y0d5
rgVnBSJRT4pujA1HlYazg+PquMyAAXPj+kGtEcF+fYWJY2yKvPF0dmx8hozybFtY
oiaPIohypqOwUFCunOpzdm3m99So3/GzbaBgt7VijerfFN7ZRjfrxGfctXdaTCWo
mRfugQya81SCaIn60pXr8YiKekC0RUL41feTq1s67aFTSTCZvA91H+W7/nZZbZb4
EzE41zEObtpoN/5M/hjpIsH8by/IO4LgCiCQL/mCZLNvTo2C2MQMmVORssh/yBar
beRHMA1LNkw6U5wcFkyOf6kFztm9CJ2japJgNVFBh7pnXjsrAC7bOMtk8X54L6fd
erTtUFKNeYAb+SNYZqigpLd+qjnYmw6AmuaP6OZgH5GuglpQ1pH/2qFxU29YcGVJ
HsvWOOLvld2y8s/uvzGlheseNjhYh59cJ37R7l4TpmzXzYkkpWp5n+RNieEieCeZ
Sertg84Yrlu4VvpYGnWfvETS4jIf+aWkMmH7KF4hF6AQATaNKLThSrBoKxBLh+56
z1LcBZ23Zocz5QQiu2gbPTAGCuW9qewgI2MxfkoVJISXvS446UYgjSn7pWOWiST2
kNEUQj64T3vPpGqjalEnZXehXkmTEpSCPpLMe6mWcMC6VIwhG8EUH/khH0qct8IN
iG7nAALgvhlsLYnbNygRdYA2qPrqss9HasjUWlHZf+MZO4c3DmUGtSOhkbuqfrxN
/JxsfXKPWmWoxyImB01/HnLCDRA0WnW4BHVQiRULBUGdmmA1u9nbh4GxWQZv00D/
mt6/CBptPOKkgVBpjSfW7FbM97KTm/jvlp1ILRredjozC4PnnYD+pBSKIlgesE8S
DcQT1PDqHLaSX8Rk27Qi6jynKkEANPQq4ZnRkQCp2pP42siHO3GBmgbfqzYRqeOt
+KIcvozm3IOq+Kle+n1IgpFOLw/+Gr6gg18e3vYNcKFK1WIs15XiSZn4Pcy00Rz1
MOhbqhnvk83S5X+7U3L8j2OytexvMsyXIe5kmdMKPwws7jOYAQezhL5ac6uI+Pu7
ZEaZhs31EL/+VNennXCkV+GnBshOFjCQjKm1/OOFqPT17wEbvDCfs/Am7xBuqF+r
ZW+Jt8XX+cccJcS9/Lt6SWEMJongx4YkX068bIm4rooV3trGahyj0oMCmUvErn+H
3kR19RzLrOwknoRF69jLCaOdWs0N0yiM0YjFrmgkNd/wO8TX/YWbDIDxEpIeZqk/
XWB/lbNZaN/7MJSEeuuvWXvVNab5qIrg0MKju3E7vIVOhwp7UElkkEYjX8xaaXxB
nR019510zsbKdqHF5OYrREo9UWUMx8XNTAoIi/TTlhMaIDNJLAiJy8BazSNTlIwa
gy54CP0tz2Iyx0QHAej08m7dSdL1kJaLXRzhMbydUjz+8zU+MKNp2VeHD6B3nPB0
VTCqSjQlYZZLdsU7MhuYM0cmxrjwhmzlSOAIn7r7w+4iMx+C616GE58DKmfRdUUf
0tImxhy4JRfoNcOG8erbtiCTtpZ/I8tpAZrr4/FogIsKfnt4Ae2AQCXsxYBlGN9K
i6ofeIgj0QA7/Ghh2Nzo3nBq0AyaJ9Eo/cZ9/9wBHUtd8Yob80WEZzq1ZCudV1v0
mri2Wm+XKbv0mLJnk9Pt96lF3eTGD9P6OnjuJX7HJ1ZOO39oPi2qS+O4X4/1JlIe
T8cnvxVZnCsqQ+QIQTgMSNUTrY4BI8xep1WPmDmRKOm3nVXmqfuk48WYA7+oxLE1
7DYonYGCpAGTN7IdpWj1z8dx0Pm2KCc2z06f6b6qQ6yQ4nEKj0GqnkLgguUQ4ph/
dK7OsO+cpYVLvPDO0az8b3rFzAvWK991wmJrDDeBglf3T3umkHgOqsHikaaZzB8O
NlcfvTexcq+PZwV2XXj/MB9yFBNbqjgZ0V31L5KUZXC7g9xhkPxE/TySGSZpawMg
VHBs5EXE1rne8WiD9YZdww97UKDKRlR6czg1kmXHG6z8NGgwIPk2grzEvVhpjQ7t
+kdU1CaM2s9scyDuJHkH7kIR429B5ffkY9y6JAnoQPWnmEbdDu5wMVd4BdT1+RZa
BWkrpAlNWX0w0SvVlS3HD0W0ARXfbRpEab8ZF5p2Y/zx3LjR3tYvyRCb/um5DcCd
Y8fOzyin+mezG8mo/SVhuNoZtFLtYETSP/Bm66PatT2c3xF7x8RvCmhr/ICZO+Mj
alXUKxYPvPrgclVs/sXUBYn4xkTe3qnhuJreUz4wHIbAFWpL+RmL2xqYElslFmwk
eMHcXuuFqLk6hLlx/ewh1rKQJL2LsvwbQbveEqKjcufktqN5MZ4nz5wWn+f8ExrK
hFn/eR6Ky2bZosdTMMcz2GaCQoNDwBRONKKpQ3pHLX7PcfnN8kcQ6r4iziZPmzoG
uoxSXgmHRtU+AChKsEWpoClIDcluSHCNq7AVsZVI1bGP3ODbEQa/mj1OE/vkIIaR
M48ilud0Vf4PAslWZTkRIQHocCaiqOdHLuwBTJs+5Oo8OqhUcFAhLKb9QY84xRLI
WquQszoGM38x2Jq9soVyNIH0MSJG1ZtNmjW7WMnPAWgu7kx5G/vGZlEodjnZVJVC
r43Po2Gjlcdr//8ih71BWIAWg7mxlX14plfb1KwIqUMxdmRhR3ZEHA3ojzqjKvmp
cPocxhZ1j5JTgcR9wDCfO4tMhP/k1+ey2NNORtJybQCH7pNMQboXRPtVthcCWLPX
ZYoab/PHm+rhKy/NdQ6JsbCcopasNbaGtpTxg1U7b0fNOKeDRF4yybrYrqTA2tAZ
3JdAhrFx6DKgg8OAkO2zvPtVxtxssv7B5u0nPmTNcWKF/BaMGm0YCQyjJU2Dc6n7
VMRDNwLgvEpxbrbo7JJNwoy0zAHP2i+52476/+ok9uTCSlaRcw0k18NCewD2pDBr
R/CsWJffZIlGkAHQrK/ysqSbe5HSdg80BNWKRMZ2/d7RC2QpQyEmz2qqtaKtCD1m
d/IuFvtD0ddtRS/YploclZXSBFXMMBd11fW9u2i8gwldnasN5b77FJBgH8mzNaan
gF3HRQr0Fyd8Ls16mql/57SeKK9pvOhTQsyMaKB3ZrhmhMLBQl0f+wMMXr4AV9+d
RQr6jwD+yCxMcDRjElsU45qH0YiLCcjZ4mUHaqdLmpLSAZsEAAIXewksXp7Y+Inj
f9ciMURIT5d2depJnnckXDr9DN3GTRLD1EPIMdSWFsA5HwD7xJduPGXzRIMJIuJF
Z5ld35FsGNPhd09/SfALJBbB8FvZFCSPFNA0bOXP+XitOOgJATGctSanzSON7wWR
0CBEKir7cYu9aHvx0LQZ8MYx8ghqc8WQciahj13QYgfJNo/klTyktAMiM5SdVAo4
EBnLu4Toz1RD1K6KwILJF4tGKUPufy7GT0MhIRUK21ngTCp3KvtSq+iS9jzE2qFl
2H0CtdwrQaJqjJ696yOu80+Q0x/LeFLWjHK6mR8421eReNBJQfS7DkI0QufehvxS
8QTzc+Jd0sSceP5Swti4akEr51OpoW9LY7Qe3uuywPUItQK7iogOFu9uZZ0VWqTB
5TwAfYmkVD6vmBLsj52aq4fwXnyG/7NCNlAshP7c+dKFNG+31uFb5Uk2xvRG/bAs
vbcmIM2abP6ihldY/gu4prG2/UFRDIEe/yG+u1KTjSPLs1n+mWacdCD88lRDR9Vl
CAPGeUzCMgZl7oT+TfhSqhaq6xy9ZYTutV96ZhweKHdeDijjPtKQbUZwqzg2xwW8
Cn2gBhM5Pd0VhiXdlplUcu8T7IzxB2c7XVklUrfU/ekAP8pxpGw+1I1ZKEgVbZfO
vHEErrbllgbpgZ69xXSPON85WiWInKq0YvAjqgyMo37/srMpH0ohiyDDeTef+CJ0
ejFuJRiks5RTdrCLKo7cP6S6zVyMDQr0JpkRwEq7H2SWdeN/lJWRgaFaQ/IoALM9
HxsDb4EWanYlevvpWYkoWGO8oENCV2fn1EH/bbK/Yro4Yo6uOGeXcagi5UGHkjA/
p/2ThTryy8LWMUXPj/d5gype7lwuHBZTzTLR0v8/+OtiA1cGA/mdAYFiA1hJEmRQ
zNL32mF3S/INuHll458EsuvsySB8lPDLMAKYUzLCu82Aas6Wh0LaGBArHHKKAACF
YhhaqfA+enVbP2jmSPOSag==
`protect END_PROTECTED
