`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f6brl5E01FagjVO7tcX9FlELJlzldVAxDuYdO4zApfQxZNxbtrv4xzGO0gCxnsD4
/hBzaeuZi5Tvj+fnZe7Ef2vsdt6EzyuBMtHpIEheFP8fuvXrLR8ez8sRcFRCPgIx
hqcmphV1FS0T9/2lI9dHtQDpzon6/X2mLipA6PrDL9RaX5DSBxjAUJgbbtQYaVu1
I47jiE3t7x3Cqj8/rweaekSSOrEIjKpDlh72YbmzcEsGfu2ZEl0lxW+/6zmzR5zn
kVgPVVrgKegy4RoXGnDt9gmdf18z9phjGC/MhXkNbNsiknrqeRqbGSCFxsdw+3tS
z2iY5o/UI9sn6r6Nshb47lWY4khsjF65AbHaWvP8vua7oKgZ6oaySnWgp8qqcshZ
`protect END_PROTECTED
