`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lWFQzOLlltlgZVIMYAGofPjRbc5mUlRQfUXj5uMza9IQ+jvhyXsHM56MyaLBsh8n
I1vShD8/aZHEjHDrGsaq5WBBvNJXs66BEy0d1E3MhHBdO5By+QENk7j6ol7kZABo
CHqPLWdG8eHjqkm7SSzYlaDBpuyDIwi7PSCWayhM9rSvYGfRU/By8Jej9bgAsU0A
9qjLLV/ELqfv/JCnL2T1D1kUa/QKd9HjVwcyKHsIARstOrpTdFz1P4dkg/WLe1zx
hn0U9vGbU4EqAxCUz3/lzdEIpzTWCv7DEaTwXgksWgHnTL8OkhgJVCmGehc/3fVx
OjX8wh1YaEpUKZUcZv/roxzmOZ2hgVJ9UlwQUi6RvAz/sjNESEToK37PKsyatMrX
2xVBZZhOBzp6Yq1RjFYBWg==
`protect END_PROTECTED
