`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l6xLrDiB8MAmc7bxWX+uOslo1Zoqos4sHuv7kZq0gY/IMLP8D3OUyEQDcojKeW5s
aQpeUVKX03pHeIstsPdJd1WGZafC6bFjmKegMxg/DHcehzA3AmqqWRRcXe4VsJNa
Q6BlXVxCGkiaNGrt8itccipZuF3smr5V3jUTeMIFAg4bATyd/WaSUUF3FZiDhYFZ
jVWV7QkEYnEK1dC0FhtrLFofhvZIZaMlZKIYskRi5FdHFRvEn2+GrzTM9UfORVvy
Td+uKsEHLJarP66tJPXHEZFtSu7LqHAcdUTUO5NSBgqBog72mqJCzhfUq2abSMdG
7hSkOaZVgsG9uILAkBgwhz9StjEM0m2JNeu8ApS7GCF06HfUZSKBUvJxDB7xqsxU
WV/A+NfGLVzxnvqXEzN/2btvnP0Elr7M/mIuzMgkm2uN7S3Th6zvYS8N864GJRiN
XauuHD7UFJ+Z+C7FVtd0yceFOleEeWHPF3xEf6N+0wQ/P9BFq7q5W7rz1OnfKYI5
9/n1gzYRcHVM9ajlQjhZrH68j2Udfycakgi3mubcp8U=
`protect END_PROTECTED
