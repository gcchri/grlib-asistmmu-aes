`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JkcNmDKA6eLAw6TnCL/wnLJDX7lngBsWZBITR93jISLSPH/JYyqDSKghXzxoPGDx
eK44y5x6ittqGPxU2zsZK8i/px3WINNnYM+ATbjHYkkQoOkq7FABomiSaKpSLy5p
KmkSFxqVC35ZiKorcqHMC4/0A9068MvUMKmH1idwew/lSEdru7zvOC5nzA+80v0s
M65nuucvXj+dRVlLX7336AyfIOIYMDH2GzU+R5CFKZuyqJtYQplsii2W4JZuZNKe
6akK+SnlgjPQzmWKCRdsiAFI7GHdtVG1qsQLPB/6g7/qHD/z+imB9YMXh34Z/4zf
zL41ieUGEepyZcN7sx4XYt10O09fg4DOB3iFkSzvSWyYEvNBEkLpMFGQOWhhnSIy
aqWtF9bTRZIurf2fXQtkUwex5q4OcWbQvQU2PjQKh/mwGEtJlkyOLce5K17p5IOu
NgmqaA34uhlo4Td0ocvHIrOPQhqih2bFvk/Gt7AM5Svzy9sMfLUnC1vPfNETArfD
9GzEEVSFs5OlU9CYOazgMuWbsqm1XixYao+r/J55nPuTr7augKcxPr3wX33+n2oj
36eF3+hAXN3GlDFi+3JfnMdVzaVMXpueymV8vgYDyWrTYBVi/EEjw6k8LNr/Lp44
`protect END_PROTECTED
