`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ZHWSCpuwCO7ovUssw3Ng6o7sX6H4yl35B3gpCZc1j8Pok+RujBCgzrTSg7WLoqY
GSJORLTvI0oAwZ6YQCBuKK6vFzPyu2S+u5Ojk+CRlTwJMqOZt+o54tUUnpEEOTsX
bw75CdpEfhBWoxzhVRqaW5E0pBN/fvAXAhpX/JkWDzvtYAU44v13CfP+iPoUUrQf
D2zKbSLCfXbwZRkMYIetzSdATAHZ3579q5y7fOL8IQ0lEsLpQRwOeoNoQTpdIqo0
d6etgJ164TUuiEYvHzHj5uuKXwBNJ9W62RDz8L4b2zWBQ9V0nH0h6OV31iy8Flmf
KELd/OuxNkP1C2S0XDxOZxAYhcpNtkcvGr2yZ1vnlEnJLokMIj+RGOeUHwlNQSiT
fR7YKoCNlbnaR3zuShvHkNpn28jkVP1XG0Qjg9q1wgrOh5PRP5RBdkUYPzwT7U6C
anzCSh521HCS8TcfnegYC/xCG1YUoUOEX7IJDwZy95ZGdUPXx9rIVPmJUSO2D8D7
iNXhrg0Q1xHh6DeqU0Aaec8tbj4ISFCQl90T7wH+1pB+SnrEDtj69IP520LZY2vy
NFe0ZDQf8EvXhpofb+vwip/u9yPRmDrMFeGuJDIZFSo=
`protect END_PROTECTED
