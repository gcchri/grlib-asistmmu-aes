`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ewtz1o8BqVE94q0q6ldN5T5uU9p4Mp9/IOvb0SMoee2KFCZsjSzsJGtmbb0sShcG
ZMKDg/uPR4SFOqOFFdHSnrm9uZ6aDn4vxKz/ZEpwlQCmFp/SYCxmGDKeywC+KkC3
eZdnuIRBm2pTSkvpzwTKxW/zL9c3XlFdezU+Ul6jJyGH4NfqFHzXMsc1B7NLQ+If
4whCQ/F2+vmZt8r/BXLELmrJNih5O5J3Mf2KDcEJy1+367tp0SnREDkhDntAEhQJ
2udEcwLbr5TsCkLwR/DFJaDYoTQgqG+gLKsDo4vJRnC1FGDfHSVHz7OyeTybQE/c
jLD2oCS8WFVqsNTH7Sn6/aFg3nURzJe4fKm8aJuhoeQHFg/l6K9tKPDFIqD02w5/
M0qqae9cLJ0kKE+UqcUNcQ==
`protect END_PROTECTED
