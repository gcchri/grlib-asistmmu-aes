`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zlY7oTt02zgRBAmsJG/OBugb9ulvwudBB/rOQpZkTqHRbdkbHWtTxG45gKnW+Zjt
6NIyzRXU9ESpGLdqAFcT7kqWcwWrbNMcuMnXoxZPp6q4gdDb93qHCIQpmNfeCCvh
MUuwGycj6k1qAZQOe7A6l7MO+/o6L3GQ9WIuciSev2ySpYpGIi0cBtQ64Dsef/yH
WOA2+gPjY9Ja6ldTFxw+OZvGFRfMz1nDSANx88Do1ke5G7NdKJF9+FV4V32Vb6RE
+D79exSg2NJpvZucjTNyO6JJaMRA5dakutEdxWiJzrP6xaqpsC8K16rMoZPG3ZJp
qbY0IoNazwNWoGQjqA2PPQkkzRVG02cVGZWc4UvD1sLDxz13/qq5ck8fA8Lf+Zp5
nMaqG+1rmANBvMK9HyTvtiPj/lnzHkdqXTyKikZU42eKsSPdddALohqlRbxjNgp4
eOdYPH98JMwaa7dIWX3zuvD++wyCv0nw9+rC1qX3SNBjFlp3l+u4AOaRi1DuphZ4
`protect END_PROTECTED
