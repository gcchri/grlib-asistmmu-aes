`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M0qXpvfdHafjLzVrFiMxklVJFAtkgqhflHe9s7D6mzFQ9ZJauYjDkZ4BpbeueIr4
3k6SAA7KWpiux67E87HDWYtvCjHFoC1aekwdfkeqqbpN79ATg8zXAHQ+fGznNcrh
nQhP39UTOXRjwY99Che20agFIGT4huYWrYGoAhLTZqDzMTOewJEUqcXAxeDN6KrR
wLpuSsX2lXj6qCjE3gXZmgWb2IjVSfiRA1CB+4WRfb1YxH1s1fDRJJJL38GItSL9
1EQeQtmMG9xLyShsIQlYOBESrTdCmNuatnqTEHnyqF865AvuHVayvPFIAjEviiF3
samXAD+HLBwU7j51my/vKvig5QP2vXxmqRtqPrfsjphH5r+abQw1JG++6RjFOUcr
C4JIUz/XYwar5mYJnrAM4H2PPdAAlG+Vvj4a3Hd6UD4qJYPcTfhgs9U6a/8JaNxp
7QKzi8aq/5OS/jErK6lztvZUBWATFo7i2PuutIkA659DVGttCxI+Vl8SFrARe25v
TzF7r9qauCJ9ouafdLQH/FSvwVC9Ese4lCGSiM+BSELQ4aBqVe3DObEnUX7RIFyd
6y53XCXT6Gl6DyrMAD957w==
`protect END_PROTECTED
