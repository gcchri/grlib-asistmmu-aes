`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fi+y81cM7fAdcOQenX5ZgL3sZiIbcVFP3daocPv/bjVTWwu3TZev73DzZs07MDpq
kH2vn1FwOwvSYj93PdZQSKrD6+K/8qpFEOncfZ+1l68WnTqIDqJsv8Ne4CXQfJgw
W7eaQWiT5IT6mR6t15fTo0Z9gzvmJLWwejMYcsaOunlltzlXrEmg0xxJSdCowdrK
2QibTUuu4YOw/BQIuGfdmS3QZb22VX7fHb5MLehXQ1aRJrA9mWrhd0uZ1YysW8Ah
F3Uki6xkyCJ4XRH1OelqXWfjTdt6yynXRRObBYxh2avX/TTFUhbH7WlG0cC0Ygcu
lauvYdhXo7yOiFuTEbG/a53bpzpfTMWl1Nrsp2CfaBob8BL4RzwtzJbkgW4/w8a3
Xbw36nHzYn2TOHmXQrggSg==
`protect END_PROTECTED
