`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sm4DPC13fgINAOdteG+b/41r/LqUd2zgyzysn6SpgncDP2pWJyZKyN3+sT2XOng9
ahLTitfCn6cwgFHzcJx2s4rdh4hP8euIxPR+3LgJ5yH1B/ykcjgV8GHDxDbtdaVe
qZZl+P+taR+ns/dWMsU31P9qN959V0WZhRNvMvETxS/v0XIzp9mKak5loy7xraYj
lSgbORt9HlVblwdgEoPWqX76IeNj37N2o6cl49SXHtiW7IywMPBEkNXbcQHKlPt4
pDOWrIW6OmMvx1PgLzVyLOuRhoAPgXamg8sBA/oKWkxhlUjGJjbzyhTzqfoaEQ5M
z6/9sTEwUknBwqrckdkVSaBuHbOma/qWmIoavH6c9PSbzHOu6zYuvrosa6HLKw4x
e10uYfcWPFICbL25pRZUU9EBSG4mzRm5njoHFnIqjT/yuDso/e4dRUA7fFmuiKew
sEHTTlWg/KYEc/MYO+7zR4URjyGxuBbp0YdbBIyVkPajnlZYGV0TImKPzDJvy4Di
3XyEeps0vUw3AUWnzMJg/r17fwFR8YO9roKCE7y7P00YdXR2Y5WROAcM4MnNwaX6
39s3W8CvQL5KMlhYHuNpHck8kzHyPmQU21+CgwijxYh+4Sgf/Uy+q/DNkG+SM1BL
WfBcCSBqnurXdyMe4f4OACAH3MoqyF042RASuW+RAu4=
`protect END_PROTECTED
