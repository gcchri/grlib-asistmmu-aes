`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
codn2JR4G0UOakkbKTnqUrqhTDqRtiQ6YMvgwWfzqRah4eFjGK1pshUb0viFho6g
LIEC03gaMSNOJ7lfFoj3XHPx/lD8dNt+Y8jWQNnxenfLKWqUIL46QwKcCNCAhly+
hCOs6vkgEGoV8MXJL8WrhxOq+YH8Pwkh7ZH0Yd29tYXfRsRvL1G6saWopGF1Gcue
m8wNe+0art5eu8vorKCS54s41n8NIcrfIYFHUlUebdAkFtYiylzlxyj42DnbCbLQ
P7cam/NklG2vHpQC/AXDoi5VTMvwDclyXaeoXbq7Zgk=
`protect END_PROTECTED
