`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9r/nPJrboapgW/WtlL9OxjNGvBSDc2d5Wz1gOfgwwGPDKJF2TFKShkgxQ/v4yRpQ
50u8HaC4xXke+b4XzbZlR3iHcmFTHhU0MyhGYuGCty4/BlAoS3JZNcHpeYsYM6P8
sN/ayUyfJnRdZVgt30DGsslg32eIVzlHDojq9eh1cfU/yRZCTIp3SH243PfBVa9w
iANidWBf3yz/Xt0YQvo7s3THlRh8DKa61atRLxeVDogu4dqAdB9lA1tzCtu2O7U7
rcIlvp5dNZvW8xw6xfjGtTMHCAFoFtPEwP8DUZycemLhbaXhayxW3iYFjJ5dUrsF
195OqYVEt/vcM6wQdlfjRFl36dE2g75/Vf2TtHYdnunyQBLI1WNo1RTUKpWQKKCb
jrHamicz6FWQGpPKtVxSPgYdQjQqYms+d8ReVQzJVii79x+G/y5a157ei1/wvzdq
nae3znjaYeme+HYhNQb2BVH/QP9TFE0BFDqcuOoDYMf7sjPanHH6kL4dnNPuWt8i
`protect END_PROTECTED
