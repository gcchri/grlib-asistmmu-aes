`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KcDIiotYel2zBelNtDLXzqolaO9+PIL+oGAt/fuIz6BfTdfWhSw7GKslwf0mhEQR
w5iEOij983/2X07m1LOMQYemzzCTKsrISMfWAIrkAOkh+qT0pZ8UiS201T+3lQGu
TzK12WtVQNGpHujbnfkbU41XADclB2JZsl5ll2qG0nse6lbfYkzjCmOVWyXhrZuU
l10u5/1n1KJLC42mcZsNeTh5uJBmTp84xTmjSKXxP+Fib1JY2lOHEKymZb8I3v9F
5+A5HdSsIMGv0Wz2KamqSqmlLCklDJ7dWz1zDy8EH5cwRhuJ7+mLqIMp49a1Ddyb
A4C+7PGjpFEQWPo8QeWTZLgTqCRHnTh2qvO+ql3QA40q5ZNfo7gzBwCB/xwfqPlf
aBbVWWF/UCsDZwFglSbTu2Y2poNhh3PT8qYsuMwQv7iXWobS5kljs/2jzgFyEBQG
v9QxSGEOAeDjNTs0MIB7zRYeLJKhJtN4F7CyABDkn7kLtSPX2VDLOeMYrDOOBH9y
yqaxl89WcMpq08Dq4nCMb/AO3IRavlSbkYnQ76ahZZ+fSeg8h02HGkIyzd0nJcEX
kl255/ACZDg/lIz2cctMiWfw6QR51ug8EnQn8VJuE1LhZNTD3D1oEzCSC5gMaQMU
NQTX75BtSttHOgo4TfxbqwZ1EgbNFxRlNeySxkAEwQ9/8hxTZCzy8rK8xCkJ7rlq
ClrbcN0HtGSsEQ1mRXtkRKbyD+ZnplBBohA6wFvMADEnll7Bj+v8D/RsKW94ChF6
+A1yhTuUOuKoYYLAp/vUtrU/4bbzNzqHO/y59lx0q+j+ZdakZQzveN4StseyjiDf
nQ9/mHcrcf1tesJBrg0Ucbz+ajWxwbSYZiOVwXXBDOy5+Jy14OmJDS923opp1BhD
ZxYA6B9bRm8rj/jkX0hxSlVyU/IhATJKdcFy8mletCH2paMWZvBDNhsM4P2TyCZ1
4qNZaVis5yyL7II4OwP7P5hO1Tz2R1LhL/H6ssbLsdKP/IJwgokipVSqg8z+GOFg
lOOEVjr0fxD8RhsWhg0Jq0tZ8rK40R0cDwjfGN+2t27nOFJ1g+kRtsNeSU1dDhhE
rL4BRzQcNr64zfpkN3vG+f+d33+h67W81eeyZR4SBYEi+aGZ1ke5+2WvbZ5rhDpz
F7DHfVNgj/MKO6ZlWr2vUbpxNGoGrDLcEPDJzStzHnjJ9/sfSXaH/i9xzp0jggBq
glqLYex1LMh8jrrfVP95ziIdk7SMKVwb9Yb5rm7R5NbMWiBbzs9ieDXBGomZgwsn
MSE4jK+1yW0gC26w6OVAe7MGXy2dC/gSfbHclVrPxefRZOwenKbI0X7W8F39a9l/
YQ9vMohWTukRzCDsFji+nLp4LMolxv4fsmyT0e2kPRQo4DTrf05h3s67zhgNpda6
t7m/ulpBVRuOgcinpGBCpVn2ob/8TCutQjqpWgxX0rnlnrELCUjOVFiXMgqT9aCT
wdvPFlLBVg1ThzZI2D+/gVmbf8dlE7lsK2EJENZbwBAhkJK6/SX+9zBehyEZ+UrX
nsHxlSNJ+O3VFFnnYoze+rXjWxQil1F8aQ381DoTuV/UFeciFVbLX8uTXwSi9Ywq
m+mawNkciCFvSzNSOzhmA8SFXUlYMT34SwyFgXiXmMTSuHWaKRx9RjCLGTcpelzu
yk95vaZsdYvT/5//B4o6gcs/6lQ+wIipGo3HyExBO4nrhHkgoV/i6/UU6wG0dk6r
XsLRwrnoDL6+LonfIZIwHgO4Z4fxL7Q4eEtYiK1i/L0iS6ySeJ+52aRpnaycHSYm
0bi1gda3vNGHKUmzW8lTreov7O3250g3I2BZUJ9RhsrUpQiVe+0G4M37rKcNBPh0
MotrckDeaSQnsakRb3LfcZ8OdE8aoFAWy2Sr3KAuhjyKa7EBjJ7NwmL7Hs4nCg/l
/kcfWoHu38uORFUVPnn+WduoPtwH61uiAlbKtsh81+AtahySWO8smcvvlEfuzRou
zCJzeIEQDuOao9JKyltl0KZNlkuv4nbz2ut73mzSsRiOp49DdxRReqLzvr/JA5zw
wmZd7pYPYfCZKUICtH/PzyTu9lRiDTrWf6gdeDLQbEz1AjnHI++0W9/Y3Z0xJTjY
dUE/Vo9W3L7fiEl2BWx/1PPc8993hWWPusRJzrskk3x4sgZEorfq/nPf8nsNChx4
Qh/Uq2RiBTl5jI7yaYww6JoXIK2juNgr7mcmQoVROGU9HIELvM0RoipRW6TH1fFd
NBhOraXuK4muJwpVGWh1imdyyAdepyuuRxWMcIJ4BaHFXowGG2DcsKGEV2C0bLMo
o9ngOBlByNmCq5BPcr1ZfMX4pGvFr51kMHp8+brjeBl5dQn3KI5lxDRGKhPTJazP
58TXSSIKVr78jGJlVfGG5XrHtCq2B3Zrhn/ADs1nQE8KE95/rMgInCCljUJkZpOS
IVt/6DajDDzwoPP8Mqgk5YO8Ej2V5s116ufhTA6VrdDKEt6h91XIkaF9wSP1Ec92
2JCGlLrTZZ920b1ZZ/S79QjaGepyajgCx6gCy8BKGYe+/9b/deL+Zlovhq3CIgtG
htU2DjRb19CWrngpu6UoJLFWBejzQZVO7caoUQRMpLYCC03MYw2djmZZpAzZwwZd
rdV/cqZhCk8BUpj+4O46VSZT+8hRVS7se6I29Z3x0uuw3fB3+/h+SRbSu4WPMmqk
pSpqMqNQyrAN3dmlkzj7MEE6+njpWFv9x2NOJ4XiVrQL/lRdIxf5EP2KDxBBUCDl
8NWG5zoxqqtVD9kcVET1pIIkkZPKb/149KATcdnB9qfguqsp2yxr+YDHhbIPJQJK
kAKVEC6g7E9fJBMSkSIHd57D2m2RVSHhA+pl1mmqAhjmmFwMjj0Fh8967iqJOTiV
tSFGWlax9o/fDPaTm2ic1IBRLDWfRzmNGBac9UZ4IYzC7F7cMBF9ZZnfw0pV6kpx
+q3IodFJFxZ8OtegIb3bD0j7sYlRdYyKG7fiCpqpS8G+j2dQ0PkS1p4Xje1Dyvuc
pLDCRmHVqacgMAUlZnvv6g3ZELq8ECWpFFTsvSkdrkEewSt4kKtTI57MfVOIUepd
KSpW7XcrC45047oU0QuOl/x4wuv82dZe6M84gx9bWh0zcB7YtfrDiqiEGjXmZuTs
qGXXPFwUdIi/06qE+WBy2T+uBFnv1Z/foqKRQdanJ5/l+xi/Ipqz3ng0yhepNYNc
`protect END_PROTECTED
