`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cc2AYLnXZp9Jpv20jKM8xdmWSeNGNi3kUFvPnBZx78U8D3VoK+UMxVItJNW+4ojM
qkWKo6HM4UKG4nzkmPszCKbWtMMKKSWYtvrf+CDz0x4nct3za+N2ZXp8sFArd20+
4o/1010Y7PNAaOJi+nKyPt3HWLj56TrDUqArSa19Bg59k7u5aD0E1RKnV+CnuZkH
Ws8hWYL8FYq9ijo2dHPBjYYIxCyWdEjH8qDvZYyFpF+tBKNQ1mFOLodEPViPsca2
HoRXFKWGbnD1JDEiBQQ7hl/zyrT/QEgpVaDhLCwQLeLKdxyg/T52bDlLf4spAb8z
CRBcDR4cYLn/CypC7pfP8oN6vn9bDoskeQ6UGoUqV4ydqtMKLuetDq1YXzXX+piH
vqZYn8uHsr44Mac2w1TsBg==
`protect END_PROTECTED
