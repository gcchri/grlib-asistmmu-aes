`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hM+UcQl+uxFOX2u1k49Ptf0d0q4Vp6jWyBSTKzO1TSxJdS8j0/nPYFB5Vlo8Memt
cpRjurNztzXe1xr0zkB8UhafNB/e2FO25hL8rOYNT+54PvCmbln37zZXdl300FRh
He4FnF1rTxL3c99q1M/SgxaIASI/C4oybdjOvk+E66tSJDmv/ylUvPBdwJUajY2x
EGGU16AVDQVK2rZNsTE7uKEaiTBh48848f9VE37atPcMALWySC+OMzX1hPoFVfZP
+wEww7MVZcZegTHfoynCI9y5isudfQg1MJFEJ9NB91rjKEeOK92Nmil7nV2zqn18
h2kQy32jxqX1XBU5/shgKzTny/Bz7xvJUoCDLL9BQJf4m6/j/hHFldceeaecD2i7
3p0c0a7g+bjT9fvkJJrbWVZZ6ZJM0k9NwmCXL1DqrUk=
`protect END_PROTECTED
