`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Hv1iIC6lfgikTSBmGMR/rFIfRh7J2A5bYSVCbzD5S6JkTCzkwNYfIRDsPXrSKeF
VXmHZfiyWssj+xRdBbushPhbC0QkywqBP4nBe+cXtywUyz/ag+I0D0xiPv4zgKXK
G84PKGzu0XymnoeOTwMTiCLINGwfcfkwOdCQ8Xuq8ILqcRnJ7nUrSnwu7R4KuoSg
lUUfA1hR1VygIW8nOpzWG8Q37CpOEwX4WbvZ497W04+aCc0gu95nuZbi4kBt4Rjj
LVIoJXwmmFgvr6MspZU6PJssI40gfp/4HQpbtVSTk+hmOu+kmaP+bmGofaEel8U+
U5/m6LFWgETnsTfstaLDEku9u02q+RC5cS+DeQJVjJd5EX4flrg5hfqJ4RMXn/wD
8Mlb7LHEdJviIb6maS4aXg==
`protect END_PROTECTED
