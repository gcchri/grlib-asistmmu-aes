`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dt0WoMOnQO37OZeyZghuZSVYO6aevqGkbeQt0QLBy1qHznTqrZlfZttOsrcLCyUM
M34HMfwZd9WIxNN5Qm4wP/5ccZKQP7K2AniiD7L8vxNSgfZi+PIkcHTG+F5d6IrC
TWKjyXpjDGxFJzETBGyMRl8udw7Kd2cye6wR7kBw5GwaOz6AQlCl32908hHMyQ6H
05KWMC2l29voISyBYbDXKMkiq3IvsAXXdNvwuXpBR7arT/IvNa9Nva0dc2wROlwF
XAanI6Z+mj1Tv/+4ieKYmiHEYEnLcgP1m17A3gZn9YYnfXGHkFAQDHR9v7Y76xMN
iCuve5lXpqkyQGrQpgLDdDoFFEOdyy+zs0fnXbffVIMapq7ExK42A1RBqyXDPcFx
Xc5WgG7z1RfAYQJGD398SdKMpFyMtV33/+vsE26gyLdJN4ffGpRzd2PpUmLY+9nT
yS06svNlF2Bs9fVedXBlsqGMRichjB0GBqTXEmyTxVExpY0SppJJ9zc8OUSTshGe
QnEkdEZJudX7qWD8hHF1ReihYMw/NuTIid925kOTytBChw4g3g+IMcDgbwdB/4Vi
cghkUVygcpKheK6D8k/e/+fRu4BFNlhM4FmrhGeVUd2u1rqp/a8N+t9bItHLIENh
INqQKy4pX06ZoFkK4M1VMBPyUhudbBD2bHucH+CwelAC2w7eDNwUpLSuTojUN4o4
Bw3Fshoh7xu1vrV4K0X3OurJ9aKAoXb1plHP+qauZNzTZ82FjH7PsUJESuA12Ulf
Yx7eBKh5zg6b8p7/ZDUsLYycd5zohqvDP9UC/Fs73ZC5vHPovKjpeMsXPv3pTPd2
PoBrODDfe2Vca1fiPxSixw==
`protect END_PROTECTED
