`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PI+TpWtLaPLnPxJhZvUpXTPUxbLlRUtFWjb/D0gXDqE2QFx1UXSDKz6jno0KkzjF
Rvnh48hXD8+e4xyFnyV13irkZ//FOhhgODjO+O5mrpN1+wm5QZMQ5m9PhzTAYM3l
FwUP2RFGIhr8qnB86ns1vuDeeEonsmKfNYfgoo37V+GyKKSHriJKMEvu599yWp1J
RN9aM7Pi/WHR1aRtxrHk4cgPFnWz5ggk2ztrX1ikouvLJ+/HivZIAE7+fBiKFkgZ
7yzgoS7kbkhqN/LZvrqsSDKUd9+bQyF6j32w0B2V0O1gnJqkkrUZhYCC8MrifxoY
2M3cqJrB8GWzWo7P3EK3N4LTdwWPRW75kfEnD8CNOwBAYc7TG9M/rjZiPXvTju/O
t7HKtO17er8G2gLdyB7zDY9RAdyVgL08ZzvFd3x+Tv5i5CUEQG5gaJFNUvqPn1j7
/kCFlR1iNpsSR55fedI05A==
`protect END_PROTECTED
