`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WsepS897///PpH/CrBwTGhnIvVtjB+kOq0xyILFG4GmpkWR19M1jrT/rUAqeDUdR
rDOgUcYohRgJKJwt25ZPSuJkg+YMLjdl8fE5l29CjC0/B3ciQO3Tx96kYVGCaA5x
ikJ1aytUM1dZ94fODqVWaP1jZFhlFDuGCeH8LX1B/El3cjLwJZSN1AAEqC6VgAeX
IQvhFFv32YJjHkXjTYXLbie07URJ656ysX0QXmnyZv7p4VZuN1Wsvy/VwVTbDUhl
Tj0QT1bnuGP5a95cIQ2logcAO5rvTH1DVLffg/NX78U2G25U/6t46jJU5G98SROM
cziVaMoJa4WxXI1GynpveQq6HsHn+rlgsn0rMYdiRd4DYxXVcKOO+nTaFiYKgMDL
PvDGGif2IbDK9fB9U9jU8+zxaFOq3Y89ll3MJYi9XN2PxrFbTHXVlMkFHD/+z2an
FbyrBKHr/Pp3efwUn+GR/3KEgPpu6G3iCQDd7yUWPcxSBXxc53ZeZnRn97UhfcJ9
74JeBWcwSlFZG9vhD7MpsVy4WN3ii/q6AoS4PUMd77gBl9S1r41GHmK8IwEoib8+
ICWJISik9tYgg/lPjIgLuvPd6s/zwCqUbt580aFJ/g72YHV5r6I13RqT+eo4FsJ8
LlJHDDgvTtwDnKO1IW0KUBd1Z3gi08MwDpA8AHD1YwhTW/T4hbxfennQM5IdIJXw
8R4En6ONRsaQA9hxkIfVp6tH51Pxzb7FaflRXoXtTegI6EWnausw9ptJfzyU4f/S
q6gRZ2rMWz030ajBuNkhTsZpqCsPi0pLIgk0wiEk1Th0s37rMcNtmF82BrThbaSh
JRuVJQYS3DzfTATou7A7mawn1L1NQITz3bdrHHeBmeFcywC+XAx7gc/xKJ5e/NVI
67/7OmWaqwE9tOeLnz/6ipw6aM9ApVQZ54kffJXyS5tRPHYa1e3wLT72rdVFPS1B
0canAOdeDKwrxm7w0+YMNQ==
`protect END_PROTECTED
