`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ku2BhaPY5UPRD4VmMtCMUHfWMqGZANm7jrlATb/NHbMTwqLIvlH532vZsFCa2TWS
1tdZEeT5f1txwnyX86gfKNbFwUpZptXqt/aWfwUD/xZY+ZwEfBGzcU7Bsl4rnpqp
6uFIxzK7Slvs25cvTKVa8i59UxI/vXZNrs1a7T1rcas03NAFTyipLmWL//vSdINa
gmA37YKT/W4TOu4WLS+/98H/AniACbshrfWLkrnzNKPNCF/2AWIO7M//Jr79v0YW
`protect END_PROTECTED
