`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mrBT2MghbsHu9hVbWl9mpO7KXVTxz2GfoetUgT/123qMjqpMVsGqBGBx/z+Z5DcL
N4SbJAz8jq/k7alu4xCetqWwhhRqPEt0ptc9+ywVvTbbDli84gcDXtpYRDtEek79
eNJzI8/kkjcAtjQZBS7aHDbf4flb1CNJkpflYEVLWU2SnWVtbsr9E8Wlzsypmvml
y7tVpqpxubBs7INWe9hShvfqt8HHlytDDXITb4WC0C0zAGkiVB64QOnRTSgMB/an
iHK9mnuqxuI+XwY5bLcxrexM6zGX6GVxnLFve22V6y3lD7cgHCwf475A13p4tZBn
hKRhBjANV0EmbJO6EpM3JISwhI+7ifKI2tb3rho7eWFlQtgtwt+TC9vLpXsCUtJ/
zqzWtrWgAS/jrtzg+HVJI1CRuNRXhEAT7YC5HM4G5lgg4C1wZnuTKQxzwiWAtuXl
Sm8DyAQ0XJ0JsmlX0IkCoeBfR6tBi7YB5TEsglWXvmBS9ba593ENrhx1cNNz9/Fv
itjGYj5vufhYD38i7m6g8fd6qHkogUL9VSchTxe6AUS7c22vHn9lwST1ebd6dsNk
HsmKKmL4u2TJMBDCYfai3FE6g84wfuiZWwcznaEol8e4IHvoUtyCXpATdz3cYarb
wn9rpPfOxT0EbClqJhnYwvFvpD9rlyjDYo2xOXM+TdYTxrG+4FhM8vZ5cLfZsuS6
uG0JzQ/ZS5ogoVPZ2GcGlsPu+/KFp6nWyKbyBlh9uQmjFGh1Lau1xFroDu7QuuEW
UuLUBsPb3xpLbBki4HaJSeKm6Y2eL8hETbWpb/mJd6VzSQzyjNoXkWgvq/fuigqK
uej9jPcQOw++W4TJZkYoM7X6e/Z0QLH6ZlabB/tDWvc9Lmak3Y0RpI52RKz3rUf0
8YhqV0aLOGgLqnF7O8U0hB7nOO+xdWIaXB5ZC3luEdU07QcNEPK6m6WvBE8u86X3
JbHMbVbaERrmhWUN1SoKaKzHNs0jsCBb7IzqFm+JJ5R0x78mzY36W2CkKyw9j5AP
GPcklh31wt/49Q6nC7X7BK3YtT6POHEP+uowCMh42xzU7XL0WX0Pb1BhIK7MVh3t
RBHMPYewbQqC72xJDv6IW1ZqeyDnkiXOGQiQQu4CZqkuuZZXbtH5D2wCA+it6Jq4
DbnU5kCi62FJSJZOugql30S6pCSUu/Y1ftgsm6RMvwbOiF/zb725TIYxSDP0ExSw
dSEvHocsdOPcPhuJfHF6Y5ro6IlFr5PVRJS3F9EVQB+HyKBk3TJ3vAxVs5yxUUIN
f02GZ4Y7l5nAmE9mBTlBLpWOcoH9e+f1u35wZ9VUEA+MZn+pyTTml3svUPtmxbXf
VUtVtZlqWGIBi8zVl+3W8WPiq7CDo2BgPoCYkGtjT2f4bXag4nypP/lYciSOi7dF
aPT1gKpVGz1t8hmJOeEwTrO4JPkpPY77VHbKMAAAxXt2D16OKFQqHxkHDO7kLVw8
N0IStxAf8pcCdZI6dXDL9W/z6hmMXkbfk27Nv2yIvEWaPCkrD8oxz6phu3/foioT
Vr7Anqt4tahpH4Ci4oQIvhtqRCvLzrIsqHNdAmPxaI5VZD83UXnZd8xe22u50iei
j40qGXe6Knio6bDMoAGRaT0sbl0KSAsdP2GQDUCA7BfR0HHEm97vbmQEDp/8o9nc
16/0Z/zkEjbJJiPrBM6gpQ==
`protect END_PROTECTED
