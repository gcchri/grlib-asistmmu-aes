`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bRgV2eKkXcConIePz+yIbiL3wxswU7xmAq4DB8/FJwrdWRFhz+AdiWdlAhsBvUlb
oc6lD2n11FcxEZr1ed06O4uP0m5nOzqNYuqaWjm7ZZlZ1p8GSEV4iNj/cZDMUYc2
P2Dvsv6r0H2I+v+mxv9Mk6U5KjlgoM7KFnYidoNw56mU6nY5/2cANz2iFMNBGo3h
0zwzUbZxp7imEnf/9eXNG43/4Do+nEA5ULpViSjiB68vSOHgIH3BDLQtuh0NH7OO
X1jWslfb4o1SEmpjYv4d+huKHlIbrvVccsggfHJWEjQrpgs0fQ2ZpeDFRltESoZn
utMHS1aQZ9vfLACHY8ysZfK/k3nDhLSDL/CqYKoN6VDfjhCesXWXJXL/Q4nMXRqE
OHsSpniAomb3w2Jcx6hmk+kJWBKrP5kCnTLwhtiUc3rC1BcipfVpQSliJeTCCPz0
Wu0RzxmYl90fPNUjLAv4/XfbiC5SSiMMMX352cKM0l3LHMx0/n1LVlo6oy4IDFqr
sOCNPIAdplcY3mhmKkJ8K6ivbvHhD5o4W/ic980ttUtXWlBAXEyViEs1pdtbe01Y
fimBdbAitl/HclxiqFUJ2oopDhPG0jnCtnRXfNo9dXrrftaesexRwOWrKN7iLk2o
0zzvb+F6kZGQGOb9OXbCoASY+sxGzezl7XZ57WMwOtc9yohI0XygT1zCxKHJwRzE
useqEY5l+2x8mSXPeDUxwDDGkb/sGnB13N822oHQCHkBwU7sykQnm1mLnRtRvzXo
1XViKrME9xUgZZXypXc7UpmuzS9BOfpQ8f0EifrSK4HE8slnCQwJVen7wyk0Tf/9
5BxCbbr0DTwU2odxy39sia24UQeRawnYemoRkKIKWdngvkDJJZx/QGw0ZYphYhXZ
v9LFvUKey4CX7122KHrgsy2BN7pHbr5+wourl87MCguYdzigO5jznhDjNIKpgycj
EZ5z9eV9U9G0Ski0ElaYZIuAl486XR83AOA5imUMC2vZQqc3E2GBzZahXsTygv8Y
wp6iRz9VUzpHAqB3jVcLlpBMbc2Q3Mzqn5BtzKlOmZS0dt6gas/hiDqdTVWXc/Rd
JHRSuZj11Vx/biWjVj8srLsUhpYULCKUc8dOtP6trIKflM9PB9qufskJn61yFTJt
Dvb5wubV4FeHKgdq1fenOLS5ZJ97C7CqGS36zp1y6ZCFu2BoQ4zsw6dJ+vfVxJU1
ogQvrF+sLK3J83MljU5OcEtdqMMZBwx02KhqGfdhBp6/T/HOKS6uq3BkpuG2YiXi
XZ3zMW175NSITxvqUkcmyWsy+QO6Oxbvq7k9bulpE+FeXU+4eJUlaGlhijn3RkFL
hgaek6T6/ycd5lCn8KKrsRmpHpSMlCAHdopEFXZqmfe0ubguYoBY+a5T/zmdeUhY
q+qOz0qwNe2YctI2zqRgus2wqgFE5EzYhxShcgC5UaVkzfOCpoyXRp3LgIskSIvz
`protect END_PROTECTED
