`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KwtMNUy3LBYO6Kn1BvD1WyvfNhTGYYJQusKQd8r8B/+3pGM0wg0OcJCfQyXBRFp4
HKTXOZzJZayaYdyPhIwdkcEBtl/T5MvHVbtFzdyFwcbXiLkDc9r2USxIgWedzHBY
pQl2E+r6zi33CZpu5z/dikjfAdLhXIhLxxh+YYZjlR7SzaKklO7ho1B7eoVTocpc
vvWa2YLv+AnQydIbDKuxSjo5gztnalKGvQSBiQ8Y8s/ZWiJALHB4wrpuktVQxCjL
OrPlX/hnwmwLZiPAe9oA3mjJ88hU14SHAnfY0JUG4RunvtsUFXv0VwRExrWLssYa
fQl6JgjNcnLo+0FkCGszjUXWDhJYGMpqqBIS3ZSXyjCFeZkyCER2QSER1o2vj3/Z
3Swx1FeLBsV3ZV3i39RhuD2sm+xOYIc5UAxXVkTOve+ex9ZCTdI9aT/nDe8ckS3P
`protect END_PROTECTED
