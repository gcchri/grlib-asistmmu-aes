`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mpsGq6bb24T4hSt6fnu2aSfZ53xumm9eqURIwpQSlhsJd3M/BM+kvHPTGSMFDMXS
zC5LCq2pWy25Jsy59b3ILOBCQim+QhL3NxGuihQtc+THgWj+mjnT+QDDPJGFKsGN
zae3HhPqHifSCUZ7HTPqL/8QIyMQ6bheBpvAwAmUxlLjHab67Vdqf8RC5PjMm2ml
sCyLmhu+dAJvnH2/0BeadzuEXEPXXcQnvQD4k0lkISQywG3Xx+Zzs1LdDGPRYBLa
SxotLe7ucvUVVuD/ZgvdKImQmYbewMsPMK0PNbJ35e1FQMaV7M+l9A6/s8++0ML/
ndUOHrLM2R5fq3hUOW5XBOeVKOrKfAAe9ev1GiF9wJX+x9FGppSItnOM7MkHPLUd
tUX6apXoY74n5hIZ4PSW6Q==
`protect END_PROTECTED
