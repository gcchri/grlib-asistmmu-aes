`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qqCSJaLXP+P+kZ6/ENNgXpqHEt7Wdz+oVxUifD8dHvj3+tS6HcpTM+PxYX3zRyX0
VWLnNztu59fP5+mN+iSwwXajRR9krx+5/8xjn+0/ee3sbZgHfwtS3T/uQJCiFTOG
HAk00Xm/ore15oUOndpDuiI1cJyzcGmP8UVmzMHVqhjvQd2zi8+gryLfL3/2qdBL
83PEdO4cTTc/iDh+YTs1AqFoSHBUJd7bRHJotduAn87E5+8EQC7uj16BZTKle2L8
WRnq+79Zs764r5stFnpg2g==
`protect END_PROTECTED
