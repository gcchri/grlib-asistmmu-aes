`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sI+SrmLSAk5dJi0Lh0YOIWsSHbIYPaJIOeZuBTefMAbV3IIFDphrComK029ApBe4
yzPIr9Op2aNuFQS8IaLQ318MQlvqCFm8Kh3WhE+UN3cQ+MaJE49wgLpKuql/X+ed
aLLIwcx66KVlauxeA4Hi+2zXrIRbYaCS2YXi2NpaKFi/iz3rxZOFp+feBpy6gDN+
dKOwIo9UN7Z4taA0erFUgYY5sw3fFABiKgSmKtXZcdWJjdbzCldbReDP/+4fITpy
BDLzn4xf1diXSn9svv73y3UTTwocERckCP5NCjfM6Ya3/2rFj7PIJhQf5+vXKvkH
WYluORaf4pP3xVqKjp50DFOhAKfY++oqvs7lbOC33ndRT3vpjReJHy/VjfggxwgK
9pnNb+mRQj/mAoV8c5zn+m95QfO+byq+UlVmDOxR4wz4gaI4ZrRYbqxBK00ddzG0
o1bIKtUb6TxYaqhAa7jitRL6JsxI72aNXWD7HMpIZiA7j7SjhyKCmGg6xMWgrs5i
rWWUuZEoKG95HNxVZ3z4hAiMi0f26djtwgnaWR6pgqX4x4yszW9vSjLTbV/UhY1w
Op3c1He2uKHvAzVbFZtz9BmsgVawuVgZpuNguJWobig237R6ZpTdLOcoDj0D+xIx
bqDzvSITxHSLW/9cnSgmtM3lUzP4sx7T5UrAhYzi78cumOUIjpbDIoAMkzPLlTWP
FLXx2bLRzOpnOXel2XYe98jN2ly8C+nIk1KSstEu8+nt4vV/R5Lo86OT57x9/+Eq
7KPmkaX1Eeh7u15R6LywUH4RTLoXpSK3tbLXlAL1igDhAi8hTW9hpvHfbK24Ex18
XtNl7X/8qSHGlsLgxWLknbQWDZ7FFRIB0KYDFDqoA7M7fZOVM/OMKEaHJXh7GXln
oB+l+5h/xjf9a5QayX23TT61w7x0ssmkwZpWfZfSd7QKvYjuVLlNpEShU36vTPWh
vFDJR7l5PYM7V/CyGMtcJ1Ue7hBKl8VZQtcAUmDWh4/kBOuaIPP7/zTXB3ingUvH
EYBOSqgo3y3eWRPmdgPwKtc+koyPU704QmAqztRT/ixLv8oaa/vO6EHQRWJ/1ZCq
wv2mPxjMdVymhOPHb9j56TqKhpLEPG4l3ingpN6gXKH3xTPpJQ+lkKRvAnXAoIpj
0Xt26msiyrz4VnYAk/2de3S8Qf2TCG7Ak9ITKKCP9kCDLEaJ0gqLfRUhIiR7jf0Z
cPCAUj0i+cfmlOerC86+cpaN4xqPSu+sjctp+RPQBI0KcJolwfCxx9p7/TU0ITnY
kcJwD3Z+ot4krfNF/Jq8cjKx2VKlwQSDE/YZj8MoNEk=
`protect END_PROTECTED
