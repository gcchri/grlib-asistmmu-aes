`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+fjAn57QJNhmcs1/nMO1Jic3Pt7PX8FvwtBu8GZwmVBG226GS1ZaeevBX7IfpM36
aXQda7hL4h67oczVJxJ/E28J4BCeR00Kn8h4Yn57/sm7lhNEJAcr0hH2FMQke/d4
9C5NAeGEaBTzjCESG5a9DPMelyqM60J9yGnWA5trT626msKpz1IXXOSVyKP3iwd8
GnzQmT/ZndYPGgyIQwf365cKw5YPKZTRENAprvrqEilDgWuNl6krK8No9zieJ0Fr
c1t4pwUf/ROL3mpqvOsxBLdg/UISvPltxU+UMb45anfi5R/3eSoCne2bPbg09rww
S+Py/vSUhZwPlOkne6rELQ==
`protect END_PROTECTED
