`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DwtaOu5lIwar42NMAlfuOIpgZvYd9AqsbNAmEj2OuEBwF69ElSKepubR9iqhhKA4
k1gixW7QwJx6diEpzzf7xRuMzAinaimPstyZkZbv8SW22/RPlr9TkWum3nO1pbCC
Jzadcbtrkk6WHSharif3rXCXgwo73Fji3oO9xU2g3UzPL0HviLsCnM5xPDLxBTAZ
XTYqzH/GqqbBdK9DlSCCxedS95luy2qVKNac/t/s2YfWIE72zBLwSqYVTsShhc1/
mEWteUsR2WjCMiJJ59CnShU8hBSv+bz+JUqh5R27Wbmm+e0Mz0zA9qsWCiWlZfB5
PMv9Qz7lQ15NpwOPFGgksm3Nwzctk5t+oKea2RJsYuhJe7RVgSiM8J2Y8smL8zsn
gDc+a3Y0piY9J+GrDZFwcBNdujQ+ubLtNb7xFR3aFqEiruw7202Q3mRZNFBn3tMK
jiiigajFwpslnBxKA5B9Y5PVa3j094xJiPCkk58MwxttXE/HEJPGDNYiYsNvRk0A
`protect END_PROTECTED
