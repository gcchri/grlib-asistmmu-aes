`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cfY6HTo3/7NIFHiee0E7rUdpLo3UREzjHKaeyNtueH1HB7FxNF/pjWcQi+9e4xUq
bG6MppaJspHdK0XCx5/R0PqkMAVibh4GOendAdIXDshKb3s0ZqUhefYrw5L/w0SH
QPwp2IURx/RwggDjZ/TgmU6RfFbiLEQntoYdMf7my0lPSVcrNEE0uBn6PfuTr39h
9NlQQTbZwFCjRpLgLz3ZW9kt0maT9Mr+vRJ7hvfdvq7NPogtKC3Hhe1IWxQeyqMH
ZOp8smAfQhauMPx2V0HE6XRBu7ediCJywjgbAZklsa0vYjJDEahYz8EGJlVTr6EC
ge3jGSTn13Yi9/S1BxpawN2udgVvuqAv3XFoPmTME+YurqslyuVqrEzQ3awHolcT
zg7zs2fULjFOKYmEmO49Vueqv2xVukOyNb6Pg03N06+eMkLCWVNAMtxE8Y/u/30N
Liy1I5CpbVbMqZ0x1elDdA0hbyYyK9nH113KNXImD5cgZuFqki8anh2mj9vBWiHO
YMyriicQPl+EyH8vF5xut7+hY4PnuU7YwqX2G3BdxXqJuUnzD2GJTnSMlNd9ax0c
xXSiPUqL7tWc9qHV9TtVDK9mN31hcI6El2iGx89pHjFYULtmbBwv4BZK31+M6eSs
PJ7B7Hl0BU9kt9OOtAwhTYmNZYl1viLTqn351PKTPjde/aAYgGCD7Bi9VLphfOSY
0YE049p6bQCvpaKzF8CN6FiWb3m0ai+RzyD4GDu/0+3WrgGMi0sVgMEGxr4XMyoO
DJ0Jrp3IECO8SbSXXZCR9sVUGQ83f20ZyofeALBpvRuWlIvgEcGV59CW3sMEw3Ar
jXBz3RZBVkE74HtONX/H1bi7tf7pbUrP+UmJ06CeeDZ3aCKcK2JuP3Fd7MtIIjsy
LVxc5OhYGVtIO0Ykbv9ljMQkgSFdfrUGmDTvdiwQvw97G9JS2wMHZpAyw3doqF9t
x3yQktrCnOJOxebq8Ltz3y3Eez5BcsVpo+y37IJK2iYpgrdIFVVVqygWII6l4q3T
Q746FHCSdTuNaDskoGC+qB40p6FWSMV2wA4qHsaSroD5TgIM2CLzs32p4A8vtfuW
bwhMKkkuTw9HuudRnaYGwF7xQ9ia/ruLEbhgEILBT5nQmBFIG7GJv9GumdNF2WtW
2ho9SOoKNUdEUMs3QRZF70Z5NjkDY6zk9qNZ0EpotW04xc6+hnYD8X5TlFi3XBmJ
dLxNj0RO3JBh5r4w6bi5zdAdoIe9A4nfCb965biMcoK/M51+3ddnu1mztW03U1t6
zm+63LDGdJ7mRMzODEJmtTJiZjq2hM/8/sU0mM08IDqSPzWvyXAU5UL2fzIxQiNf
iVuSOYW6LpnS8uZm5NccUiLXLu3FCxKwMirmNb6uZb4QtwlPbx2Udn5NxGtOCZWW
ExZ3P8UJddb8AfB6byQt69KHPxm2M6XQqwOFg9YiOdR+RjcIWR9wjpuQxqxgrsqO
SvoXx2vJb91SohuD6kJtFdH2D5/BIJPui0/wk1YS3tidkIy4P4IILHkzDXcV+50B
6ZfHEiRY3UU4Ph3qX0RWq0FZnjBpvVTzmY8t6vg+jk5WrZK8hSb6XOsiiY2VLIsJ
1c3Z0gWdmHKpTqq6ePF+aYQ5MSj7ZNU+AoelC1xsvlfJlQnp2G1XUQoDuBDcJFGQ
+FTOnBTdMaw3lMSBtDTjt5XH8GLVjqKKUgBfriiW/yuiTTL/N/UsGD0t/ZXqPHgx
POPtH+3JSjluVFOKXxVgq00ByYo7x61OsEmfdwq12EWZILLAI+5hKPC2wzKWoElI
iyE5cElfhKZfF9N9Y5kvjXKehgSTWLcYH9oEfaHikfA=
`protect END_PROTECTED
