`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9A/RiQD81ovxbFZIhrbllMVKGQPbcm1e7tC/xe4u3AENw+9HUjdYcfJgCcp3PUkR
+A5owqKQ5JmGGDw8bAd2rKQg71cT2L63sizXrCjv77Hj6sqm7sFUSUnMw5POVDfo
h+ie6mHvvQ0hcRLPdD7TiscOqdtuT4F/JztlyIsCXdr9gw5eodtE5rg+YwIPBEdG
HBgTMOFWJA6aIwXafvuM5+mASVBByinl3nvP166z/29YDFQa1QCm125H/rTMKJae
dpDx/GHtImLCfxFZ96cderxZD3CHHU/jNl3K4LjyBw2WJBHKfHeAjvdiALwcUTYK
7HqL/dCRleOwWRhgjJ9TRk7iTNNJndVBZhMhU20Vblw=
`protect END_PROTECTED
