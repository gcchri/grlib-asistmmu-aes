`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q/2XQ/fpxNoVoLKfc+/BLchWiN54R4SeU1UpJlwuuT3/ev8aOiWsE63yk8S7fesF
b6kZAYJ1qDctfXEI/vy6C5fhxwDjS5H4TNcWZGIlx2lBEdOg77dQ7XBRYQvX6o+M
psi+5eOgil/Wfx6Pfno56f5iqpgKJ8YFm94PfTcexNgZKMpEIozk1pwfhC78iFsl
tOTW8M/0QbJVSn1iAIVnv5cwin8vYO2Nzk0ieRffnoOOvzO5/hvjoyCJTjFYimyS
CyhdWrXTaTwJExivruNICXLEuZakPZuA7o2rSys6jRGcOxYewcjdbWnalbJf2/AK
ss7ZdakpXd06qk4ys9tfZdZ4/kfSl+VpVPc27Van/4logJupKiHZs9RwJBBLsC1X
bd5NiKlweCTuvKzMQCLefHJga1BHA/GsJNsJGSkJ224qXa+W8Akf24KodNjX/5mG
W6iUbg9o5E4mCB2kSCyAx/JQiyJAJJ1T1ebG6H3kEx7kUCcIs1dYkRImwpRjtpw9
J8yb8IHro8DHmHB2mUtQKg==
`protect END_PROTECTED
