`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U6+7xJD4jgZR8o9eK+Yrcls3KAcc7gMO/CfqZYQlELbAuVWfz0BUCFJTSN8V3XWP
hLB5e2GGjAbx7EWD6DwugSwW/Tbv63X01sqj85cyaO+UrqXkPQsK9bLqAgY+aJl9
+8cj8RN6E1JP44UVQwSxNHBIwUVIMJYc6m/hcfQsiCcdUHr602+DCNPGAph3SJmm
iKb3nC4VXZXl+Q/Knz9qnYs4LYqj5MCNZduf6EitkylcHAFZsSDRnz1L1rXcCgai
D+G9+OkgR9X8UJ4GuWdU4IgMRLPsgf1BuiCbEyNVq+lhS/H1IvwzHj29561pQfWl
2JIHFmgGiuQjRovw36EVuWPCsmfc+jecc6ajihc2ppToeo6CxizbFSqnVqfAhN5m
afj2vJJfvlKs8wsQ/3HTV/oaJprWQ0grp7EbOcUC4o4C+h2U1vgKBH+gimSRIXph
q0QUuFTvt8vALStSt/HBwM3yCYS1Z0HxIZNjDhwq/Qewyz65kbkVI7qFwhFHvwXN
mniBV9TOZyfKB2EuvS7HnEfsxsyJVplsEHudgAXi5gs=
`protect END_PROTECTED
