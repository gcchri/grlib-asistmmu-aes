`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
naqMsFay6kZFh0dqKJXAjcY29lXsDI4+23Cqht8i6G5bJ9APHkK4De5q0dTvzlbe
/ZJUwG4fa9pmZCS5/+AyprPtgFY22F/azpdvvR34I+n2ZJwmz0Jq23MXLVWwfg1B
n1qw+a2SIUY6QR6sfTMc73zMeH34F5rg/NZWhxKTEUQ9ZMi2TW05D7NjvrciDjkA
YiZAcK+OhGjfGDPpRJOLuId20cup4xP3of7y2/c3U/oNxnbz7lYpk3sy49aHEu9f
M68GxzgZwbP2hNb7V9YTcdIkODdHbIUaXVKXcCXaF/wcK5wBfLxMWGmnR7AP+Gdy
v52bYp5LHWUfrmynkxG2eH3gDZgDuZ+2mLVwpJG97Gja80NIqy24Han+hEGskDjX
Db8nvkNebkp/r8pQ7EZcVsi4jn3murHqoEYwEprPjfkD/N9SSSfson+kyTW5JlMm
ICvhLqrnSaPJF81N7nquISdEpW92q9FdLZW1wsF4QcNl/Z9bB2uuu9cCfmgwvDlI
op3XTRqSgpLsSHW/JMQzfUqtOJcLvi7nzUhZdOibhUAMq9SkDim0ixbhlHwDSgp3
2I8o9MCS6hPNpBjJYe3uv3xAtq+ap+vwXD/z9ireIkmmOdgW8WsNX0tyqkhVo5lX
iXpDM0l1lDyGekJUWVFo3FZFM2jgo4XDXJQtAyCguxuItPmUUzQAXVM8FBHw50Fb
`protect END_PROTECTED
