`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FISu8v2mK0N4I6qsNzOihjqdpMdz1ixcULFcsPJKDN0Q6QknLUeHjqYKqawb13sZ
LoT2yhHyHhq2nYxSGzHGJgSQBA6HZDT33V+vx+hsFcVdIUn53VRnXS3uEC/9f5am
9riWYySVwvkc9CUAsVmMxzy/DsQ8ns9WoTyjGpSDPImftJV0hO7NsDw+A0z0V2OI
WDvlc0MzVNblE0YnTlI3AT+yptv+3AJAkHdS2R0ONy9tF86fOMZx00lLW2MdZppV
5EJ8Wdq1h8opvNOA3Gm+6EWCKVGRkoJHPuk9mCK6Dt4fUFre5zQvU2W0VVf1gHGa
GX3T6rYiWFqWXaoq3m1Z9qhf6Zd4B3bx66pUcsGwHtjuJcEou6N8eaDA8zxHmu9E
c/5iuT5EMzmTi94onJdPxj9tplIkSoJYTrIWtNTWpzNatOIjVL8jW419fZu5BWTW
vLr9Eyw4lCqLzkVtMke/fO3HQ7pUiMHg+jIM4Cw8DM14c3NxSMd85rYSSMuLail4
DIeYvUYQGte9EVy4FFLJMoTDrAYd7td0j6HT6p7IQbb9RvAd+8S5NPfev5e3LgZV
PHRzU88pMvyzWAXyfuNjEw==
`protect END_PROTECTED
