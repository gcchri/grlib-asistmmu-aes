`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
StHw3xLHGmM840iHhvjEVN+xQs2AWQmxZBVcSHQ0EFgs7lKgnRLKA/E4LU6Ih1ys
UQMiVcmzmcC07gcazv2T68GGBuRSPM81K8p19flUgaqSxDoRgEBs4rBeYp/eJeQT
2R622mFB9U/Mu13Ul2nB3hO+OORCUU5OgNQwRec9e2NylmjJEKhoVYdhxaV8SlF3
HKlf0MzLUdqN6iow1BKzm9bDAHgj6gCIcxlkVRhRSmMUuwhfHQu6WEW2xxMZlCAB
eyz65D7Did2IXlm4Ys/xEog9UX4MaUvXiPZBTZQcPZ5+ZeYhOoR6bkACrzHIOtR0
Ax9PKw4udai94taMrNkuVMe8a4gt3ooxyr0Wm/poy8ufyJVLbqdV2bSIEYBjTx0W
zikjTuX2v2ZGrZhoMdmQJ1B6D9Iudrlqt5CK7xjiPZJBls+WaAZ2R1AFHZ5qz3gV
V16cwJ8luj5hXG/g/paSQDbJtpc/6mIacxN/TnFinBK5Q0MQPLncJ8h48pE/7+aA
9+h8xqD9Of2fCFqOAz4NXeMzcUnB+Wva1wA5gFrcUv4WhJZ/7IJ20aPq72nme7kf
/ACrxb9mD1XEHmuxtCP8QSHNdVVxHQcZxTrymhNOWSzkZTiJ93vghvkaqraeKAJE
5SJwOB7+ROsG/U/4dcFWnILiFPrw5/Na6ahV6YDUOaWC1ZCWyrsNl2q9q+gs19OA
MDLS3zUPhwG1HSUGKTJjkMdAzsN60RMXDJOOkYANTK485qV7Bcb7dXa1Rqx3wrBi
48uHT4ozwMU6bWXL5AwYPCgHnAVt5fq3vOUYfhY+29mYnKVrC/8mBSPr2Fa14Dl3
yDFSAN3fZ9QZ0z4KuPZIMCyBts+xsopj6Rr6oA2yPMLc5dt5lkAGqWLe+vppEtCk
co+JhE0YIs5zNjOyIJWhk5RecfdGUtUEpEN5ThkdmuTkBqep4/9fGRcuF6ibfDoG
BVlRfq2tMjX2bt/4MlnlzgZf2+KTwG2RUEiWF/pM4SLJ81rmTDmljKJaUNjjw7Ye
GNLN6USg15SbQ1zWZ3kbvwkxAyw0kBeR+HBdSE5FNWhjJuYwHRbXsG8ExSvlPcOo
nEAPp54GOQZb8leGlA5OZ8GEeSvB8HLbEWxBcFB+CkjJwNMyhyCpUv0SpkIybYDG
1g7wTEXWAZEgWGw7A+E2LAe43mwCMfVGvDubpQX0QjLXpGnLWMUei6klt7IXPTZE
i07D6gavy7d5wD5BowBlJhJzlZ0QJk+je0exnyEY5o6munvl8FNTeP9adyE6xD2U
I8iVgpp32LzoIjOq3MYgVwkoGr4TdZ1DTK68Jw2l9DOv1M3anYEw+YOphxM8yUve
DaqVm/lpm1S1BGKqJz1U+gxp50wKlOrjFK7ucRqPESTLbxFn6r8SDTI8Fg3OskxL
VDKmkNtRymPOBXYNwUtSwdlE5XHunN5gFq3EFR7hRoVfwZdxsapySLQ7XBbvzWAS
kiZuDkA1+vRsPe3pdtQ6bYzy1PjminJ9BRQcMIRvnsSlcls8IG6YwfFCMRZpSCZr
km0/BXLHwsYRgceQLK8Tbs0QFwIc1ooP9GVBTsOziCU+4nZgWPuVZS4nFLZmXGA1
JfpPCrkzhtvHwAnrc6PeeblAkVach9HdJw8Z2ejYtlcGjD/sg8isx/PLUvrMh4x0
wOx+vHvwAnW5/CPUTD26yk974Vnjerrxp5ulRi97BRdoADWiE57DURqZj4+0dU1R
QqWSV5GlW9nn0HXzngfAvzzAo2A0cneQdRXl8q/99lKI6Z2i7JMM74BHWPWPDWwd
JZNCjt9QN7OSU/zrQj3XGJBCzUh1LffiC3b/xFfL9XsFdKshVOdWyTaLdQDa0Hb8
IIuDvEhuY5ooJjvypiPy5b30O8xM4+lni389e/fPYTdp/ua5Can9Vwk4JFrtqGyN
6o/DY2JGGR9D4VlxuRsvJCxIH3vUoTzlSKj2Cvhksvyw6UdtRw1vEMboU1Yc371l
/ds6IjNuZqsEYDjsxl1f1y4AyPsZ/NeD8tX2NLtq4EISVsWNGZb08V8/YHbRCGpC
VE2qZ5LljNM/luwY2JderSIeOVw1UEq7T9PVZhsZ4lqJj1F2Ni8Ba7VuCjZ9iY2m
sadipbiySC7lcqxITq9BmfXi/2ub1ahbiVySaHh+Rmuzs6hsFeywKQ9IojnRa1ZH
51a/7PmmsA5jX6cEAwKwOUKMTXZGvkio6veSrHMg6TfPvaYBjXxcyt2abvImARsG
LRemoTZTwPaZGCT4/GfX7OIFGHx4zrQS+PBkp12eFXcsafp0jv/gQgm3Be0wPHyW
GnCu3Rywa/B6JGwpj1b1TnG/f1AY9BlYMw+smcIE2e84PnT+bzNBxPiQpuKCXb43
HdKprNp9WDPhlWVRlXPTLagF0sUiVhNoU2/VZnS/8LNCbcetDXHU2dsolX3pQpca
tkAQ8AaYsS+FFEG0q+oZJSQ9ahz6fQblv6tJ78/kAGPZmbgqNmxril2j1vxKgqGj
1p67csnALyk40ylVzqTxlX56sc3DBUq9EKIBqG9j4qO79/26DXneTHSAzreRZlHF
XuwcQ7xhKtYJ6fPJvwv7p0zPeiODa0E+BUxiNGIQoN3iMOgBjwVkIOOr25TyOuvz
YfiuG2kElI9O77sUXRixwBu06tQQjrA1Chjqra5Lxvf4Ikq6sdUtt4l9rEQ9GfLR
NWEizFOaFE6T/KT4NskLeJaJAugTUIDze8xLk3Bd1Fq4y5++GTbfeRd1AtEZZ1Ts
0GE9rDQ0236DgDE7RpYFdtuvFBCKMZ25BL3oZuHMedl7ovYQJG/RnOPqTYUSUiQ9
rw+bIKp/POn25Tg0nclZMsfpYBlN7mNSjPw57kAAFwbYDOVMzkMsSSgK6aKSzMR+
8SW140d7CfOdtUbIK19+dMpdGasm72Iyf3SKycUcBU1rSyMYsYJYxEknPuUALM+J
vN5J0OHsZFzMkHtTcFdOfK0ek72nqIf4Au+APcv04y5G+MjROe3lIX30UCDM8rCJ
mCc6GskB1EDbv02Kcr053OgHsgrutzIHefMGuGNJCt/Z2kqxadSsK6MswIAJMW81
6PlgrloTycNgGA7/nU4JNKLwSTBwhO5Q8qqHFyJHrCPlsh4G8Ni5aktqQG6b6fzc
hxPtSgCzDFNiMLCyBmW5Br+EzyibpomKmNKO0nW63IU1KhnZmTZQlReIa+O9Phwz
J34Asw7K5SpVPWgeCF6gmxETIxOJTgThp6vfOdPxslNuECLFzptJkax2yKu06wyx
m6NCm8kSVJUM0YmHxlo8kU+BwFxBFwffXqPweb2ucHAyCIeDJluZAiiO4/IMlQlL
dzIp+HElnncLFVS5fB93EuUVNxl7RZf8cLLzkNnmtS3Erd42pMw1seC3sAINQddi
8HwqqvJ0CK/W6v7fjVMszYxkp1uBZzY8QB3O4SYpZ+sqvMtMXZN3BCniUAwdwkbd
iMqo/n1H2ijmzQgHod5HACFXt2bUlb9OiCjsFAhz1dIBzTHO4eSVzkplNlT1/oyf
qKD+Js4ZrkUOD6dAQ1MwiXLzRWkcay4PY0yWDHcwdj3aRYgannl+Mdi9ZfwI/EtH
cjWW8wpJ5ZeeeM3rStJFFhuXvxamsJdrRCGFylJ8AyreKa1uUrWGLn7NZioNwvhb
mvQblURucnpg+IhWtL6V+3sfrdhph2GUfzkh4Y0aC3U51vfBI/bjNHEYLd6x8avN
6ZMh8cxQQi/AEn0IHftpv+a/woEZvXrJ+e5JpzBBLFqVDyPRobF4ZIjxDX55CT3u
egjKU5aUhvjcAdNfmkzRU5yt1iWGUMupH3c+mfRJpt/6OWWuDLrYPiMPV81oio0b
Bi7JtNfSPlj7G2v3dtN+QXNkwzSTj6WOBCkg6hkHnlQwniDI42Jh3GHfsfXwsRmF
JjxiqwyXnvuyPSa4ntl+OKFWvDXhHkI6CApZs/uZaDFgpibkjF2KiE/VY57Lf4nd
vy+bZl8yUFkwK1uSvjoplakRVGtQKl+YeHuqEmAbNlQMIzV5Y3JSE267wqhzxna6
JUFWZbyk7sTeEjdtW1nFwTHeALPmhcdqBM85/XgS/lW8/uNO0xJTV02z3o5xkdcz
ZVHbIV2yqtxrhmLKiV5WBGeysvH9a7dGkYRjyH2Q2t56rMpb1x4Xf9tCXyYu+fMw
jDKGAxgHonZE7U6pnSDEMOx/Ctn2pxnp0rfLlJiO3yhL7FTkCih5DhW7Nz3tO1oC
Mjpbpxq42gD6CSLahYoOGGAWWsLtvPDNsDZmZYyp7/uUi7848TaGhBoZoiZ9B8N6
AxEJeNXo6cvVxMUVJ1Q6a114VeDsR2okLjTdEkA8brXhANORIwKVJ87sXhVSUTMa
GacXfvKMMUq3iU3VB1rcXib7QXT32cak4J0uv0OvhmARKdRJ0y4BiN3sGWaW1p4T
D8ZNsC0Gi9IuG1tL9ran6T9ocHoF4AiSNsf+DpPBIF7jYAiEBx0/2IAc3+2LCNbM
nojcvbUDa7NU+EDLYvejM8hQSFdf66o2ppy12zeSo6F4xhsTvVpu8byiTvgYKGxy
CB4TYi8meGYlou1D4uiaA6hZoFrW7L1MrMNPuH//GGzOY2C2tv1IRTaQWt2q7sco
rSjYgah17MVamsvnhzYOFjSK4oOzSiv4kL8FPUeLAinE3Tuqo6ewpqv9IhIFCf5D
GxcKdbV2nho4WGcLUesHvlDN7+HPHIGAtaEBxeop7XegglV/Oe7vm9j9Yp2gW7C9
UXJSQbMMXJGgOMxihEXZxNAVG0oNQ4+6MIo1GdEcRgR0M2bxl+4g5RjW1EIZtj5U
N+7ZFFWQISO2MXRUSn8BsRi3lW0dUmGFZ5fdQ7/HHfZn/pRGriH9HU/TNOivwe/0
ep1P4u4mOcH/9ICqf8F7YcFylV4t0gobH0wHxYJOPxsuMJ2I08BGd39WHa4n9K5M
g2XIqFWu13GNIYFnq2q160nRMXNnaYpDDA5nd87MQB0r15YeHtg/JhOp6akPntHf
26pJ+89SkvD4CstG2RLC0a/PvEFBpnP1KGfbObhYf0r47bp2/GDogplyJ//z8oIj
gZMPumYSdHnVgxfVlLhRIdyyNpp+UPhEGGMNJlUV45F3IL6NL1P+miF5+ssEYQQT
I5JwjF+vIEoQGGmbfbwD1WHlAHWWcrpAbkBmmiSnSv0vJOu0jQYqSrvNSUmD+bX8
m7H7Hk2ji9AvantDyi4cf8pdVnSNEFif1TI/uuluB2DP5y2kr7CsKUPAPwG9pW/X
ex9hODQeOm29fHCa7WaEV2lR5eKFRqHS67KS5ngPb7DlWgatoqDEoMxxPs2/zVjT
Ee3evJFgPKxv7AjHVdDTjXs+flQ5teBPptxvLulReyPLrOkWas82pEiXxbJV/ffB
iV5Tjc1woQVcBOdqUrKnEJCYBsTsTyBmoEE43fiBVQeVXw1Hr6jHIl5/uK9R4Gvj
SiiFWboBTXbJAD6GNIpJ58RnEdmMKkrSsPr50B94UWBpupFLZrU7M7StsV29FV99
DmUaL74zojIzNsFmOIo78g7iBF5hq5gw8HVJOlFgrYT3uxbZauXUtoDBQY/kgXSq
gn47X/LGT526TAKOZL+4v4DFnvNAN2Ee/KWskFA03SilpoJ6TXIuAzyGefWIxRy+
G3/M4btH+N7LYY31b9MCRnIXrFxPr9dM5Ag7D1gGnzNHzdyak9yw1kTSerFZL4zQ
7t8dYe7I+k9uf4kllQoH2ht89p/snu/R2rU+NWTXFDP2FkEc9dYG13Ot7ChIAXUZ
+dujyNXA7BxGDsuIzFsqNAtorM04cr9OBXmRaUm20D+cuEaSpFyjwQz31j/dJtIz
OFQtJvYS44jvsosD4JK/8COo1MG/VchDK1/0U3jXbFx0qFWEhqTM1I1FKoyLZ171
eeGgP02Nz23JrQmsv6mP1A6WeVGbqjF0bKjJ1BrCvJ+oL1oBV71nunQZfYgLHt+s
0o+epDcAFbPFhVcsVRWCj0O0c5OV+NLp3AoZ5X/jlo45Gi0R4CdOAn/1I0e7IrvB
tdfXFX1S5hiEK4uL1KLjtgH7gmqQLBtzQM5R1W0tuU1Ei8+qEUkCxGqBSHaZhhoe
mhJqaFy2HyZhSepWYCKsnli/XbamTi8C0Q2La43UIv6T26fkzU01uItKaa8ZpOxr
dcv3VrCR+h9SaOZI9sf4fgQ1Cd+qHx5DqerxYFSolVDNE4jOpFQ/Igd/pr5jR1+4
3aFtXtMDEsQQ6L4QIRyIjX4q5EPFMVSSWMvSGPq/okB1MMgs7vFgiRtG8LHf16RD
rePB0bfaOu4gciruFJWvVEIBWEVtzu1Ybw305WdymAg1CEF9sDqNptnezww+TYgX
Mo+/D4WjVtQpVtzVX/TSewVqEtrSjfGDs11GAldeVFbO2FB3ottseISWp9MhPFG0
MxY+KAGrTqPNzV7Fn0tWZUupFCX45Y0BgOQIbQMgXuXqpQKNYMIeBUqdeQNqMcYB
idiQdJ8ehBPiiGR69tUUQhB3Tf7406nOIhIOOQIgm4w+hMN1zfTLDbywd1XKExcc
ObYH38OhYdHRu/02XZqkHJX+OUgHWPV4ItWGRXTIOYBuX9zSQ0gXkpZLWfHVMAqY
7tvHhzx/eaPO59iC074QOK4mXSnHZ7c33XN6Bibpmm+go5wc9KwjMnjOZSNvdP6k
z2AssgbhuCFAGVILFRcwtq+KJ8oPomG+aRojiA69K5xN+1uMj+PwOwohopfUKSpm
0saIc5I5yM6cqfApsy/PmzgXpnS7iUABGpcJ86u6FN1NAFi989OAbLZWrx6wkIq3
hw5dQDGEfJiwJvh5kbov6zPNWi8pfiWfl2YCxPX1Uj/iySSI1ACdE1sAVkJHOZ18
OBAm4glN2oM8alMbpUNugSVYgWrnrHz18Y7DBulKJGw57KxsyiWGUlQcKvtYQLuV
Y9VGJ9U42aDzhuRQatqM6Q4cqtFRH7eLyibgSKYdF61mJXafXUV35Z/uFm1Zn6B+
OxqKU74z403BE+cl2yej4fVPL9IVddP0bypORiNhjeed/PYp3zrdwp+wMVNEvScv
JjFV0ytMikvW/f0UJEmOJtk7XpKq3ZdT32kpGAzCTrXqE2/CdXY8c3HXn1FpYG8l
WJcr663NSWPbdNrChfZWvtQbJRI6hJTW7CTjGinlOcOuRxa2TJUapg+MbYd3YDEW
Yh1YR2QAzAJd+dc9FDLJI25RSdUC2PQKekWDX5xQ80us3GVgZzAP/bEeV7OnDNig
v7aBc+gWIvdWO0e+PNsV99K9KDRA8LvTfMgYKmT6ay8rH9gmUnPL0TWQ1kXAlY/S
/NafzxDn2EpDDO9E32vrMAq/T7Cwvh8b9coVhesfdtsxnWj+vfU7zAs5KX9LtKMD
ji+D3RfrcVOk4YCqbhwdS0bpTIl6huek5yif4TilYezVGAG8LKSB2xVMYy2ktm2G
fXlCC+xkAqPsqBHbi08rXttpT/zMrDAabPuLztW+eI/BS6QxYaC2CTIjzGzyDZkw
ELPnrVzpf8EYHribZH7gAfIIw5xlo6u5d0YhhieIMLQK26j9hdmuYV9NlEqV1eQv
LNCEKP6PEV8/VIHfudk6DF4NqVd1PClXQbMsvPfajQG44A2AAqai64KVAJ8E2cvy
UPmfM1lLtdjHc4Fh52EbxcQ5IVzglWPkqjo+yImrSYzB+QeD0YkskZPB7UxzkbWH
sri/vMOuI22mLeC0+vcY6RQATGSs1RykwaMllhy+wSad8Npuhon6GvLl5fytKDQr
CHTqh99HR0udPTg4TpfVV/P7ZEuQY5B0SVxLxSKE6QMCJvbRukMAw5kONdcroZ6s
SyY9XL1F/7gMVQLn14TeD+kCj7DQ2K/uvlTT02qxyN+kSaNpepqFO30kNaghgMqJ
CJTtlEyobcmxlBRcuOvstRBkHWlLEv39SOKAqeZV+ieKaEHCDqwanfhzjOT2o3CL
Neam2Qx2UWaTJXKe7KxfHtDfa55iwben9xR7J/8XxQ5eLOaQOdXftdGNYHZosxOI
2scGLKAYOsSWji+cFhITLtQUKsNcMfi7enN/XwPGcuh2FKaHCDD6ujBUZN8OW+Oo
3P0QIbwIo00+2T1VP9ksZW4Z691/nARd8u/f1WcZP20hAyP0FJKYQtYafBM6oXxy
MHWyUGiqI4QxDya0DOG43W6y0FewIvDQRLYJxDT5ZcL33sz1uAnka6U97zqgMvhT
j1Y+luOoitWm1eIjcfBTFI+e62dMfWSE20O/YjP8c8nQRo0fcNxx2Jyd1i3JSB08
rEECpuYBcX/54tbFrA0I7q5ihHTUWy2UEvTh1uRrg6lrGi/9HwQz67f3/02ohjYD
cTzdipu/7KhKun9p+2NI4FdEZIGMc8PeT7Nw9+1TE1GyMOfp7HA0BBUsDjEJ7tOe
qmDQggTyMtdB32WZCrPI7rFrR0oDLCClQFIO4JTv5hsjVTiGdkfcKt4f1TKtDq5r
t6ivaPRZ9+eVnblYSaGyU33Hj+IynU2aU4Dt/6BHpRqwauMX/hYtS9ZvvyPgDOgC
xmzE7tKOart4FV/iu1Jii+ziACh/fZYlbAem49YMVTkaXtLbQ11MbFJtR/BlVQIp
Ya7SVnykdbt0vA86CHfpIs3cX2dYTQXxOyh8rm858FEz4awEWxUkwq69VNlwTg6s
rbB00NC8WWLNN7GwGjt8bi7o09x+rjnn+vTz0K0FzWu9h6cUPO0XcizmJ8etUtaw
M51Z+xuSZL0VFHKaMZBdcC3t05DSLLQIM6TJJSF8vPecXsgmetnyYpsNbTYmEURn
If43p8lKgkQ9fswq0aM4+8WygDsnPKJ9nTJ7tVK4PvmwYy/zrXkuYJV0OGcGgjBJ
8/d4lrmxfC+gnqUCn4+1FFWRquFlMjvsuYA157C+s93q1AvUmG6f6GJrx9Ytjd+G
1aZtUnmaV6dAGBrsjgHAqQO7fL0nBqvrdwTWAKwNoJpe0meHKFhF4jNKA4dKjsji
On3jyWTMmKOY+tZgCaiOQBksVXric/R8xbHNmZEgpwr3QF2098vgpFi7j+pzkc/Y
DXW5aAAvvEDY9fuTZ3znnZDA26DiWScFOitfl/cV85oA7BNZ1ldhazpJFK8/Aa56
3FPiR/QG+41QnXEL7jKE8SA0Uo7VE2DeguZtMnQo/rxe/wWBWbF/mF7kxbp4u/mn
vwLnpicnGlfKGPw/1/tQWKN3SV8tAPd1X7R9YALUg+Lg+yVUFBnImS53S/VJouBV
YXG0iHXsar/bMri8Esuk5Z4mb70pCi4Jyz3NHHAI1dJDW14duhsIfLn+lPmcTLP+
/B0wFbG0jmmJKvMDKZCCHpXPnmu/OS8qh70vuSbw9Z3/15GY+UNmPDeWzA04t3NP
7Ep+Ybs2oGfxdmHKbboTp5iG6i2XO4ON3Lh97l+8fbvZEAhoKDvy0eEvvhyO6eMt
WolIIy67sG7pypfPZiHYGyYb5pMH9Ymx/gOg/CXePlnmmpqEbrdba06ZmaWeZBZx
TKBZgLpLgP3t/4Z8Q349s+LZ5g+Q7+udLL0VcFA3xjUvKw+Lh8Lujx20GpXJA6SC
PmZh3Fd3Q/yED/wyRdb3XXn9TV5ahNyv1h9nTbJPrRsaFQVYhC8FirM8g2lvim+1
Vg5KbLcD6SdZS1lAFBoJlD5f7CqTQTtpsbpHa7q1Mt9EjODojtQzzaJa2MKlmS79
gU5Y4pveF6N9jnxeECmDhY5IuldsaQMlJuIzSW1jQByyVLIhjXUDna3bADR0GAXP
TpAaYBYLPMi85rDkssrdQSLyhFrEGEe2R77xRsj+axB/Fgk9e89tvX5mgENdJ/oz
RxMpKN8jhSeYZu3Ead3wKI7/z/3pOi0i3tAhpmrzAyHCbsSXWK1j3MQcEpKx+GnT
cr2FjgFonYqKKiltdPVj3COETl/LGYmp1wRbtI44Do9KrOTgPN8y0E1E8IZwmeeN
Ju2AptqZ9PWT6AVw4/j7+MCb9CBK6hOv4wKBTg8t2a9IGgrP5Pvuj+eFyifP5afN
JAXmjDRG7R3p99RBfDTFXDJQ3mGOwsWOJaN+/n551nEcxF7yKm9fxqgtGbPKqlL0
3+x5L3r0OLF/51TButUPh+BmelByD/C4mlxIHCcw2tmSgBeFjnPNlYKb1E1Lu050
aUreWBznMFcsdoU02WLF6KRBOnRkwHUxIW5RNUXfm/LNfz/e09yoBJXcGCO4k7/8
d3WbQEaYwJNPL/zMlnEeQdreSoRCCtUgdFrS3ibyojMNV2f0SFYqx1x9/CqL0X10
vfhn9UbyEp1C8q4mINCZHnlv756lhveghRb0E2WaEzz2CPKLXTpPcwS2hAxjV0eb
LKQs4mFPYdc86wSg8Nq80la+ElZoncxwu7MUsQZw8OtlZ89ClcLp9CH/H1yyqNq+
4BdavGMPNCiZbmvqYsYPPv9MrFMqZ3IojMh2bzx6Yj50MGnxCo6AiVLAIzUP/YdQ
mveMWT3Wfg735EYB2O0Nxzm6giAw2wPVB62JEyF2v0FyEN/VUKaEGOVIdSLl4dyt
ItIoRLPEd2F/nyyCUAjJXS6WZr8m0dGDAAOZZVUQgbl6IKrfW2DLSYb6N5kWjxKR
D9zTTILkgmONjft4Isa6sOh9+YXdGU9kCYLuQbo4it57nTVAVenxChps4cDvWwVu
eKAZhnvgP+/ddCOR0YyauaWkk3CVlYC3z/J8Zp3pMIYEVe2JRDcH/dT5zQp/H9Py
XlFX7jCMQWKdz9kZkIkxDQZgKT+vUDQXKkrSsaQPleEicvRyl7jDB/leFmTq4XMK
IVjP1xLYRm0EgHW1zAAhr/fLt4jYiBxdoXMThsa/jgtMjjDVqvXxKU9OdRr9yR4M
w7TmTvk18cJA8wEIJRJ+ly4L8jCXUAckh8v+VcnxqJmZACs0t1D+cXP2kAyhHCng
dT3bqwg/GSBjtvOOz9J8gC0XQDxb1s/IQn9A/hy8bGEXbreSDelT48snlo4h1X1o
HrOGFUCfXfqVDid7S0cYtgcGfXeIJm09i0Zrdfu1SFDaG+Otux/ZsCfkvJ++9hfr
56qDy3GlWpTJI0N6lh1V/n2nJq0+kIMFo/C91MEyb7Wi0tLgaRGixjSrRFylyBVY
kuOjdd5MwlJdExXB3BHWAOpj0TUlvPAlxIcmU4CJpw8RcCVOLziChPRYQ7DpzGJX
4tIC2jawxpkCiOTSuxqIGHlGfTT15GHsaXEy6aFliuOVGKQquassJBcDqrpXJ8YA
9ltlC6z10+danU4tNyLXtnRjqatYMLeoR+eFMZliRR7Ao+01/xnH6ctteYxu1n8I
kGeOANVoPpDbELDwTsHYVOGiwGEX+NbQNrUZ0jR8tGfDgDbEy0dIITF6Dej1Yops
jNul2RU1zpM1kGDNEMvcV9IQuv1ACmjc1lIu11o1KlE3XoqQYqYywD4nIUp8VPo8
+4938SltjwmM7mEtuZIyBkW/sk85QyUmVMJ32tAdiRhokPwhlNqao59/+EQteQW2
fdBFu2Y1ZdcH6cuIoZ7tpILh89JzLKrqieUnfqDaS/uf2/meTpib1rflPge2kqSU
lP6E5ndCwCs4oUwmfVTje7BZHtaNWBV+Wjn1iyOHvKqkmMR4mb6zF4Jp9ITsPHfj
w4VDk5rgI1ER/1rqrqoVIBltPEqAVTCE6upfzlfCwtyLGtDkwvTUGbzz4jbZ/DnX
eRzyS1YD97QzoS85iAGh6E8ZD6GTAjMj/vO6Fe+3NzLzFTi6Ll7FxsgAQ5gtUsWl
eBWyYcq3KDbRUX5iAYz+OBmqSsFnx5PjdInDbArQyCb/Ypwl3MqgzJYeknc205au
JEXrC4cu3NklpyGLPqhj/SAfdKOMzOqWzfVq4u7xMtXn/BLGH3A5oOPzUquBFBEl
gMZdv0oB8OAuq8QAklkc+JVd45D2To8NJKJbVOpoqMHnLewY19dDAMYwrGONp01X
e8P1G7bRS3VRDQAnHX1vmoTcSHD3bMW0vu9GP3Gagg0VNVhiceGJCGgfc1Zc7BF9
4ayS+YKu2qeJNhmL9IGQmAupRZjK2spP/JiCF5JlwCbLtPq00HNoUP/M09sZ4Tu/
la5iDvbEAzGM7LsSqP4T45IGyF/gKgRpS8J2LcRVnjxVr4AtNyu1rM4z9aiA8TxC
KeycGRS/JrEt4Fp6uDakXcHrcEh8TvDfIybbkZINgEDGRXq40LNJG3KuxoPwTJlC
Wvn94mYd+3bBRQByjb7bbpTlqD0WNliIVg1j/cZRa+GZO7/tULN3GpK4wLAGDpno
flRlH0w/1+7PWA0VF/Pm0kClT87aTZa/zad0NNu9qkehc8aA3zPCOqBm1IRsqvyD
`protect END_PROTECTED
