`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zYgF/y4229czhTXoMs/cPSiXQ7UJpHYRyYi+PTTENjilhEFCtcG3oQnb8yFgbis3
LTZYt844yiygEL1rFQierlJ9YAhLzGB6xl/N8ao4PAGRY9wqXIf+UnssBgSp9Yku
6IN0gtqgCOZSt3/btZojvVWBG9yY/XRQFCmZ4iDRp3AYR/x6jIG0lu1Yqj8mGP9N
SS96iPv+t5MoMKstBr1AkRKYTo1f+KhicNd+U+/oTwg9WrJcmdEwWEx98RohMJ6l
dwjvUxmarjtHD6V00niT5+KxnCAPI/PhQL+gfg+0uHGR41WCowygwVaDMfHAWW/w
sao8pAOF313ygWgkMlBHU3V3fDL/5OyEzJd3+dOGTxSV+g55DDZsG7+hAIRXsyfA
dqNeK62ZILgVMPuNtX1JTV68ZoPClTRFZCsLDMB5NVswyvW1nECXe29vs2F9GBrO
v6wCvAMHvqTVcjuWR6m4zfBUOrqgUVn/DqGFhHWMQZccyIYVntPj/HTuLFoCC19J
nathChyGWRlSiXLWVU3mwUEGs2RWurYWiVA08w2dkmZ16pA0Y9bz2Xwh4XcL9iTB
sssDJszXg/BGsBt9+/1rRKk3gflBqYYGPf68vXg3777NQMhsAx1SRe2rpzDidcst
rDbASrboHhBTdwM4Y50aVL10LmzTFUiHBGC5yrKwYEQEIiMp4LUcntlIQb93N4NE
TVl9y1AkYzsvQwpoYzOPZhcmGw8dzLthV7+/hhxz+b0=
`protect END_PROTECTED
