`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kxZhoQHSrJ7VxbE3Cei4cX/QArKpPyc1QvYEVrF9DgCjPPSHQcQT893jwypkpQTp
OHShq1tEp+NBrO7MdY2JlogSIa44Nzh5gyJ0ZbEokZRN23BGBD97g5gKyGUpLcHH
uBUqkoILzX63Lijxq4EkXOWeLIlN4E52ClLuNt0xOirFCyce1g7qXpd2UJIr7Nj1
9KlftR/hplCjqsRvauo2YPLXR/ky8ipvzLllIYuWZmZ/Nlbi/8BZAaorymPwrep5
plDd7Yywn/R4a5ozr2pezP6HG4LYuZ3E4YHf/NeAIzcRlL0zuCArD9K83ZsOrQxU
UYh9woaPiTXp+aSkUandO04AHVWlGvct/hhhdJoyqwyRmHSWycfOI5EkYRLsf9AE
Uf1CtHEfu7ouQpdPUgFVj+4b68KgDC6zqhX1qtQ//z+J4wBsx0PfYHVHWkNzZRMb
SJMav6+okHreSNBp4RTP4aNfqDqFp5zHWbRZYNvrertMyejAY8uMvKsTam8YFQzt
VNzIWRAH+9i837Inc1gslisI3ZggdByrdoYbUscXiIThx7rsLz1yHhJao7T2aFi8
A2LCIEwRtnUCpZXj8TEaFm1YRQGI3x7h29GaoAW6giRfTGt+T3qekeRdKKicORRa
iIXQ3Hjx7nQzgQbJnt0UFp3Og/GH77idvApS4c/EKeqmi9248Hk19LrPUznkitig
x0g9dpZSF6ovclDPU+P6apLwXa+AOGYuOKtIbHhascmrJXeIEq6YzUKFt9OBvpyJ
H2g7QQDBgGmz8FdP1UWVQoZwqF+ADncFGt6+up7trjd3K5O2gdX7j5pFeBE406Qe
1qWZf9DEmUAHDjKJplDwvFvxI3EXRp93XSmvcy7sA2KBh1oawN4lnZ73dTsTfLtf
NsMf/JWzV/ZKmVmaJh5d8Ua4aJ7ujJ7lb34FpSB+NJ2GoXURWUdJzvLpEhLofira
1gwsln/EjyHbsLIB4+rgtdVtcjYgHGYPdJ6A/2XqTgMKKqjizCCLjZZJybN5ouTr
dl0P2cGUaCOlaZBF1veiUDJ1DpqqL3jXXlm8hu9ZR9Q94zWzYVxl85ys3vcCaBaT
XV4B2kXNPmIMkKt450hIaH1MvchHtH+9KJFXkjdsuwuxjSdlhVy1o4j52tD8O1vA
EvjdC9d/5eF8luWom+EkczQ44d7YDjVp+S7wnke5HBtT67TXegcVbZdPWqxxPfgp
y4Rf7chSlGi/9gCvlLOuNEnBSpwP4R+7OQ+LfsVPr3rERluoEPw49oVpJvpCI7hM
IGSX0VcT1rWs5gl6HezzPPLzaNxeGcwEyI5onMivBwXMM7hMANH3q8wZREKcvCEG
OG0XNxVIMfP6rMm6T95MH/NZ4ql48F9d+yfTOWHqNIXdEWYMH0RoYcpXWa1i5mJC
3LpvxHk4U82IbGOBmcBB6MrBYrfE5l5ZEArxpjC9xkPlbxAfnWEBYl0Rce1SKiwu
WH6CF4CW6ZN65NF9+ysxx2dNWPDmWye4sL49iK1TlgAXSM6+CJV8LsMz/bvAGQk4
XzJ6wH1Sb/N6/P871ANKHVjN+JZUlmI2E/xwKsfyW9h7C+A6ub591WOyEJkJofdr
3vgV69QrXTaQF17ws2DqBRqG6ynv6AOVUcpr3ZQam5oeRhNqMqZrsKMRS3x+unUG
/3Eqy7z6rFtUKKSMVXysyfUgz3QuUCnzB0ul+KhnJCRvUbVTVAB4lW2lkyvMm1uB
1NJV0mTksT/jUsOFfG8GT7cA9nnRI82od8/AzuJjNh5VZYB2ORbPvU7/yDWbSAVJ
5Q8UXMsFUsyaQJSWHM6bJPG43BFdzlo/sCUStan6pJBCk55+kJppPfPx7+udQmq5
gb3ebM+5LqrziUmLrCDC85NuyQ6FiRRalLMoevXWAXDU8AkppYexd4wV9Y1o+YIi
coagPtlONOcVvi95lFQq0w==
`protect END_PROTECTED
