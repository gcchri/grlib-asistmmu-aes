`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dGnyndtS7S+sWRy5pdDVJEyMbAdOH84aooiI8lEAfC9mbnKdraqjXlQjxR95goJD
U8u0GA5+STxQke2KV0drKhZRsBseR5f8T+zaHomecA2b+Ji3G1mor2PoGnN8GMQn
v4iH1Uj1wUHKQ0P+o9EJcsVknSEYZswk6gKxmbY+5S/7KPTd+gVg5GzXY1g4Dxzl
R8fim0AXOVLlpAJ4LdJhlw/ky/+jqCmwidghVW2ypfkg5vLZ1VUrnBsXrdtB90u9
Y1DcK1DkZiajuWJD2RhZdxA9PU/WIj2rJF1CnO9bR+YMhviLtTwjLcvuktWw3RAV
GqaFcMH83+RE08LDfC55kcAhKASDahd9CVv9JUOdClMPQNNDNsbHs5cRHfXX/ttI
pH4yau295SUOGoK1ugWgUNHw08+sxJ0N+xpPxgA3gf6csTxBWlJzoAPA346n6fvH
td/2Ow+LkKhKRLX+zK4gJjV3K12tEBPI1Fe/h1Mar10Rr0xk/GjQqAv/4bF11xD4
8WL5R+Sbr4eaHPoklvQ75FpiMCGyxOYVgW75hEjvkTNtD2feZO0B8aGa4hRahn44
nwjesNBfD82CCaWrHluGVN+wwB1l4XH2UrQyKIqyPiODz/kAAVQxONC9VMlSv/6e
IT5XFSiNZkx25tI2T4CNeOsEE3NxXi66UsiRhH6u76/2JpCO1h7sC5og/60JBM41
Glc6gkWPE0ZR9oNEx8kEJcfK5qroFWgbkWAKPLauXUhDbDcY8G1iqaO3MQ4Vm0w/
MZKK6u1lpqg/gn5SgbouswMuRfXnY1Gd7CzmmdxN3slcXgOSE++NQTH7kHD0CKB2
Fo3bfxXUhXlrJBrO1ND4uzsnIn/gmuBfGEWnsso7VFs=
`protect END_PROTECTED
