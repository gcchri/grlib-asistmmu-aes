`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gi5LNOIhHKKVINIWetUYZFEYrZCWhLQfhq1PWgXDifrb4HdpnWkYZTZ6TfuMhPA+
z4fWkkV4iYDpzuntQ2aa2dPGXO+zPWl8ST7zShr5IFnFv0+Ua1isFZaGRjMXXOMp
wSVwwncyc13cy7+nMvW2iKrV8z3Xi8coX+4EQLI06QPr6OHSpRZ+5j3PFJBhHxoZ
V7SzAABh2aKLw1Grwg9MPjoxy37FPzO9EsnvS7CLGkRJjbCZtZ6TN0j8oXRZuWyz
4IsNJGqaLThIA8+tB0cDuTvsTkp3BVEJjnn62aTiu81xOAGpz/LvKZZfelsRymhA
WpqdcP4mmN9gDik04sOZgg==
`protect END_PROTECTED
