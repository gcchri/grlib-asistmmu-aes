`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L1bYayt3dRAIN8Gsycjfvdo133+2ZvyO1yJWu8SENoGlVbr6RhAoLYOINFo9W4d4
e0XJFrcnC8qiEghtBaoDBCyUC8caRVN/JnWJN23mrt11rW03BosbWoX23PWgNFKl
lxjoWYDuwmfWkt40nXZP+Zlfz3gm25/FDTv3fzoJjVYPW33w3fRCEktNZfNli1tR
HV95WsT1zMwHHuThvfa1ZqHlxV+yUwBagqeCr35h/VU/a48q8bPuBhj2IumEkGju
Yz6nk1inigjzkwTxsWvFQz80oiEeBQIE0XzXiPs8y0jJfzIaLkD+ubeCGqf2sJVy
/zn/yT5N17I/DHpeLRpw1uGfvFQixMCdfUyWRnhtV9617TsWFds9V9o7x9yju9kO
SXz3DDdgUzo6jjxPGi248DlgNHZ3/yl0f46+kcLndG0=
`protect END_PROTECTED
