`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y7tHpYFK1MxDeQ/UNlGsjORSdBs2fFW0rFWAVAaRbMWFiVgpvlpn2lb0lBewQMoF
ih0jnPC4iNYXptiilk3WjUCxd931gIu60NnbHGguGL6cp9MA47ntXduLBXP+ii2W
mqDid8bJY2Y82WdNB8T3dyzW5VqAX8qksNJ9q/NQTTUz1ObZErVB2CYFOfw2C9fV
wzoUBdmFaPclUfu4dcsQpLJxAHESdg89Ph2zARqR7h8woAxUCULGq+4ymdaHhSa9
AHSPfsTVqwsPlZpHfg/JeE+3Dpn6yjh470Z3yObFItVNNVGCfPKQko+ev+/OLTXN
0tLZMKmQNxla8qEL1MZo7p97iREj8PQ0TgkBjUTOQJJ5eWqqY7G2GdwFOyG1A9xY
XvmbZ5EoFOumXwnKN6a7KyedFtGfK9eGpzUjxP48sJIwZrm4WNnRKQGArZce4uNa
2Bkj/xZf0N+hBEf1W5gljw==
`protect END_PROTECTED
