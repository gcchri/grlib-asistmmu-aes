`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OGb6UIIkuyqRdlH4st95nE8HN4K36hwH6WyvG1VIsA4kJfNjjiqKfCKpPbmQfB2r
zZm7+hQZ3MDHoNkANUorv4vxDdN8+GFog6xbQLg4gyQbtviiCok7JKWLFHgvJkgU
v9i41hLm3Twy5HYNcjF2neJe2K8xCJqe+ORH0HGkJtTwlmnxmo+VfmuD6uWK5TC5
tY9G7CCM+7s2bXWg60YAK6h6gPENSvgKkQkWk7T27dCEp74R2WkaIaqNYWvc57NO
D/KUiucp21ippGSZaVSnXg==
`protect END_PROTECTED
