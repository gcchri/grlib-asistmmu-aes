`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ugZaVUIerL5Of8Y21nYB+ff9v7w7mnj37SkvN1oh6mjMbqFkxtZmjU+2BFUsO1vX
hm4mza077McJgDkNNMOQgJ0p+FgB/bS0uAJXfObT/UDinr8reLB+m8mObcPGCR4R
deGovRDJKG4YMmsp6s5f4ovFhGaKTEQ79VqDbq71S2+yD2NzIqjjbiMtgQex9JZI
L931yFseHUW9a2tidDb9PpY0Tz360prjtdzzZvZ6y+aKoqMApNCTBXrPW2FdveCr
nm7PPAXKtThrCdqpiO2xWL+5PwL8/+eSG49z98KORIZhbVf8TqBrKfzQybH9CcrE
VEzAaXZyxEHAP4XN3hsy0fVLSonK9ewwdlOmMEh4z70kN4nveTBMwtZOyxeTNUG+
e7pYqPKAOeTdCOH5IPk8Q3fn6Sef5K+830/ScQWWdy7AGcvwTgn99FQvtjaH8Yuk
iLQ+ZwJrauGBLdPqvJ3MYQ==
`protect END_PROTECTED
