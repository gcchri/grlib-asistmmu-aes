`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J3YaVg1tDjzEpryUFUt7ch+jc8/ZqohoktMEaGqTw0ZXoC7jO2Q5DjS2XYzUDT4M
0XIjanC//7/pELVIrbYgIIT4iW5CNRIAAVRIq7a4zp5AKpF53ZKJQ185Q4FoPJRu
jqnXR6QDv49yFOR4Ci/rd/Gt3j5iL2lPKBCOGy+SiuStDMPy9TfhqDYe2mRHikCC
YqmJmBOczkVyk+iaySfhbvb5mRKhFoKSBZtRPexu3A/jMu16kOaR2qfeSTYGXkSC
b4QnmwcN3uRfd5xHPa1vVsiWaGKM+NFeEle5xcc7uutOHSnXjOCqwqw/HuGGBwKg
Pyk9aQANO5G+o1G9USKvaaqrxRhIjyRawmQGPZNKXqcb1LvAyw9A7+8AORoz/BuX
lDXb2YJ1oMJVtwW2kfkBv9KGooCfQfhNY5alucMSfiBotle96YtfT7nOnkDI7ibg
qL+vfdCJnFve3wYIwg96iwQPaCGRfjh6fMZCynIKdzfMPj3paRC8i7FoPGazBIqU
GqQNla9i/d1jvnwKTk//LETkKLUTIpVHxjYofhwTh8c/BOHp7vXDTj1V6cst9lbT
XIGutEZAOz6ZUg5Skkv5C3koM9Np8Kp4flKCyymBq6uZ8K4zmQeVKraTr5CulMot
hmW/lNr4009roMDBFigO6PwcwfzeXKaRmdVd+yZ6oa1O1eO7MvES3KOk31QitZwN
7OGPb6wzuRN3YuaTa1/SyxVHZrQRHhd4TBp6CLZruzekby8BxCSjg7U+Al3a4t7D
45D7ttI8lzf/Q1wKszAQSRV+Z21kpgg8PRsL9II8S+scewHi0jUlIbcM+586oMzz
5F/F/+xsigNsHbiBytTyLYbZAU4+mXdj8wwY5GsdeMXcb6HpEezawLiRst2Zw2jp
8qu6fuE5bIrXjwjvNkxTxRPCyZMBJxUN12nwPOfTpSJr2odLA9SRHRCgP7jXUQzN
wFM+lXlqBGlzan4j7fu70qWFgiaLLd3kL0KUZktwwPsUsWcr/Vgf0sN3RykkhlOZ
e1GNCgpgVvZzQhkK89xN+zlIRknWRauGMVPyO0vuYEmHQZkA5w0no0tHJ5RLJ1wO
cpDRnS44V5HnuUF7YW2XUM9eI7g4F/RGl6ZYKjD6DrypRwTE4qXc0rdLsM0cCZMU
myOS041SFXlkg0jCjxZExK1aqhYZAJhWEZ5/7UEm0rVcEuNAHjIjT4j4qnlajsra
UqHJqPh16Tjgrv/fRMjdaIg8/Jvzqcqq3e3pAuIX6nTROFIQ/gcykOoRaR74iu86
qdryspIlJXUz82uh20V+Z8ZTsVZTJwCliCCqXuIfWjeilGcR4HwNYdmO8CdgCZTe
hoXXiardnNn0aheUoea6TBwieH0sMTgIFnrTQzELvrgf/OtsoAgECvxqvgvbDfFC
t6L3DKDAknBVai1F7xrFewld/nORpBEmb93pAPLJgG29YtQpARWXLDVXBiWDCv/u
ULjWIZZn2Vka7YRhmze2JWl96pkoVlIibcxP3pd7tmy+RbLdS+E6NjHu+lcs0E/M
YXg1C66AzRJQKBf2b00VAn/yoH9Tm7CBkp6TlEF5BR6j7V1Zv/nXHx/rv0O2OKji
OcPBzlLeLMlEZ7ZWqB1PrDX3i/n8rhb0ROtfYVyc+StfRqpC4YZNhm2Ja+yC57lJ
QwgV8DsfzvZwXmmbVeSNajxobMB9/w5oy5ufywUAjoZpLHPaVfj8SH/JjTH4km6L
C12SAnOSh/hH/x3l8gvxtPHu+MSTcYx8LGgejLLEquU7PtH1kHYXFxeX4IKmOvKy
oFuqvioGSZgpk02gg4ZPOPxhKVOBYmBAIBRrd0PIHgsz3sws+PVItxbv5FrDzfZe
pYfACSMUGpG15uyb+32xc2L1uTyTMrv0c3fkO45P+rqd4n6t6EY7UhseO1um4bor
aUAs1/zrYG3G1t4fkaFxeyb/xa9T65bRoQNTXmI+oRTMqqc887qYd/xTvuiUqnwA
fZWx1ac19bQdyVQ8gNSR4HfcYo/CGp9OVN/cjINIggZ024wt79SwikDVuV+H5jQp
A03/5mJP/5FnJu3QsUgpn4l6qqXsR8eIZWLvdvcTmuo7D/AllTjywrU7CgaBJAW1
zyW6yCOAQWB/hPEpTN5wsc18YIY7V1RUCJbWphGvSqQNzvvemV+PLMGe4O7H3Bkx
FNEFAcne0hPtepEGldH4vVJNxr55NgH3sB5tzbJ8jjP6nUQn5kB/fsao7bAw7zDh
zIwmOjhpyWByfmxysLwcdU8kmADXTi4AMWSQNyVSdVIWIOlmrriOOdz8f3IXTsYx
nHGk1RRMdkTyLHdSmqAZp8KmayfScRy1oFRBw2gLObX7ANEf4R4x5RP0MeGFm/XR
vrvO3/DV/rhxsKr/yPRLk2/qR/KllZZK22QjtEGHc+N43ws31kWRa8K1twWA6EPf
1eSMxCf6RL7W9CecT2QwJ3BunprdYcgDOo0xENi5furZHFZgpzfxeBNi9/YhnAQv
PzItxS+BKV5oO2APjWcxoi+SbKFUZZMxKeRfalvDug3KOOREKige96KNIszSqqsP
z+hObOvprtXZycjVpdJXyTFrlSOhjJHkemZsI2AHfKCGm02db2kLJIKrMYMMoNrc
+2KmRw4+OwmeJEGmaCJiCGS/uIJF1PyghN0MAz9gfNPZhaBQ2l0HeUyY4GDexJ6M
WUzsbqHD5y9Rb9KaBxP2P290NT7CQfDuV8hTIQEH/Mw6wg6yN2hxcqxixotZHEKO
MO9CHbRCq4HqPTdmTDjowgkeRvPb4oNYw8CA3ruRBDw6SKU+ryiJD9ejk1AZkK2w
mu0FdaP+cAYDDJG4Er9GxkbWlK9r1+UXWddF/ILHQ+l/5CCNvxn/8rUNYomHCwYO
FEfO7u/qG3kd6LHRh/rB48oef1lJFEaCMrG0MmUrNtRpBcSwsPwXCvSq7vXPFE6v
IeFUBDCedzP9dLm2zJfCP98ghsEorpFZSdNVOSAZMlInS2Q2HeDrdPL3/GA13uFh
hC6guEnXzIwnJIGnegRQ3+O9lFpqy41Po+LMaIKa37WM10gMC7sI5Qo+oYArHGVO
loKoGbatrW3oL4FnsSekxsDK+KTnpNmmYLVTUbZe7V+kf5Uuxkz09bcLBLr6Yb2q
3v6O9bq8CyYR83UJ93ccF34tYC8oP/f74WxVUiAwKByVwOk+o4oVDgTPaOEx16jf
P/0wMwIVzo6Ko1Thm4NkrrizRDX125H0wa8DoX2wDvScXtF1/YMWPbBKtb/ZmDpY
dzEABagjE9uczgtcHBD0uFF8powZPE/fbyxPB36niZSNLDx2LRgyN0bqk1x1kHIN
tPO8oCtXKve1r4aqiEygZPnojwMacDTJ2Wfe5e+uHZSRgKBUyVHvMJ4dn6WWKPJS
XhjvdCzUzOXEhjs9p/jCV+jMQozQ5loYgkWwcemjy1Jjhk2Be9YNAjnV29alK6HS
iOhQLyjVmPI3rUbErA9oM1ahkvN/Nc++oZxYjRljTwCqKaWxRTUEKKL7XRnT7y/O
C6qtY5QeuHAHwYAI8N25pRiqbp6lAj8l5LylhbMD1tPEIlkMT2kXEl5cnham9fyM
Q+zjd7xFS1Dh4EPsz3gKRTl8mU2jnAcdpqY62FqZgRdkweZ11+7uZHFcgJp50h0D
03vv+cG6rU6S/wf4d/xhm/Lkp2687y2vzPkd2EPPlgat0i0KJkT8gaAyU23AhHrx
YkwVfOXJJQwthUEOCUVbnJ8S2bK31gkwrB97R5tWl3ZOBZJjwtGvGvBrJZJ6GCGa
LfwGPnW3b2nXWYrEOVV+ltFFnR750IomN/4MvD1BFz/+z2qhwYaXl9NrA2O+6hMU
+XLm7bMrs53ybptz3PpwASC5Cn0ScGcsYK8dERHp7JMz6y6VKQq3cH5U/FFHWNFy
nH5I6bMoRm7xHpA2m3s26dxrX4+/PNkPkr/6acXUYA8ZpyGQGirSYDAncGAXi818
zy0K1mJeefWQg7iqRiJlwIHx7nFrPCFx+vHr25EiYZCASawYG4Harfyy3bkAO3hS
DD1HF+eB73490JD/5tePNJBdAbbBN2kf22PySv4rYCluzWlgjZzUwXuMsMLUusAs
az3jb1ovU246ZgDaQSfEIfAFBMnrWxOaTHzYmK0thSkJOPEvkGKvtfUTgpbECk9M
b4VtvGkNCv2pdJi0OrpC/P+d1vRgMyR/mPL4xaQunPTSSpjd3BpL1Kyu5Mosal4m
mXw2uGN9bm+QpS7XImY7uftc1AwGDiYzG67+hRXgLTXXZmhTQV3rjK87GRdhLuov
FzATYIaqeE9sko5nE0TKLBAtgKkm+rjMDApNlh8KcFNspQk5YEl9/Up+/7K9ZfXK
LSBme0IZwmXEwrS2ePm4eSLEsgQ+rjpT3ZANvzwp26rOSCbk6fVTZ6Ge9JEHSivj
Fr9tbTQy+gTT7hXJ5v6pJs3oaBRNOMZNoynh79FTYJFEUZOF0Awl/QYm6O3w197u
YsejyiTgB168nasmSriSIjghEHq68L5EjZ56AAVIjSOXOto41tVNr7MG6SASrKaG
rPrnOP48tGDkYEBxtk7Mb6R+fPJ8uqohiTJTeI9z/Zu6AMSIQK3EnoKz4q6xnG4X
GMojR/P8l6NGbuSzG/HGQAKLhhD948yb/m9NtGyjJCGmZkEylJWNTjC99Sr/9X6i
aOQdg/2LsZItJmG2SGVwT6rC8pRx/rjrQXVuyeYvr0NfqdzOalufysdUEmirupfV
oJATlqwfusTC2oDMapKUgpScDNm6ALpqy5sdPvKKTGOTgwRgydopmE7sI8HKM5PB
UPg/mJ7dLstnSYXvknhiHL6p4DzShDoo7Mz62VLhy3Yu5ar1uGUr4/A28S4d192K
p0rDTqj+u8+w6i+/oPhAlNit0jQPojse5v92QVZ9W5BXU6q5fNzNpMvF0JJLi5um
rAXWTAIU3wqIf3xt7nPuRnLVofZ3ibKYVJzW405+JK3+BLmTBgvmC7c2FAvDsvrt
ozD0EXvxGWkmHoNQBkxZ4WIKPQo0Rq2x8MRQAutv2ylOcEz/CQS/k9m0SeBubrVy
IUy7g2nE/rWPNGZOfJpPL3E9Be/ejUYnFv4PabDBr/pzGdMRWAhEYDtCszuSUxmu
PUGP2WseDNCaXt2M3bgMA9sBLsEGnJuRim7js3I3Kd8zgogdjWD6sRUUOHeDugCA
XZcBVYI2GI+ZVq7EwhAkfVuJUFsqfqc9u+B0h3CZmni6O1RpTCOR9YbMwhxxcft1
/j17z1u3dZGeK9SFRAJAOQ1e54pX2USTJQIYLgdXjctAd7qYkyUaLwMe9MfXHD3f
qGh3aWkJ57re22Zaud9m1PrJ3IymVVGsQbeKjy8J0dh1PxMKe8tICgS4J7woFdyg
Yz5wuDXcUMq0AkYxlfsJ+hR2bsa4PSZ+OsD/Ug8N/bklU6u94MK4/vlQrkYipoae
FiRnsmhQKoVCjtNXzG3jAfd5IFR049We2BeT1vbMYVna25RVA6KCS7w0BPAiF/XU
uHo0zvr/mimK1xQhZ82D/Njr9LiUYGgth+RWvFN3zED7UYp/R4YGX5axQc5tqJo7
p0ibb1WR/yg9jai1eVSGrbdziDKpPoZp22YhqRWGPb9EbDiEX+4nlG8IuQKTbNPn
5ComLuMtOavadrXf3UuJTgAyCmcv13lYijHNupPEnoKb0BAvpAosbt1Cld0knwYN
jP5U2O33SVhojZhQIlZN3g2MDHMereyWnMS6uBoX4BF2iaZFWSf8cI+YKHFhqyBb
x/BvVCwu33XQbYlCtL+fIxId0Xq9f6hfNoqa8VaznLrkRpbh1QIBiH+yJ4XLUAQP
EU0XLIrYJh2mKlIOJr3+rdsb1R7JRMZMiP3mUkYmoqnI2WzhYAUnGKlqkp97bEhp
+sINfbOB50gVgvEdWFjDP6ne4IdGkfNH0rha2YgQ/YKi/qsT6WlmgjszS9hTN3Vk
q74rNrcaEGihtbNJ5yQYXt+5+5nlLCwA/6mX5bwY4OGfihobtYcGZm7jHQPhytxg
2+MrI4pQfkBTwCgTxTtVclkQ2k/Tbkte9PyrZz/lPM+BtIJR1YugWJj3Ne9WvIYN
tLg7YnHLgCjyXitIdFdzQ+DnaCK60JR+oe/O4lBcf8ogIN30UXYu2qnZOdykGLAB
8kwDUqRBuJwGMYhiwbAdjrlGruBaOpwIXdql9XNNTTfyPgrPiKNxurOODSyZhgcG
qChR8uoX/eh9XPUeBHGPEjD335Q7iS2jtUIXu/83JerleYZQDcDrtwpPoVKWv/Bw
fPf04ygrzYVk03FmeqFfQkwT8cNklz+ZrcIAHN2i4LosLzCEvWmjF0/Loy+MTPUg
CU/nwuYXGpoiNdKxMFMv8EgExEA3dV5v7a8Zi3rqMqMuIB0TqSQO2foH9kBNYYhx
Q+5qljFaIbneiU/2miV2uoHDpALAE7XCNpgyivptBFFpoiOxRttwqz86qOpwS/1/
rShDrwYclc44lg5fvZVoY1BdkproArBJL5AuDxWEwEgWXS1Paz3dp0lur8Mu62uF
O9yOdyVBDg9fEob989tyz3gYCkDLZVnFS+RSlDJBvG2MnoeDQvgtEGmPYonxLOfX
BylJVzUkt81DPQeVJHzLFCuDVb4t8K7UFIUEnqmCDoKsEkMetM4Lt0J4GnAATkjG
NtTc3mdOXNwvdkxiGORkvLlRpgcgCjnDSY6VMMS/QBqP2ZnX8TlV/YRSJXUzDHOr
UPPTAJi+nE1XkROF+ppMgLXF1CQfX/Dd55+vqBrBWCTs/zb+MHm9tDaYFYeS9lZu
a0/TOZ4iQqIdDsBLpi8Q8vnGhQ4YL7yKfDUeLOLzgARgKhoGto+kZ6VPZ2KP2Sep
/2khuAXta0ol3KmWpPRQCOA/BrMbZ3GjsS4W59jGA+9ttSJ9FMIp1e0OaCEQLuy6
ly9KRk2UpVdfzvuPJt5iM7374NnFfW8AKakI1CiWIu1j2ZQ/doLX1EErqXwPBT/k
jL+H0oe0wWYoEbYrzK8JqD5IZn7ywc0PfuQbM13gIY218Jmmu9NX2EpTapuw0FGz
OIHV5cP67RznY9xfixpuGQAQpjueO2dIqkiX6hv8P55LdGiLAtztDnNz7zR5a2oG
JyqRPpQv5OnFjmV04RBwXo0P5xOVmtyBqoCup/1tSqiOhoHGaCx8VPDK8Ud6BOvl
BjvG4cLkDrNYXFfDF4QSxwNTk+zARaQ6d9akvk7ienKqVKkyKf4IYFQS7nxTS/4D
Ox3Fau/v2AGReLBdCnn/Hnk3HvbNDgm0znPD6HQwzgRzmpr5XU3hLhoFh34JQr9P
F8OHLO8ofiC+wVU3HxX7Nnh0wpwFv0yBklTo0qhBI0CISav3HcS1WdT2B1jCaHIp
Jg3v3Na7/tmdDjkj45YR9Q5gNL7LeUxepa8XsoK2mz2v18NMeFF9R7820BiRY5eu
heR/mlcEbrxgiitvaOe9PtazMBwH6mpS4JGTofG9+1wr6z/q5kBDkNhe9qAE82Bc
4+3Ob/RGxJpOIvz6DBtZsmYFBNnDWU3o23pj3/3f7oHwFnRpzimPUHxucWvQubC4
wqWPQgt0ElzGTk7r8crpaMbImJrItyJADtrrGjDdCDAo2clNgxHap4quqI9oEu4R
pByk9lVy+Kekam40lXhsjXzW7/+NbmVpW5OuaGPXSQniOv0DSwurgX/9Ht1dU9Ad
arca1SGMAny6tHATxDiUohotwG0Z32ZfCAjMilX9V2/DSsx6KaxCHTW5lZfr3Bq2
J2ohVrFP/58x1jDwFLWoNaLIwMUOU9FbE9OYxp2ZMYyMSwj1i/o+1g5poNl7k4OU
XuUlEar9vFZvICk46+LWKGVI7nJs8wC72ToZRyNQjtr0mZZRaAotDBpIN08hSBab
6JbuejS4+EvMkppvI/QFltEQ9kohd6RyvvF/NFSYtSs+cNMDJVvHzRklDWUl40vL
P+ijel6/DpYC2cz/xfZEeN74xy8GVTGuLmS3GTVkrF2e3qgXOFNe5/SJAhXSDnbb
y4z9wCJqzDhVzQwBvj5G3qX1vruPEz4linQPJYzeTZn6Y0VZ2OIdnaKWfCdV+AyH
HqMApBuWh38jXUvwhyKP4+Z8n2PcE2p6IFtBU09slsLDC3iNaoYsftW1nHip4Gvy
VdyXcxRM6wUWBfItLKL1Oekkg6V9NUWJS9sTLEVaJkpdyLDRNZwMTHvZH8PwQfR2
yyjhqjqCi66vT6XGjSG7Mu0wA5Zv7fWMd7OqMiXb9RtGwvRHfhY55pifiljD8lsF
QL72QY8OsRht6DsbnLReAJCI0VEUuSANhNAFpoVfrKG7hBdpCgpXleXoE7Gl94Z0
6GMX+v2+XhfFYyFtbQIRPSbTFj30hZ8+G4/VV9uG6IrfJ7QpIRHvetbPA9w8W6Nn
Osw6OLxXfFt6S+CWCmdGNhZmMqoH6EOrdYuLLBrG5iPJidjvCdsBqcCA/ALO0rG3
zMyXuDMXLn9Zp8gKfEVqAIdAWGC44MhnOg6D0e5IfMDjwhixZEkN9qEm8/QPpDqD
onjw99qXcQpKVH9iNBPLQXqABU40LnTAoGXtafpn2Kfl6Rz0aUAyih2Q6BeXY8Gy
r422FMWUOP/gxZ9vnUWTE7YUDuWpVM8581S5Wjr8rdE2DgfiU0424CvjZx99qQcv
FoPZY9CEQrYl3itWJ2sV6lVBNIPPjQVfaEl6uJ2ky4T9B0t22wyGamrPznFL9EfU
RW9fVgKAzKqP95/VAFCFrolfWgfnw8QQ0yqbQGykRsN+TtzqKDMWgzxc0l+Ykrpt
qwq4fllMWYbjiSjWzciEAxiLcBidDX9nMXqxQUqm+nUnjltT77YXRstBoMklJoBB
rKyFMY7ds4SOHuOinvvPqbkyIh1rNrSicYKckpDjp2jLtYYoXZBaDD4fmbY84oAw
RzkrtbS5ZII6qYPjvEFWIYNxoQNO3m4Po+hg+imA/2zYFHfwUab7dB8AffuN8Cd7
88y6QVdOQdITRqQazQzAGVptx3vC2YqqNs53rVKyvel+LmgffBOiA7ml1B5KIU+s
6bS3JOTBwptLJ/078SpPg0GhL7Hn7zUoupQB3WMMfjC8woT+gHXzzEH3GGMP++yI
x85MGQEsbLWT3Ahv74EKv+YTaVcWPYQHJT5E/OTLlg4l7s8xGM9Gz/kwORo7YAaz
it6d59omb8rqapKiQFwLeS45Gl4tlTIswsnwkJFo7f2Ddd/28Cewk2e29mrxmVzV
C+Nf8CBaHSVam13sGujCbrVpVC8P8wO/nGlHcC+NW4uWzANzWPo4DeY/4viVl2fe
KGfe+KXTRX/NQcYg3gnMeJQX8KyRSSnciaEnA9120it5/eq0YUTIg25JluxCax0A
7ZJ9Z/xR4ubnxkVvShbQUaHSD+5Ef6k9UFL/yGF+vBHcYuuaxb0DNrrYFuEHEdoH
FgaIGzKGLEYU5fNRfkvcBOwpRnVzVrsZ56IY2Wmzp9OIs1l2CfwuNbZnZlnsOJ3t
qsA2IgXboYFTmBxM+PxMJKgTleQ6TNeOivRPIoN1qlXtbPIaWd7kflDSei7lFu/K
ayqgStAdmAn6l5IKjWTD9+5c6LAUxEU+dr5yew0b0OnaGY4BNCHtQZsEpBfsVL2S
JiuJ6ANPbByB3Ca8Z4I/J8SadsIdC58ThtuPSvTd9sUfWyrDWtMpZTTeJmgJP2wh
BSMB+as5OXOn/VUWAM0ncNkRjrT0OtG7BcpuDwOCU1JHR9yzcLFFVVUvbp3Bot0z
hfJu+39fktJzeNzwaM+3yzpcWibmopmJxLVRE9gCXVIjc4wXYdkqFK08b5hvY+R0
DDC8MdlQOM9H4alS3bghekZmoaJgy6DfUa7zkTADdWSipoXwOQ19zFOy0PO978tj
3TUS929Q/AFtdM1ZM1UYFOP5uTLM7oMLekEF/LKY2pCfIm1VqdRdyzhOEdvNfCe5
8+ZwMYYurPRJRF8XXya8DOJPJnFv75Go9OuaRQLRSLQYZiN43AJlMz7JkOcccEO0
FFQWFy9I6vq55XfbQ76O4xoSHY70/nxGsZCEtI3IkWhx1kfPxzC/++3Rw/XBHF90
je/q8g+5VKg+9O0vFFPF2LiFR14l4/C8A5VcFOFAiQZyI60LGbXyDIl5dyitOotG
r499FlIvUDOcNVSZjs0XfAxcFKCyrTqyrXRquPbEsWJwYtgLf3NoAqqJF0dVmBsw
lieS7n4l61Xx3OSN8m5BiaWf8SYOenusmtJklFjUBIpcd1SiV//kpAi/SBh8yJFH
WMaRUp+yu9C7L1SNeHcH6Mt3D3ANIIv85BL8uWwrL2fMkFOwQiY+mKvpNdnIYvXV
5eOb9MWeBwAZ2NOc6tMvud3XZgzWL6PDltiqAuM8Xu8n7IA4JVIUjX2TlrPNrE9Q
2d5/O/i+AIwWDLQRM4vGmxDGj4CT+lfzTHHkIg+tJuXHwBfviUwIV1iWDLWs7M6n
/TdmsFIJyIKA9gxbF9IjjnaabFsGCmc75gv0Lc02DqA1MrJmOyTi1pAHgvuqrO6s
1Qll18/HxLPtWvKXEJs5Pah7W8TatnSQdEfdl2YQDaW9NLXspmGQIC6xti2J0pVf
HOtfk6RS1rGtCSBXfOt7x6kmwEc89Xi3VPlEQ88jbp+4TQj5PiQmYZQTnF992i6i
7Nn7E8mQNLUuF0ew97jJrxAsPoE85VmNGp0VwHWevIFjjomhwv+4w7sSWehXs9xx
w2uN/e8gDhTv4BfkgLRwuMcXb16bwf6D4DPFtf2YQKOg3LXXRHmi1csinNdybyAY
qAKSENhpZkbUsBQJjeA0EqAErveDwE7s+oJg9HNshQfQbhEi3o1e5owKntgU9JsS
ku0plbmC5IQvBn4AceyDjnUYQYHikqDaA6iH6tEO7Wly4fVWWzK8sozuot6N1gbn
EU8QQrtjm9vPDLbPnI2W2RTDAz8ilS4NQpRpvL1Bf3GLxcDDpJymxOavx/Cw6g4T
pDtGhnR+Y7ClEHr3hzymmLvMWuRbXz29Uwlinn6D0GDjSboL7w4lqfmrr+V3raBp
OVS899BO7qJGkU+pqBRJ87Oy9ddgKZPh7jpGjVSy2SU0/BrlWciHsystMf/QIEy9
SGB3Ahn7SjQwBs3z9XUV+ubAdceZ17kMIVk1xyN7vXAZ5zqhGcDy4h9hxILedGBa
0RQTUVasC6GmcMUoJxrZmCIr/wYhiFTFwCb9ld8p0t1w1utBmlC8OSd12i7oE4Ad
E3NFzBTveL0ndd+Od4rMUrt1e67nFLdCOC+en4qaLE6zT32qZfJ3tfNrQkEWzKtF
D1f1zbXiOrEiJzCBRFBD+MwcnbOzBvi1OS04hUeMpXHAOF9NHs7SX4yE/CzfTY3N
/sBnpTJM0Ft3c0VLXqg4JGtY3M3fSXJYO9Hks50/940B7No1AFyjwiCmCfAiXTjR
aBNj9EqffTk7EZEYLXtK5u+PTh3eVsdX8V+KlKzGkWR5siIBY9F6i+amM0BTsFfe
pAHtJ4p1GaVYUgJCFr9j9mAlw/qHPIglSb72M5SoiGpKsPg04/wyYp7qzTy80/cW
VCKRt4l4UzIiOxtKL2Se2pl/sVLvT+gzKHY/4edAK4CBzu8HgXPoLt+YVAQ4rpcw
J6AAUts8h9Cdfrg1kkXDTZ3v+65d2StA+GqIyjBkpM+vFEE3y9FSBrT2om0LSVzX
eGEy5hDh8Cy685bFXcePfm6KCoFJSWQXsnSLl/ksCOfFT83AzO8kiw3ocawVAi9I
ZCicN4R0cJ2BVQ3ddVzATynCJFWBtwVYex0dpv3g1KTpZEqw55XbpRIw/T47qWqd
W571PtQ//2UtilaruwZLmf+h8jWAC21MfbBATalXh9n4wQs9Yj2hjzr3c77E+w8k
Xxx5UoGeg578Js2Us8A20sUbuVngy+2hLWbXPbc7LkaUg/cLzufAszkawrHft2JO
DCLtr9jIpYdef5kCxq6tMnlddL1A2mBjAyomdgBoVlnciZdbBEv++hiAdGDwC8xw
JbOsEwixLLbL4/Rc0qEiCuC1YrLOjmWuGXeGrUYmfwiwa8WsRu9UPR0fpZWVaEDD
pCkx0aUeWNg6D6BVnHk2zGg5qkvHnld+TaAxNDQ/rLUOhnLUa28fe3KvALkvsW+w
3gCBUet0oPLTXSehY1fo2HrbLMDK+08xDKER8cS6ZA3vfAUBCbjQEIMg1TyF54Ks
DeNOXO8I4/DSMV2vmNSOFa0FAItNgCJwxn85Nn7JrhDVggsspZPqEhx8nMzrfCJ7
SnsLFInys5auOSRDgtolzR7StdAacUcsO6PO1qEp2YeqgOxbkeUmkoFcMzrAUlcw
nGx1bBL2wBqPsd4164DPHewRDUSIJOT1NCvryJNP06Lb6T782XtmJiQpe46lXe+M
B7MDgq1Xxw3oQ1mP7IjJb2LusES7qJQX9+u++cGPNgZinMVR5vaVW5NV7let4tV/
vsusafdfh0P63AcNpCaO3HW+ANfdu6wLyuEitWkDNl5XRrHoIVrUZEZw/hbscrIV
DhRQClzBi5sWCKGaUOVL9w/oQz8jajlswbm8jd/8KHrbbhraQWuYr7M/9fZjAnoH
IVJlQIon9c+JrRv2nkpfbUnYN4J37ykPIzPvqt71+V3pkjGROT+4ummhFD5d7J5I
YI4d3fdoNIPkuMIs+oFr1JSmdjltWOIU2+PmHaU9PF5Nn1Nb/g9ko7auyrF0mBE5
WIq01JXvEd7lfFsjubKbO7uHA7X86GjvjSRqneR6x2J/Zw1qvVEn7mUxVlKxt1eJ
eLoblWvmn4Zwg/sUt9JCoCVg4NefSg3M6EvNXfmmuhia+ThE3c0qZWaOxHmYdOqW
g04az2M35wkZoFAPgZ5LYlPoN2TQ42MIpgFFbGL2eaHQRjQhZ0Jc8zPoHxsB4m0K
QXqTOU0d0bpw42OEmqJ2/OrfIDF6muFYNvmgkLXbf7x/rZF6ldNvQcgTYScNP3E7
4ixoiVWlYVUorWr4RE5ce7YLQ9UEzy5ggI6PQhXskLpjaRV04+ICE+7GNcUybmvX
LWNDmnxumMVhNI3n2PDVduIXwrFbtYV8fB8LyJ9dwZCLMBwjx1jqBvo6RewGv1E8
kTXz8AmLnPoX11RSoH85T9E7BaQa7e4a2KGEZTLzNYx1uOg80tWlkw4fmDjT3zJ1
Ewn3xz1TBHorHRI9CgEV+rV/04X6cWwyfkdZf5lo8fGSQIqXgJuAsbgu8y69RyZu
gUfVDsO/2z0hYDRKzHkDmJXxCkTOnMc5uHWZ54XPjNaQgAJuGdRzm8WWR4E4f8fV
vei4lvjaeuuny3ssFRWKPGGTNl/OxVR3ehFHzX4ecWU=
`protect END_PROTECTED
