`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
leMg/jnzFrohZdsjJn513q2Tlz62LnuOWXVhfOht/ZkAEPQj8uPkNgIT9gw3vRLn
9hQnDPO4b6VZByt9wEO5+gAlCUwoKOggOaU4cHNcZ/os6CoiD5NydVOgZFAnu2fr
jFy80wqvMsdHs0/RouiGaBbF/44/Pka46Ux4pCVbSUOGkVD67aPF84h1RR+KDe5q
2bNfe3j7sz/oM/S9NY1uAIwoOcoO0Tmr1hWav5ALE4hIafNpmFTV0YEqNK8w34Q5
ASLN5W2NVlTr6afBBzHdyodkW0oNNxCBm9oxBCpH+qInWBA0GhTOxAQE7URNkbNc
y6cPCQbv0arZUkuW1etVw4S0b+gO1a4BXYqxPwrXvbtxgXvFXUkpotAR+nM8s/P5
bqvKkPKzXgRxjAHxP9hfUevYspKRCYG6Pbh5mp0kCoj2QOp1cOEhx7T9HKYZqBvm
jmJeieHPpJH9pefSIgpqNM+1KTZ73fh5f0sShaiWkna3MftbWakr9x36YGxguQyw
PGlrLNqCFxznib6D/0esRekq1LW1mlSnqdzKCUrsIuo=
`protect END_PROTECTED
