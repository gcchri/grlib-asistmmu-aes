`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OYsnx1ZkibEUL4nllXwWuiE3SV0AhxZ/mQYNAedFIXZ38Hb/q4mOpxmAahaa6ffc
wJgiUxgGQ9/NYJHCBYJx0z/wbs3fPsHLKjfC4FVlcC/ySIUXkIVcOcEoQMANH9/h
htoyLXPzecvhAuEg87DYCi9Pl1aBjM5ZEuHUDd+sMUI8754g39TwA4iOlO/ujzdD
bvAQR1m5mHDW4GYyIpGtSPHklHAtDLwPzfvAKnYyoo+oAH1i9HDZj5qg4gZqkufy
87bFZEMkNekL7G3QGEzF5vxSLEg+KvfFh3Addifd5rPpfV5LPA+b0wk/fzFld4/V
xrxPZTmt6f8ewzlvq95rOGjOQfxggN5Ca2fiQXQM8eMdjWxmQNXx5H2wDZf4Mz2M
4l5cI4ndClHbwiaBpRaDMKvi3TxvnHoE+XIkqmeJcmAQhhwMTfYUoyxTeE2p2ObO
UmmKngp/HcjKv9y8i8iSTY9yUwpsaIqLMsq9Z/g7xSEN9chHp0AxxTGPantIM9eD
x/aGPTmo+QFWMocFggzjRcVr47wfP8XcE41tvj6iHvgiysu90ePcXrbYiDAJC2df
ItecEGXjDdLf0XtKr1B+qavEpd1n8DZnjbpgZorm59QK2d4PGAU6WBHSdr13iFjG
+BwllW66F6OhoFfJe+Tn8celyUQDBa6mBZCSn2xxeyA7z9zW806o/+vFAh6QNg0x
w9vgXyvRt8WfD21IPtLbo9LK0hhogeE3PSBHgYosBDp1UU3B8lkCgqBcL7lNZcnR
yk8CF+isdqvLs6AP5tPFhQMzMoaGN9E88MMITgvKQznvQh+aXQDP9+j5r9ek0SXe
k3GDDYXCNsnKNLDY8/jQF49gIG27/BziYwfTMFSTCzjWNU9/Rz0HJMXdqNhdu1XT
gTXANYrT21jPIv2z7Kp6CcM2j3Jqcgm+XVJ4NAOSWglLZBuafNZ2Dz4SJuNxL4J7
Ra5nPjbkRPdEBCUQcEOOY34qQwUfN3CH18cV3YRRrIPqCJ6TAHkKHxyGLNoTZ7MK
4gpBmRPMk6J15P3LPA14N3t0wlQhPDRJ4I+sq8KMGDz8desAYNdOQSdGAp7aCug6
UTL9kwEYBPocLEJpjmfz8J/vMR+Tfgx2S43clvObDUYHyB3V4HlViERx7WqMJC7c
+7SFo95dkkIzFaRg7IQHqzrXkeY5wNu8TQEQZfdOLEGU08gR2gm1CkPu4gbuNEVm
BvAQuFWI7E7JsfIciJFpFmeDheV5DkvAE+kQ8HYaqHMb2n8Mgo2xvoY+snIy2BzU
dI5qTWPicDEuGuQzjqGJ9CG8+TSJ0VPnr4KanJv2j5VAdKSsJZm7QeZh2CdVjlIR
JFBoIjbFgMj3bqXVkFq33k6G+Ywvo9y9+FqOkKCBztubeCyFQTn9R9JLtvwTSwn5
2LFfm5n8f2mFC3az0DWZYvO4iT/Jzve27p9oLYCK/30ekgUqisubpWTH1BkS/1uI
UuLwIst5NTdhUAD8R4xa7BZEU5E5Io7ivH09JXFMGNvJdLPccv5XRcrghTB8DFqc
8OVP38+UEYBCY5G89rDHt01fqrA7ZKPscy2Uv8Py6X4+aWJbajQaJNE74fvBYOw7
w4BWZQnu41bVBRWE2vS6QFZsIAZ+i0jPKdmEjlWFox5cLLvYxkWOJjmbnojv+ttS
iBiGiPPDh8g8n5UMm6wahoe3Dx68hryBM27aOqj1gN8Il6ViQsFJedqLdiUKqdQY
VH9OkO8Qdt3GTzYjHz+z+MaCc4JupT70EQCcMfUgN9sxuq+otcg3LW275CqYlAct
+C81HFV2M6c99SBfW8wHNQ00IRfhDrespprw03Y0SMvl9bAgzbC8aRjNZgpuhMqa
7hxOZzldePcKxfYmiLAUT6WCerT35CV1r2dkWeZVSRhKSbVNrwOckTi9Pu8Vg/R7
5nmp/7zAeaEZ5WI69m87Flp85yDMs1L/JAwX+lvAs3TERX/U4eP169DRA4nWgtfo
J4Hqh4a6dY2l80Vl4Qo9QHbzKBmtvsOUr1yn6EdOY7EZPPjD2cGwru770Yr20AaZ
4dXTLCIZUAOIZeOtDiCkk+f3UrkQeVVA0pjzuvwH7T4Rj78X4v7/IZc+lXbfzm1P
wMEhEcjgxgeiSDJz03xSEMwEjI+XHwIwEdSpOMMwvnEd/fM5mkXrAzwhzq0xKkgt
7JjXLDNd8+yEans7apU+gRMVrEK5lf1Y/oOB9W07Zek8bXflKSHEaWXd3PrwEF1Q
fZxDNkBPT7pab5aZ+mYejFfT4jAYegXT+zWCl19MlrYEmkx2wP9LHlSouZtlb2p2
l/a6wpaDK0e4bmF6aVQSJMR/b7vb9fqSS+Pvb7utk1yoPLZeO8kXFbnBoRtOz4ml
c9dpiEAZ+uSG9auPmHuF3ravVqiNF4dDUG/Ud8LzjtGZGL9J7wDV3tTmH4J5xtsV
XKhuqUAt9roIoTZYgmaUGEhwXAX6FNfL9+4ryRTQLRqKRjaFbNV6tgMSlim8fn/Z
sj68Zo1YXHM7RsVBIcp5bPaFS5KugFABTHY1YPWnaAdp2QWlskBQaeuVD4iH2EeX
ij92ts410mL8RDSxtwsyNd3lYoGHx+0Gm2M6l6XYaPGoFz371vQF2kvEu+vnMgdB
RYUopD1/alDBLwU7ocxAiPrZIsRa2bNNmSK68S/WuIg1nwCyhKRPp1EIN1VhTmjQ
g0O7dzEMyE7OIRQmJvr7xYKF4+Ix064FpG8dj5/kS7X/jmDTk0AUxyYvXISbxku7
ZoIt1o0+7M53J5nf2DnshV9kNW2qd4nucURGzm337B8Bm5OsXvF+3lsk4Q100GDx
1c13bpw6dAEle56FCRGAJHiSvJ8aBIRxOro+G7jU0xjuM6OhyL/9RAXlwXQKpWUa
8J5fVn91PvWPeOurlfI9ku5JFRHko6NpcQV0u3QSGXh1mUU6/dudS87AKoG7NP/W
34zMhvSVsMriEt5cMEWmFVYojorUJ8YqdWNc4bjxrg1eafUm9MM3atkchL/s05T6
F1ui5f51GStMi8HOt8atLrAIWQiixYSM/FxuNl5a06WI2MThxMcSVkSbnzcrN2iX
iN5UKA9SkRWKfgEzIzC668BUT6647C3rdCG1KZHkgBLez4cvParVvLvNaQ7YXTju
nGVcGTn0cyhPzVmHBTnegMg4gqv99zWrcbOc3Gao8SUEvomOPY8HqfBj/N5TVJyt
Notl30oxBaVbPrXVCJbWVqv8xOX1MRPIuMru/xZ1MxeYO/xv+XAo4AYLhjE9wu5y
TrHpplV85wsvc4C0KmxmI+nmHOVpJ9Uzh+Q+rXjvkd2zOFsW2MDeGKNf1+5m15zo
bMICx+U+weRZLr+oWQYD58EAUtcydJ+REpEgb2p6t+XCN9hWUSDTvLR2nQTZtL49
qjc1Cmkoqp02HjB+cEiGhMUMqnVC/4Sji/HKKIGLGUwoMvqZ8tVTJ0rxgxDUc6v8
rIOgw1biKM6uvX7kSJ3bMaKfxp59Rv5iuA7N/7ySmcvqyZ9Rxjr6iRL6mIA2xw/k
7KuCWL//MB17SFasAAd4EUhKJVHfOdiBcpvcQEt4/eXBfM7yZD8y9nm2AgBQRDex
kI4KGfJsORvmKAVyMv6ghRrGKPm8P5DJ2tZw+pT+LKNLAD7/jv2fGFKsvModn9Tv
IYEKvR4G5/61RPbRP17a1i+mDWfKpWivBsxRgSL3Xjswe3S8/lr+gOlgY0tYqkxB
1xWBVGVIRQFPRVMU3iNLJUFl6PdI639xlsEBHydZJN3z+rx9d8C49WOZf77kOdJm
AAuUoJ7kivCO4mMhjtHwtiL8W6dnuG2LwtTXMahvajZT2mAQi5OU5zStk6e6vZkG
XngJPeyx4mq38bYRPaEJoJ1JQsMtppnAM6Gs8/AMaPGCiixc/ih9TU/x3q4wvIiB
imS9pzWRV7MGrVTS/HeQ6mGws2gfmviKodllVPFGfLvLkeb0HM8Pb0zQl+qerImX
RR9m0IFotDpxnAodEA1n5IVdD6GTS4GhfCxG58ZmGYiJKIDm4IpSQEsvxoRsMVgK
UfvGBwXH/4hnMVJzqKUuNad+XgWA434FhLqNB9u8qR9/d+Fhr1t52mk7d2UUWhIK
N/g7w9OQ3eUEKBseWIQRcJZEvpjmys4Hon7VaRGc6ZY2k3na+aUdclWM26d7ZVdw
emmMJMmQSkGu42Epv9fuwFTdktVAWN6QV25Smp3CxrCYK4jmGx1DBH5T4hYUu4HW
CLeC9WoM+xbo8tQN2Jn9XKOwuAK6NXgN8+MGXVwW+qQ8RGFqeDIyybCOJ8nUYuEH
hcdDGQy/kBs0yaJAlKcd+v41WtvTtWcPLNz6n16W64kIEXbWcM4NamNdvp1ArJg1
KqMw1+ULDhGdDpZpjaKpOoXiGgbaAFS3beKi/HntFaXDz3dXD3BcWvDq9WBOmrEC
0oINGiIow7WjYwvPK2hkGtdpjF0W9+UQgQZARno6E20pxZtrf+y/D+//3LLJpn+p
2ljRf4QMLs+hrWq5akcP3FNTiascUlJyXFU27HixTrQIsvI8oSjpwBmIeWQyGQq7
Xvpce9lL6iAHO242bnxvd0PeIzkcmzjFrONNAFNAABpYQoW/JDwDu8n63G5begcV
DBEtKhKXJfhcIyhsmwfQ4n50VIXjfiK2/clMfzwtVh5OFsNIP4xIRUIgtlneScU7
yheGNbovbksAFg8cJC46npI0PJ+en8zOWrGxEOxtw8nhJxVkscaLZqSaG/vfyvCt
F5kPbz5xHeBcoYHtP4EfLEVdxWEDbDA/lFW+cFu7UD3xS6MlTdCNmciDQ5zs6OgV
6Z9W6lFWcMZ3U6Nxo/MMxZeW8RUhqWJJtbd7rgbOMNNUINaUj/QprLeUuqjloTLo
/G4diArc1RB2OlTDt8hJ3dutNR3bk4cE8Edic1n+0oi/xRNCSpJNZIrxKDTZ3bAg
wuulMqOh7FAbkmekDA8oNJy4Bgkw6HYmq1YRiyHZMUf5sSIORG9mSuWEejJ2JC2Q
25T/HssoHICf+QUNk72DqAk9VE+sFpEP2gOQD/RUNVvT1H23CAj+ldTekxs5yA1X
fKK/FPf8ZLPHDhXW1hBReXos/bG43DhJuDKxdQRTPeAXPER3BtI9zfHbvRK4MWJq
sKx7f0qxwhtf7Mb7lZXFMVJqOKngyLanslJgr0kBCBzcXrIqNjg0H0Qd/P8klo9I
zSWPCnkXjqkd/xftgWgtEi8T+g22iZTZwthe7aQEubbvVNyL6Rv/7wlf28EyRHd2
p7prH+4opkAE3e1rQNoilg83ZZyrfliS9r8KF0uQ+Ie48/q6S0bBjOPNQgWtecqG
uBAyFHePsNPLzbDf4mh2IGh21ry8xmfk4ygatwj1YQLHzWqFf8EixeKdy7cs9LKp
iyOvlNeb5L0CMyUEyZNpqh8ml5E8kIA315Tpufrkv+9O//64ACt2dVrxvaTmpJ+A
MG+stTihYM9ljziCKftIdxClTO0arQ0YYCdFOV8Hu0DF3Pg7gPmcY+eYWlBqOzku
PWJZBCd6pccUUhu7hMRgmXtehALtj3elUE65yIvF05JwYgH+jMtsH8kLq+dsaYLM
s6BBP8FG9fgEb+CC5ibq2GG4ZyoVgF+weeaA+huUTjzmYxogM7ZuyxXLwJ3PUFHS
gBoiIMdT9/V4dFWqamJRbVNY1t05jXmYMrNa/+tdXecyRWegjwrh7jRb8X6Pam6R
POQXQTeYws3FiSxLWU8EXFmc9JcjoHw2r7TBgJ4Im2LwZBPXOMSri4GzGwgKBM1k
c1+WWYNC/fzJ1hQbFxmbAC+yp8nUZP+ooeys3wA1SCZUGJfLT91Lt+j/x5prXjsP
CMwEgz/PvUxrCISqxadn1BboOVKkJsep82iWHslJCsw0aY6lGvD/zju/xQVN2owh
n6NbvmFAtAVwSZiDTDzWOtSFXGzle2UDfB5TIe21x6GyCJrCoYwZCkK5DbGLxAMk
l+LBWNx95AkV6cm8rXtGJWptOtYJb1lEy683PubhQhq/feUH3lMSLiN9t6xbgzR0
Q4XlAxqc6zw066s1DwfISKUUhHuuX4YiaQBgrH985/ZVrK5U5MQlyB9Lqw+iOXEE
grCU56Zzq1nxF3SoXWxut6eo/aKv8ZkqpgCzHUVMYbjcWtnp3pG6ehqCNH1Kfbf6
hWo/POMKlmn+5RtfIjBFNCJVzPsEVfBrtH1hbv8i61Cz6sSTtM1oFIlQasGzYZTV
XpwXLFCPEXDac/LO1f0BksW9JjpgnQH7qI0sOrgnr1O5r4bpELiSKGhTTlNGFZG5
lmVXXkpZla9vbJJt+QupcWAZ3mI/tCxGOIutRwxaTgnVilMnA5EYvkdmHIrk3Rz0
FKWKz2PmMMwxQrauScX0Ge/BerlSOOayM2Cplclf1BqEv0zmzJF2HoUUuqwl8k+4
4qQfQDCqUG12O5UKxrpJ8OS81HLwr45TnQ8w+OGEv02eoxNICozmq21NctHN0fM1
FdsrIgS3qxSGrYKUR3dROPjeV61trG26VIClsBeHP9fs5WtqpEKkz8vyrP2IvSzU
9nkHhOZIjvSWA7dTCvQu6XnQRRQ6sF/yNoVDUeYyr1/Tm80tNpGbeKQYIfgde7UT
I+Q4O/T4FUx7dwo286uLLJt5vR1dmXfn7Nrf2jsNad7vAB1rniX1BMC8camDEPkl
IxsqBa26d2faYwAZBc0jrSdsYM3MQnraqxMkkbtyGCpGX8vZcRz1JsNdTaq7/2IM
XbruBNDZOqfuDiUedAmyMEuV+lDrjoWSQ/9chUsbagbAw/BM2Y1fUjhhKJhY0L6K
eP6H2qUR3lxHz7st2BwS1mao3xvX6eJDRrSbepHXjlnoR4R1WVmWYPnjTSs8svq7
UcglYukknN8cq7faJIxkMTHQZRYn1s4Ok4o3gSMeXEk90nDs7Ps7BMfkjtF35x4O
5Zu/9Ni7ym6dGk46h8J9v/T1/xUtJAwEKAVCgjanfIfhM8tJJ5LMO20YQOslN3bl
RwohwHxmm303PYAg+XrNTVx3LCjsgk7VEGqLGWF4Ff+/d/tT+YOtwzyM6UQ8fgpt
trLVeDSehhcM8bh1rmmXCJn44x5dzcrnVPhilowvXef1YFCPfMk3QLl5hVV46I3B
f+y2tcZQyOYBfqiQ/MJgz0W8iVBjms5Bz8Amxv3seJzMIfB9fNNHw47iMNbjme0y
cR4mmoJEXVMQYFYNg3gavby97XE9nYzvVTsB3oF58KtBWU16F5IyuuKVr04fz2Ku
8+H8I5T9zwix7OSFWB1Ds+pLRI4PQ40EzmpVpI82C7RgG+DhL7oSMnnNHKe0gruo
rvTowOkONJ0tzaikdp3a37pu3zfZ2LGK16rqzJy/4UVmGSInRUwxF02qqDbOfwfJ
BViybqquy7R7jZoZAImYeYPyncnqwwgA7cNzbYK6zRMFV8o2O676UM1PzNX1mG51
960tWlyWolBfomqI2LUm3AwRIiQc1fShkJJkw2ZXQIkGlf0CU23QkvEqtqrBw4ZO
W4fx653MskEDWNkROE0Ull+Lx/lKtx6Xs5k2KgmdqiUa8EkbrilhQXz2IZB24i/4
CC2u2SDxK10Nt/YCqHB5KsKKBZo1nqeS1YQNdCmgDd8TQg6uLFgBKpc7CeCSTYd+
1l9Gs3dbD1yomYsWWl9g/Y1qWDMFN3J31AO7eYdQyGnF7qpNUQHrg/DWB7V0gcXV
Kp/1xQsS7xU6qHm6Y5Mj62EB+zz100UU4vBFM7qcWhX5qa1SLyM0OWoh1SIse20m
IsQO0EZ3044YWf9tD6nK2Q==
`protect END_PROTECTED
