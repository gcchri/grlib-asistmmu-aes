`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I/ORl3y/n0fvaCMpdRBX4T2016AitUJFtbdLt4rZ7/lg9HtXFM6OG8qgjrch3JPv
O+2HXnP+P1uJzjayXE+kZtFwxviukRbEF0KZ3DasDeMMKoi2xvVKUByDoHr2YPRo
SqgnE5rpIT1zq/LjZ/tiuVQJ/WxwK2CMesJs2JsQKQmWhthjcC0wAGPRPbusLX4/
MB0cq0GUCLl/dIjbao6sZ4Kto1YYuDFxuJ5lq5oWva+Hxn44rDBPZ6O7L8x3Hace
sU4vMZ+PGDWbYGIT1PV2hhFreeTXtJF4sNEDhLCPtpKZxSrcxqW3S7x4sRSsWbXF
rAIm2+4ru6Cr9ogI0M/kMBEBYUNCwst1KYXa/8Vzi4JLSd90CDtjcvwvThWIur/r
OvzfMCRYso+Dx00pnp4JkGG9htJb8MaX0kxm4E3Bfq7xo7FezzfvWkV5jafBZZVJ
aS8guVNlB4Jkf8b9Lr62tItKLdrq5eEil4/aCW/6YGePK61ZgEl+w4MkojVqqwYg
kVD7QAjS9hwIJ73jRf1VJemGaIwLYFbozbJWhRfkAjFWZBd4GYZZSlGwbkLyd5Ug
oiCycyRG+ZCrEbA5XuWj/59BQ+oWkMAGvJrBvS0vpmDp+ldGjWgBCX8aNp8ULFVI
lneFu6d3HeTkBMC0Z8it5zGrEXQvQw/TtMA2xf6rYe0kV5GpXK/YiLZ7KOjw3kKy
sJAtAh3tCQnnvW9NkR2uwammZDylOPyQYR5a9W1wG6pvcqGjDFTRwRxHyDHul3X/
ZJ85pZcvRP7FfvvufMefqVRpomTOvCwk1FUxMuxUvTKrnazBnqDimOeaQhN9Vl7W
wLC4YSD/eknCZSxm9T6Tezypbcw9zK+Rk5CApFfxTGI+8pHhpktuFkiwJhDa94yL
zUcmA1O9AGES9xde0Wt+76Mcgu7ueQcmOAFzVTT1R1F+mfp9emgGjLkvhDiaSWZV
SmoEqqSJVRCZxgrn6KxWEotRwB279lA3CD7Mn40wEDNXd7Zf4AZ8dlLkKLXBRBFN
u55PkG3i6ySvxeCdTX9g6Nn8K0M0JQQjegSyi07Sshf00GYPoj/F0ivX2xMeJe6k
`protect END_PROTECTED
