`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MdNV47Cvl7uGnIdvAI0MARbvMOcGa6Nj+RPNFpr9dYC5gNrhAqhaXGaLS0xoNdr4
2K6nwAUK7iIxrtYEqpZZj/JIhmf8auOmNg9zusvliDQVLcr+v4oPm6ABvkRfy07/
jJY42pTEM/1QeshyfvBIr69Ymix7Ulo95cddwAGNWG7A7ULAqDE+1XN5mDMzekjc
cFneTZaM5Ma7+Y4f/ROgpOYOilNU4w0uZfsqk5KFPbDCpHBx5IlgyRccMF3SNQ/U
szHYMesB9dXSR013S+3y+PpuhJD1LL+679327PXUFxL37KhRNlioQLUhs45bWPJC
H6QEEAc/T012L2jHNwdcHJZxbbiNsx4xxA67NA7DXcXLbnfSMl4AL2gQx1CzNo6l
tIinqk5lo4w/Xlcov6HL5A==
`protect END_PROTECTED
