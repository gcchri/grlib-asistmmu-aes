`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T4wv/6URVzHmNnuGetuP8bVAfeqjwE9CYUXkyO2/SlMEhFMyxTM1Lfiglg53SuGb
P50b7DYpysZ9roalApI5cXnTS3B+/6nJ7/GaWl9bOT7hlocKQn1BiueZox5sJilq
lGRzYYDsJMYpW71PuBUpbAczUrJKtdXHyXOp+LnqVlJKq+xhkZmFXB6tO591H0+p
CjByEcbOIjvlpgOmwmPN9jr/8IMVY2I3XaBnUgJ+KEzjYA7LHnXyDvPsMS6CNTNg
eSDdUo2ifMx6J1R8LA2pDUL6CMtcba7aK7mpmAXsQtFuqMlsWqdTsDo0cJ5hmm/m
Mrwf99UVcBTTtxlIcQ/+EwAIk7Vi662rC27R9jgqK08Y12lplfGhqxPeLM90HsO7
wkAlgaS+cVIsZ7v9vk9CrD45RbQ/24Usx/Db+n3cILANLrW4banOwmqNwAGm8TWM
Zr3m171fDPdE+WrBz5J7cYojFRVJHlFGlbmROZjRPAVZ2vX4nRIsSAcMzk85+qpS
U+brjEERQJ13nS8CIhZId0QiGxUGVp+PCoUyhIYVVsvB0lGWAsT+pnWxkmnYlGDj
b4YPDVmvg6yj9YpAxVJv8a4cQY1LviMz0szJ8TJY+3XvSET50QXZAGTAiNe7dn8Y
KOCM2k28jp+fQ9EELSHU47BYxnojTTu5Wf5kV6hO4lO9Vx/4UOgKyS7DYdKF8RES
YdYSezE33PCGcGGAr3J3tRmD5iGXWUshWcfsBqIfrvvWvtE3gTpWb2fjeyK3oCl0
f7oTKlXbm5d0PxgPfwQOwwHGOCV3jgHk5GpdPne+UKUZx/ltQEOEK9v5/cktA4kV
pxvcJlRgsPaygP4CwB/CEiQtXuQu2T2pRipAWGkD7OfJVqmoRxSaWPJCbJu4ESb5
6ntZvc58i1wh+m1Q6qpO1OpGUMkE6ItjKPSP1ndL8J2CMF4zmIAsI/cCGKUcFkmp
lTix3SM321exf55VCWoq6HQxK4wUouLAyi/HqF/m3ik/uR/P2U2QDPd0fmWnSmgi
ExJ86dZ/HVH7j5I1bnmGU0LlkuPgZ+UVm8isqBI/jGCNjroEbsBV1H1ARTMk2t7y
rEqUlMeVlPDgVEFXY2ftYAynDzh3eD5bwr9+nLf5UGfTGr4gPtFYx8Bv8/tklmBS
EHOukPpwWQi5PUzS+uZFanL230Nc/Gbk+c90ITCo6DKKD384hEBz6pkRKE3BXNHL
1mHAipAiab+z64d2153gnYgIgCA8gdhNtOEbxaGH9ITu8u6baSI8L0dCTRKeLn8q
3wVM/JZFm1OFNMNfaQeHJcjfGXBtbGRdYqCjm4c3IKTP5wt8InlpQRp/yT2w2GBQ
vb3wptHjxf2kOiqgOXeoxqPmZ1Xa7ZZqyCihVUdV8kwYrZ5TaIQT+hcTLDxc2BSF
xoOeUwDOl7sd8Vy1cqGWCieKmDllQlDvF5bNbNiJai0g6opgHfPer1OEmnzION8O
3z9NW4dSX6QJhXZbqhIoUaSmsFI4zb+aw1UFKBwqPCNQHyq3sDoqWvSPS7aXyDkV
uw5himkqVk4r2k/d9RBlsG8K0nwmG/X582Ek8bC3KgPh6yVs7KObWaAaj+NBdczZ
O7M/9rXKVBwYVJqArrlxfkC9Z9vKBhB91FINpFIU/04kxLA43jMovuxwBRzuhiOE
qpc+7a1C6jS505bvKkaNwfpI9V3bT+F4w6lfOHD6q8Fbd3eqTyEf9WCcQOyxHBl8
pUPTd4IvfElL5N32WHBBMOXQvt5CrXgS6tLBnNdoFk/eiAwp2cBCT1BWbkVC2DUD
jWIKsUVH+yTGbH2RwWJr8IJ5TDl+URkcKDXzTJJCWGSOOrhdyliAyHWlCzoiEsXS
WPN/lJBftijAZEToN9qUJEWlCpBkT0CPQBiF5ji86rRWxvQonRxmij0Gwfk6aYd0
8J5WF972Vu7aKzTnxqDBaIC1fquUXofUF4MFXdDygZooPG2n/mVTwrV1MzC+9stg
gMEmutcyEOTqCVwcINe0Xc6xFLF5Fo7GezDINMlP+CmVVog0y0NXiuSB2pFpS8DQ
UYZx9lJPLYkfNk6Rn6BXn8BPwsh+59UBuuCVUAhS5hexK7Lr0h86uZgbH/5wMcnG
Po5T/aKdiViA5yHc7vWPSTWvN2jVNsE5xLduH4jyTy8ZpjXlWrBINAOiKK0ICO80
3Ffn4xx8STipNZMQ+2Dl0rP849rMY3LHGhUlllsVOJHwBD7zHw9flnUy85hD9cpq
ZB+DPsw1Z6aF5zuPmuYtx8emOEUTuQcDJVdD9737Nj1JncytYegnLfQI+UtCB9YG
0UbQWBIl33A0lzosnTypT6Lnd4xzHura6+byqxGMVICIh+cs3RGQzZJds5SJx6l6
N3JcBrdmre622pjuqUW6SyZZs+2RwUZUD4mMf/CH/H/uOEA3glVc+JbZPmewuo8L
ss6fVexN73UJTkBpqb7/5kMJSHOvvtKqTLwteVfyc6OceVQ61vSR/YngujtcKw2+
TgZLhTudkDj3a0XR3ZP7tNG/tm8DeS2b0Ikmj6ZKw1qgYZAphwXCJT71i26LKd/F
wHYuRf6qfI21EtoqxA8y3c7cNgdHQRn2FA2UtvTFoxULyUO0uIPqXP8hzIqWOdEC
TLWCkYWXnSknD73JSvTUPdXMDUdTpubueobJsqQoFPzXPwyBuZ8QijJqNGxOUu4Y
hXfATNyVAAMpxa8xScFHdjfaHYvKFLNmxKJnOvUgAC9epQ7nXGDrR7D7yw/6eQhe
iIVVv6BQjLZatFb8EUQYawEHLxspSfl/Rtc/Egx1IjalbW/MBiBAfTsnY3drKfob
DBqMGFb4B9RcHnQhjv9vEIzjcVxbg3ZDAEXMB1+pTMhKEWKIH1vTwqJ/JJKzvi5a
F8AS4yv4An9pc3c0M2N7TdKqbLYMsS6i5pjVbCm5PU9eBR0mHKwuoLaE0/4DPxLj
fODBRIJq791V9Cxj+pG9eOhZj3AFt7L+wn96gkJx7RKleCqG+lMNUKq2Kq2XUp4D
LTPnINnLrDwr0JgU0BkKZy5z6qD5Us3w11/eOxlQPkAJqkFmDUYSQD5/hZ2rNlvv
V6TdRsHNczQ+nhlbMOG6XLKHB4FfGtm/QWAgHHUbHbnw3yJPmbnHC76F8Ncte5xX
YBxfhAGTW7cVXlgAdXJXAOwnZos4IrEQkw92T5do8JrI4b5e+WeXa8jeZ9NaaQ0j
TflMizSfMYPHOsjF0d4MAvrf+FIoYsmFp36tV6u+qh0KtlO7iWas3Tdk+jxMlwIu
ZJgGlYEiuW601itqHJutfi8bPlYU4YYvH/hO+DrtCaRdbEGSHJ/5XxZHA4EnMrSZ
rWSyjo82QK/UIDYRuwI3pqb28/SP5imMvueyvvo0lka/kpS3i6+rE38gxEyeXkxh
M4UnSIAHMiW2iky/yReyWyJcPVZgOVZi+n6dK/0izcQu7NC+P6eY6MuPArAq0KMS
CmKmyBgFpMuVtNbnwUxY5sge8cYnS3GACarb4iB9lBU1/tvZ5ZPVgg0Iv6NomBNF
oOXCeIfRVufUqxcTxnSlUqICEoKZTR1hrlQo/OtpxU7P6gMKCUnhWX3Iy7uWag7G
magFsq6e/fDGvpWhGazqVRRhOqx3nmKOn2eQyF/aczL5wEe/GmAKfwx3D584pWoW
kUubcOU9l/H59SIh1iGQD3PnjV02PaEzEuyh2x1M3j5uBjvoKcroFVVEpPVKF0fM
cyt572FKTyUu8vAtgYbXdwuqiILVmtiKh2Zq4FnFWfW58fp4BcsAgEdVuOzwUOsu
vjttNuzaqW4DV5OvGWEbg+eit6uzxWJpmXcNVN5xJu1hE+crTFCv5cxrraOLzPAv
w0QX2qI/DIx3Psm0xnQqvcEHeCynfPQPXyJTi2HQ0VXNKoXQDiVzRr9FO9VnfhOb
VULTnhGIpDly7Ghqa2JObYyif4B79VWYKeIwcuNvT8Q2yoB60rmtf2BNSLzn2xUN
qTcfWnU6zmL/D8MThM0daI5eoEedFShS2qkmtun+N3MZyTMGw3hVk7eI48Nt/AoA
wXpmUTbQyAWAlQv8pblM6OVaRvr+UsuNskX+E47WtMoafWHuricHULmQ4m5dxk9T
nyqHWA1VA9DB75AH0GIv1DpAS2CL8ogoWGjHrpf+9kzIrXD6NvU/kv/yq27CVfmC
gLlTtiMaZITN2/zluXaWZdBWyvzyie5XzrQEjvqqDjaIy4PuKDGTBgVv5wb4hR5C
B6B3UNGbRrqS/o4hTb2fS7fPjE3k+BClxQ3t2dcC9qiB9Ba6OyuJmiXH9QHlM2Bf
76eln3RJAxebaFgr4Ty6DiG3tBr8BLVJbZTy+yMPTBzhac6AZ5IYew3sPCOLTRuQ
nUmTlH7db5wvVM+e5QEm6z7TceCURmbI4cv8yX8vnQyF0kUdOQiRwffU4s6WXdNj
XxjTIvdQcv1oS9qGrgXmU2p4FXJBmipwGebTmwWhGmgEl7oT7XTjEqzMOBS6rqcw
U/je7dUhNz0EJakmBOG54LFOnqZq5MAp9tY63ukEsJJ5xbteNqvCLBsFJkcSmuNb
1D8RzOrikQ+MT9Vqhdm9crPe4nS6ZZXvNCdhqsBBknK/bCbvI5M5YVN4yUgAHyn4
l0RKQusbwjZjhNb3fnMYblxZ955vLfzwrHBM7Rzgzno+dQ3JwnBYDvi8DQkeQvCd
a+UZdPe/6aDRzq732Tq0IcxigkUoVcWcbqLsETxP305A8my2ZZckgE5R1QIelWKh
EqusvqzTJjoC/9b85rVcEh3iNT/RNjST25zNZVVXshIspl6qWZPFK9aDZKbQhkHm
S/9uT2BcHluFxyDbw5r005D8Hlx6y6Z9E3n4yMNSVoebr0Pb0GwT4FQN2EzCS6n+
pmYmANt9nLN2xUjCCc4Jz/DlNGZPFXrbvTVTa3qhId5QdnQ+dJjTAAoJJweV1m45
3lxUODDJnh/X5p4/K5pMCND0T0TbKPtnzb08uLu0C7azig/eKZHUabSisqCaLPaR
NN28jaQsFZDZXUs70wJe4LA1Ene9I5zg7851H4hx1Ux/8wmA2T2NrcWL7TwI0eaI
JeeO5wN41+5GzspWUwM+AHKjcpiHejPu0a6TA0fMYL7wGlVk8hUpz4zrRPwo65OB
w3R2ro13l/4YzqBjvkLhqkNFF83yBwE7MozQNEZS0yf/gYOE6YjipOJCocsjE5OZ
QVZTXVio7/rmiE2d2NO7JUWV2hoOYdluCtu9/mfy7DL4grxFv6j5dD748zvyF+Wi
Wt9YKvn7i9ih2zu+t/+Csbfpscfv41ukDaela+wEC7KEVgCsMGU/bfnZLTnU5Ly3
a0gyvGmyHvbpgFiBaeiidlrqaxb2/ycohUuJg0QwU9GSRjVMXruay8GTca9SYU6F
Nsdc7WKpfB+oR+3f3KUbOA4se99V13pmLy0DdLC4wOZU4Eke2d/Sf+QLj+m47WXz
6FfixC0TrSxKBJok0T7xVJSQbvpmY8sKYp+dkeEZjP8zm3SC1s8kDov2dV5JS8wO
HPL8kJeFzHxHg2ZcIafGui6Cq1xWRf4fNYSUWts4hDfNdznUGUZjykO22lv6WkgN
CbpGUMLI+f94aNcoAzMHk0EVFiZ2NzSWaUVFq53znDPu6f7YVuTaOce/ZgXa0qnp
YFSYczD+Tox43InZ0jkYxguw44rRwOIN8jKFM1VpHEDla0DdNYQdsWiCtJe+giyP
apAXbJEjH7hpQdYDKicmuGJEMD18SxR9QvfJ4bFBYwkPLpwSF4RnVA70lRMboy0j
Q/XpoJmnj0mE/MTpfhfLgSgWP4J5WyO9Vbvk3r2Jt3KxexVYrCJzyUZH3RJfUAeF
j1of0n7QTVAtuYV3HKSU2TRviw6PXhiqykouqEimbp6A4DJqlOVRPlrvv0CbptdM
mBb7yqQmM/ypiC/Dl5XzbdFJvL+8E8Rqe/DalYTnMnpJaWn8/C46PdXemu9IjUus
DtyYUxcuSjpiY4jTc5X6ewrOxk7eHGksRH0gHoLrMf+nUyw+DMvX4j/ZGNw+dKmU
eBG/mu1cPVIVrDD2FegXseW2X0YriU9Ues8Meo6BMUnJBmABT0ClvPD4lmkHxiMP
9TcUFofLspra3HYY6BmWHwusHpe2/QeSYpXruOvpWEVwN8+xaO0G6SCEDcw/f/Fu
59wbK30lHS0IeukruVz+SyrhOWmUEuo3fKbeBXk/+OoBxp6ALAibdqYiyGEgkn3u
FXqq6+iFp4WAX49EMtClXb5eBZT/XNn3D1pCkEt3w643JYr2BhTg1kAlDuz2Bw1Y
N0SXAa+zFXCbFbbxltpg9jc4nuUwKbF7BtVKmx1iYPxNLRPQlJkvfpD5ChjaFfp8
Wm4jDNzoTJUDufXvCJpr/ZsH81dadwkdUZWbRGBn8jWPUGEOmabW0/AomFqa5TtY
bJrWlW0Nx4zIE1W9sIdylrQWrGxLdnLXqM77LDkt8EGihkpV3i9a1sw02x1gY7qH
ptU0f7KT0++A0vcaJrtVxbLWYNk9js62fhcarJPCu9k/2jidfMP7Mhm6VoYdkYfv
33fwNv866ooyOK6HE0lSUJpDy+aPjOD8RpzC1qUtwt7L5ff3T4y3n33709xm2EYr
aOKHFTnKFdkR3BRB4ggzxRqw2lVAmEJ+m/4ka9uVDV3Xcf4NWNXhDaBNv9Jz6s2p
tdb6o+/Uips0xjnN3lNFiVo+gwk95JnrZn2LYfYM+G/IP7WdIfJwekGas58j6XLO
cLr2s1dFMgJQ9CnC85Xnz/OlrDRxcS+BMirshSuDWZ7hwZ84MP73PZsjsp+CUsLU
zfFSicvJrVUidJBq/230+TEhCXc/DtViuZFzHjktqYVI/otle3+ahp/H1Qj/VAZl
HLs9GSB5Y+JPChaBgorsyqmr3n3YcDLteoIx2qfcWmGjuFinER894CBUmh4zvAg4
yBtLmzyn/ThDFukiD/yKI/6J2xVCoJ6a+cqyuImkEpcbx6kA509VAY2iGWOBUFT1
xNT+NLpsK4KEq04zChiLYvvHXHSys0zp+DZRK1EAA28t4EUOoX0MYJkjx+3AVuk2
QjQy7wOXr0CjQpvPw+EVhvb/NsutuO/JFZaLAY0NWRwqVrglq2oKXM2jYuNglgH7
kT8MKWhiJK3D9aaz7+9rCOHT17iwwmkAC1RdfKkNrOcYGHL30qrRZ+RzCJxhWeKn
Idp5gxyL7mBeVFI4/gp3DuvCt2YC7ykYFbxNIGfWiLmdZ5JW+62tl704k4TlM4bK
jxu7bwccFDUEmLCNsF+9w0F8IFuKf2G4Ed8+SMX2O5Ppe46MESe5XvpgA2rLck63
qu5lfNxiAxK9suU+o5R6ZXqbn0bUame30zPm/iWz+gqtULIBn9Qu8gGHMcD2KH7E
cPB+4FnbsrILrUraj8pjLU5zBQxjs7FBFY29/DLiStHyvg7kFGZJXs7F+E9GfQ3v
BmC3wriGX3o0v4G0fAhv4TxsrBV/9tZ6r/ImfTBUJcwyNQcIeOO48oyuzRRwDPSO
P/CfcHnVojwKq/m9t3xBNjsxUmMp+FkPHU1Bo7ojSp1KqWvsCq4kQQ2O6cC6eOSf
gGxZMniw787ZgE+ZeT0n/vYPEIWArJ6FwUbOO8VnzoHuBTPXzk/DaRpCSru4nrZP
6cD2xOiMIuXL8c9YbxEhh/a3iXtcUt6mBx+G5Hv0VxwQBQqGcwUnfYkhr7f3mjZV
TE1cHIPcjOng6C8KKl+Yy07wsibnCJU7JIlsR+mCsfYyFxk+EyS9Efpksb27riXQ
NReojNEDOcub8ln0KN/jsb1HYQmtyBRxnwPAmLlm4hSKkNls+rqjtxmqoxayCa4s
c205+GgCitpSyxXdT8pioXOiTy/PVHTPuYFIwM6JNm+bmpSzYs7yMpGAq9hyGVo9
E8e0hm99vmGBwWap9bUzzCKDEyAfwhblTBQ0WKu8BMeFTKpQYzSUnOVN+//ytR1u
iq4+pbrhFWV2KpR5SUmsXqdnFtYcNe5wVJYznc0VOcXnQN6EBEKcyZHkrgtdlaYL
JvVkznHZXSuWXPSxGE6k4wXjce3drbff0xEsnhS3NM6NGCTT3PTOt8lXT3tCtdBt
yF/j/WlOSG5ZYlkHvTfEFEhW9EXiGuFZdLK24EF62NyoyJ4KnKFpCE9Y3/aQJcZM
PiDZPg0wN0/TvfplQ2HM9teP4QvayLM9rclMFnC7ILp3ug2lgGzljf4Gww3RUznc
7/DFhe76W1jOoap5TIDAwi36LG3uwC7btXFlqTIOpOSIyCSnDAEZwBgFxCSMQaDJ
kz2s9OH3kZSEK7ayFNbXwkoWL3ajattF8Zt4F3fqeqR0lYP7VKZ3WJ2SOH3Feg13
MryPq3n1uq9n+yUDx+eUc3kLfrvBvtxuo/SRZ0Q3IYKM+Qh0IhWTGraBNiIZCgEd
skXva7X97Ob6Edxo5GpVtCejklt2Ybvet0dOIyiRkFa4FFM/giKq4LR8/jgtnLud
4xtjs+/OvtRbSOvfJ2ZMX8tDVyY9bbjzCyc3yBwA6r98JfVRs1qaXTSF++3KJraM
Bn/hs8E7IyipmKIdEL+6jWdebfGIqiY17gi5gXTH390LFri5QfEVDy3zsCOgLiq0
T9It7Omclc5MTl6M+Cvs115vX8xCEAuT2ihomdutw33vczY2D16PeYWAxcBUnini
sMNebSAeO1ijI9eJEpFsu5RQWvoxYnYL0GJQ5yJCBSg2jBxBOXvIlRb7LnVyRNmb
DtCkl+mJlfr6LQW762rYf9i1vNYyVBSOoCa99gUNxko00s/JcT+k9ade5CLWDvK/
mBxeNkUUurZ9Jo3rXD5kxsxc2QPnHoX/bC98eU0WVXnyQOZvr+SNgXT9WsW96a42
pUSxz4hfCGQwQIgxWxrrv9DdmnBf/cvMRnHI9K4HNsGSp0BdWqz0npjo22Dav2Uq
Dp0Xezn0PBNPRqe/SuBivBprtOzbu2Mbe8umo2iPP9bAQQuZ+gabiaMcC0ptbI//
1ClMlBGriAZ3Wnux9xFWeNupenSKuS0BJWY1fVBisyte9W0C4pcOq/2H4rirg5q3
mJG7Sm8DS5aHRJxQF2jABDgZolY+AVH3wRo9TNDDTzZz+eGfD6p7OFKwg6gVsiRc
jsM04woFvTUefWu0+FtKgUmg7yo2C/LO+Bm1DAbdQK+K68xYssBGVmcYtaOVWFc0
yoYGWpX2Z/LmR0YtEwVYzfCmc4fWoFYdyAZlg3ffvu10ASB42KH7uExYn6MJ0KyW
o4BhoX+C5dVb6UWt8W47XIlh2AszXNrn6LE7VWWK3hzBoyWPhWjKkJkQ9mkxu7OI
ZV+m0fcS1nLajJjtHW+d6esBmrZlS5WF7/pf5dLFI0xegihuwJUf+OHtFl8ZasuG
0v21y8gBSST2+ZCCjFx7Vkn9f9+HB7DVZG9p/RIdwe8bKWY8NrBN2cSZECwvv1Nm
+07hpM8aJXxWDR1wKr2wvgq2Ew4iiPhrntniCb++gyUpUDHoNTZ/xpLebVT5ACVI
aiX2wlaKc49TBeaJfAUhCLmbZVmJ6VP6zrHGSiUl1fC1ZxZex+BGCCERPqmVz7zA
yloAEdADiJNXrHDyUspIieKVrciE5GjQHEq0klvOH15jFje60T326QlpgIfrAaKa
bILYZqZX6i+wvi1xBdvsKOTr0IgxCNDkdv+si1gaFm1U0+hCTSogmM89rrqbHlo0
FQ7O2Da8IRID6bj7+0rUUKo+R2MVwdhYObce69VExABnCHrKiBmGx8hu8mkqyBHa
wmUby1HSfOSFseOex982EUPpjDxDRyiy15uCSHN5bu/qURKE6CDwjbGUwcIaCTE1
7bnUyHX6e2oRYjqXHbS83dirWTw8JhcgDlUtnz4nuTuqWePJ+wmHZe/dBJBleaXB
dAKkxJ746jzuvcplAa/MO/2tWrjlbgY36r6sLYPQ24jS8wm5VTfkRzYAp40jYkH5
dHuZcpaGP4PVHbDJfZU6u4qOs/AppjzXgL7+fzSiE11gjLdtSwUlNSwYqM6E5dYt
CV+3Gk8cn6LtPsY1t6te1s6ngWX+AogffOg9LC2YS6C0YblX4CjSo69f3KX+4aOL
Yto9VfkuMkdilVflr6nlkLQokIkJ8IMWaKtUHlD4noWlzptZVVTFGU3HclmJpf+D
lGcC6bOP06VBmtX4AjeYkK8lHwSpYkOHKksa8EhjtDPKQgY40wENHs5s1IsgbPMg
pYtl7R7n3Dsvoy72qAGMfzvpitxtf5EnhXE0DlyNIzmjHk5TqHx4po3eU5IUBK2u
FnVU0OhAOiP6Q20tu/UqdF7yNPQPQzYcMMi/bvWYuL0oWZU+OiEx7NwVwzMfD1Kk
GWxhzdDNPJHeA2NvIA/fhU36naipTEsQXNNOmSh2ThuLd6cxiNQcAKnEl3zuC6Ux
2+fkacfgpfxFxYQlyoiqcdC6S5FIf4ejt8OLobCzIZ2ylxp33XyD1v1DkWpcTDDi
EQFKXtSNENMeHf6P5zsyiZAReCDMNPRTsZ5ZD4Wn5opPi6bbNWhy2ClLdwoeW3Y3
wN0nS0lT51RZ4weRRxuwfT/EUA0NVbo0Xvy+8MWyKUMbZV27Fz8SBlu1jy3Nr4XO
K41z/OtkqeBxq8i1bTzlDy+8nirF76p8ZXezQyujBMjpAfRtLS8NejKSNjoMy3qj
R/I5uuoZj4u+nzptRu1I/CE0o6n4kmdg5O7yYHggQbVIhDwo++wfoOy1E0gEEZ+3
MkbZB9wE25eGJCjrMGtY8Y/AuxcKZRZ5ySr/KRV9XkkloX62W19NeCeA+tvTV7q/
G7ogNuOUt4V55gLoW89e/M/30q7LrQZyGaE5syJJyH3tqA+uspPpmmodcUV+ZwTe
NTSOAcUpAy+Oyx6yLyJ7DAnVe7zdFWhbZfzhN91D6UvxFo5+pDxe0SlJJJwRXYeh
BfdLKAa4lFqzC169eon0Q/gvq/7BwGsQOXfyMmHG9tdwF2IBkiJ64brI9UfHFcPT
5tyzU/flUGyacTHLOQhERQ1x8YtP4J3WFpJsI8ltxtGSqjNJijHIYpXiifkWEUzp
fP7ZE2RbeCRH4HVBWx2hiIBDWcydIfhgbuPGHal4X/JwVxkEPeVTFw13D+ovZsrc
sBhfY66g9T6Rsx8HfMQuded4vvLqMzP1OKaC39aTGPkvR/oRf3N/7XQbSrt7eXUX
M3WCk0siseW/vpyloV7ynk/xGqAePe3NMiyY/YgJW7UKtCSZari5nJHmK+Uz2Q2/
D0tik/a12ZDYP46ERPumhUvIcQmTD6nhO865g8Pi347DCChfEA9LkhTi4hEJCT0n
QGqXUd6wBSnGj6gzDLXdPnI++ZAkQKll5UZ4BqZAFek5ilTH+8qD1cE5pSfcw0LK
YhfQdtDB9hKVlbDCH3zDr5VZjUYpbKg0/2iESVa1zwWBjkjNakfHIlTGWQn2p/lB
m7kHjACWFUjCJXUDz1UvfnCkJym0baemgeBR5wG8o+E4NGnf0nHaiobP6yiqjZwQ
SU3Yz0Zv0njycIWvNn8TsV9RT+5BLex+Jg1H5Fg6vfm0sR6czAeyywlLLcK7mts/
Hda1onqsPof/fPtB3XFxnrseI0cg4obmVuA2VHCkwoWTJvqBRI85ozUPdoLILSOq
kKnoBYvMAXkWNxQTG1stSdsg/BFmyYo1mSMdqK5+ynfTVt/BcJMjINkx7xxh8gAw
1l4GlSuDkTjnj/nEA8Q0pM3Y/9pJUQlQ1BPAc+iGD2DVS7DZB3veTDZ2lEM9/7sc
8WicZEQAM8yWUw0KLR6AlXZ8G6KTPuJgT8GR4XMOe0W1m5ZfIpGK7sUWjPyyfwoK
gBGqBXbEgyObJLpQoUU1Q5Pt884PvsFbei+qzzFG+ZUBOQLo32tng+yKPjB0di2v
6Gv0QB4XBpWUS86zpzNA/av46HbEM+OYsz9eDv5qYjckAfBDQ5AB8oV5rk+ory6W
9n5apbW2Hhb8c5MOU5sIli9TLjGbyknVvtsXQ3XwiD5uunhE2/sIRo7B+Y82fjzZ
HqYBPSpxaYPQhNyVgKyKVN2PZ2tCKxYXuc7NyqywzdRdMxLKhXWGZdee7NB1POHb
r++ymXnB7/rEdAqmjhd8/+cAduvQ8lBcsOuIHPobaWR8BrSxXalaMw2QzoL36OMz
z9TMXZmz5YhPbJP4PUUkmJD8d9pHUeVxYVISD/bheW1Ed/Zj/gaQrKRDaKJ8blbg
dw8u05LlXXghkjR8EbGe0dWZpkpYO+jZytUi7s0dzPmEiZ9AMIIkeQ3fOpARXaLT
TIfVnAFNzJO6daRMNjkQ4pydjtg9kpZm/MIUCJZaoaJv4riiQ4ycG5FWkHjbOdIk
oo1uTWWdFq6HVjc/h54qV+1eShAtZYSGlpfA5R4lrPX8U+zOE+6YoHtf+I5YMdwU
N+z97NQ5/yVjCfBWE0b4ZShhNfRana0bp0c3WN5UseFgRUQCwbemb5E/v8Qvk34+
iHM+51FK6fxQYztlC1/QcihS+9Fe7JhyWNP/kB+NbUoZWUeTS8pdc0fK8+6UXIaP
F0U/cuUeDM+cBRwiGAc8OaRSHZNSinPF0IP7+huqEo1Uqwd8RtYJpo95F68eIPrL
hYP8WT8tE+uUA0cn3zB9L0SDJJqelTdIRzGa9tC1UHJX5HX1tUFWuYCLqRfAAOID
Sb2khxHTraqbaBUYFXHcILR627uoE3TOD0FvlsSdcGvcyyktRpIWURTTaRr7qKo+
Q8JQAvJqtqlZYjwigqiTRNI30418A/Df3MBYD+uD9wklFgnovc0zokgDFsOJtnm/
mcr5lpYmX8+BGV92KbYE35R5+7tp9aewz+IoMrb8pGaSTszOOgUN6E662T8KASp0
xeYRlyxfJJ1ROKXYEFDNvtejdTkr1BNvv02ZBUu9vvZ122cV/AV9TODbGwf3exZG
DrPZegrhQ+L+9OoFP8EoJQYRLFx++7URCC2Vioup897RYHPpWGMCjz8ZH3OT7nos
3L6rCuh4EAGzTbpSB9RqaskZPNKmXYoiI9RQRVMDeSiGIPlpXwZF3Bzm6TlqVrv+
khjbLIQbMBfRdphRVySOfs9kxOBAgDAv82ZHApUIC/c4+cIFhSj7UsUkHcjlllok
by73Q7Kjn7QOMnIAZzEeX6P6TClPHScQbGtM2lFcC3Lk3wDJLB66od8iT8luH74l
E270Cgy9HE25lWVfkcO73ykpNYZNet6ApxdmKxFmChp5/XfV6rGooGbqbcDTYW2G
+O0QOsfHkAjjkHKfFzjtb77PpMHSZJfbGEY96SK0bHZQtayR6MBC41XdA/GRV/YR
l8bQhP2C8QWQCTMad7wwtrGcjLwchjyMh85U6INuw3wBHdNziRbI644/G9jN4j5P
ZP9CKU32GBqekjl9X3eM/Vjz1QNGgieSOLTq7Uch4ZixzTjWoQ+rb6zij3r6qMJv
gN+RdX84S5iO63BAGDqneYZkqzoG4xXLYBFWqHrCJ7V4J4AdmNcigA8sgoiLtVYK
VI2XLcwOCTM81Z9mtPmtw1LGfw532hUmeLAtmOtXxZ80+ZC7wFH2jyETI7OamPHs
xsc6xWzEHtzDF3Id3xYEATokSj8mE+VVzx0t4ahYqCCboMLO7hYN3LBqgQCfj9Qv
42m5w3pMirVlL9RLAT96n7aTh5saY+FIuq3yClYyL/5RQYKzZ4n6wo7VYQ3KNUIt
o8zB0jUdKg3SHniFqMvZ6bOsQuws1zMAEq/NjGtizeYVUuCLEp2EINx0bux51pbG
Md9GkHRVSw7OEMddO/gE8Hv6v5PhG6xIOCMbBlJPejis8XHZuxXUAnYcMsspViC0
DQ2HDqcOJc/lUY7daiKqkPJIg/czepxVdd/iGg1mxvVvgc60trSb6Oa5+cWmzwXu
Ec43Axqzt4UwcgREB04poS1nOGQKIdDoKOhKs4ho/eZbxIfxnRCPT9IQ7BFLXlim
lt+DbWve+vqcnM2Ri4JFnOmMP1CnexlGLGMDvzE3itEEWWZf1Bo1Gq57vehmS6Xc
nVY9Dg7wu2cdJ7vjKfydc6MGtK5Zt7BdRnI/UwnFR2AI2PK4LRGUR1gEIHixGyQJ
2ioYFwP4pmQu4HlF2bpmba/LJFmYCaQ62brN7GIByc9t75K0N8Ocm9hTOzy2qaFH
dWTe3vsO4lw9/Mo+d/LCf44fQG5w2CIA7ts8r6ZcwD7/5JwtZ3319VdSRKx+6iDo
au+1GQeIB+80wQTAIQgK2VDDNcNhgARYMRplWKDPVIpPWgmJpIS9ckrhm3kXk/oN
lQK5tFy1+D11aSpnDOX9Ci7GWO359OELotxZr/LaobuApRQ9BZSOFhmECqmZGTre
6eEAFxwgR4DoaLcPlQiQZhzOMLIMMayyeNl8VFsDFCrOEs/TEp24UfntpB+YQBel
R+AvIOG2YAbOM7wcjPHNW24CxUuWavE2ahdHUPRxuBI6Tzn1LIZ/NevXDP7JDZf/
u/lJ6OnKgk1xnC/y8W87IT7Pgoufi/7mm+kS4Wqnj+Gj/JdY3ZNU6/1MQsuUxD27
DE8/lZO3zuIcMTHGHX2caR02rT7K1wma7Xr9pi+Vu0dPqJD6KNoJNL4EBelPFs/9
T4gmiBvAnXFDcpE5nmNXexJ7XPd9BPWBahFuKfXHp/k3Kqlz1XjbKkif3SsnwLC7
nGGpRc1VKl4KpX+I8MsLfNtdg+8PZMHCNi6emDDAaZkeMhJYXGRbczCf4F5evSKt
oDdUhC/6X5aMs2P3NoLAUcJZGGjcwg/CbdZ66yAcoxW+MUiDDZvvLiAbTsGcQ6EE
CPGUY0mBa2LH58c9qZEYkkoidePyxR7duLKzXDkg6Mr75q4MQYWguK6tvYXScdWG
Uf8abOSH2PTX42PtIWGc6SrP4UTLNJINSWvWZ4pvZFBoAVAl1/dpd1tuyBXYpCLb
JueXBYrMp3IcF0GOZ0XuDeurecseSmdEKDLdQT14qtLQlB3cemrLegLxqOJ1OkOx
UjLilTlOQpbGHkNzksdrYXvLHbMrzmzj04lTgLDxmwD7Lc1azykoIkHbuq8WAbZy
5ZzKlH7HqoWNp6D13/ZMgPaaYwjB98dr0eTZ1tJwzY7jI4nSFvwS6G//tlXd4HAt
pkwZAQ8XM7fRxy2kCbMDIXg/GlyM3G+k3bDWzaBA5Bs96hHbKOrFt9gPtwUNsYf6
iFMDPeBeC+7aDbRxBc1+nV78zINgZIkVYly4fxNW8zF/qk5DF5tSxatsMxvvknWM
BKNptSh3jNUbZGpn0HX+irxjTlpUd4bJwB+OBaErLNNiy4wpA54+CuhLWDZYSE3C
R/IeFIC/Vwi+BCepU0gmbizOb4BXMxLZ5IU5/45esHpl9dGh1ZQEl2uI6YG2OdAU
PspQ/yWVJhuQQ3Z/iv1+UVhTFIiPQkIkqflG+WM6gsh8A2XWiahtxmHaOZxcB1ro
MAB4PP22cOXwrL8qfBdxpUtXIbpGycozwTVpD9F4DtTAg/77nDCWf+09DGSl7RyC
qCVrkPiDp+84EXky9WWyMXvbfqVKL51cxSEo9De1MDkuaRgycm44wNGwLUvuQbvT
RVApKbkcZl1AmP43pdtX2H20lIHdqW4/902joe/W9CjH3HHsXjuW48Lx5fW2DtBD
1xJAffWhJbC20zWSn/tCn1Pp/XPMRffMjnNhEKMsiqhFrEAtisaC31NZj53P+7gQ
se3cvWzpN5aO9ungEMNx2FcMTMxaDBPpaP6Aj9HnHkEoIBcIg0eIrT3Sut7QelB7
Nun3O/0lOkmg6+ZnwD86XFaW/KITf7EbLQB7Fnh+zqmyNlJZ0PZbo3MnXYQMPJlI
vUz/LQDyOVQLy2asYSa66hWdAAZCMVutiSaQ8sS2TcW80fRdndv2gDDo+kd38Aki
KR8Mc25BaFfZ/bG2oRFI6PgLssNV16CqCQ8/+HNb5PMe9WOpb/TagFb3A8kHxSqK
xrSxDgdd/9cQCUR54D0kec4MJeUsRIXEkP7yIsugaFILxoKEi3RZ5Rx1vyxJzoF2
Mh81ZOUFKKhEYPH6qz3BqN+367bKWNnHsJ4z1XWvf5QQrBoD2fKDgOeQV1TTx+Ub
X7gS6XUQdlbnz/3VPhmu2cPNlLVihAAkREA8Aw5c5IAzlfv5yRLDjCLzZs3fhc07
npoIkK+DMffJu5+aL2gKlcdcv5Pe0tC+A5uUZZDK+IYFvPp7OheJPIrp0XbxUan1
5C8ifujJlLkcP8ONdehlL/7Q+fwvnFnCFDIARnbpkcTgURMeof4mo05B9gHHO/7F
mump/BlzY0UyUXWsOQ9VFcKnvYtdqDreLC8rIMSy0X837GN/CwMQQ8EHv/xqCXKO
tFuhpklJipFmtbEX3ZGxoHAdNC/3i1QfAxsIel0KEQ+6mk+iR+vLJ58t/UvLjGgQ
7YomNcLPC7uBK+BGauPHVzxWUCR/2C8hYrDibLWKLh+/k1Ga7NsNMrFEOcJ3rT2u
Ly4OadH94goQpXYsMd15eQb8nZOWIh9MGI1UJiETGm8HRS6ivaS9j0N7PkrA7kEC
AIS4HXpzTzrxHA7hQczFJg8A40uSxfYGMz5mJTLwNSwi5k+btDT6M+VYTn3SJ2e8
u1+P0yxFheSSiACq6cFK2VA7W1VgaECtWxDokfHi7sIY5Oxu8mpqCp74yz1USCsU
eFvRcc4vSDqGmiy1wTIJLDWuFFDo002oOsAo2JRfWP8QDtdvfXdxSrNwe+a2Zl6S
YsYpnNcu1GXSMSKwmQf3k/Z6Bsk9nw4jybfpNQZo1Vltac8XjBqpokhy5SO2MxHK
AEvsdiX8iy8mWRAGp8Tclh/2bYfMzSWeHDH34PVN5Ma5OrI0/1szdlOigAPxv4ah
mQXCi+gSVcW8hByFX4GrEwvB9OEzRHHeNP6S3sUTP0sg5qaSxr7PgMfBuE9Rn6sw
7hB/U1/6sr1BZNrXQZCvVWRrqkGKEy4vX3IUvc97l3sK1l4hkl8qOGVZvqNaMCIG
sldxFh8+Fnq7dc0MdGkhX5yOjDVT45P0AqD/ALrWA9S7XU1Du/s5LWVY9VYZVCy9
Ec4VmUb9leGviFjHlu0AJsZadSJvm9bPu9OdeqR/TT1rMN0GiNsQ/PwpOsDUiqyL
j0qF91bqGijvOuQRSYZ0GOPZqGZ/wA0j0vsVpy4ynb+k3QKIb49UqoKg+B/y0g8D
VTRsxuhIaWO6AKH4CqIUOhgVo0e+Ralrw0ny0TFLkDlTBRh1bXeJThK5WPfITvXa
ZW67dhxrvkxyb/yRT6D8UNfQKGFgs8Y5lpBCxRzUVLo4ht8CRKid6MD2xjiKJsan
YoLLusUqqBmttMEmFzizUCfm5x6+cQ6M6V2bYUjydYIT+M22yrb5ASvuHtb9dBWt
d+DhmD2fy1m9NEj/FQqRE9cbbTpdxzafAk9DkyZW0F1H4E5nPZkA8ygfOANuQW2a
tb2yfZ9KqvoBYNl4hiBuzjmgKgvNf+stZ5xnO0agAr4oGWdy2e51PTOUT8T6vA0p
rYnAMVG6aFbttjIYCrxbipQ5nrWVY1LsMa6j8J5gDqM0KqQPMQBdb3FFbQqM9K0m
7Xbuqq8yIKhzvh14irHMWqxI0XhVf7DRisZV48GYiJH5W8DzFI3AlfheWqvaMUBR
a5hPshRFH4b7afKUv1zH6UYec9eFdj0Pp9pnQ3hOGqfoFnvaSivvbEav8IYi7xyn
6tikVt6qMg9Q5AkAa9a9I5dlXgEgZv98hguwTjRLnyFiLJel8FaXz3Q1fVpP2PA8
vvzvyGP/Atnk/sFAliNoGVcTZ1z3KPAHSUv9H3fd4CXxiFBj12UnQQDwt9KsE9zc
ZcS6CQvcO1s8FQh1qJA84hZJrIpFAwmV/EeEdni3foI2czw0DKZVarqg6ZsCmP0q
613LP2SRcEgWbpL9gHyV/g7YzLcnrCI7fQu5ZaIWX1ubXwkl8H+mq+ZT1d0eNwbw
gKvqvv+VwtQoK9Zjhh3jnSZw1/jrw2B7gwEw7fFAqs5cDphoLUZ06GjEFX8qqA5r
H7sYebOc63cBbMsL7POp8iY+WAVqakuPN/mRDDUTMWSxGgmleaeMpmKr6WfdknML
zDQa6NQ/c1PUmfPD8wBa6LYltDuiRs0zSvDeJwirnsHjPqQMsaYb+Fq/7a4UknMx
zMNPplnc/3g6jh8BuWox19cxfEk2wyXyfxb8mUk7FX+9BxAsSrFoVEo0zxZ+J+rq
SpvlK7GJWOFks/XTvMRWq0p63t89gCjT6nYsIvsHN9+Br6eZp7vUEx52Nxgzkxrf
i2+OLjW7FJKbTFOP/NI03yVUnx5x4m/CvkXn71ZBnHLEo3QSwh8hq8H0CwT4NJNd
Ff18CjIxJXcEwig+I5pU0cv6dtRpMQdmCv+awOo6WuYbf8EIlZ/OKmJaYwnRVuY+
dXJPKzPMsdoxZdYysymIV2P1hqXy3q4R+1YoHm9DDJuAh9RzZNs+c4QEfH14S/V4
3svMTsf/pBu8wub/siefk7pSVJnWA2ny5o0HqFXKnhUNG7oKOSAopcHgxSYV6cKJ
IEqFVVcHFg6TTaZucGLwvaAeAzsKk9L61BsroIFWE7H2LnwvUYjNnsSMT1OnBTUG
PosxiBlcXRLQ22XVswao6WbIU3TMKhm2OV02ffVe6vNMHrHXUAmh1jzz0Zxqa1oh
nOIyvX5leyCAwmkIbWQ2pFUMMK9xg5XwnXWHs1h4OVgjw3HuBIYbvW4RQ2NozKUN
xG7jzpdxzPk8zC/zJ0pwsJZoAh3yGIXGuN0B6mzqFaCoApI2wo8yO3cumi84MEu6
9BzIDWAjuldagNaC5NV2puGO0z5RYzVKsAaLNr+9fspt75odP/Ferv3M49qgbTo6
arrStAWX1LFUcvYmk6i+5Q2KYVmVeSnSHl74ReljK1w5YggEZaU0RZgl68DpixKl
CdQX4PkPuIs4JTaDg7bJGuBr4220xXmJTv0lmcjL4/W5EG1b9PjbGlDHuwN8b81b
JX06s/1ZOpaofCaAU1jmfE5bYo2uEJYNs4nxxymkeKG/DoUeGEZ50UDKbDgm6512
9lHnkeurcV8mWk4vwewbxgmkdHKH2e3u48SXmWYGQL9TP6poWWnLqp8fHT08uYp/
hWbsxEVkukyk7LQqkLqVDcdII0bt3Q4y+fiTROTLADlkgqiuxquCycyZx1y0aiec
k7QJjIfE7uaTQJ1XH+WEJybeUetrBO5VyiV0ttJr6/nZL2fGBHh+lZiebT8x52Nc
oUwzx93HRwc1tVSCDKUqRcS1TWdbE3MefyoAdMWJB5xdiPh0Nex/NzGWc/L56FxR
eCCnZAHtAY3JFOtztSf3tySD0ZYZ7e8ZS4xJZ8SJ2gyd8OQVTHWzRsZVfIukj6DU
U6XZwMrTksKI8YfLmAe0a6xT2/uVkzBFMD9CBv41/vIq+/v+3UdWQM7CkLofyVxI
N7LsNdJI0+S1WKO9XBoNw4bWsz1WWIVnY45RYwhf0x4GcEwKh8Qu/Q8pfhpAL58p
Alfu6aw98c2iYelzKfUKVE5nlpTZFTHV2f6V2c5uvNSxQNvFi2SZmuYrnvg+F5LL
r8kK2inPgqhyLjczs/8UJVcY0q1qsc7Qi/rtyBAywEMArTjhIvBRT9yZGUzP+Ym+
e1tnaXHUAclX2M39hGZO5unFWL9XG7pcvFoVlbEnXX5QosegMvXEPO9FQTuzMUff
kFMkI50WUo8vNdL7hPF5Je2kfwtzVzNpQrZ0HoLZQ7MAmLcgVUBdPAVKoLaK7Hao
mQtS5eeMfiUlUsqlhs1TsgrY6lqt2NtuXKyArk0P7pHMV6gD4nz5mGMKp9AZTQ/9
RGobIKmWxIjA7rT8OnJ1StkicXs+ayihpuXnuEQlCCYu2ukaMO2cFcIM/sCn3/PL
dRxm+/KH246M8LoirEGcMSPeu8N5n+piE2dGDXFC3jH+c5i1dZjGu/r2ujMqIY18
znjUmGrNF87aG6l2jkTbpfO/6WcL4pjkWWXNi2W11iLhpSHBEGnq4kjDT6FIUw4V
1SdSPOIATLHyOH+ZwrJh4A65D5JvtP5urziN97NbBYNJFlav5SFXnZqwzkBNZFWr
2atnEMaopnlE862hbQO4CLqZawZM03flknMK75k3kYXRtaRN9RsgFmMBZ/5CtkHp
cClDwjssHF+mxaYRAx1cb0G0zH2CyhyWum4pocVRpO+qs9LVfHkCZe2JNvNiQ2OX
rXKEcedGlm51h2j8B7LSRlxyAGJF5zDKcT8BPwByLYFNsDF0WhRAzNnHwgz3bc96
9Bh0NUeCThGV5p/FzqWgNC25M2vT8s31lkyguJwx9bDCsscilD3kgWC8ZImiJpBP
fPMWQGLimz9MaFColAs7LcfSralcqXgyktHri16Zwu9/0rdXwZzWPcRg8NRFy2lM
IIb7DGIQK9svbQecAT5jr42/ypheHnwdt8/EytjYevIwnAjq/Gvzf8rQ2WqISMgt
0ycnCjBOAC0XEuq9Z+6GUZTs4hYaP+Jzm++bTbPKKUX34VgCeLx8SOu7REbbYKPH
04PRoi/FzzVlQG1I5+EyPXG1OnF5N3K5Vje13uJDLlAjmL/uLkCFDGzpFmF1gWWJ
npPCkn+s3vAiuXC8KYJMlaPzu9hY6vgTKCQRqBSJr/xY1dX9B+Nt3LqE/0/jcMF+
1jjoqe0KiTtep16y1zXDBT60wCHLiYChqACUSos0M2rmvRlTwoTkKLNJVyJPapoZ
1KXntI9daFgygLhjEoSYhLDPeK8c9eE7EieJwdZHx/oG0Db7y6QotqVnYLSIl/RS
JXgT4tzscsxuu+KLEi8x75j3AyJ9CPFoeCT0wbGvXGJCSRT2zoMboCs4yqoE4GL3
7vA2jPU11gGh5cgTblsev1UxS6MiiMfjMiMM4lzfrOTJLwlRDjYle9DjkgLplqJh
TWFFAIInuueq4AMgmankdA1AzpOA4kL9DKsgW7aQgWs7btm+C5zg/DfMj3zzf91L
aAPd83N4kUivZ44Wlk4S9mMi50QEjB1ofUVgq5ei+StAn4h2bSD+UqG914pu3xvm
/R9A5dH422cVt27sstUHgW+eR5GU7A8zQ1OCHmbPMhWB1zRYMqorGgSUjgmwp4DD
N3bxjPO2jAqeGx7R+9V3Q4ZYMI3FKOFb4f9u2WdHF9nsYy4DgPX2xX6Bjp/IIqUt
8fppw4ItUgxWKiiQASRo0uHlfxaTWSQ1730nhJg2hQKb4xtnp/KTHCEL+CK5b06Z
m0vQeZz9rDzl9ObvRrvZayUnYz3S5D6PXMfB7amLClmblPY62iTte6FtfDJF3o/8
gnUMqTSZZAfBnP/tKrp3vf5bJxRskmC6C/KQBGTDiTT8CbecPFB7UrkRZA3Ip3b4
pxcmhQjFMGzUyQbj/Z5GVCvQzcPzpu/nHKl8yZGsXfZyQ+STIfBjckiLWTF4FJ5V
KDsMJgBn0rTjd8xuZ95uxCE6aSRG1VoNVTn3pSYdnamIfKBqszjRvCMy9PuslrCJ
oZSh5AzBPOtWxLTsSD8chYa7Wtc1b9MYhUJcQxx39ECfTaV7Vu060RzRd+woHYxG
GsYZ0PQchfu4GTWFjxM8Su0FuRR/xE3aEq5JZCYB4dVxf0Tbjtq6JSldSg/lym5P
nqnkr6tq1HyjaD0XDwfSJZXCex9+RdJ+KQgXQ49pspHO0RGRNngldeoERuHq1W60
FerD+rTZPPuPJtrIJeYcFstCEJuW2/0Ik6qCesXD6WV/3WdhjuViA/ti8bCMprnv
kcPPcTO0HXT4ErOTgl/1IDGKDX6zSMONjeFENIZuxZII1cBj3OzF9EMBPF7H19hP
i12VPy5AbI/RtDmM+6CkJknvlldaKhZOs085Xcxv3sqrL2TCOZNx1QthalBcW4lI
dLjfDPXMroEp4h70UXfdA7r7JiGn2iJu14Ht0EVHIvPL711a4rSqFxX5f03dqL64
fd08fpzqqvj1BCINq7vyE6rvdKlpSPp7NtXY3jOvy9GCSAQmvzLTOw02vwTAf7Ai
maylSk1/fSf5YaEcPGnVIPStQqeV7U8mtDVhpoZlt6E9NhmsNAg0NTtPqoYjMf8b
jOxBbdF7jYbhT9Wk/lYWRIXFMZoFTNKL6fsXsTpjVL3h92GFLFkbNy6yMzNZf6j3
05IBDhGqkgpsU2fzLf74nu1Ccm6n+kZSzxdQYQDTrllQxwzqYUWVb8tKcc0OytUH
TS+ororWSfV8tT7BtLbz99PJrNK4IBTqXWoul2TKmPMJ6lrTZDeX2lOaAzWFRKYz
jjA10nxEgp+SYbMWNvnxZWJDzuPhkOUa2SWmXeZUrXFIYzVTEHFCiAfCzMnUm2oN
QYAwrtdxMTrMUOux6PgPziXULn6BFbDXJ7AAh6u3Y6ZbQsupRF9ZHPrNkSqOeHHC
w8FeyZq/HDdPj40SpMbg6NdXDUbE7gUBaS+OVK5fAT+GjP6Rg/pNfqjm8QPg/myb
AOv5GwKjTYrfY7B8fyq1zDFEcH618NtL3iiaSISeVaCrUn99mgmrhVaPIhjdKRNx
NjHgHCMQYwMMo/D4hoAxAW7XVK/pRcwX/KyIKFT5twR0FAomnbQTb13oGkbO7PAM
CH/q/Rf+Zefh8bxTgm5i5jW5lzQqNUB1apDuByjtCv6r4TdQ5TvC4SBdTkGBWQkH
I63Zr8VhD0mkZ5C7SVHz3HRlFTGxzriKbxKVsdzPtM25JQZhjHxrbsaL0EGFFZzA
AOpdAWmry9tfMF5HECy8uKbvlDCkqIEpNceojebvMyMoUwCLLFCyTLI0b5sNfUr2
ZxEo0GSWU+TK+ZbIiaLtMs0qYqh4oBll9vnr2JpWhW45Dx/EjjE3st777fU2xS5Z
gbaWyQkQP8eFaasRbcFZM93GJBtpj845bfVcIs7DZEnrpOt+5LkytPYlb1c2GDzL
zZMt6EfNvREOFJ+ayMhg3qzEmMXFKUpkBkkwDeXYh3B4w44PqYQyIXMhbuKlSfut
K5tdfhz9v0irJdjYjMZTpjzd9MYdC7lo+LPXCAvzMzLpPNglU9anhu6F4Z7UJuik
W2lkz1OVhxCRo2Yvc7oL1omWLKZS0R4TjxsLJXb4+jJhvVJaM3wkwGozh6L70T1n
tUWfVKoPG3JwteSi+1dfDEH2G65ijKIq2rlSQbglTZjPj2/6mxT832EOOIzjWeBU
49CF66/WQBTJOWzMOu4EHL09oGxjhCHVUaTWcTRkCfM7vm8oCF03Z9C/bNkmUAT9
iaYB20wmHhbTLW7Wjv3Shx2NutZovKr2UMNqasKWxxW/q583QKPO8zzF1ajfYvII
nWs3rKLww70yLo/bSkFFLgDuHnymqZjaGxEgrpHOOqeDOTWSOR4OSxjBoSbL1rhl
n0i7pGVJJec8+jegRnQJfZ/yVnhv9q09PsbIerzuT3TyrxoCbQQAAEVUainKA87b
PeGF13Iiao4154OEcS6bOwbBgRHMPOODzKeILprWSbqpEDwRK2OqzoVwlgV47ApM
tIcVK06eSy4d5SGiKW5OoEfZewqtpQ9a1u+Zd+mtrcch8wD2hgRGPwTfemFaNK08
VY0VTimN832219DZzpl2k88Wf8EE9qHgOKWvBGX0v1LP9IIorfq9jJPfOp1lNbnw
3rutdOYwZAkWveukJYiUbSV0feC+g5AAfvEwt7ohLxTGOCOXjDvHmZdeYoegThf7
UdLvgZo5yyOK1JYZgjh5LVCg10maHYHpHteYzCh5NFyfdOXu9FHLQBJc+rB+1USw
r5nzrzXblpsMQp9yAAWv7LnOyWYhRqYbtxA3OgTMRPa0vjElONxFFimHEmsiQktp
FwocjVwXO8Qw5KFvbPGJMXWpYkW3zt9QalZfihZC5R6v12BO/S3Fvw83KuEiZ6we
L5awuplFZQJ/lmgZXqLXhjhEO1AeQg28CVXXQvpiDniW8W4V7eM3pfMMEjdGxBRN
a6+5nwDSCZ97anTPlfSKU4BabPSdYkLxt6WTrJ1HzlHhK6ns3la4CKIlt501dyAS
xqidLSNecevJZJbgphASopxHCdCmow3+V6IwjBGUXsCMTmF5PTi0+VKs2N9Jg6nE
6dlgn2d7ShaHec0/ei2kb0aLAcVRm5vdAJmT8XoiBXvJZ3pvE5stojG2jHHMugq6
qwRtfc6BI8jQ1npnkwmh5q0oDEGwzkldFxQFxiPqWCzplvhaDhDepkWyou9wZxAK
Hdb6JGJm+wRtbjCvwbu/7ZIIofTfJE25AV36yqU6cQyBNkuG57TT8JNHWgAJey6y
PzUxeeZCwnJUnJP8cz0xjJ2Ui4gwqLZe9vs/CR6Sj75OkG+US25KH0MK5ftZjwCv
IU2TBTcDG4n7O/EDves89rUEGVdM6s4EhCElIOFV4hTPewW9FKaZRkecrqI8CxNK
u3Bl/S2nHtRbNlkKJHNTFoKoPCH3/0eabsCO3TDEu0uPxtwudg9MsaOeQm33e4Hg
+c1Qk3fOhNupG1VVxr17gzMiLOcQz6bCc8PfncSCGMF9w4v8Vc6v67+Enj8CF54Z
q7hAXwde1yyWOMos+qbq/w7tVHehuF/Wg3HjXza6q3gx7jKlzYcfClGeA9ppsSlH
wuWu21U9nJ1e+qiM9KsHMCzaZwTi7iuJnB8TDMCI0UwLPggQ09ZuMYQVRV4yAZqi
ubbyJTwbbfYigCTCKY8MDA4SZYsTx27JfqHMHHT79fLmrq4Tgb+uALIMGv1xvoPn
somZYe0ISA62hd/eb29a7T4TutbvyTSH8dKVYhT+M23d7tkIWn4o/F2zakmxVa6S
R66iMKHz7busk0mZwU4CJzXjMEC8hzNEHGu2mAYpNpTDRvo0UMHaS8D4I9/Xrzqf
Sjz/n1fwXhNQpMK4aUqjJdES2JeVAPzxsAVE19JgPVYCmD6ocrsL9gvqiH/++JlR
CO5iLpRqRhh8I8BTYynN0d0IvAje73QbZVREgQ5jk/zRp+Y9GXelTcORiBx+MrRP
tynfJkWEBmXdQf/OIyBfmj1WvGY5ILZe6MZsNYiIx7VP2iBsJXqdRl3x1tPb3zD2
Zds381Ept3PF4Tmqfz3LaTqLS97+84eDFFs57iJUy9T0xz+D3qcMQnXIoNfjfgmT
88n7o2awFiIOZNjHCq47b8YW9J4inK1W2M1MOXKVTSjgB8Sk+wQUPv5Zuw177ddd
VPSYJqA8WYbrWreGBPIQHWrNDOAI8W8l4fBvDlAlgtsEH/GVCARguKZuDqw/4ECP
ynA3KVt0XGUJxkoX+1Xu4qmAhZqxV8EHxk22dCOBQ14YJV9twT51dVT+o8qzAyrd
XI3LcMjjRpI7WMmXY4mB1vwDiMGB6YCMjFOrsjUnuAZS8qlTy3pqKL/DFssFuGi+
dhOQhDhSVAcG5EnNGwfpvTvfdyf2vbe/Xm/6hWEu0EaSKKae6OaLPboBxleBPjN/
oprzD759sOwUB0ZwyCXEFyPpki0ZG2HUCAI7F4RTBDR4qrT+9W/7AObmSJufm/Y+
8kXW9k2fmUt0tMFkeTGmA95QvirmufKFSaovFFiuE0kMtnscU6xJyosAJilfC288
t9L21p9ezJaBoHBFCG4iF606mOGh20yxZSBEWXcQX+6QJ6lnB262/m1e75FWt8as
bKkCIJ/HmoFikIqrdLLigg0spFoEDUR/fWhqSp6Alr6grym0b2W07VHIoXY/5QCp
jZHPtTob7tNQeis2GLDXiCXGafx14N+/5xqAzZz8+cxbC3cAkh15Qj0UKpC5TJtH
q4OBXfp74+9VPFjkgUH2r/qyQ2TNFjmZ2LT0+UFmHOV9sYZUXleShjDiPiT2GpXO
jPdMhqU8fS45XsWPavbWXIM1v6P/JnXJzv2ayoUikAcq5OCMDybDgUxcO7DFNrMS
C5vwZG+MeIgqkhFgsm4Z/Qq8cQtgyFM4cwP2UPtnc5vsetLuK0j8eZZPaNt9JGd5
ZcTf0snTtBfQCaJbvd0U5X7CwsMpdWmB59nhjchzF8jP3/Uet5a3JFkFe/snDVXB
lPUwwPOavSMha3agMqD+C41vyogeSCu68WroRAPzR159zxoB9wJ6r2L120AG7RZt
47YW1JktL6IWGU6e14FTrCfsFYTvYFaHeLAAqVy3PPyISBcllvXh3wHZ8lfwBmzL
lqRJvQ4IuxwfCbCDmvzUjiN4z2mOwn3qqkM1NCFYQg0/66T2oM94/+DMSFdbAT36
OZH3iPAKtFaK35G1UNwtKZKZyZm9Nukc5xZnLsNSvkEH9tsoKzZm1dT2E1jnOt0T
/TqW6r99zxHV+cnBQ4TNM/KS9jT4W4HimpUs/VdaqIEdFx3btLFu04m0oHtA4Ow/
QfvAY0rhVrwY1Hva0WgNJjbtklRas/nvP4jrZktSmF0MOSzs3YCI8fJsD81gdT8E
915GdBmiwlsEuGRiKRGLf3zZ1qnuEBxRUHmq9At+XPSN2qUYrWH/43ZCcRCIGIwI
4rofhN2SOeh/aJ0w3KxGqJ1AhqJ32JtD/q7dpF5Ol7F0eDcMIAHfO5VckYzEsVi2
wUIbtE9+08Sutm8gTP7VjSYJxZFwdoNOknYWwxWy2MNyqfroSKwvCc8auUi9ejme
yvzXL3f/cxkGHdPr6bYygJxg2aCHEOAj8dm5fBvCJ1nyCNLigWwr92CDfkYIylq7
CTljowGpxysezU7mFkxfPlTcmRQJttud2LL3Zbu+4l9EvSxAkciTfd/83jPYXB7a
D9FhhOdbUR5m5ExyoaoRxhvoqd5hEhSte5LsTzVDrg03iKoDzLkunJQ3RoOqMdC1
tu62WAlzHPClo0jcZu92ltg9+lWgqA6TN53wbWhqKuKgF1kYOxIwNqdEAQyqM3Hz
hpe5so5OcSM8EDe/EjyS/eKq2LMbbixeEnLaiF54eEbwkw7EO37RNDIC+MJxpA6Q
HEA2EIdV171/hC2+SvZimKS0Njs422CKl5Gi8jBIdK0Ji5JRsUNztIsWOi1A3uUh
1GGtncK2OLyu6sqvYIUnTE53MYRNwq36f9ySr/WMO17A4DOgTMzOd/GmMOiAHzHs
BYPUKoVSUkdbpZsEbFvb5/3DfjVqjKaY5OvroZkvC3C2QphefAwjZGLQtEw1RxP9
L+zsbqz1DBOHR/oTufrD3eHUA8FozQHAJnZQoPF4TqW7AL0DnEsbOxB5O9OTiYs3
wX4RYCQHrDzyZqFmNJm4JXUClYaH49vOeXNLUA65DSeYiG9BRtRsMI9rx66uiX5v
3cA1daIjw1PBGz8rmqySdZqJoXSAdap/IJn+9UKVdp7DCxyCZM7BCGF9fXE8kCiW
1HvA/Yoz0HcYMOc+yx9Az0nlzZtTKdK9f37dTcBsD7SebB/vgcTSYVJbKnoTnDur
1QqtQ5WknCS0cFgeLMYl+NKo0FtJNhotvyvjdquhIlr1sf09dwEdjuarqCFPsX41
9oEDABX+BhUbcfKFhsu0J2GAs/y7m07JIwfPzbTwqxaxVtXUCiVonMYG6ojAOmJN
pgPVWw70p9+KvixKLmqlMSplb8Btzylfdj7p9ogrjVi53JLPU7XyXcUdLWa3WgGK
L7Nn3NxsVZtq86Ub8NK4dvOWM8I0MKIsOf7SnqOK1/jHDMhYjyNy5+bWKgE3NlPe
dFaInAoj7AN/SKn1TtfKiSUOuq24/63dKyqX8sXc3a28UntVE0OmHDS0ueNKYbh7
fPC/8HLHLtsnVyh33Z9O1v2WWoNxkFQayA1anCQvMyGMgEyTRdNoGs9NFs8T7FYJ
XlDxQsly0Cx29F8F+G5t3mkHWKvdeQWp1eWqOYnKLTyggaP1m60DqTssaL0vKDvO
5TcbQAZiiinnW4V2b5CRbz65fZ2IV+9l0/WTFjeQUrXLCVotxf5GCJKHEGP4z+YU
X6vmcqquz6X/QMfBafY/nf7MfKWSQSm/uW5Bl3Y7AZVue0GCZ0jv0EUGlV/LbJQk
I7Ts62RBl3G8Cz1+sou0xq336tzshhB121Ijis5PDUgK0vJXhtjIHY0IbQ/C2YvR
Idbf0aO8i4xZT5TozLvSFUnhChHECjl1QnFcC25WUuAsWsPAsmoJip+s+BgwNk/A
rknGWn0MkwX0h0R9zZ5R5YNdnFPMWLFquB24aoi+/4EKGYLdJ+JodVQX+2+mIQBd
R4xOQPaoFIzte4oqnuQ8R3pGDGmQfjhv5qt45fBR9iCWIz9n+sNwttAJmyukV9ss
0saTLdtFiGPGFwNZ88WOjKLkfM//ER8G5mvEofj3BmK3hFOmyqeFr2hwu6Eip/o7
aUZIqENsEw/DtSftsWemIYjslpXzZ8mFDPLTEQEW3POZIRmsElZsX7JrC7K2Lktf
WVhwCHI++jAGbRRG7sbJqjpepKhYE+uMMgSiINXpt5B6plWXIJQzyiVkDFQqdqo5
FpqdLqOYgfGEU77rOkIEL0uVBQgB1x+yvck9nNJvojiXakF0dJ9PO9fQXxWkIAxZ
kBAeDW4G0t0QKDoEkUHrfIUiDd7c1AZ8ieF80Tsr3w1HNBMs0r01UGuvS+mjT1K+
Oih4ouSomB1wiIZfpd3+C+AIX/A2eY4774HaO/NKi9pC5f+pkc/rlVhk9Py24zXY
EXuTjJamETv5HU5ykSvejT4hjnW3K31WhHhka3Ff0mn8UWGvRuOuuKzeC5vP6H/0
Lk1fQKMZ+WY6kKHi7EI5v9t6XcWq20niAoiiu4kmHFjjszDdhy6qYhLnhCIYhE2t
/A2j9uLFElsjo7SeioyLrveKTc8bSN3REjfZnV9CiQ70aRA09/eV4CPD0tHHD0NF
eW54LNNtaiR5wRXFNPcIOlNtZxtvxKE7l7tobdVkuPrIbKow2LvrtZOWatC0CW1B
DOd5OxjAbpYh5D74TOtj8neekTf3FhrLhpn0T2rMwm35Rz7eP42gVh+1RibNUtj2
fM4qCsT0FZMMlaLIpKbXKyDSIDWkStSczSJnyYryG66vgePjo+VgdLQ/N032A8/i
vw3pegqY8wH/CtkfcN8OEVOYzcL9TYIrcRc9TbKmfcI3TxdjYNsxictByB6SwCrJ
mtXVB6qxUrXLRl4jbT8HRHxNKUaI+k4nMP/aXesFY17XNFN8gqn4QjRX03X7jMWo
mCCviVV3241VIVh3n1/M+Kr/izjLBJ/QcFvWvknv7mdnb8d5DgUlsbxzvnnijnu5
hKD4YXNg6Jrnwd+ByZ/jX3eXhORAJjXoLe6tC9p02GVJfGtltOoO5kQf0+Nl4uB/
PF6EVHoSOhQnNJwKDT6O/dm/rOwY4dbetpnyRAHyjEg/oRN9GcDQIHY6X/4beuiu
Ln/47gtouxN7cALaNXiAoRB/2VljQm0EINGkgiUtTqd0TV7gZXf13Dp6OsYVXmp/
Yp749N3XhPgs9O4+apIDqLn6IzPSllNPsPsKaLoxf2rzRfGvktj6Zuxynjwg2itE
Dm4CePrj2jzzpxCK9NBvF888WHRpXhfjrb8lSExpCdC3I7fsjitgeoTmN/gFbaKZ
FRuiqE90hSPtSgDnHucxCwq+C87/f5wr6jqDym5Yl/kozY6JdMkiugCTw27/aVW9
wx4GGObgtgW+YhPwwPRO1a9+iJm+rk6M26Qex0u6Ufq5HI0ZDewLikg3FonYRHvY
vJH8udgjbRrgdhUe9QYDMIAPgkTmkUOhl8P0LKsC5XBzUHTNDn3i7kD8kW8GHH76
NKlgNmL0ZeoXXigdw+Mq5WtCQ9OH1HngM8Xe+8dviC4fBdOVkaoNaTs+Vo2NzlTG
iRea/WhTI3DU7fkPk+FIrdfbYnyAb4UrYqf4CyO5fx4GL3l6kTg04SyA7/LJXyqg
xtCM8Xhyyn3LaaqquemtnnVRenqmsyjlO8Gda+dyE7WIjsxA/up7E+/VjfG8gnAJ
jbkbPcQLFZOoZmP5UjXI/+58kCu9q/U2NDnbzIpamQpkAeCRlfKieTedBxLMxBo8
OLumRPiYTWfAtgF/2xAFJuxcthkBlpb3j6BHBCXhs6YNRMEMgASyfHs2CT5f9SUF
O/Ui1lxpVAyUQ2YzjKzDOj6yHSwqSZlG8ikMvBefPQvxSfqqcrhsqvx2VeMO0Uz/
db8rt8D/NjXRPHncJkh/TpKy+RxT/SBEH3DfWcM00XSkmtYOx7PbjDfkHFGF3GFn
Y6N+CipledR8TP8Pxz7K0+E8BKOuQNYPDhDUZIKfj9BF4ke5JgWM7t5Zlr/0UcK0
60Uo3L6Ruvpfu94NLKzNuw==
`protect END_PROTECTED
