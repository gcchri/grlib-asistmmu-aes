`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FxVyzDDX6/f2ESSunrWyYfRQAD+I9kw/CIjQb/H5lrb+jI+h6AVtlTArGYLtpkHx
LoiiEbY6kyz3/KSzKiuYWrw1lQC8LorXU5H11vfrpBWOx672/RYoFJiVsSt0I/bV
6uSmlKbRMUMUIGPIVpvi+v3oheMNHPCUtRNuAqpaW2xOTjo1Aa2z08BfALXhBy+j
g8aBcLys5tZtWUGbTIwZhECMoQ3YfFIdw0JZi3aHIlrpby7LBpBCvQix2AWmC1sE
upW1d6fAoJJ9OwfnjwsebyaJr/Bu9fmyWlj8itXYwSA/yWXl9cLVkcrezZefWvNb
vg7L0WWTuQx5cdYdhUOOKig333ndVedG5d7XAtiZPur8newbhxhfB3fJSNeXk/iZ
Pruof2OPVE5TQWOW6hBQhS+kOZcg/50l2R3HgQOxNNh4pHziC6xc3nitR+3FGo84
Uf+spQ8AuLB0EUyItppMR5y3FXDjMFJJ2+ocz5dNlsT5+oelFAJ5RwnfdO5uvsZg
s5Uvn0glqsE8aQxPAPmJIWOmBMWc38BjrFsQS/4p9a1ozrqoH5fiP0kfzRT4L7OB
hDx++XWkz/o+gRrprWNykKqXWGb1dR8Z7erCHSC0jZkAXcYoJ8D1NkUTub5afPNU
lBpWEYLgaq2XmTb4VIvZsMP6B1LGjNav0Zb8jETr83yNhlnEnxzvQAmNg4jyOHaz
Gk9h4kPPJYe1tdlUPWMW6mj3005HTvN0+c6JLvU7TEgyzK6ORu2iokw6ajC9zO76
HuHaU8k8F8O7LXFcZ806AJUbakzqQVGhzsMj2lZ8U9AYFCddMXPfTc3OrsEgwf7C
uL/3he034K/O7v9pG6t3kom6BaI1rlWSlNH5Xh8OS16q/5OG3kG4CRwKuEm2X+xj
pEQWm1hXETIwtd2SXP9Uch+VNVY5uxol9kdc7mh+7ydjV+bR5XxPmF56oVdpkTvO
gME/s/eXSdnWuliJSfSl/NuS6KchAnyBY4FLvqyfiESVAQ57Auzwwwvsh9Ih02AE
iA5m65bAoyLhADGD24WZCGM64ImqpIl0eD2zkGiOyzxFXFU5J1xpK1D/xuE/ogod
nBW7AOYICSMROY0nVvHM9wi+xmvba+FI78LEDwX163L2HtAjTJXLu/3b8J8kHv6E
PVHAH10h4NfRtzOJq8VLcA==
`protect END_PROTECTED
