`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K5YTYU0ycYgKeeofphT2xk2RoTYb9es/bdI5IYVhhDNXiYjQpcuZW8YeWCq345/j
ea+IWjb4BwbOI9dfscvBkFnXp7iV2eIo1XZISbUmTEQA/OC8PH3c/HIouNarBAU3
JmBiBJ7JquBmLSthK6LnInKwBwFweOsD8wDBrO99+bQRHPuhk2zyweyEwimeXF5a
zEi2KefElnIRaR6RwGdU5E1Gm/urZYwzw6tuSQH11erhwstI3/7KvThJ8+akis4o
IfZdw4Zis3XaluUeILzDGM6E2T6ZBZUFkOaLnuah3M5RMxjDjJ5IqYju7ZC7zSPd
B7+DwtDFGFMA8LCw/TF7Hwa9K6jehqYtUopjR+RCr67qdfsV3AzZGzJBv7btYVKi
x4y3z5K5+yHAg57KAzXTN/KOUxxHw6+hmAWIh3fg43iZoVOWNTS5z4jmnUoPbjlR
t9pyvJpvMMLmlHECoGiBLHfeS6+NLu0C8iE/QSfOKKgVabk8SI0mCle6zr5KLKIr
kq/BRYkW7GDP/qjyDRH4Yn+s2ed1vpcKdNXF3chudKwTtV5APKGuMfxT9zMitVGW
iVINqgT4lnPqD3VJnFi/9/c3YwEWVHVReVnerIgVI/7UifKfdJXg8pOZ4VbfpCl1
exZyeP8VuNSILiV93K2NQEFxnFeE/E8tg15EQOmozfFvK+NYpSBgRVexarzLb535
txaC+Vg1Xx8qXpckyJsF8AO7A1gK3lYLr8sE8dskfOmLFBNjnL2mUPAZOYo86NbI
9XJAo8I5MxW+5IjBMWyzGeDzyqv70tELd3L9R4QVaedVSHKn3TsSKhdMhJRQTcTw
PnLNCF3YsdLtBOtkfuk3Wv/Of2dT8FmbfA184DfWwQXntXVL0w8YbIRoggjQnQHq
wNffXot8+AIa181Qw7mBHFg26R1GzinXCRw0AJfvO2Xiefiza//wkG51KLtrmLY0
WB4IRzBE2DK9j9NQcZSwcsFngHvHLdT2KYnG4c/ST3B4/5hBx/xgPjWqi89/lhbB
6s1yXg+x6plfGtCG7nwmSToJybnDSWJ/rrE6OEILEgBYgUwAoYO7XnT83cnQLA/W
uogyuWhNi+Q7FWEwWJmZDDCIH89creUegZI4Bpl8cveq5aR0Eb3XcJuK/Ns7kDbD
u+U8Bldv6U2qyN168S0QXAIASPs+O6qwX3zKeOPUgESRyB87hkKc80VzW8DkFni7
9PJhdPOAR2TL3M4vMLtRLxRJTdE1yK1QynVyhCjT1FefYD48WLrPHXR05KZpaas1
30O6IMUlUmJzPicrbV/7x1D9zA4Wm/sCKz/+A0Q3Xp+P1zSdOh3Xw3n95+6qSggV
FEpCKIm7jivH2zXuGQq25GzGFv04hqBgEha4ZOnxewtcebBxkntKKVAodrDX/Hnt
wBpP2unaXnNC03oh2iFlYq4BwqhVYAqR2p3Q8jyyDz06VrbuuCcD7+qMLOeN9gvP
jIqk+dZ/S5zJqlYiM2yDAXxh+/JzABIKlZDwT4RF62++5t4ICe+33zJk7c8Sul5E
ZFoEOaYE1vwcaJj+g3fu1kwcPbMal2n9n9VkmugD8VCXy/HPWmgRg+fQdSIyoyAC
BY5f0DeVSYEDsjNbkJYGPTuIQZY3pbwo/ivLoWA4mvhfAO3LmjVdxMAX6F39wpps
0+unZipPlvomK2biA6Vp6oRFT8RJ7AvenYn4sDwqjVUNEr4z9AW/Yca9j69u85T9
qntb6rRtbihkkVen0zpPXBcJBptnzXFh98i6zK3KX58xrVJBooeBhCRTTq8gVfDe
MROEiqmneTm6ikkqS7VmRRi4cDBTCOZ41DXLX4qelXq8wsuaOy64Cl9xVuD/2H/j
54+fLXr4wJKn6FiDgBMoalaNZAELD3iiF5rcqAyTBVIqTtb9La5MqSYiYnXDPDQu
Y52dHtAdcSCuLMnRcEHNWi4q4ESoCManODKnrrluzaqO7ZRlDBRbO+0ctjC+erRK
ZMBiZ2NkyfmlIxE2qE8rnbee04KSCysqax9DBCCUhxFOophKRB/OxnDBNzRHmuBP
2+1gUkP9lhzNJqIxMidkXQ==
`protect END_PROTECTED
