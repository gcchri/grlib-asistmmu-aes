`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SNcDL2fyoJTY11p2RIEBX+AXyQu8pP+5rC96ttw5dk26ju/kqBOrr7DWEfJtsaU/
xX4TJxwySO5jGazNNXkrbiS7AkU60NSzi5lEusqT4eIh0OVuqHFhaMmruRmpKj40
aivgevPBI6YfVdFkqctgBmDpQsLb7IXUki5dy+ep8GansuVS6BZSu1wdLjvmbCl0
ACxtXHY7ttMkv8wQWyo8TO6kcWR8U4caVqQ2DR5VYP9bBCw/p2b6VzWnCnvzn7x5
RWy2BKl7dTHPod4YUNPnH3iIzKygp5DWor6sQFrI8QBK7VEdYBXil4tvYlMhqfDH
EjnrwhaNbD/aV2t7lqBy7ODRDiaXiFcDUk/PgLQt0XOpcp0MAQmR0EqUpZuHbML4
qfuRcKgDQlGTx5Pnfp4WgOmQHmitcO61jtI8++YI9v4zRpnDY50/n+939jjuGmF9
Y3r2m5tOt7rAw5k08/PyquNqQN8ZRxhKyIYLL52Tv3JvxD64UmDwtyZ3atZJTdxT
XvijrPwuaTAzfJVSf9kMqHymGyOMwxnNQmaD4pFDZcksXyRXKIC9kcmLfXCleyGN
7uPm5G/HY6U84gTe7GhB9muKblBSVBcZ2BcuiwKwYwXI0V0RmXbQa30HvzSSovE4
ko3XS0kHkJkryeiNnOvnvQ==
`protect END_PROTECTED
