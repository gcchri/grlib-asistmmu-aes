`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
79n4pNmuX0uhkElxJU1BC8cIvd+/w+uPUUKSbzLOsfiWpUSuqKMaLJggxTNZfBWO
Av60a3xpKZd/DExIJXKHLryxeN2vO11ZFh1CGl2mUh0D92KLUaG6r0hWaDRmv8qY
XB1fe8HQVIwGJhqf9XdjolrGHFEVVN4fsyofz2yUs8jsvj/hO6BGhfLHpuHa6pWx
+fPgsqx8xSVB28s7JFfvPH2UzipiLK/4+ZUM3cWnBXaKzpgEI/O1Q4Qgmd4d1z3W
FZXs4ul/Dng4HgxHNBTZEZxqiZkS+X/kngo+x+Jki6P1YgaxRTI1cnzKIL4GwykX
zd8qvg/n2b3TShZFa1gv4/yDX3eqKMjHwYffnsr09Zf5dvvV0NrFvuszutMgAQ/9
unBq8L4NE1PFgRVBjOCypQ==
`protect END_PROTECTED
