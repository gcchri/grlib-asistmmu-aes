`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DS96HmWECg0uZkDyqI1nIGz6b9l20XLIXtbJhpsGf0V12T30Z+P2AtqH/k6YY+tv
hA8+9B8np0n0CdCg6va4Oz/ete64ySpFmkQoHYKwl4JBJyaBkFIDCGW2bzjePoD9
/I+kCj9rdYCe9zA7+stQsRctztELhCDntcdgaSBXc9RE/d6hyuGOFryd+bYNCRS0
JKIy9V8sO+OnaL6H9od3xsvwrzJKnVHzsozw8B8SJtHdkap1MyXmqtCaM7CJV/rN
sqpdnJieYJj6BHVj7SK7AnH8PZBjEiBhHEqQH5JMm37ZrDvC1pguiAGoRgdhUMLo
pwtYQLCPS3g51cyeoFSqKl7Kh6K+KH2BiU79dgJiGTjBZv8LRig/wyPMsPWDIV6i
WgBTTfWF2tK3N0pVlE+7Bw==
`protect END_PROTECTED
