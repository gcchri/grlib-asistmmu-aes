`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YrejXRNQaJhnOWDHTyqpwagPsffEAi0oCGNMsk8c1q1IPEd+PM65PE6gqGisEwNU
PkkZ/1R2Rl3apqRcAX1xLWLFEkGjviwJ6H1ogXzmV3reCe5P6A+2eVEX3OztQIBY
Hcmh/pDsJoxkjUDrTQ+fm+l9yfat7qK7UcDvaGa+hCszc5OGr6pMRm74K4D3iIrM
eIcQRt4lHkRCOzpBdd4+hCboa/YH3335z8Y028OkSbQ4uq0Gn5mHnMHvD/GKVpIF
uBjX+ByawKty+BrhsAKFMa705jOOVRwlMHmIWGjo3OaRnmoK/e5So9A/qsyp1yV/
+5i9zuYq2MXVE/o/x/OcrmNF2EVuiyCqlM/ZgOcHTDFdtBXvYvRvS9xGSf2uIEFW
tyWOdL8vdyrfywhWSwgj8ZBQ9GuWjURV1XmYBy1T2YidhrkVM7tAWbEo+KR74Qxf
`protect END_PROTECTED
