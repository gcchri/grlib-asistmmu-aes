`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FLdsYVzK1lYub4PXq86W3Duv+AaFU6T7KIGZX54DvjbWl17Ghs7+vxJi4FY40kDj
J1Q6UqIDA+KHcAcF0asN75cMU0yyiffG2ZWfiuMYajmehYKmDOa70C/fMN1zSPs1
4JSw8EgWjdliEZmsd1AMKutj+8OwDfdV4vC7kEuW+wWV4HFZTI58GC5hsQvw22lR
W1uSO1bis50RY4UkllVfuBH0WlTmeocQqND5YWbPdr8ClRqx4ssIBlNXW+qiBKvm
/iV7J7kQVhPbZdYrkF0IJbMkoasby71ayoKG6Tf0iWXi9us3whtZtUvQkp8j7xqw
PT10eNREPYZgkbulsWXuwOO9/P1EIm+N6qzduyV+sKWssXYU/ncHNY6EvK3U6FoP
6vDjh8PwNESn6uEd2NY8wA2R3HTW7bpzql6gDjxYPPI06Ce7zWFnB8VZxLoWlcVB
bpBptc5raLAN2PW1HCrfENKeJFI1qjyPKPkrh+HpZoLsUBD5N6EJNHsH+BnfgGfa
HJsBMzkundJE2I5UwVTWQsq40dSsVBDk/nWEq/l68YXm4c1bU/G4ZYBvrjaTz7XR
W22shv3WWtZwB9Wdoxbh9E2uTlcCLwETfL9YNm82N6TzGrqVfMJCJBYqi+Vn8G4i
UxEQs6OK7KvW6girPnPp1S1kz6fnJSFoX75dnoNwbOJp/lGVohYuSCUDOM1GzIxP
YWxqnpmT/KjHZQLNloi/rwplApa6xJ/BS1IfZj+9gxs7YEL+3FIR8YRfQxlKddD2
UuSz5GddNunYodG8M/XU5Dnp0gAfa6u8iRJEitJ4KMNOT9kh9URZME7FAxx1yTya
sXluc7kIdYrhA4pb10klt6QHWWiNXcCEKG4y1R7I0MEnD4pxR2w77JWgpIXVLa1K
Pee6cl8CX82p9sDxSQ91KGwhHbNsYWcQkaXma1I8baup1csMOejSRw9MLu0vknKC
sle6crBwvK+G9CJduz4fM3J9P08mBy6IxrURqAeWZJSzOw7kElnH+wX3th/xU6z2
mVuiuKsu/Zbw0nMfL8ndcKoM4Vj5m8k+u7PIwVaTZ2N2KQiAW2hV2l+G/ie1Q5eE
cenwOx6IIPdDGD5HhCgLJ404eWtDyjsTasbp6KXiInToYvt1ikIot9W07VdHh04q
0EfygHOnJBalmljPcMi8Lcmp/L2aeKltgfKYtZwtos29t5BH913F8t8iLORrt3QP
9nCDHu4It/syp2XawnubFHMHr/4+ZT840UPZ9SoBj8+N7tkWKsHwehOOz0bRDM34
qN8EAV8VDc6mJDtLBcl6cXSzCJbF+wumKU0qNoB/znmQ0cK1AeZQLfsOV8ZxJZOz
pPuXBaQGRQwTBlAlRJLkjRaid+dz/28XiYuTUFA0jxHwz07zwuIfpLqSnND5zSiY
H7wNYHvEvhZFBZHSF+QYzuzBi29XM37j4LQaui0haQGbf9jPpNPS/1cAxXulHKRU
ZXszhOin18lLdZbl6dL2/EBNl4d2uSCZ8q88/ci/3zl1MXqSbXXq/wJIM25Lrxa0
DNzrCciiiq0yl4ng+MVtlBUQH7/ciUffaLtcy6bbn6q8eA5tjwWui/ja4UW8cxPb
3H7qvU0Iz32GYMrkMp0NC0LQK5P1CZwVqSO/nwam03mKtxfzhC//KZWDfus/UUba
SMLm/UCdNENVTU55WtTnDi9BqixnEdzroiXoP8p9emJqK4UJVfpUKjOudBekHEf3
ijPfKBllejuWN2w7hrUOjxyClCHWYB/o3ljqSP01b2uEzExRIs6RpGGAlQZIdYJS
nedQntjZdCs220e9v/aJLPm7mh5179w4q04NyC+1LnvErHSFwqFq2eLgkgzp3rHf
Zl3oM5bTWl8z1/7vf0F02BrWDyKDpezriFlpsdp1sggOYjluQQQebFYRhshMaCb7
VhYHtEJqTJbgOu1waZ0uVNWxzPrzjSBi45MbDT7BslLgKvfwXcDZLgB/J8DauNVX
9/mAXMvVOmX536e/T3dbXzBmUONcgRcbqJQAZFU/gPMrVUN92PgXynEvUguSwMAH
hTEzSz+KwubvkUqqGmwE/T8MpdLX7nbm/VfihrARNZBbUGNlIMc1/zbB9A8VHHcm
PGLqOWk96R3Oq8c+3xlqEWVfuzfW26+INzDL3LEvGjIjcHICif/OF2dBm+88+nw0
fPGRNAhVLO/vQPWjwKNHgq6ZJiMC20hAKIjG5DXrbmAnUov8/oCSYWO6TRlhuGCG
hyMEZFh/pzg+1VrElzt9a1qWEHdvUpA1C2nmvQVuUxeAivLtgke3vOdwMA56uhtX
eLeONJf4uQ5STRKvy7rBgbr+wAyk8b+JSGvoOtshxKpKSQU27Vq/NSHuRnONGVgz
GIFaQmE2RTIu426ktB25OAYH370bxRya0HMjumqSK0h1j2EE8uVsdHplVL+Bqm+R
mGt1rPcR9IvblWA/4a7xp6dgZ2PCLDHoIc7dskFg/daI0GVMjaI9jo7matN9l5JO
Mw1fb/gwiwopgjJedf3ttz9QnH6VDc+LWuABVu+X/hWLC/UqWQ/j0/8/Tbv8STR3
r1DiP8WU36U6/G3uAJUEwW9uyBoelcpjO5dFqN7WWpTHg2M1q9RaAh8XOjp2y2TM
/xPL/9nZXZWutPnhRSl/SHW8ic6CB1rdVE379E55XQUYH8qd1WmRGbb3sGf0Bts1
fVzpJv5QIf+4TrWP60GuFkn4ICSXonSUBzGBu+LO5Zw+Q1TfZKfSP32cALOQ/AwO
I1hkHBbPMMdAS4EoRvMn9CAjeGRekN6x3DG+jkddyI1drKykE1zBXM/FK5v1w+V+
TPC+T8RpaFQkpimkTukNlXKbZxIrYooBEWu++GF2xAeWTsoAv7Q+YbxvEUzm2zGW
oOWBX7Etfk/9vxjuvZI63C9NF6rYkx4kkon1rAJ7W/K1ZLthVyFJWKOF6VnXP7hf
xBAoAkT+hwCIaIqIwNfKTVVcNx8L2yS2pj6hsT4tMil9rUoiiRZMK0e7fCpVNask
eZEYI7z85BxmaWrk6/5Aii8BfQPEyKeU4UBdsc7Pz3a0w4tVpXL/ySEsc5+BqobP
pP8299MeK8Id0rN7oGqfc6VC4oM4/BYjfsGVrGmF7JVrn0BnWOm4TWai/uJydALM
3J1JO03T7grxHiQSdUIQYMBpVGz6fw0xnWq1gLtIr4IymVmJEl5mvaR1lzeqowoP
4AGvnLGnt+va8ZR/T8nUVFQf2HUIaMd1DHiBRhSmkQUa4QWF5l+9bf49d/NX0iVh
ggJp44jTdA1v3n/E/rPIgyZ1RAPkYrV+2hTRmklRVhfecL37X3MbrMBoTJ5HuFnl
8hYiZ4UfHnJt6HxYYBNVpXkZYgNK+xPSc946JGF4YQJtRvZBTgFzoAXBAGKX/aE6
9Ov3k96eYhCqlnbFeJBD4O3tqUb7ptclkXUFYsvIoFWRex2PdDGWl5PCwMigQvlv
v8vwRNvCqk1T1Gtp/N5nEFeH/fd/KXjoQu/mm1Vl/ZxXfohlNXTSImQN9e+lnlkp
+mmH1nPcIpAI/dUvD2OxvJcw9rQycFARvj7srYdKpSr/NaId4+NerZsGbL1MkBSS
AeXzkrq3QOr+SfoTYk9FTL93jaVN4OsS+stBKJLgZGDkL0wuvwYt2kwqtFdFT/XR
lyR9rEXnf01C8bPd7LIwAEWAw1gt5DBEDoyHkeUr7VnJVs+Vx2hbPSchFr58HbWw
AIVBAJ7iMihTBqkxjor/tF/zh/kUL/qa1zT0RP2nnK+v/5RHhg/CDHGatsSmxBjg
lMmdw/zOeGurHF7g+ca2fWWn5SF5WxZrmwko1Qm2O6MZaQSduAJCHux2dof7iRIA
3uaOzuiQodtbsEIxiIwskyPArMvzQ993qRI2JkGHBrUsvhOqSDM4UHqf17M0RA3o
Q3Hnz4lUzENMt1jhRe1k+chEG5yfvf3f72aWFhcBZ3ACwzKJuqOk9jHxVyH1c5OE
oDb9P1U+LFAfMTnyAimRZmUI09KLPqJaJZd7idXN/PsgfE594pRmbSufYQ1hKL9L
FyVCsj1EggItd54gwQZCFP6OdwOul2oIXvGSFw7GlaWQabpjN+aPhLNuQk4W0T//
IJ8ocbPRU2uvp3cjvcGa464hBSxfRhSmJAOlF/PLssp5laXvI2M0KAPyn7ny2ZFt
EvnV+K9qRh/REFnnlyKpyrnLYVPzSLVAbQRUHHNcrdf/k798rkl0HWiitQg3Fg9Y
pU0XkPkt/MFqG/WrW1InX8Pb6J+C5Bcss4KEJDgGzfANKbdKej8p02tMT3ZebbgC
feRoYXSKOaLmME+tnxEJrmNyIIhJCJv9+RGkdM5H+eGykHQRa7WBr0sEttTN/4O3
USgQBHP3XqIQPRXzKVUSiCtOhkgfA4xDyQX3I/Ahurf4bBuz7rPG/Fmt/P882jnt
tuU+j5aZLOGiCR3Zq0+EI+RWXGf9kUnxZ1NWdgDmdfv04g5IoIS5r3dQGDFvU0sb
RhgVgove44OQBbzipiT+cCWUNhsJHYwqQpMMJ//kfthy9QW90a9aPJengBj5ZBeU
agAc/4igARhvGVeZaU9KqI3Q7zmzhOXBpYhmywJRAQBblXfRzVtLZA0YU6GQWaNb
RxNNGCt4c/lAAOmyjrc503NETzXBuspZtDl5qUUDjDUk06RmfHIuiBgxOT+aNIxh
2q8M0sksFi4K2UerE2pQr7iuPob0uk8O6Fjo9sVtSDP2QhgNUrvAjR2LF/5Uohie
+NKEIFHTcls9wb2X4qEyk9gNqShOmAtsWsOoJW0CXeKGTetJ/3onOaWhKf5dV3D2
OOopxNgr+asv6sXweV1SAdK910v+zHWD/dsRi9ivhwHU4F+hzfgGLTLtcbhS+cPV
eshAZcl+iDEI2oXKKA6ckTIVYb5IaCDZ7VTVpXpkq6KaGbyalMcoEeI5T8DGFcq7
ic7Hqysz7hBJzdwXZYk9hPx3Ov7Dg/4UBZ81PXzkCfh1oN8n+/lRz4bMhHqO3wp4
y7NadqOOGjlyQaPAmQWD8I9gK5rWLa1KucLqpuM+AUm46NBm/C8iao4j2WGTwz1v
m16iaUv06vmBuR8Zmhxv9dPsjOgisBAsr6Ex9DMVdTZiG6tIGlfXu6hs/UZ8wICL
iXxOdFq5XRYru943pPTRqZipBZFKdX93KNRQ2MhqoHEkqHriVwxUB1eBZyakAKUt
JQUimohpGJ6FxodIleqjdwgp+U9PxA8vsGQZn0YINRzWBhjOIXDuzRMSobv3QVdi
hyBKshzwQGgIqBdJeYX1/zKxsFwXqmFS+2jdg7566eUO/cjKZOvPF5fMRGrd2LGK
MDMRF1XDZPeE9QiDfl8C2wdKkPR3qGHnsvlOxfuEYmLzgPo1ZwoHex/YBRb/+5sc
tl0HECSgvu+ALv0Xq4wNO6v2LUyOpYhno5RrnfaQN+18O2NLfOIs1YmaTMl3Rjx2
3S5bcRem5qyd5BK64SvDkqa7o05Pfbincwdl9MMCW0T5U731hHTcMPUl9bxWWSvk
EG9luuxtTjRi3goGFmweFZ0E/RGVF1owsAeIFGdaGiuz5MFQ82V8r8twJ5tKfuuJ
p9czCMBegJ+m+mXpmXBRBdVGw2BgD03mJfQJm0i/ucLaro1ivYsZS8X5sQo3NLGV
br0tSI2Jt1cxWh53QCbzcyHEr+1MyTrxk69MSROa9OOw8+vLpD4zUioZTuR2aDWX
0l4th23l8ilO54hXVTfAHRVDP/zukNZ8VeuQPn/QFeEIPBY/gfH59sQeCBDrPf2F
7bA5NUsVAiuzBVvUVmzOxq8o5ca8MnsQDtUGvGtVBvRBVUtd6hi+5i++/pFFDM+r
CWFDrKHkfGN28jF9P3XWE6MiruKpoR3HetDNLlFejvlcC7gpEmjqPz9ewKBLpv8x
xSuvwt2QzSwIxvH8eg0f9x/2kgv/yZvhtBucHHfj/lo9J8Km0GT8NYbrNJvnQ2nd
T3i9l+Cy9yM3k+Lms+xIhcfwwxTvIGQAuQorJdIvNkI9Fw0XxgC4jv0kfmw/BFfL
GId8JnzSg4nUGYsefnfQ0dzMd8LvEwfeqVja4YyrD7Qu9HJZqmHlMeWaJuhNphu4
gbeUPqVbac+myggMclxEzCVH5a+TSmqTc9eVLcV0yTWK+fYUwM8syU0uBH9Qe5kr
vI+VZCTi3tgHnLiM104zVKkHzuvD6F9l1s2RjMOy6O48rpaNJvKGApeVd2xNHT/7
MBJguxEzQ/VpCAwC2D6QlH4hcCAbO8bPDoUhI2eTmZlnLpbUHneBtUlWlWBPhsxa
j0aX4Q8A5MkkLYRD5e8zjjuLCoXaLc+0S/g4+1eiZ2sn5vYR3VZtPH8+DAxY27c1
pCsmeyBpfgwmCiWXAzuNFFK0fGrJP6Hru2hanbYDZWnohoS2lDSXfN4R1hnOJ0jE
SSXXxZdgOptQ/nn6FKMeQT2PFn/x5RUodudIhT+QkvVdOxOLECso/V3Pd1A0Niiy
kdxR0bHAdv8SOdikI52V7qK87YDGH412vI6M0988ilM4PYjVkC5PsbeM6mMFjRNp
x6W3CYfwuhWOG/WfXH/QLcac3V2vFT3V8uh/f8J9M+0oCM3vbR+WoerD1tPCsa1+
F94xYzCU8VN+EZBiwri+pFh8LoOiwYQb8cMW2HlAc//PJLifxw9xTIHPvSSFC+XB
wpsAH1m4yjJMRznYJi86Z7JW7cb00StpMYJIRNkSPaNf4OC68odXlXl3Hr4Xo4o8
fo2Cd7/7k0fNM9o6vvQTf44Vd8FTjCVNxLihqTbqMCRz4dFSlElQ8j12oYjSxylY
fKI+XuMYb2UxYwnDJn3q56+uHFU43CWNSmKrMrinTK8WCn4j9jWz0Sf0tzI66gXd
LdLYlzik1PJDlhtAgfv3jpQ2lJVlxAykA/zePE9XbOtvkcBHc1/flgyld+etvjjX
chSeGOXNQvcrZF4xmrV+hoO3+Lz8msv34w97FjLjzQxM07l64NFAmOxQyBSS5JiT
ey5Zu7lpYpnEK5pgK7KKOgvKnqqTonI3fB6f2MD+Tpo23V0sF8HshB+H9h7zJVTd
LpQWmB8CFAXgYBOo1sSUIywETxBQGq1yc8ILT4atLAxGb2c3ALA3OwZOOAcbjp8L
kGqCoYKpeEt9XlJC6ogAr9T43Yoyhc4S1Js3DbptXa1D/d5eEQHCCth2OwOSLQ2G
vArq0RiRFoeFzBwt0PQZD+Msv+tQ+LUgIqS6UfFrDvX7QuyYzpj8YlSYyeJiCXNe
fyEHgZyxVzCbscOSM+SLyrZNRTE9Mqn0GAzT6mHwoyFtoK1HDG7Zrw2jnOiYfwpX
5n2q4O7r7DYt4ljHceiVbKOHNK4fd6dbUDcevXjTE6U4GCaifqGGcELI4qidtCBV
HzshjrZuj90RkukIyX7J0+k56tyISCebeRLh9RlPU3z0iJj7ZE3Ni7m2zpzE4lep
2LMchZXGCSlgs9NMBI9ItqcKJ8mgDWb2ox2TZCLs18IRDE0cZCFdujtgIge+nY46
u7YpIOBpnoeoyGX1Z2kbJgDEP5aEOqAAlFFVqMmY9N5XwLGyynZZKBD5LaxXdxXu
ZIJU6uYr7T19oxrWNu3RNuIi1irGSDvuy2AQYzddmMwQGKKhuFsq7dtWK2XqwvIA
xb24RRMqRK7vOgD8OZVh5yAZ2LeCkKepcvHL0QG8QydoJ0Gn4wUjItr0xw/Rhkiz
doSXV1dfi6UrY2aeHlu5QUv4io7PV0a6mRhW61JxK1BikJLBRnDkVBV8GBvDrgYl
JcElrxz1svMLYngY8CQ07W0xRKAq0Wfw+v6lHsY8U3hc+T4twdfNH9+GrjsIs51I
Ee1x8S/7xR3gfSlblVKHq99Eu9SyhXzR7j6XObYTC7KeKCAaL8GL5J4kGfz7wTPr
p9qeqcoGTngy+if2QNr/BDIWkHDX4+sTQUG0TQ1YXmJg/CyAF3kDwmR4IMWKYmm9
Jyv/3XByLgZ7BdxIWnGMCstrhuptbAkbzIAAVDeB2jFTRWST/5g0AMAbBroQybzF
ke55MhIYThvaUJ7Jypu4CyaBufJIy3Z3F1Z6IPsrOLd+BPJPzm3ytlSasf5wlsBr
1QkrP1E6zhTwq/4RivD75bpN65ldhO+aK+spWb9kB1N3ixa7KNAtbqjn3V5zSaz4
nu88T/HcqvAFZul8bPPtup3JNxBzMDb1YU2gVbchpMLWp3pDLgC72vSIJcqfxZET
XsvurqJJKUqg9AJD/cm6V/E3iWaZsU+uv+b1WXpNe5QWqvDvMCptZmIbVvu20wUC
vKNoCdxTpAVraPZYWv/L8b6XPo3Dv2Hv8pwDyjYUaJyBg4Gpep+Eja/Y1AkNtXAr
/R4QgdmHf/ktC5wErm5gmBzi32lbp3LikgkoDZZsXGyTcrow3W66u3n3guDhxhnP
XrT7SVzzKX8daidpckx08a0Rw66beHgBFN2OdptODjI0SYiezDANi3QYinvPHw94
XA7Ghlxtrpe7iA/7TNAZe7hkLK8h93MASC0jD2gzTZ5dSlhUIHId993uhxuc49Xg
Clo+jmg8uSghzwYygIMRRRKFSt/BYo1JVtSP0A8m8u+q/UE9qOtq5AwdWQRhmbWV
Y4Q17bWZj2TdaOLi59dNQ5t+qiwhtlOa00VlhrqHmx9anfKyIROINNIvPwPRRpyG
oyDdb2Lrm1A3p+VwJeV/4NkY4jkO5fJtwQpaNdGgc9ijXfuDpU28dKOFN4FsPA0t
C9s3o5GC+0aSsXM1cTzdGcgXPWey1qXyOEZSTgw+viMpnszUAEBN6ajFnciBxSon
N/zzEP1C/3QWB3Em9zAXafkJBHESptR1Qu8m3cRKtVzx7dmKcyWhTcsrjvuePGh7
G6hwkMjKqc/xg/iz/Ffnzn155G0E4E4HNo22gAjGJcWOsetwitVS1x1xzQ3H/j9V
NpX+dAiwJbpGzGYqdwMB8J9u/bEvy3a4pmvd258hUCPV8E6hsqG2xr6Hdpbo1Brh
okGp7VMfWNYqbBY5dOadDa2RT0LXoHM2t5G0oIDCay2SK5LTbFzkDCtPxn5xtTXN
Dbcvfr093zOOxXUth5TgKtMGNlikYF8iAaTDFVRWeQLTFQM/Y2dAUmarn4AAWadX
JG0233yCTZrBR1xNj04aoMyAdhcaSY8Olo/1bXVy5KJR/poZhF8MHepAOt08s9dS
+4Unrq9Fl/ullqedWHJn3B6J4NDZvHRROj2LQ+cCx6Fm4iNaetBzfY0lfmuJBOXp
YNHWWbPjsAVdpwjs6oaYyAqDFoVgDlf3TBsfePa1m0FoR9v+FKIdPt6wP2BtkIfe
e3eXAKBWb7sVxVN/eEMvWKJmEhC9ms2vwfGu2bbHLJaistJzA9eS3HML5/X0tuwC
LyW7yVofv+Ik+EwMQaCPMdw9hfbGrh6ltbBj83Eq7dHNwbyZyd2GbBtn47ocls2k
ZnrS3JN0YVvJDD8JCcP8/zs3n9ro6st8w9vav4qi0GpBCL9rb4Ii5EV/pB/59/Uu
scbWAWRLkfLZz1Z/v2iCnIxHNNgjbuFm39+rl9975hLSjEdje/HWzXPZYXL5hlCo
Dpn3nBpokH2kQEZFCe5xPK7hH3Cj4SmvKa4v3sUl/YSEqiJfSLQxxFkcRwZz+iHq
sVnI9Quym+YXfJqGyowzBcda9O6DOp5EUgvhYgnE04PrU75shxkYkdVVTeB2wVFZ
NYjl7AF0cUedFeb/2thRtw2KJig9i/JjafUdV+lgKUzvAR8Vocz3zGfBS+1GTTEg
zu6/Idb4CUlVkIwNz7XOo62BUKTycVGEF3EtMrvqoepuLC+pbTnkZNq84fQg6ThT
A1V+8Q13Pw7QsofcCX2hreMCc5Jq4TAFWK1isDV+n3gUIKtRcoK2lRw4w0hH3Gp1
KzlrVG/MngbOsnoObAPNMIJ4DCfa8mHnyAXKn2AsZ+7bhPhZEv7cZjPylz34RnmN
DHr0aF+lNg3X+wrLQPKG19ZgyKra6xpeZ5yIMugJ+6PMgpCMovzNVZuj31cw2kvT
k0ZCKDeui1A9/VrZOlX9vtgRpWsh9MxmfkkhI8iNR/eW6soFhWr13ZmEFADsvi1w
x74Yno/nmXsQNVxJWpotNfsyD1jrOXkqc5UAGOn/9VFWGu47r6coT7OuZHUho4ib
m4/X07D6d0DRxhkWvZi+LCDkO9UKZAd7Mku/rqWWC9UcYaY0aHPCcEKstxYrL+ge
Cz2vXcmIJg8eNUvTsT8RXt1EKiYs0FJbfileoI9gb1yUr8rEjh9ilxTm8nQs46w9
pe1gOzg3f2E6UmMKYK/XEGlSsz16FbNAlA0jBvKaTluXu5oJuH70SlCVbDT5bJtY
cSCT/NjaVXRMuS6kyxRJBVl7iysDvSzdF66f0nwzZGkzrh44U1FE6B8v1529SiIH
2DYk7qodZRtvcQj5BK54DtOZRm0LdokTE0Xv8e8L2SXn0R9vz9d5hK866aFLqz3f
s+apvydKEDgU4GJczjTiqBZnN+C132eu51moc7/DpjGpx8a74/BGTKc/CsqFbhd3
5/WjU6ebC4N14F37a3pOcp2sO/5WZEkvU3dPz7QOiGTYGaxqgIbQOsinTc1LDPqT
BOD4PtEc7xp9L0o/uEMXsCNN+I0omwQj0IGpHQg74TNsJp/inI/nHIOu89aGGyPX
Mte6QTQ8b5Sppf+bSvSIW0tlmHQN5akCwZrtB+Utr/GXxw4V/PUwC4RBjqiEutUh
MDLDzamMDALevJ7PXjhC9Z50INyMVMNOexMoRsYUVL5YPP6YryU5lEkiakeRu78y
s96eXEXGjevGTn3f1dAKxN+8XmPxri5LgNgac2j1jRam6h9CKlhzZ4yaSD6alg+Y
Gca7pfcgkV0wX96Ie+sJrx5kFD4ZdTpzpDLZWPFjtgjLefsReGck0iXByWD/yb7E
t697N/L2aZyh43TM5rYxsj+MMZlqjrIekDi9mdY7lY2iJmn0jPUD/Du/3aJ74mmQ
MXlAaZmsxTot9yxXk8AbOncBteemDpcNhMxesOWB1LgkH0rUp1kchn26Mv+VybwK
tmyqGoIHyorGtXUi+3xgvFycuY44IYBA2fK770H8PgPcSNOd5eZAOiZ3ecnnUFly
IBKKY4WWiqdvXhdkcXDXOIWeRvJP+cgyg0ELyAiNELdSaCPLPvnTNxiikxCCYZ6f
zw4N2niki6GltEHVIWtJgawqep2pr8412LUYM0UJ5qREC/I8x3e5/Z0gZ0nq1wXx
eo2bMgDpCjGBaT6vVc8XkQUY5If/tS6VfkQ3JxDKloGEmcZKuZn1Y+V7XiXrJ7rG
bCSvNbORszER/OVo4VP7EpnCzS1xR8r6S+xzMjeaQeWoejyV9nFREhdRsiV09w4Y
UTl4OoplmLsR9Hw14TPtdWulJmqeH6t2EXaYllQpdJPpBEuMNMuTaHmnV9/2G2xY
v2Yfro6D4oTbv/zdABpOcXYiFXohxuML67ypwVTBkWi7F40nvdj1xEZXpsAJDQK1
CyGyGbFlFhDmlzqD3sRvu635mH74t+M1iB0Ru2bF5ccmsoal10yTtAJ4EtXxdSQd
33zdd/EhTPtLpYOV4/AuoV3SEQqrrqQiYnN1IiJ3UD+jgqckyX96JD0QHLVIRReI
zFpjmMKLOen4L1FTN+ZKGYRUNGBFhM2WVo4TjnKa1xch1+Vwz9T65ZplTiCMxMo6
uekY5KeqSAxgM0JQLaSc/hHDrwET6aqkzmICrYouUds47g0SajpXDg/MtLqXfXOt
alQ+TCxwMlXcjxQNLmDcgBcEEyUpMit10S3qj5jiioYm+xXYrh12unkWMONLuCUN
Z5MbV51vQ3UVhzML8HL9CmV0ftIMmqvVAJYq5maYW/JtpsrJu9Uf8YW1WW7aRJrq
eW9VRdEW/l9IIN+nNK57cQGARJ8SULJ3474jOurDn8emfEx18VpVXTMGy2qxHEpa
vGi99OubOIX7RVkbID0gRcN6G674Jo+RPGoWnKWkV5p6JI78yebaZDJBWASFnu92
bo9cbFfzmb6rpmFKngEO9YAMSfKIqBVHmXpHIdHOJZ7Kn7sHxQOtQkGQ3wRWIemj
9kdQkqCxbPA+GmtqRSScympav+PMbWzhcboYgjQ7zMETDap4vCujp3tWkR+QQTzF
UyC73xFCrGoZXa/Lrt/4jZzzIL8Lt3i/vKvCdAS9jCIwKwXkoBRlq1bdHJZV22xg
pPY5SNeJnXJTOD0SVQJcj4h1ZmbQ9Z3VGbBRvQQ54NKBkqaQF1xH24gZww7Mqelm
YYElxrkzE93GkRpplxZeki+4KFpH3eM2lQzaBjJ6EwEd/i6BTQhapsN1Foo6ikW6
M+h0JhCxBkS6b3tq8wwe8m5Dp3vY37P+A1RydjP+fuiZhu/qyd0WM6Z/hrV88yvX
BJeZNH7AFl5zhbHUWzcFI1QglKMKsqjl4veG/vos8l30FlTr7Xi8IeW9SZLZUQJn
ZmNHpVR3c3xgDNaKgbu/rm5QzkbCx69OCrac1zaflURLVcgSici3huaROLe6DTHG
GwNk7Dinw+y3oABlFx8TR/4Kg4Vt4Ik+QO8cugDevg8aSVnVC1ur4J8bc40xM7bj
b6BBbuu07l78ZhMXONXIYsycvCYgAoysfPuqrvWdyHdKmGjnLfCVe6gT7DSubfi3
Lp4psC5uRhcVNOC9KvG1PbIUXUxuXJMhUlkhXzykhmYqX0Qbse74CgXGFCd+0yQO
+v/TYjGRfL8pcJVfcpyUUlvSWOUbGL8KDIWaL2SVWit4AxVm7nUE4CVa/Ujz9IoF
KD3d/0OoL5SXmEJ4NvLwvy1vGj04GmT9U6iwlF20bNDf0lBMfmf6yE/E2H2j82lP
JfzrPBiG0X43atlqTRu7wGtj2UIEqksgg+sJgnVvr7m6IuELrjvGQEPh+AZNZC2X
yedDY3ECvunRkkGRO6HR80qYOJFz9YQWdiqPaNFZjvlvULIRL+iLvjmbEzdpbJnD
MqTOBM0/MSZrL2ukmS1Dzjf3YhuMOAOciy8kEniPNGHN4hB+P8Y1qQneXiZgf4lO
mReorRv4yW+COBYQDBDrVwsH9CYowkp9KK7pnbjA+RvyECKieZ7vHnX71702vJz7
QpEricNSZOJNFRzyehBDT6St5/fy66DRFk7Z9AFSI9nNiU8K4iIrtH17r3J8bC5m
gzlDJkPUH4SPE0dteIOn3uB1k2kZXf0Vp0BrDEnzrN2NTPYfKpxjz7hiJL20he9V
VRInzR8nTRcsBrbFzZJJ0fmZMqbExoOkuFGhUXUosqGZNDY/SEJU2bK3ihL1knlU
hi36DLCK0hTchzAfRNt5iGFPvriDyAVghguGx3yCl8kotoX/UN7QBIFfcZigO5MS
8K9QuDtOgaz3uPPYS0syHIxLUnfYHd6kiPwbnzP0bAziiSbg+o+7cxWvF8sZdQjN
BG3eRALQDhL1Wc7+eGN27BHbi6Hh0siFMJf12MAcJMMZVDGze2WBArxBM5pQMKJp
pyTWGQIyD3t/kYN4SU/q/h2u3KnVOCy0NIDYY4uH+/2b/ENSLo0HfqEXBqQwD3k+
J8yQpl+LobDnBS+bfQWGdCMjjRWhqilC6t5/BkQ/XTOZheEcQEVfGnc+Nf4u+lP0
19CoT4ASoC+dvVsWBHXDF1AnHbu/f6bPJwMNtqIfPKfTUr+2KDlUCUEFigQZg21E
MnBsVKTgbo9P5Y6rbbvY4pa9NTqqU0Zm+NMpanln0izmZIya+bqzaPcNON56h18G
C3d6iUQjl0AOJVqhMkUuWZaOvhes29J1hYxP0fYx12Q/n1/bJMbD/I86acuRn00r
z/Ekw0MyLIBkg9vwMNp969uvbxPFqJyDdKUybO/yxIav4BvuhD68bPSdnOGst7ez
jE8rwgX67FxeZzTgqWTIsI93CvP9biNtd64Vk5HgM4GzGLgd6Gh0fJsWXvXJ0yRx
Ra+okI6ibhLOTeK1x9n35XNO53MWLG5bZI1QhjOWLGyxxFI7l9wQ79WQbqE6MqKJ
r5VKhLshx7r30Om4kM9GO0RLn504+suU3E7FYnhr/obWXqiresGYwYCCjuockpi5
e2jYUB0DyEzmiZntnG7x7cVy0k9wrRQo6V7oNDQ+qTAcXpwPH2ODS5W0XyakfmCY
LfcgVKvqaCFA5kh6cFeFyKsI+qihhHp8LwZiNFG6DIWrS9o5M6GJmuQnY8UV4wAq
QAmSN7TseTb+wO7fdHZI0eYQT1psGd7dGqthe1Ucz9jZMm9JrB3T4SRQAhzyL2+g
pn+xUkiqn0Glka79SB/4PlEt0Oe7UVyjdeue8vexR2llMXFgHl9dqBsWgdA/mqef
3CP4r6odsprPiXt1lPxDKn96tW+jv/m5F8wvkH/JLAaV1txoMjZo+3WC7+Yu0Gny
uya7nSHlDfevNHQMFP2WMRUFcMtG0PRB6dhXXFOcwCYiwhO6ybHIrPa15hQJWyGs
dbqCpzxuZ/YB8bYZxkSjP6CVfynD8lOYGM3NvUYFlgWrOgJwX9/VrmkpY486rBUL
joUAg6BMhZKbSjEARTy7vL6e/EZSyphCovxdovzN2FuqEWGgVc7kL+Qa4qUo3TZa
ta3pagCyj6mAnIIrxaeX1YB4aaJQuU+BXAfu0ychQPlLRmYghacSXt1KGNDN8lOQ
fdfd48gjlWy5M2L5i5EmlsPWa9ZkxxWeVmR668KxqGzrAk9VEt6b4OJTyFsegz2j
6CP13Cmk9EI/n9X1ce02GY9RHmhmIzX7yu+eR2HeInBsVG5/zJXmTuCfE4zqiC1+
a//1O0Jq5OYJVqmN03Ave9i+lcAqGWsU/c3JELuV5bE7fIheqUKNdNbNOtcb0RtF
xh+IuQvEWSWWOA0+icjw0yeHtXBhJu/pO1LDvw7CuOD2Dxqwcl5NKPRMcY9Lqklg
YsXQwrThAOl78iUp/Kz3hFlEXseJ6qhC/dcFI4mQOkxotwhpeuPzCTqVI60bNePx
s3pPsC80/84qGbofjimn3+NHCmc+smX3wEye6/pbRkd5YLYgBwfg0/OvlZkXnbPu
xGpZNWBScHaPVYr1PIVgPNnDcvmeyioAUfiBd1z69oMCDv6NbTDWTxNIcLQO6qqL
5EPsnAmpX1IwOgM/RABzK98ynTmcTiF3V1mXUYUrXQGHR1+PsnUqeVtAmWAMoraz
eH3R7sM5aWYlUt+NEFOFkyB8KVDBcLvkn42g5JZ9nRkjFeXaVX/Ih8lZkmZ1lffp
KKizxSQsLyQWQ7uW5EB42DVZe2RCd/QxeYrxNyUQeaDA8hE5R2iqnwZT3H5fnJqQ
ACJoDREszyPqh/VzUHT1c0ZB933mgxKTWyQXDDPGwHfKxYn6+NDrU5toQo+g4WQl
MkhJ3oCcG10ys5opeeK7UhtfCQkRPOaHAWxeAzmrmUzDj6k9OmtirLQA1nLjy++E
tGe0+YSEP7ea2K3xzijQTfrEkTPBAf9SbTO60Vd4A6UX3Ef54NsmY418X8zHEVyf
FLsm8SshXh2qPpsIZv4xpsHi8C34umw4HLeVZH65p7pQ/THiRldX/gOOOKYeQMuJ
FyienxadVL3kZH1ocQjbfUcwA84QDG/DXtPwENLZU2aMXYcRL7EhiFABmQvsbHpf
aeh9wlOkZiTsbQpSBZfmy/aGSwmBt47kEfw1sPQl5nI5okDwB+Vg6Gei2AqyWl+m
DisBVSrHYjSHjunKd4OQe6E+su8MuRhHvVuWwDvqXa+R2Sb4X31OaqFkmMB+EAfX
UZRMHjnDMFwtSRNwQqtU9h7ONx9OPII6i/ro0/eXi70Tee0sUEZp82iES4Af9j8a
bxL6CSuCahjDsmMiaXBRWrnCsVHu9bfndhI866aCVQbcPA1E9qU5JU/Sj5s/+EgI
QeIK+7hdr6s83YX0VB4dHcGnzefelnk3t1eh3R7NloLj5W+aTplWVjYBz8LtQ2bL
bgNM0ZbOJE1246q3WLFfFpBA++mlyzUk89+7HqL9SCJgU6Lh6yeNTJcgydO8ZzCL
XDyAeygU2d79Pos9eOxUGOMmuPHcN7f50pJURMEtddHcs2v+F0BvGo1zsv+L+gWU
SjEd7BBSFtiMSdvmuldHS9wvV6Y5l17wu98XzLAPJrK2PnXGzvSJFbdtYDvgwam3
K+pqgShd+RDlGxSeK7TnX4wiWI9whc/3bTxyBECGnkH5vwtttemDI6aOYBWxJhzN
otgDkB6cZanm0NxVAcVBdFL2b/UNpni2WJv+D9+/8jiCaZT7ZkiRktVby+IKkkjK
/q+gp01MkeWAesaTA56F7HL2kuWwUlV7Wr1/RIMRjX01ToxcwTdeAiyPDiS5S2sr
+xs2GxNUi9fSCtSDgqLKRHc82f3/0wGGxoJiy00htXagboWOF9uIFlxE7SaZvyPC
8kjAfKXQ2LGU0r6/Iz1KrIWho4pDXOzX1TWYEge3cjNrrwxkKomQK+PaQZ18q7MF
0o8sFWXvD+OjglBN/ml/sSSuMGZxNlZ8gUxmTkmUbEpRf4p07lDLFPrj7M5RjLhl
Y9AEgX7hdEUK9OoeNVtPOOlABmn62Zu7x/HhcNbjP1Erfsa11EqfyymxCSjk7x3c
skKsTSfprmVuhDQGY9Oa7zI9zAxptF9V2NFBv/yC/rhMLn5LZbSW1eVFewCo531D
iDidQyleQJc6RxCKfkOSmQgA60s/AA7Od8Dt7Bd2GqypQoIQymMsu+qahRHkR7zh
DcLbO7WLgKM03aGeAH1RGPaWNq87wnLc58NitGR9619fhXoIAQLQtZBYNBez/3ae
VlRDlGGsN5p/uF0+HTMQj/5jYNk4bdysA50Fd1tMxpvcYxtxOiE9d2W8Ysfu3jxY
lZYCjugYD5IHHK2s/Ezws82It2JjT7jFc+F/Ho87IGXtkAdTgLqEEo/3D+eG7ZZE
wVf49VZ7P3r+90mSdg8UmmoTDFIT0W0DBHnVPMDlP8I0DCFsD07EE5P61Go6OpHe
2dJdW8xA9TJzQeSHDWiGQ+1MLmP7Vt5qMDedgluBUCOALkTljlgZ1tBvdkRYjvdl
sUVEMZ/ySHQQc9CjAyvmPQyhFhouvHPnk9DLFc9g2AhANv/JZf3IjluLnm/csfZO
ndAP3Hw0l4GNHw5PIKTW0J2j1ObG2e7PSLKcBqG9CnkXzs1MAxlPdjjyDoL/HmNO
/tTq9EeAMobHWCigqCtkxA8Y0X6mLG5qkvdNGD4gb6pCynFRSR3M0rCK78zgW5P6
eK/TsKmqHjFsUWePyv7TtQWR/6BAt/9NMEpFmakCAFUZOhvy0y3eqwED6jhDNIik
JIn8HaienEom26D6s+AQphet5345mC+prkznWUUq9Kgler9JnGKPVohacJRnUCVz
L2/YAPt6kJLzXZ/8hvpn9KVIbExT6UVDwNfxvYJ8l8CTqK1cnUJr5LF9NunhNSTK
8pWOjvflrXJFjdArEeER9vf7ZFCM9S713fIbX2dEIU+t+CHkIJbqycC/1/zBjzxH
w3SexpBaT+S1iAcmTMtrZWfgstzFD8VgorLPIZoj+oH3yvO01bbTTRhvuiM3RVeX
mOq5bHAWBNEByHVYqiLhLKwgFW5qJfb259RsXYoDRMlbXu9dyeb2NRtwm12Mpe2d
VHGxO7BDiX/n+BfPMCAP8haTc6wqWjqZ9t0uLkZtTVH9OHJ+HGVf+OeoWLBEEqxY
BtnmhoSYK5NvwzAdPQThIojSpoI4or4lkPBsgWc7JXcD0QrFmHOX1cWtvd/Spbl+
8Nfku4cvT60KXLJI4nXwv/OaKOuPKcl8KeFxwHYcJEtiVVtZhUBvg3BqQMWg4Pv+
GJVyZtiLVLLqdPh/zCKrCOZhZRFd3Bfv99NVRv2q2YJTx69NQnbv6ZyEjNb1d004
3Vu6bGTQM1KECbjO7kucyUBF0y1q9izSSw9gPgEH5qjtd4pSL6si/RtjaeuYPPa8
zJ2B7LF1gsiZByiWqbHg9R5s+ZxTM5Qd/SfXD+29rrPjH2cRrClEjYpaLfjQcsid
Tnq5n8OeqPf6AgQJVqPmaddp098xsyXS5h9Hc8ewvuo2aGAXY/apABY0TvhGvfJ9
9i9EskK/4q3atHF9Dpr/4Mo0UoKHMPlZjaOF2vAhQMx3rs65RTR0nw6h10788Ub2
fTCWXZ8ihgzLENJABV6UdrawhXEFqFgrcKegY5fuYsMAQV8pyePHzzjL/YeH7xPx
dsveSEi0LevCblIdFTfgjc1JYZH70HBESr8+8+D0nXBGtAoxcNAlfq3JiyQPhCnc
NBOaoynIqoixO8bujGDVZ5/olgbBmi3jYWNDQDPaJAx3YspOb5M0Lg1MTZ4w6T3F
BV/7JFuq8YHBZV1KNQfLsX8HHhPhK8iQowB5desGDuMtlR7EWNNzQXWWuURtSF3b
E3gGKIrnSSyn9RY7YQNhBP6HY8uUYbPNkqb52WxVF0u/SzcMkZIVSUWQHTz+P9Z+
OaIRaXO7YZhtOkEdu2ePhD1FAb+NB0GmJG8X9dD1MsmmNRdawjZ9aCvPGmfrdvnZ
Y1W9seROVVu1ijcsd9YWUzEuVM1MSdMKo9VNIUd4ZWVWtrDkiM3oSXEdgw2WU1kn
HjqLiBOuvYePUcu9uJdzM9sfqV08ur5ynO5Uj09OLKZRHMiIIeVjbWGTTFVAS82A
s8iMLvUy/C3Tst07oD5pbL4/y5OEOtLWgyyCGGJC8bnm6vXBdnaYq7iHnc5k2ZH1
moo2kMoUCLTmUeuhAZBPD8XGVQEWJjtM1x8nx7dmbMjkammVqbQW9nlT2iJidGD8
H+ua5UD1vx7j0x3nX6v/xspomM7qBn9VDabGKVR9YNyc5srLHDZDC7bKZ+zhKq/z
TCnVSc719kTreH0veJtENNOvNJRCRjIs5aAzsda6Q9l9QLzZW7cd8lKoKn47lH5G
49tzY7HTjAeJyYdY+OJVeAPHNaEFcncX1zLYr3jCKlGd5M3hvBoo2XB8T1AExPP2
O6Dk10k++cAn8Fjh4Po06Pxfj9DWDMli68+zbqrjgsSya5YbhPBCX/tp6r7uvrzs
tl+ThGhJdzh+VQMimcdF23xUd4IJ8AWv33uQRtAJtPvf3+uZXDVB/fJRZKkhST7O
YG8uQJPyXOvTeA6eM8UaxnYfUpC1xuoyOBnd+TRw9H0tAGdLtQj0OQp/Xx/be4xG
WwofGHGOAy8K0iH/OD5LqA+sB34KoIBTUuEUCdVahUZJATb5VFgCe1T2FETzWIv9
7QGJq7aQCYYYyurRhBTuaahiWhpdJixnD9BAATR3At6qFybl5DTtd++FvnOtwxOk
ypHk5YaxbY4dIXL2nRZDovmPvz+noGYrvYKWHwK5vDgEQRQvGdwjAon9y8TvW5BI
kMpWwu+WjuRiRKfMWHSASixJlLfGsHbIvDaegJjLM9/1aVwFRY05Y2EgUBfWmike
7WiiF2ymAw658G6yeiuD/xex/jpH+f952vch2kchoTaV+OYEx/PD7HqZc04S7Ogp
pH3J/XGEp0Y5LrhHVXEPo4Dd8Mmn1iuQOPM+XKKM4Uc/t1Oxkabh5CDIWd4WoUv6
o0MAvTNKMsjy1BrMAmsQLHVIc1h4yyhedUifiKZAvVuBGmVvlSjXsP8bZt9rvKxo
1velaZQrY6ANRK0/XlNDk5wGDCu9Stxoks3nKn/4JrYLsLSAiUt/uCuDqQWDsf4n
fYNkApFMHjWVbOl7UyGCnrw9ocxnVtWSKesIf6h0Lpc+zpFKpv5Do/P5zNdTj79p
RKj6s2AV40VmwF3K6MNlv6aCb+Zd+UIcTR4GE0nALeBYYbTsKE6VaTPX/yaCcUZA
6ssA/RVLNPzJM4n4Ao9bvHQSDR7gtjpO85d1k6wuTsPGZOF1wgj9EgErrbhftF31
bjWiq72+KA+8Sh1/FilLHqgUY0puCqJl1DaYSOOe1DoZYXeh1MM0n82Oc366LRcx
/8vQSfk8TkxD87p0VET4BX1zHPV/T94O3b1GJBuwL6sztTDdX9sp0PnlcXzC7Dmk
e4BetsFeIKzS+Kgd4FqFT7izs9E6dO0pMd7qYcmmwWquE0kfv9p3+sKGraJ4ozNU
AXoRjloCmLwRxfL/3cGEFGCbBb86xAz5GeVUQTuGNjMqb1BhzFt1QE1p3im8Cws1
Cmkj6a7q6itQtHsO1ZaqjRs5YqHiM67ONaWXeNxGpTswmb/CJwvP5dj1v/BeI9IU
cbyP3i7t00uWQOXZK6DjmHV5ZeDzm4S/XPumD6u487SGaIkbt19xzBwJZPSlMWpk
WD4jganrWd4B6bplNrkm3R0BjznLUvH46GMAaPsXBsy+hZVoISlzr8TBElu8Squ+
v9wt7v3CFr3cvUsjDhVg7VoAShyap8e1uDbGiT3s1R6reZEu94n5lutadxG/RHzL
WkOPJFdBWnSRKrKq21Q4VCltk86FCOTZMUk+rfIFAizmrF+Pf0IxclNyq7bD9ZnR
TxoiPUzcyOrbtEV0xbZRSy3VGFVzx1/F6LqZs0QHgUyPXcGk74FFPzoPTPEJlrJi
iHAfOxl7NPyHLVh6JqYSLhF8Nnx3vFG44LpM7NRgVh2QiXLxdQLEdCqD0JfrW4hF
i75/P6CbFMqI8s4jFDAJ39FGCdPRZAye1jVsF29rJpR08o/xI3LtYIg2dzpAc8yP
4dyR77J/HyMmbeS15sVa4IPM27oC2TtzO/IZXIlcFqJBA6mJ+TkBb0c4l12DJFG2
q/3hFN8zRsJkCyMSX2NxepommG3OdJuuDksquYN9wlyhCqaclwDKvp/h5SMy3hOF
P6KPtCy0r/+ieoqc4jz2Uj9rDq2SqR7lw1dkNe2xZVYHUPEDfLXcSVSB7UjaWtv9
Fb8ZvwKUS8ze7cvNW6OjAH/D+KJPkQoYnbewoXjoW5OOgWu6vbIVWIYyj83Bx367
mOQbySMQ9yAvcthoaxTrUjBQTtd9kXyEmYbATwd3MkoqMhOjQ5Q9bFQzsIbCcvZM
BedAaoat7tOvhRrDzh+y2OYgoL36QsvzYACjkHEzy5N+Vs0TO3v3VZb6Sg0nWXh4
cx8UIoLmWz6ik070pxRkPN9Hpg2XqnkvgL4a8QAba8Sk/wxSmBCvE22QV8hawgta
Cc9w71qzyW4Hij+qwxgZWRhvRD7pjvEG9+W6JJAzZN2X7fAV+uS2O9V+bRYn8GAC
JaQjbCn/xX1KEwI3mCDxRSfUayGoV6ApkTRvMF2mL/5lyq8R8RlVDB4XhniOtk+1
gCOP/6s/8StDv9Fe++FbnPMsUEsfB9aEL55+vZZ32w16mdU0FIOeVQn0T9/eAqWg
DL+j4hqDXA2f4LEfIgVVaC1niScgqvXqmhiOM/MDzrX/Vw6oTiW9ZtTwS2GK6Lp8
lvdEKPOvZ4fwTGL57aJMlCB7IEs9/n2OfpyhGJpm5Xlp8dVd0L3fy90WVgbwETAO
4299zaSATiBm/tci+GVVthbhov9w/NpuwYH8feCAUiRkLqfdY8/b0LwcFgXBwK6o
RPEDjrMUqUmttFndUmOWx1HhPWeDZ9eIlhD2ZqwFwzXMZlQjPjmE/JgnOOhpdnU2
zE0DoajtbW/DvkCjtHjlWxOOmdRsmLA308L/+oGD0uTTB3tF8aDdV2INyjRRaVgh
p/uYWmkPXN3wJVV0tvM7dOjSd0o/cxIszmso2TkbM//YsDWhBGGXn0+tgfOkaj5C
h42RRg2jJdNSXxXNbtJZBjGu+byEAqvaAo0tcxJ2RBMT8enrMJ4Sp3DqIuryZXQz
cq3CuOLFZKI2tXWIFS+Zs2q0uzMNUELtzeNcGpBihrKtcEzpwJwGg19gA0CuwirC
jXlx3Pzl3+JN0tgmrUNvYbzUhQBCQHwVZre7UNeTnBS2jjgkcQm6HrENolY4ewOc
TVzfBadQvEggvcvtRCH4dTIuEFMQWJKnBXfBCfOue9y5tQeO4zqPLk3cvFxKb6GK
L+qFtOFhRQZvu1x4D93nTpOFbxOIjxASXNQ9fpo52tEjJfX1ecbilZWQNvFxOmIf
WML5ffmYi3qXZHWOZi98TlKeyamxeY0xlG3qmUnVrHakhQmiZYJDjCZQYKmg7KYo
EjI75a1ZAbzurnX0WhmSjH4SKr5j9rlcOtu7OieTQPe3sxJ7mA13HwHralzoGR2V
zpXYseU+jrW9FCLBHxA3WqktsDlY+QoJzg+3j0aynBsPvOD0j/zMhWf8hktQpd/f
TlixJLvWL309dMWpV67jt/2LE60/xiD/stEBAIrO51GFvh/Yp+OL0WMksVwIfNsg
kVlRzPA70xAdld1HooqqsqnC7TbN05fx9BPYMzQIDyNxEaJ42vfVlbMJUF2BUaR5
klAccGP/pXv++Yp7pfffq9Llm3rcI3fArKNzBrQP7wjnV492xVnjqvljKv1tS1C6
z33IO5X98XpmivpDANF/OUo7n/hbs2wgxqOQSrmjp9YhCqOABSPu7yNU6k8PF7i/
c6swNrkYHDAK7je512AmO/3tkVQq6Us4qbqoDR74/8EaFD+npfbqAoln0+QpSIDA
r+0nFFeymzNxN4crVqJZqtLLVckWn1+gNpv7/aeFn3JoOje5Sx2QwlOHhrN47nS0
4O4vt4mcdvACMSrZUjcsIFLyzIvAXbHJQATwjho5TTaaBujCrh+bnvJtR/6meBnV
3nK0JAUlvc2JtFvoaQdRChzKHId9jXHib8Vz6wQ5LJm65+DxU/wguD7uGNNNILZF
YXU9b/xj5CGMT6KXQ218y5TkM/CB2SluVAaqtoXKAD5WtDu85bKxsEgbHYn4WBBM
21eAXGAQUtkoqVmk/74PKCBjED5qZu0dQRpykjf2shuD+7eB0/tFHEzc8yyS17pp
9o/LSJJMeI1pbeIvRZmWKnlIfCbbN3/F3KBOokTkdJUjPOHxbvseptVarc7rSkWd
vae+meRTXapDvi7t9oMqmiEIOm/Xm9YXm5grhT/akZv7RXnz/ePxt32bwuh4dBGR
lqi8YKwENuVywFqHtYejcTsezlyuMnx4jeaOErEaF8NtAmnEFWmwBSvHByBim1Om
cBXWuSngnDskEWBoECcAJyR9R830QXPYzJGpILr2fDU9B2aTCsqyU5v8ObsRhgQl
jnTbrrgWOUe2y6GbcI8cx7ZI3pKFVSvirIIzqdtTJBnH7/bY8bw8gyO1I8oDHQnY
2CPhWgwT5KM6pRkygiFwnT217U4Z/+yq6y6GfQao63ZBupjG+NDKcEbxIPFLZfM5
gGswPHmix4TPyLmnM+1ed4ogZ35vS9a144BsZznUWGYwyGOpzjY20gxIJo4El1n7
3qaxeT8QRC08Z454KXJFt4so8/HQuxXRjixYhabJmohB4vKiGrZHP+DD5leaqoaY
NjPDZri7CB+tqsqiQVhL2ZHypzHSeog/Hz1uPwDAbkU4IS1yO4CUXfvBcEjTpZYQ
XdzdVxIijkzcGhezT13JhMgHivtGXAsbE9gfbZF3ae0NFJavE9QFvtZoQmp5ubQq
PD/iPwY6UToHfZwGCKdWzZYXtU69HcNEwEL/kofda8GJfCIX3runphzI8z/c9T4I
sBFBE9S2aapM7fo7l5EYkZTOIAHwBtoALU1+Bq7Cb+QVZWucpoyvxZufYd2X6Vc9
jwmx85vYJPXzZajgD5g8TegA1dLvKVB0LGZgE2yFFkHT97N4Nioe3TDkGPlVFcCn
JUhWdF0JtJf7KSvcdqvSMTcxk6+lfVci+Pnx7J7HBvjRuVVroLFYgAw3w50fFUav
6fcqNpmU/uRsiIvLtsitE98fdDT7CU8SH6ohzZoiBmMzmrENlqASv2MQs7rYnqJH
mikTVmt9n5o1f1FmPIWq/ciYzfqYxkDzdIbAvMFwpz7OtYeWRfPt+cFaL2lCmmTA
tRk3PH8CgrzszYNXPZKhHFh4Xlbv2tdhscMPDzzRReMeIa1kPmN/xtT4+ikO+bpe
kO4s09pgP/jx7cm3dkakbCH/NMfxESAvAt1ifcvxcZ0uIV+CFt/4zngkiv0Fx7AS
teyZQzkuj3Lg82Aic3bWr7GFGF+/6RpHOwayJN3loOoqHugNN1iIo4x5IrzPeRk4
6+Dx6eUmoZU1MIiJN6TmzV5Xok8SjQGHw95lWiDEZcn+0khZ4P0lJ217W2BuSUuJ
kvOrtmHcOZgxDdcpPhGUAZeUGAU7Py+5uo2ESweb2ZprgPXMT3RuBDCGRYdsnWKK
AbxSXi4DtVwNLaPCwdW6uhuoAqPm7dlF6WtxiFIDgkWDMqN8967CCuBna45r0/+t
eAfLHVkMv99VcSPKVWrdzO2R6GPi8DoXunYiHJySUyPZ1YPLzGU1w6tTXnEYonik
q4Xd5ew5Qe3uU+3RIEID3oMEieetTOXcUdwHJ9mfRxgdKeX3JdB8vbz7UJOsFllk
BWebEugzLgC/Ed/+9BsGiwFVhpsLUc55H281PQh0qEad99KkuIX1imOQxGUAfGIn
yg2rCFVsOOIuLiQIdtVVQlcQfG/VLn6iWduuSoteTgFmXklaTBUTVIx7NbMn0uqt
H2oM0hwlJRZjPfJ+3Tm3bOwjA2fPsGiqXo+Xawfyxq7WdQZTwZDn4rHjmCgaoZQ5
h0gvO6gLRidQUY1a7lfmJ8rObS476/kuC0zjSDW67UckX6W/RSLpB2Nz5RwwkSVO
GNlrAKta1JES/KooBslh/haph7pWMFILDDV3/p970fIDh9RFwCJfNAsozIAY+5Na
Mv8WbSrMhvRIOSMMOsccXRPI3EVPSyGRn+P1YJaGEDQYGsidPvXoYdjfRzMLyPed
XfABqXmSdp8u4lAnPaaOnbRwaKrcpZcIHTxe8LbVS9/9zRacJ78UctNFqhByv4ID
3KTxjRxJIb6wupNNX2mVVqGcF0GvdgkMFkGn7BCITWLpr7qgGJfGHPg0lFl5N+08
qO2S/Xzx2Ya7mJkBv+trvZy3UnP7T3ZxqP6YR4Eb4B8FQ2izAWKqeN3Urazfx7G8
zJliK3VGlfLXOPcdhxMUnJ//GoX0Tdk7DmyCb0hk6wtL4jL2HpwhjMdSSR5FhdDB
U9/YZdTfc0P5x3r3CBkT7wHput2XB7jTyB+8l+JMmu3qd4LbON+3NViCjOcybJwx
N1nr+qUlfa4+/jpi50CqhifuJQYhbgD9+qc/82TQ77mJTvsZq4iL/HkMP8cMRbAf
ndaxSlYTP7c+2iV7HleRb0PIT5/IEBRelua0JEIDsw4/hQ+V6ThBt8RmBVaX4ZDC
5Zomj5vBqwRIyBwaYMmma1CQKbXu8qM65vScjSwi3Di4nFu4FhpTMeAIi1fx7TR3
9Iz2r1OiIvqiU7uOQTSd9OKzipWOOFn5+54vQnzgYjoz8ylEgZsWTxBA2somwhdr
0ccSH4Ni47DOwVkvkK9ULr3ciqCLolXy3yM5Zpk06QG7gmqIaXjW5rs5beU3qv25
oY4FMRQERIaKQm0kZYIFjp+RkdC1qVJLdxC7MMMQThUk2171eDP5j07Uzi9jnZBj
mZV0mgCI5/nx1bq+SS4RKSTLRw4oEym4h1Fw2cUNnOpqsqcVlWiw0e0GRx37tTLo
pUTht7b1QiUqklwu5lyMZkxSCQKPtyrnycLIZ1jxzFF3Jx44vu/HTZmRsMhK1M+c
dmnJAViwtCP8pNJkBj+aWOsc41XqI9DAV4iZ6xkyoMaCBemwo2pCLqlWLrtTcnzF
icRc8/lfAtRuDHwpx6gRjfhQvTe2cajUiY1evGIXBcLATBUacSHWXI00k0Eb1M9j
M84pAqkbB4N1McnlCYhIwkMcWbe8EN5n+cpaBU+nzSBhtUsH5Lql5VdQe1PM3UUs
r6iAJakRElGGFa5gay4X7fg8ROpEAx4Y7KMqRuV5QM1vwhhfqOu2KmEnDc022LVE
93IFsjeK1BphIwgAO7xR9z6FknoT4oO85DPnyjg9Yr+6Yyl561cYEBMagvAcvTBc
T7lIHC3/7Giu6axFwlcuUHAAj6PNj3fRjYMQlhCAhkoi1z98uOkSwNmXb42z5hUQ
W1Ovqfx/cwn6QTDNIkWXXRLl58HVrBoEm6soDJaQZBp9ajckBVDITG7QNa2v+Qs3
HdBLMTYE1hYfQ/Y9+/mTPAd3xBjZMRvfhPGq3YPqrFLWOLHa6MIkM8hk2NHczP4M
UORyMeCZ5cmhXb8351spJ7U64uuPfaYH3A4DhLbSUDm2g6pn+WUh2VK1EI9YYNqW
l0iz1tk6d5ytuN0vFxh28jas2QQjs7C+UoIChTA348Jopo3OIsGzUVrCMeWpccfY
xMkgbL69Sf2U7xO+i9aUo8KEDMZkq55UTrza3Lg66W+58WqhhG9kyXgRZG6bT8BB
wIpflcP5verp4h/g6unJ88mbGStfx6xaoJwmFzi1yPEUHFY2hDnE7wthYMARGf2h
JNKeojlqBYAzVN7w+Oqm7F+7kI58ZjAOrMVTzOJRgHv77ilc8Ens0Oagi6nzhBPe
/uiXzHfv0/aORWr8SO1JV4Uit4jWTYnNB80JgIjHRq2uU5MgPvWOG0vN6jYNW1l3
V/fJn0dTg9yVdridvGYaiP0aoswdjveoBWNPZ641X/gZtL1FDkHzA2mKhfGib0eT
fdC31T3+f61Mk3lXxJ0F1zXjqMXZ0ba0q+2uRharppKtDeEy24B3Vvo7kK7DIEY0
8Y3ztLhhbVyEQaP0nQ8s/OV45nErBsKjI0dwaLyzRXs+M0aoA8G+CXnMM/TBVIrU
CWqYepafWXcDS/H9iPgMuOSxkP3wzFIUGrm2qL/TsgUKR7qwp0ojhvJtwq1l+B0m
bgD7NOnWW6hOyDzuyTae4LRJPxtS0JoD0O7L4YibEwfrzLDmG33GMsstJGs04BFd
rzZKNN+U4fHn4syXl/PVom3hIJ0KQr2tO3toNj/I12DRPsuiWQIZwCPr14fP8YQD
mbIsS9TID3lkHOX+MwWLRV6EhAHbKfMtXXG8AshSMUIiwMXDyK4wdl/FjMkzyBf3
VuUrXl0AXMXjqwhKv1Tvz3EI8pm6yIYxc/rzDPKaQ5zqa8UWSHiWUvEMy0ssRNw4
yzlC9eHnzkJuUHloKDktbJXeRDA8IQeKkO9Tx4V2rWdAIJbma9Gao0+5zfOVrZTE
J7TCfbxs6v9bCmn0fxcnK/dyynEBu0lOq9Bv4bih3o6Zc/PSzN7Gxapk1Xq9lEfU
UD7S1N6mwvfnYVqMD6o7oyUghBHjQ817yfT2thlFF8r2ZAUmUQW0iIkrTeFlZ6GE
df6z8LWZRn/OuBeRE2BoGVeMsaNPJKDW9QH9z6C/GAyRlPyiSmglaFXRO+p3wqx0
egswqgMLRmD8vM2DAQmv0CT7Z7oiJwqJ6nG2bXBjv77WqAwQf9Xoz3eQ18ouUmq0
K5PKFAW1OpU2YoZS1cVgavLuuCkH0xUaPStaPB4XMovR0ns3RTSkhmkIMwmfKenj
GJFNVPsHC1zybIHGhtEFR+kcYznzu27QXZ+CCAZvFhfy3vH397uAsoo3lz+TABqd
faNomrb7VBtHAz+/fmyxYG58QRmz24AiLR9mFDseucbb1fM0pEyTKtLPO2efPg5+
6uggHg9M8QmH9IdK13GzKgdIvGJMWiHbO+rUAVQKRsJckJvDoV0gbCojIEcPNiTv
cZHn1dUqb617KQpHH3fi5IgC85jAIInd3T7Ykjn3b+z2vpi//4v+Dijd4jKYpKj1
5DAo/5c+M7tv+58eKhuKPOlIdENZ7pVuGlv3HBMnteghy0YQ/ez+7XdcTYX71R+c
snQtNjHrJcvdyWN7rVasP+376n/8TMzZj7R6wHICHWQgD7UEL9fw8V/1s72YpwFF
DqhbBDxkuxbX5JRqPDqs1yDg6eNWbpSlXOUfedpDtMC2Zdu1waacQ4qXNA/mcvGS
PGXmQkelPKxT36dahD7NQV5uBJiuO+VVkL7GP/DlLE3YbKRVFCKOqLNj922cB8q9
ratx7eQpR2c7+qX/CSY27gA3zw3yWOygO9+lSN7wqV7it6su4RY8JOZqh2TMjv82
dhvWhApqyyslI7vJyn0HLzD/UvUptRp7cf5ae6L0F82ZXVVwSv4uZUhWSa3OiQ7j
AxDYjnPVYtG2ohWe26C5UqOJl2Up7rMFOYKScxQLm26sCrAhtmVEeZ+NTWN3YRqE
gQjleYGiDcu0jXnp0kz1lMcmpQoPedJZVFLwX2eE+4ONVVSHdm4iHVVZwWrz0Gsa
Kr1rlwimxiHrwC2P8QVa22Quiotds0leVNtIcjD798AejeE/jSSLnzbSyJqPP0ls
jpIUHrUzDNCklOpSv16NDikJwI5JsBtyjkvTri6y4AAwDGmE+4rCEZdR8FC29/ZO
xGrVz9KO8/H3VM/JHQe9NixxCd6nXpOwCH/rnQAUMs6ZYMALH6j6swKyY3i5kd9m
0vXjH2HZcIMVg/gvEzj6+qR2MBbl9ptevq2flg0++wmYtQ0mzUbgvjwA8/qpeyqn
UkLL0EYK6Uw1W+9IuRRo5AjQ2gAqqTskX8pQeBdZyPncCHtKwU8LID/hXB8OP3Ku
7k34XPUswUF6D9x2EVjIJFpiB/B2Mu4iuNOXGStfa+NYE6ZutB+c+5kSRFziRYZL
uhv+RntuPXewVF9owNAqCSVbBsf65Z8YDIyMSxha4BP6nW34BGx6V8QJJVjT3q6l
rJMa2cpnZ0ldX97wE0VUtO26YT4qBcugYla9tFt7c4DXJ4ezd+KjT+1tWEmSBN09
GM4HP6Wr87n6P/QFIKnBwbOWYwqCE01ce17WwIekMMg4GwPejWw5wK7Wo5SUH4OV
01t+pjKyrrG36AoXZzL+DCUj5MfZ950PHVZVYGsQibhZC/9oYfeOhRv9LMF6vzxL
H5XYrTrU14rFu4ZomaOxvdD6pEIHtV41E57igOdd+6m6dXySx9YiNl2L27DULefQ
bTXsxGeK748q04PSMKmCt4eycvhesFaVoAauOHyAb2yeR86tzZSPO/T4I3npouE/
xg0aQCxLvc0aAPgCoxwMctZnkR6TuhqSBOVmrS2z7TvY0VswLNnTmQFy7nsKr1P6
QsLtBNcI9QKGZEg5TVw4PcLeHnWFkTtNBCnQOyLvl07BUd4KFa0dAwGkIVpo6EjE
DgkHKUC3EqDwi4IlHThbXM1x925xz151RpORCO459MQnd7jheC0meB3GRwnBWl+T
AE6RcLHhGuY9jSHAuWK1wurXW197ttzY/Vp2nvqsWGI2JFSEirDf+CUuUl2X1tUa
y1kUpj1NjL8i5yNQzReqqMBQz4K5q6qH2Sw3rdQNk+CYjbj6GMGOddCPeL0SJWuk
0mVYtDO5o1RFCmBO+s4gHXRyFhlWgEm0OWvSZZF/F6d6WJEM2IpN/iqF9qLaHs7G
ir6PGlil6z0HOmfmBbHvW/qg/ENczFGzbwBUYWfsM2MRBOk5rwizrwTNLYvekKR6
LefUtCvMgl624r7FpfngC3Vq0DhKXT5xF7cOdkcoppQiRtigDYVUoGISYeMhdqh7
VKxWLss4EtyqwCRGWFSiqweCF9vI31luZEulWSFo30W9OFQ+WT5FEYMuJsGwXW73
kGcaFSkDCLpnGWdHzRkX3L0xA28wbKZ7OlWhsWcd6YSmje1FUnF7mx9/yNoC8yu3
acBSNgA5wFxz3Gig6YxXARCb8WbDQGr8s1QgX+T1k7GadToP+hdmfxbcBgaiZHA8
a4/oyLmNqdqE2Us64kCBvcsJCtVMtYpmo2PKNUhfd+Epmx4Yc11kkDE7CdjoyfC9
wnzt1QpSA8qKIIJUDx/0nl53gvHaqYlpAR/y8uWp2SA7JiH94+I0FZ4TykEVskyG
kARLzHrHaoCgYpEvg/9ZB1r0C+C0TyQJvAkP2/vY7Mp7TmHWrr0E3iOp1zQNbQoc
fMfDgVCEVE90BZoQxKw7HjdgBwNK71BKVXxpY/o6MumTb2SD17LCSlMrQkbmQ+yz
oPa2fONc5gTXwOcxsuuPHsdO0/n64iH6SkTr+m+IwpWSE6hXkvtlcCL0+a067OYQ
3GF6WQZcq10Uf5RBB6Ze6PnkHPyJpwyA24Doa+x5ROYc5yrPAzSf0Xvxicc/YibL
CfuuT0xyB69McCGpCp97d4c+1b+VkHYMU8xthPxE68H55J9QHoouKVhDbQ0TZA0e
/sLJItaaHMnoGuEbqr83V92RD7buUUJAtgwY/7M05v1N7Jmg2efqcOF7VOMuBNQ8
eVMx92A/v+YBlhNAgmN36fEw1TEiOpZJE+eJ2wSXeyh/nJWiqX8Q4vnad/TyJI0r
Ld5Ahzrp4FfdkRFhW/o0f6gWn8K9aYe00Mn1+ep77BUlOzl1nXPMYaKlhuF3Xgyg
X8aXN+ID+FRBJce2jqMBa9U87y7LycWPETjteB8t2M/j0gw9nKMGfOe7UefXvyYr
li5AzAzoJ4t8kJD84lojNXav+qMAX6JY6CjdhYy7OGgft89VE4sVfNQ6k9c8pl8M
/ouq83ZGo7wy9duNa9lKBeGM8iCFRcwB/vWoEmI8eQnm/8OrmyO3U4kVK091U/pL
7Ws61XaO+KhV4vzlLLWckiSLdnwML+hNjlruKXzpTDQhwra8h2Ml/omK7NoixcU5
9bvkAhX+Hm5pj/QwpskhQSNUVcV9ubdmihgXCKc8e0qBY3bhUXkhPkAyWy+b+WPM
VfDApzbkXIOccXcBrr0a0LVtCBwtkGbPNNMHCaNDUhNNorCELDGjn/566K/z0nAY
OR79vLV3jOhwnIXAcC7XeHYLPVilBpcAWCca2dwxlWF5Fty/v2tkKa30r2pjdvEm
9E+jn6XNLms6SkpQmSzlkmWZialtGpJWefq6GlivaR1vzRcw2U1A6/nmR8McLjjc
thfsFRJPLd4x/o2TKVTRZMd1pU6GLOYZmX1wEJF6AzU5dPnR3NbnqTxcvHLN5QfL
a11aHRlDOaOY3EBV4JmFP79U9uTwbkRL277s533N+t8rBFW7RENdwt83zpeCKelw
vgkhs04DEFrajdVqQczNF+qMdFcbvsY/x6VhmKOfyUg8Y5+U9b2mjU5WlYpseMdA
I0dMAk8vnyNP2mePq9PE/Fmv3zfMISAFA9XO4N8npSkA0iJpRdczogqmCCuvljcR
P1vkdTP+RQ4E3Zaq6kTPE2pvKuup6HYSIZDUx3RFToPrHrXSXGxS/6x7CDNkUrlb
5bG0cm/E8eCLIE7kpYHSzOOt40WwtQfucGBeUDX1BvWwJ4/NS6TcVW8sicRIaO3K
+IYEhDUKxyMlUfXnY+ort/K5lQ7d0x/nGA+1zX97Ije8cEFWv/Fboxg3drqusUwh
NSv0pCSbsnFOtT1EK5NsRUjUDGzTAk4TcHLRqUyPeIQRSref/IPR/NeW8h+AWCbW
eyX5Qiv3yPbEKE1JpMUij9q3dpnG/dukhytR8drI6yaadl13zJPMf0j2mGncGADh
5iH0YjxZDyNmSK37LmNjoIVWE8hX0UY3IsvinWGeHhxjxoayU6ZuK59jmqI1GeSs
AlTzjotreJS/sERmxh4gaJgebk/OIpk1KfVNweq74PfFo7XqBkBfrum5BJx0usiY
UmNNriMqXs1i2rgwF/801yBFJyJZc7z++fu9oHxubftKahH5lvj/Q+ej2xYZ/Gje
8dnK24mN3GfUA5Ar9TlOWQwcoVa5QRgDORx61wfT/lrhCCVzhVC+/aUNVgg/U7BG
cvecRJsOa7Pmd3adSalzpeBPBIqu0DqpB3gHlWwci8nQJfxUnTg5ExnWhFMaMzJq
i9UIqH+GzRAojTSpRHIF/RLEGzeWRqUbAzKERcIP/T/YW5gbh50NJ6yToa+GtQn9
/ut3E11wx8T8TwH7LisnZLvUq0sWkSoIBxa8bINfNR4lkZAxU3GHmmANEcAsR2I1
GdY7s/LcBL2YScdC5HHWbLhhYfgRnPRPs55V2HuUz2iW13gYoDZe+I1BjJ9h2Kyw
vRZywLlQlxubLdZwIbM9WQcAD8E6kxY+Hv/uc/nvaPA0eF7hxLs3kw+0DbSzLdUG
Xdy5P7Gc69xVMspjlIPuhPU22Tvw4eUBkTPpChDG9uSUHidfc7FMgYkKXsTMHVjb
3QU4blUsnRuKs/VNb7n5Ri9BtjyDM3WzGOlR2522A7aWO91kEhoitVWpSyDnxnp5
56DEkaX6dxtjiO0rcYSpUJ0h+jz0LHckrHdeZqOVQDQT6K1D58cVIn8fsPSBPpQG
xyJyMAB4CHUveoXqtewqU2/EJmNpLvotJErFKfTz+2/FA/bDn3LOT4HHPCENNYg3
rdnBLFB+1zKdT1F/taf+YJ5hmT7n5fjRpH75nvhAOCC5Y/Lp7HLW6NfUgslks6xC
c1zn2onA+6MM+vsee20rgoZYIYkS7V1H62C/wDFB4N85h+LYMRW8nQqgB7Lq01Q3
dB+MrRpAQlT9RVyBzsxUVeJ8V/nJof1sqp9ZtdAZP7N6V/9pu6MLtRaZzcpDeWu6
AJ4eE7m2MziJxBiB6guWoKO70wk7T1bKhqCxS+DwOUkdlg8XW2s2cGbS50utKkqc
7d3ZbPwW+EAqdaqMScNaSx1m7/QFxHXPS4375vjPdRqAR//KumDFQjrcJso4ol3A
Tuiw885whVMP3XJWpZp2wcm6nuhbqGM+f5UJ/U0DAlqc8kNqrDbYl5IH1e6C+2U3
azbzuhKXFQB/3L10wWIRLuh1dUVMiHX5lt2ntvlYxAAYrgU5jWVSYoB4JPc8b/dC
r1vLZgZvEPwD2keyf3lh8QFFUKL8WV+1VsZeg1aE1loUPE0fgoGhMh6M0gFKjhva
IZrRYVIPel4QQ+T91oadb8qEZy5lvk7zB4XhfCbZkcD1uk45SfSlAC8NAZMoMOV0
jlmbJQNDiLZyjyyWovoLRs6Igb4EGKmuxpUyyv3F+joEp7/GFNj37p8oT282og9Q
6BIA+YrWULtaqae1yH4gt7bA0Ridxmip+2MWay359jAU2oHHdp6aZAOpOWUsFSl+
QFg+CYY4nhd8kB09utleJdSUlLcX/2fJnovWrk+8hFnkI/nswKvcoDbKvzUWQNhx
rXe72qBlD3PeD5etLyrALYC9uMtbsKrcLf00Voyvp7LzlI+rkzsgyqv6dAv8p6pe
XR0wJ9NtV1qHcBwutkbuIbXxTOiMjvU+nBz8o+enXRmiGcewT3/Y0r5wQaLR+n+z
ilPKRXfe8n9MszKpsM+w1yHR7wcDP0sDeHfz8Xi2vVi7ukyDllkAGuvanB47L4ah
Qr5W0I/xoQz/uiA5j7tfCUtRDIdGAWUTEQH3mUJ+0NtfZYNGBfKrYLw7//016s5r
1eM4Gb7RTdvnJ09VoI0YZ5kYoUPbu7V4OOxtvhXGLGOG9gqeXwSI4+iuKJ1CjZ3c
HtjMUay35TiWaajnQpi++Ttjt9+mDeLgUCFFSJxPwG7JLDXuIWCi9izLh6UZCPPd
NqPn4SG4QQIrbVeV61n/TUH9Dtiw5l/U3y5tLxlUZBI0eyDBC7ZRLHEhH8Y2/1lN
H0R3to9rTy2UWDseUVrjTzi+pnFQzJsjqPQyoXHqU+Il9Te6t8F0pF3eRRmc+r/Q
hpDIltvxjKA9HbXzA3on7oTvufZeaxSVk4yZMe6RChjnL62z1N+rKDemu6qcezhm
jBxKsOD9+c/encW2OoRcknE9SOGrZAplkGSIUgrH9r7HhBckVzt84ETuIOLBulaI
NGrnh68vd35qklI3OtGVTs2qc3g0uT07o1xEiZlTbt1ipCEB/RiMavRa6Jhpsr0N
pbGlqwv/FcWeSUv9EI8ZfPfPJ7WGW8CTjBTqGJjeN3w13p/dAtIn6+nG9R7EnzxJ
sJAHe37fyiFFA1Xho3Pz3E9YzTByBAzUHJRUnc4XoPhvk9k3ZNfJYZ0scxf+ZmPF
mPJS9uCpPDQ/JvDHYmqfcBUiJJKQz7KaXS3XkIV0GwKBQzmsOWdSWI4WlYbZAQQm
l4A12hjRhuWXUBMFAmBL6WPk/KzLC7NTEWn4Y8rc63f8I5vtU7hnpvEY7Pf4Wgzm
ZE6UVM6cjV2DBIC4veoATnpTXJ5UrQVkoxDMRpr3PqJ4TsjDSsTHjHE+3XQFKrGF
/kYYb3CDxN4Ep7jB1QMv1G/56v1pP4KBWUWjxEr2sro2vSc+6soQogeDyqvoMuiV
kzV+4hEO/Uxvw/k7g76ZcTliVCJqVf32QjKr7O1kPdCJ8LObR1t006Ei0HSApWBe
PZgdpGBbLJNJjUw/fKEr33RIBPqBKpbSnhvlFfDMOXHGUpPVS+6obiQuGgrlrDHe
mFr/iyXATgPg1NkCUcDWjb3JxKZxg0HhunVc+/Q6DDkFnO/2NNh4HbLGn+3Yt1Sk
SUKxt5DpT5pswOac9OSrLlyniptn2wYlrGRjVSDFCEndBCF2HzJxncPzk84pE7p/
oyRq9THm/JPtWKmBzJJAvrQXefZe3yUvHYl2dSZXZaG5pOrAoVOc4rGGuw3VQ1+z
pKE537bMLdOe/rxmUcp8nGNv8vMB8U80SDfAo89/ddMERjxptD8lLJpFj4gakDXC
ryu8nBelqS31C2RSBXEuLNGDdne/HjDRWOz0m7wchSjR1XP6LCw4Rzn8kmVzC0tl
Q+2cTJdTBfrJ/ZORTBZairEw4cQb4AhcOMm/qljsbufODoHwYI/QSBpwKpOgTEe0
9o20ZnmXYoFDwrVFYjXom3L8Q6OgyEyTvkZh5eKJ0xe4W35HFulrvsVqTcGrH6s+
Uf8i6FTgoBIQZfyS/s/HJHb9AUua79ydl9y/W+nk8hsxjaV25m1Ezmhx6K0u1ihz
8azQVwshl0gaOnDQCzJY+sPqw/gRDnaiZyaolyNhmKSXzLVQKmKn9Ueez+bdGLs9
ZUC1vyHYDneKCT7N8rtf/QxySIrPrB2SmiVpC2/1ArMQ9f7p0mRgBkJShhB3Ftln
PhCgb9SJSvz70PuPIoZhECzgn611vAwFZ6n4OQkyBd89HhVzIURefJyfpNlWdcOY
e4TO2qhl4xo64rjamv4J3s7P330EvpL4r6VH1Hg/z3DU5zvSwJ1dhUhZgCxk4jzw
kpmZQ9V2v1wzPnlusKeXTrWQbAq7kK/GyPJdWW4USAj41o536n2odofu6X8PzCxk
EcRDv3rMzab/VpUkw1BKtee/1+calDYp1XPnPiOvWYLoFTUPf7t5DNhbC7VNn2Dy
AaeVAhH35BWHLPblJ9gLWjCqL0EcbNywtCOumx24VBjAXprhUvx3hJSOWo15hUm2
mUaHWFOnUPo0Wf0+hO0IBlBSRMIP602932W5i3cOHXry8CcJaLJCNNF8cfF5ANaT
ePqzHM5hTLNu546fhr+sXchx/VhbU6a0npwFLctxYPeZvbyX4q1G4oCxuQ1dVMCL
1WX1XcCxrwAhz7iw++I2L8aQ32e7j01SV+/D0Opv+rqBuJypjanksCb9NBBNSWzz
63WlQAmyhuamLa6UshQPsXZYDfRnRSoQ3uD1cXF/ZScJQ+9uvL3s+berZjYB6muG
6IcEC748Q6DZ/iamPaGpodWTpEoIW1O1AkutpkI3u9RBqOmtSkV39LceI1X9K8Ir
phmugUnQzyO7MU0CQ/ROGLe47CruZbxNYj/p3PMS0WbrZDon8julppVUJNDdJy9P
kIQVUV4MHhtSQycGM/v+/AhZ53nLc1OpKHL+UCS53Aqaezbi2h52aYBGnqoCje76
Y8kPRtX6KHj6f+mKW8w/V2UZDMkYBMCJ7+vLJEjSnv4f4V9hvegjacbz4x/j8Dp9
/dSAal9dikm6HQMrOreY+R28354sgM1UL3dwDQXmf/ssQN38+RpVuTHevIN9aDWc
MepW+S6eYPgtHWHFdKr0ntG+3/lfUeEZj2d3+03x4c17NwkvZfLGDKyF+Sg+O6OM
O7SaFuyOQO5pLsU//bFf5lSkr5+7XGENqSIy0UNatICW3xl0iJFfsStSL38U2JA2
HYjDv8ftNRVBwRayFeGH9g4Utwdbtv0bMKO/ry2w0VCxdKd1omjO++GkuW5T+g2f
hfYak4FB6R8PPC5PpJ88IuLxUjGPFqM18gxaE6PXKLCpFz7oUXDBOY379tPkGsTd
zha+9cIMArstDUPoB0tGgShZ+RvYi70K/fsNMqqZylynRwLiTkzUSwu5qh3QzJdx
WSRuEZjTtKrlIct5kYvVmJgKNRRvNDa+NIdGiBzJF8KlX9qp1zyBIh5LWJZ8HacW
iQEPo3y5EDxqThZXUcOaofGlrBd0nxf05tqD8hzXZDPKjBxT5Q7VIvuYnI11u4g0
3f81a7prUy5wNgp2Ykk55hAw61Bp1r5o0KQMhS4rweCMXePQLDHGeHLDuIr3yOLZ
v8s7hFaBoun/bo5AfAwbskIhA+LiWLf9zBm8SbyInK0TPaeAVqETL0PBgQW5EHMc
ZHGmYN7Xv3aWA5adijCVTIbUKa9tWZD+eE2mZskSwKrSpPHXlU4tsiKQaYMifo3O
TS6WSQRkDRCITJlvBvd1A8iq+bHTRsmjIo6jBChWtl2LJH96se28mphuevvOMo45
r0uo6IEE196KIEZRhh+rppeOPfoVgCoHUjn+QRGNW6/xuYbAiYjBuA9CxiR8PFcm
uo+KOB1qyRhWwh/f8D2G5XviuyuUXLn0T51W0z/2ukPyefKcrDd7i99R9ZAdMzO5
tereCt3cmVgukCibVVBRa0n0HetyWRhIUDRXdaeVKljcbHtWtNbSVJa11WW2wLwW
VWmO3yGxZ4lwNiFkCezRbwJyWhpV+L0Qo4ht51bz2dymGDpSFkSFg7IebFe3SWHl
oMqtITS4uUnMqAa7kaWpbMIqmsRuc4zZUsaPSEei2OLaonLM1iWjcNHJV4BN4L/K
1yh3lbGcIRmJv1C1t4xfpqpvu99xaUOdQppRaZR1vgeiJJt517mmdAi3A9nZ7ih8
qw7w8AJg3bWPJMeoeexksqs/lL4706s0LmQ3dDPoLwLlyEGJXdGaVltnoal5OsrT
H1ntydiV8gYziNP7qwUYfnV14k3cCHw+5AtWT6ha+2NWB4DHPZRizG2XMOoTee5X
6lPg0fHaZExDtkwRmRs3ylZPgkn4Dm6bD1COgvA4uj64o1AfPY4iCKHV90CdhJ7I
/9C+BLiSa96HrK1PlsJ2Y3wXuc3JqMzD7UdNfuNW6DD6WYalzxQOyoO5GpfR591r
BzAy8RRsraOCIpU0I5UybLA+DEenhiGQmOw4Od41vgc5WQWhM3eJjUUlkqQVNUpS
4BKQfiH1cZoXrn3FGl79azD8bvCfm6T5rS5bEzkvaMR1yXeWlVbW9nXfTaLeHfNp
Yk+9TnxxLCuUe3to4LF6k1SsSY0SxpEwQkAr5+GmMvjPRSqDbdgTut1+eYbcWeKC
TT8/Tlvo9dbJo8u3xxEbyeOT6129a3mRjeOYEzFT0bE6CTKP5YxZDmMIcWraBHSq
t3zXtGZYfnnThpZvSv5+McJw++pmTH0m31KPxMcgODqXUuwKgW1hJTMxadopjC4G
UEJO298zCtLV/tPwmOmQbd6Yh+kiMYL5uARll41+Vj6uYB73gXDd5l3hf09bMfSJ
NT+g6NCKUXqftTfIu3yyxRNMKeg79W5Jo+xOgXQYCCp04CisvwQQDi6/FkWjKZyz
pzlov2OSsusDIoOKPxgbWgP8DN35jPL/9QFYHzsOKLAVLlAHe8Bln4j2INj949nz
rKHIscYlNVCJTfdycCPkZ6rDF6fiVwex7Rxjkf6URHcBax1wyywoDWbHMgB/1GS3
qYXIPy6T86i33muUYmQg96wz9EElveLSJHa7njO5etifFxrYHijpaScyq8y7MmOl
2HJ6nWrexUv5OiWtxAs68DnJe/NJxjV4zs2JfZk/pIpgDCOh1o81cAW5ea1e2IYE
6yTJJTobo2kC6LOHIHvtr1FrkKVV6cT9DSftmLXbd3Rxnk06XXn73Q4U6B2pWgAx
eJrCdClfgXYXgQzudaS1TYIQLUgziL0iiyhj3OgyMsNyGAw3030Q3ucu0kemvUl6
dprIkhRFV5dAIpjFKRcHP/ICMPrqgudrcsT8ed2KNFw4XMv4kJV4BRpXFoVee/+O
oXOPnjXCubBCtBUYhq2qPlYXso+5z+0txDn/QPp5syIlAaJ1izljG41pxqW6F0Aj
2vqJ2MNEGxcNo9EFueEcWngQ4RFlR1sscbmf+HWKI9vvIaUGIY4/9UBVCcCO+kMR
UpNKky2RCeeFx2I9XgxJGA6LX1tRcxsI0PwLCZ+XucnanXRzRcRbX334P5bOBuMu
swQ/8mcG8FoJdwFGonTvAJeI1B6byph93krAjBaFVNeILep4akS/EkXN4xuZh5Mw
Beso3JTDkzv9t7rSCZwC++xzrae7pMaLCIpqh2EPhY8iKujc4gE2RVT2k4ROZz5B
g5h4eKYqRIwHOjzcy5WNYbOIqUMphQjSz6T13Ojo0B+MjuQF1xpw+JlKJzay8NyH
ZF/zfPJ+6wo4YjQaTVZtynMZiz3j2aurGErG/g0af2l9OBR/a8GnV+qKPcDbcmPR
SUeCbvO21dTDncOfWgaODCqenTbNF/laMI0bO/zh00205FsGDhm3Re/YHtB+LWBJ
mmXB+lmS4bd/oEWZOzBkK4B6GGUydZrc5zZ5AN2W9KUzZqFmTvtpugYP6+9EchKB
JA4DMSu/IawyTSvrMHndfn1kMiiJlt/kxAlFTPplzu2OvQD38NomsSbMewIv5crz
9Zfbp6M91GqMKiy0GF3fKCVBX2Pca0NZvy3m3z6nIZVSqUqKY6jVutLteJaV+UUb
TKkWGXQrbY3beA3MUafC/DNZGReuCuiGphPQTH9xq+XhoroMCKfrFjPZnieSSKzh
9PuAPgbBqp1q70RfKUUJdL/13iqE+mywgkgJBzQmCXrYymV1hXHqfHn715yMZ5Lz
dIWrRO5hSmMB3cExnztd1ozhA363MWU/xrfuY8othjrWMos8lVaY5WQ3ikERz0+L
8ca11UGaZacgC4zl88AWlxeq3Z7OU8IOlcjtdnW5DzLLciWUH0nznLcWIWRz3fid
y1Vi9g5/7J4vOhiIGGGQRQFDkvpueQy1M4xnzlSIyX/nvFB7IujSdNuO1ANAg6AT
Vir1UdfNWP9CwjOEYW5ibhrS7NVZMkAsFrGtaZ2R64uLx2DW0wDEpNUibKNRnFp3
epBA1u9EEI1n2kG72ilfsEyI5tprq2mp8Xim5QjEq9XnqL2z91EDw0+brlFLIV+L
7FIjq73r6g8MICfAxSt+IG7YlfjblYTOn/PaJbRRyfcAmB/839lJ/2dqYlPgJJVw
blp8HhMbhxHz1JJoeUOHoXxUcHJzawifwpmAS4WAM+GJNTdDrIYT0tntaJv4xUHv
Omb4rWJfR3reWsPwTmvmpUrGc7N7DWTxgGhmoW1Rf5Rv84+EyRZd+H4kYIThCI52
G8NIoJfHlQXXnk0sFSsKie/fbHG73Wf9JNA67LadIfQdlnNWXWAMvkccBpPj8Tp4
mpdgRjlm2aeesvQcfg5EtgXi9/QwgTPhuqz1WrzHXKbWwg8xJfHlgGqugnh2WRy/
LB36KTCS4xyIC5xNoYcINfJA70Vp2dBZsT/sSSuZ2RkyxUazT9+R6O/bUQ9iV5L/
yItnkqUcNV2GAjFYo4Bdw6cQ5EQnHXa6vb4ajkOEpd3EI2migXZJDmIE9GwsUURg
fXxDIxefzbFUpJ8rbHQE6+cg4BAKqBrXCdR1aPGgRbBcBLXA0iQ/ZQBV0wqJr1j5
pQu7LVUdJDWhL9LL3nr9/WH2zl8G2LFAAKLDD9nQeGZXQWhYNpDRBz+edQ7f2Mr/
kn3j1WM8wztyrybwZlFfVn8MXlUCI9scjdX/rf119n60NXADUx0NvJ3E+QUbJkdO
T6E93Zu9cVukxpzCCRSRE1GPd/0kr/WL70hmJgZ//r3hMsZXGAJOFob3RY6hCAZX
eA46ByAltONRav6gBLhOeXazz5F1njVD/EhczqPlOGabkNB6cHPKZ8OfKZUQRshm
gPLNKJR2qN8lGPEUh7VH682tgmTwhWNb3a3bpdo1jgnjUuaeEQux0PwHkVw0BbzW
dSnbaJbPHX5IphKVUMytmpHn+DI7O/HgH+p3p3aUTeYL1Nhl/S5Qhe4Qki2IWuzX
AW/GzyPmrfuGKalJX8E6b6IQiF7hL9iS+UVHCmRdvaIa2FvURoInQb69Rz76hba6
HW+Pnim7Cy6AAtc+St7RtGD4l5NgVLt8SZkMDNJiuppxKuZggd1aX5W/OhLxrimu
CzCS/Ycugg7SYJ4KKXU1FecCxg3EgV6mqbY4EiE+KQ9jxDwsDnu9cfg/M8S8cvM3
NSn9k/VS9QMzys0axm1CXj54avWxS1Fdix3Ax5ZVlQggadx62cz1gJyQ9bYspYGz
19YvnP4Ct2BvfxSPx7etrNPu4TUz6W3TlVxH5QZWA9BmuvqmRv+IkUnMie/UNb28
oJVFvbqiVT2QCdQfI/X7Ef1SMwvGISXFB3G1CPSegXKxzr0jNhuUyjAGIZyUkGE1
/FgtYosSEfiGA8UL6a1w1/2cYl23DlHGPq/M9PX7ajhoXmec2PAF9O25Pqz5x3nJ
k905jKLY2xZpvNeNAplllh5Us26qdTLlbTDs7t0+d1CcrVqtc/9sDrSCrfKwK+n2
uTQU8O5LVT3EPT2Iu/J+NQ+cFnzU1KbmneK23wNRQcgOYm6FL1Le0yCkc3NqwJwo
QYlxIZsBqo7RyWlNdL7pvupzR6A7rfhMhyXG/mVaT15uozUEhvpptjvfGIDmrrm1
NoKw3VJA0xXKDjPm/EYdhdsShtfJWwBmIRLzFBiYTwJRepfiHQOBwn808YpvZ42a
j0cboyZIZVKqf2uD9bz9m7fiYUOrheUyS3fq59peZzK5Zwj+SjQGw72UAKlhaevV
wVwZVhszDEeIQQL/Gk0mhW+l1sUD3otlupim10oEzwu4glkAY0J62roctmnBGmdE
uiXJL24OrEb1wrfHVsVVKJtG3EBd/Y/nHZ9w8DhEKAp4YlGfdypAAWuc0iwqI9Hg
G7k3pWgjzrxx7KmuMWwO+DC0UCn+Jnb79Y8rVFhusuG5RJA5FTZ5Um3JQTAZHyF7
42URizwqMJ8oo6+Dpz3e6GC+1GTg7har2QFPd+09tqb9TY2g6zGuB1O0mAsDgk0j
dn1mE81AsFp2C1NgmQAkPQiwkm5lwT2/i1z6NH5IuMOmRoi5Pm1SRL84pLVmbTeg
9n0UMFLJTfB9trPEoxxrWnlAX0EfRX3yr2g5w7g1S5JOb5OjVgFaBYsxcSlb8NlU
UyxwF6avylrpzYK93J6F+y6mmy3LdZjgrGjFxOOrRM3jF9u5nptdBSh/s8hU68pg
vK1aqU0dSYc+K1mN/uGcludYsrnnuNF32fWKstzHgGKuzbUxasWaMiublV3DBwEh
i+EN39a3AldNJ2jLuGwGn7GM8c0lkIZ/8e+6nTZe5xPOMvMRy+I3XMFDJSjl9C3D
nb0OU4OIUqA8/qS0E4W/MNDCdsslI6m3pAuKH0RqnMgcxCLh+ANVcXu38bYzmDZW
obvOXRD/ZdtBMKeLAeOA/I90oE8d0bBtL3dTPomUXYNsvc/z685rQTy2H0cSYpVg
H4t6I2fQirnaDogdYcjTfi+hizWUW9OT7UN5HwfaPPwnxgXlHP2sNvTB6OzLXsaG
L62CDkJZDxAqBEud3b4RI7x+eBOMS5FeDThaDD74XnzvAsyLvlnkzeYZc72kO/0l
YBRPnOLsLrVHE2mr3ryZ4vfsa9qeB7uY7+GrvRAwQBwuQf4X1E5dedMRQSum3Vpi
OkDlUzj8069z7Sr1I2zfSCAl43c8CoFs9Q8TeCbjj6XI/M0PGUw6El3OgR5cboSI
kDtSiv9y+OkQ0KCyx47g82hoaB3qmSbxv62mpO2OTnB4FzOpXoXq12lThIL8SezU
uqUpCI7XLRkY9GIiZt3m9FWnYwUnOxDCBC62aTLht8oCBTjkJUPNLPCBDWYBPmuQ
5d6xMWZWIFX1jBunNykEZ1lL8dmOMlPF341szvPH3zKyCkkXDt5qO4pniGaRbqHH
0CP4Z+WZta1llHeN7iuffON+xWawakQuasg3mxXgFSiWUqzuyZI7n2fyceHW0TMb
iC3xK9CmOcYXsOzIdqb7YI9v0X5K3iO/wSGHTmc+dDYUmkIYIW2d3Jl6xZ8X+oGL
dOAcYO+YEaP7fh1gXigQKkNp/aCKAVnPhnOakksjkzfN7r1/HJ79OE/AuMA/VNNa
CifHE2z25/B0vugp2cOvFWaE7ebuMCVOz3H2nig17oW5Phh2WGX1mFs1qWhfWa6g
Lqasb5XBKDJJAX0Ql/g7dd8l3/nebsxrWTApS3CuH/fyB6P7Zm4JMqmmRWl/2p7T
JjA2hFQBik8dPRrna9ymo9J5mfJdn5ff3jGF755amdFeFcJNRW0UpB4m3PJAq5vU
UVajfkmVRI1LHPMt/IUoojx8QOesoXK9uGvdvj2Svk+Mnk6KxtuQodWJbJbfTFOj
rwbJUxS2ulrm0SgqGlZbCe7oP0NQOqn7BdyEhybUJPYtyRtJndH4nYZfLiKT1kM/
YqYu61FC7d2d6gtbOwnr4lUTYfZH84wAc/q17Ir0l9KVOdmrSX8BYAp2yOFG/zlf
gp520M9XhnCs7nmnYOosbxepKnZ0cVKEOJNgN0/DFrQ3HFOqANSqvQPyIBeBXVs6
MVdllxsZ4phFQokK3f8OO3bVi5m3XqsGlwr9LGq1ucIiOloIhT/N7zQrMTLQWAFb
27+UcIMwta+TR04A4S2hrEL4MMxfDUDjZqvWP/M+sFi4XgGm3OXg2RV46BoTSLwL
w96X3NBXWpcRNX3zCMFOSs2k3UHbByifklEANy2uueCWTDug6zLbMsD15DFSY6JM
hAgmEyJ80is/B11QVx39tO1yLBD3CbiMGazh24Bppn33F5YD7pO6QAPaIKObiEhQ
RS752xYNMcH6fzIqHD8yZn6pU7hpV8eg55c5LvuQqzu9sZRH42XegN3YXGD0z88P
r2+yeTCr2zGuXhEKxadZa1E0ebQeo6BC/rLA/gLfuxepOeqm5xRwTiFYLKxQ+rk7
gUrn7NZGWmEj3F57yqbVzw50qg+CmF3bR+ZDQy5RIhtBrsnobf66ADRQCrklqZrp
45SaVCgoAzSAemIsEBoZvbT7sIpV+zCHfo4+KvaxJIJxls5ENZN1rRj5oJEfTMal
eCBxjqMm5/IfkTBusXfOspFKdt0dmfaXeUVr9ydBF5gPhSR7mM2+/OcTL/PCmbTJ
+TQ66pFAkV3G+7wHMraToRyX4rVgllRKWX6Q7YratmCmnJfhl46D65NQ/z7AXJAf
E7Y7CXPsBuG4X0R2uFoiXqJVPJs8HIOU0i7U7lo2A4k+ijVSqh+ps9j1oTYssB7L
gcjOX1PwzwcYcgj6fELpUAgh7tNIReGZlfrWMzZUFWeC2nNWEirnI9UKoEGxRq0u
HOOUmO3V2PVxCPbobUYMD6lCCjCrPi3dzbkCQPGtinrcGbCdN/wHNjCUalOdbE7L
D5LbAJzfHttnwejjHMY6geIdkEv/bNtdUd65clH324hsKAGdXa0w5qoJd8I85p84
VfW9QRQyGYwhgpvAl9D+k2RxWSrQY15rfp8S+pFgCqNFH9lLxnr+tofchF+PJig5
+VRQT2LJHRowQYngY70d6/2uSxkCFOAYCfQTzcY1YnGVBwRufts9t0Iu4OUILMe4
BPBI0aqUHHFAGtp6UXttGYIO1xTutDsosVJbo3EhO5He8UuOOTUmOfgyqI7nCFsu
EQtGnHCFCzR4ZbuLeIy1oorLinhimAJwVNZ+OOgaJz6e2p1Wl6XJzpinbQqbAJ8v
MM3S2ne1+iAmy56fIv/RqOjx3ryjPw+nKVT+qc/TLUDVIraWf4S0HlksFvVVjfjg
Ud8z3p/HoR2k6gKoujL15ob477PRiejajAnKKjNzfy61PqBp2DT0tKwVwBQs1/1X
Vt9e5MS8cTOZRO1tv8M0Il1snS0Zs0cEpinKal50AZTFN4d4NYAz7ksRBe8ppUnG
irLhPS40JAC/eLKvmgCBu7nTLEGW4jkGm+KS6nlH5J4ny7lX8dVTSikIhtcPdXsa
ujmAU+lRwzt2WpgqLCwUcynmjqJ3kL9GH/bqGA98mhhC4jke5dpcVITW71bp48bq
yHUT2NCIfGLeNP4AocGy2eOE592TQb5mYtsHsxKF786KGopBzfdcWZYYIeBNjr+Y
cB/U2P5H0UFCJtzmiwo2jTT0pHiOR41AKgCIbkCUfLXf9xTmw0NDAXu0AOsIVjEH
zfiNHj3VZ4SKQ5nN2yqbPR+c3vBsyjohR4ZofjKJWi4gRP/wOpHui17YPX9UON7o
ibCuIS/OfGNMsWQ2EwFmGsAABXWE/Dntt6WmcPnqKz8QIowaFwoyttM6FdxYblMZ
dR2mBkeN4RqZVZbOcEDPoqtUs3JCC2076z+P3ppvPHBQSU4ZfWRccUQwyWIiy4fS
qpijPGp8cWDF9z3proPAcGmPebL/gpSu7lOI5YXXM8FgzhTl2VMGda4MRSt8CBvh
xTufc8lpcDwxBm7/kTETCEMci5wfS6gKVFzeABrwGnHnB3HoMd+BJeMrww8n6Urg
Gddb2iqFuK781ECpCCtraynpzfRH5MRycMhwHdiCXvgQAmvzdIeZyxDhXDRSxzQL
zfy9uapBbgGpaKjvAig1x7R97nqRgl+g+SKYCvGVR2lOpgMOrlIeN3biLtcV4UXM
awyBvIszhQY4eo0dFm5BRqmFCIZCopAUOjRaVImem4WfZh3tfZnoA8SIQL5NfSHm
bC9rbg0RhXx4PnZznU7OyQ3Hd42EZ3Vi+Go/aPylB2KbdMGw/x8HNbA20HehxjCs
tsJAGh8IyTD3/5ilY47CXrPmUGKueYgAh0vFRykbaD5yKJiLN8AXCiAzkrajiDil
bNvNoVu3Pyw3gDBkK5rOqWhoN5GnLnr3krw7NI8qd+V3zcj6NK7s+RMkbY9jZAHt
9TgwsgOjk3ZZjCCH0q7hYtfn71FPaWw+yEl4Qdn+3kvtijeX02aTZ30vQAV+/Tq9
E+D+sXwPNzvwPC6PSW7k8jx1QMeF7ntIEEHv7juZt8UxgDwDJwOgembC6EJMbZRY
Uryx6vQRBA1w1A6e9ZTHrHgZ9nwWiBOkDRL1Y2z9BNpLH32WGZsswfSs98nF8XdF
watYYD4gjfOI+VGReGRFiME8EnzMePQqx6Mnr2lCQh47XGNr0+q1Np86+oW7Nt73
Wh5BFINy3ymN/qs6TJrvnILq0QzTm/L//tmljIY31bxxstcDdTD2ngFhG4tBBN8q
6Y0i8wO9DKuWRKJjNjEVUGh6gXrj5lUzWXUhTPuR5Ui+I3OLv46EvFOM9GXZmp8b
7mnIqcD9GwPzi3bhU4IB/aDyZCZvQAUJ58aZ/ylHBOe7uNNz/k+jUDMnAh2i+Ciq
BO6rPEEdOjDPpyh5vEWuHVWJBAaTtWOc0KUpl172DUwkJcBfCHSwe4PUswNR/VtP
gcEI/l4cmjjO6BVVAHi3cyWYFvVzdPYvlrRgDIF1TNfBgBFpJZG0SRqU44SdC0qj
nycvsgSSUONj/zc5/XucgKiFo4kZcPQ3wWvPiksCJHFhh0NGS3JKK/FosXbRXZ77
SYmBuW25Yq1iuKUxxlQy/GckFZEndP3zcIE+kHVCjPBelhuiJka0d8bbx9sUHOOY
LV7Zkg4KnSRsv7V3UqKGTeKtO60tXuDdaVcj8jdHU1QgGfcK1/GbONH4FQ7zgvqv
fhQb61ZQ+2eMkkFecAMA19xfH0vUOhBIpKDvf7qqWQJUSOnIYb8wR4ZsNqGSDF5d
8bIZOlYhOMxxOZG6pQwIzlMyVTf6gq7N/PYyE3vBmKuzVhRHsZ2WAeYHaE3oP0j5
X5Wtbv/j7hrEYVt+c7yOToulm6daM9ujaGSHpHYYwzy22xWticqVXyNI0WsJSwUq
NUthJal7TVm+gKv6teQVKJLdlQS+nUg3VGIhPTgr8cu8UojcbcGb8mFKMUsEVAIY
g5NC18rOYz7wvSDlVyEKqVcigJlOtu+puaNzGkMoH2wCS7ogUBK9pq0kuVsZmoST
eH06/9FNfNSg7zAT2MCGV8z25f8ee1D5FItvztkAVOpft3dejxlTmwwIBjSgXHr/
Ub4KpdM9IarIpupUzHN/194/3+m5o1/imFYfeqy3fKGxZ7Ru7NWSZvHzZ/cKrPJi
rjjmpnXWTsOMIEO3B4RsgTnSI0nUZSxwYQISCY3tARBvCqV5G+ZEIAyl++8Z0DSi
iUFVVIrOghjZZVwd8ZxVqoXfPDa7g2tGu7ikQS/3aXT4h2d4dEWTI0ZkkVCFE2br
aq/5G/QGOhULVtJxJM/6bzsPvYuQKuZbp1LeZrM/k8Wag4w8D2ydeD31OIdQGsaH
SbvfQWXU2jHx9eiYIMtE9ct1BBRj6qgQfKJ/YfYjoQ8zeNN2KiIFe5LHqC/klVrH
s7btvvwhCgjv/FkFXo/Ah9DZK5KB6+Kb8RL5FpLjUx9RZ59ILloZBnm+r80SmmT4
w3GnBeTndoIDolyhtm7OKorVR/uqzsRTQM8P9EFgXDSw+KGhD2L6FpenS27/xmb3
bdEc8JZxo1wpvlINrNUb/f/DWTlcTnIcYBkWhV4Wg1QTa95xA1lYOO7zl0C7RByE
xGjC0+8tNLPcEYqPGkbzGaigG3n/YIbzHvr5Eqk1Xq0bqpXtJOilDtSdYqcO5eAV
2tw49/KQ9Pow0erQFgkT89eQkEaeW29jdop4aLYdUPLMX1EID84l5h7i8KJlHCDN
NtC9qelE+e0e2xQHYLMqUEBOyXSDwNi8aygKfVNMJp0N9b+rIxPCZWxnL6CXySK9
uMZT7H0+wXwq4/b+wVfV8mOFEhcD+UL1xZWmgR4kTS61YZRK9sWbo26wBZabnUCS
yxKSdq4WKA1FAOtOXkYYZ51pT0zDtoU1A3SWdETHs8alUv8zmmEoZ9KQ3qCO/VSg
aSzPpxaXL5X4D+L3ahUfCh0wIBB3AK8f1wn5XQDswZU1isud+0/nl9Z1S6NrqBUp
gaiV9OSpLFmXx0GReLvAlWvbwyl5qFo5x49BFVB6WSOiGQNZbti81EI+E4w94ifD
0r9IlmpGWJPXL6b2Ekn6tNicpXzPFrQ8AgfxwhVf7UPENbTN/ZQkeboscJifVVGP
ewMUCGQ5WmnPcMclBMCrxm3Ky/ERKKb4y7PxSCsSV2EY7UN7K4UrSK8wsSTcA77f
yZkx/I68z11XCzuetomcFXwGiIV4HP2h/Qokpgs/KipffPgK2kMRgBWz6ivNuopa
tTGSt51H/w8vHxeh77KOGUDkAMdc8IvDJEZ/URIWbFnjnkPNILnKacXXujOZ+K/X
qKSvb1jId8VM7GPcvXZvllCMUiQbNMQs1WwrkVPIgyGBKUW7+8JyzNOXL54iID9Q
W1928GQBKBMJti4lQKQTacbkteupdUnt40MXj2PMpll8vuBMjU3/l7pqNJHID+/H
9AEZa/c742xnQ6mJ0+NwouwIOcU57Kx3zCuBNbJsqRNFKAdAxgFW0yY734SW6DGE
+iBoGZzfHn6Vnwt4cYczdBAtMnLb+bqOyoowCmTcnke/GRaCfziXcFCKiN7x0992
/EbStlaipBdynAYW7Qrbq5R9WZTdTgfkGGjA9ghEi/36clEGeBVPFTWzd9zl0veG
pAAQ6cpVmjp4n/1TfsUFutYlvao1M0+x5nMGLrmmAMza+Z8lmmOu7eeikddqObvO
NPrZzs5i3YdK3ZuN74AZJxpKcGqWLMAj02F8qau1e+HAyYaCTVW6rGk62LPU8iOo
G+dHuTCDoeKpSyDdMyYiTWR9qUJ/PP3iTxu76f9hV0rOj3fvyll3MrrEnvjXnh6T
BsP2kQw/h4PL+7WrX24/myb7fvcVgedBhNFe6Ia05TBmcluvIGZ9EgErUssk+eSv
tsndkSPIACFnFKjCxklg/NR7sIlquMOWajWENDgyGA4Ks5KH6f7G4RD4+SA2kYgn
TDwkAC1nI6iVZJ5ARDigS/5uI3HmOrYfeL/chy2gMy2LnpoJPPiVf4EAkbvtaJaO
sVJxSaEpy17UmmtXdWHcn16CNuLfjjhVXVnrjf7d4urkB+Tu2U7Pic97h0+DH0ss
5te/PxKQW/T5s1WpaTtAp5jjamtt10Fh5uL4Fjez91CFRIXG3ap8ZRd2w/YC74WA
ZWgnHOccdGENbb+19Mls1HrAJRy7BEeyt+gsFEJiPKBqF05bUqIcAK1lL5I9jd6s
giIUY+kFPgvJ2GzdKBtjr7tZVmhZsx6IrleM5TJw3+eTJrZbiQQG3p3jsWCu5hjl
tuwbhKy6Iw9/1W6zP3qehDJo74sbi79Eu9/i36FfvurRYcrk7ilJRLHqGiGNi3hh
E3i6Jovc93G6iYoQFPnqy0tWLENeD1qWYfUXu4BYA1+/jm2YTtlEAdb0pOVAGb73
wexjOlWgHDqqdvEDf4tpWaKPHMy7Equqi2p//tAV5SLCrJVQcfsWQUmHnMWmAbgF
fTP0vf5gCVpq2Pvvlugu0YlqNbJO5VqKQ79ipcJ46cmrT5i09JbniINpa6B+KUnC
jlZqcaoIbD7AWemj4ZP4lPzUyyG8mdCmUWOX9qUMshHbQ5pbvbCjnWY5BfSGES6N
YxqTbpmS6lVmidzeveU8BMLNqdrAav6Kig5fouIVswP6Jr+kyOdd22h9uHurf1PY
+EVAYl/AeVwNGPUMYPnLjX00giUF4BwrLtA1weOEcvBNk80CkgyqZv5uIC3UiwOs
LLBM/kwJUdI5nw1WVrt/JJD9dn3NU1YN3mkFxIvjuaLBMKPE2Aab9VuVaAQ9Q6s3
7n7CHmOoOUKe06xDR2vNjsobWxYx5C66VWsue5OXXyydRpI0YGhNLasBpWs7OHBN
1xEMU7QtgkOa8X7xOdIC6AgzGjCKSYkTcjk6b/gfWfegdP8plFl+Rtc0mMRe8Foa
WRXHppibPi8ZHDym1gbjntpTbpKJTplPhb8DKsSoj2Ve956PXKtGmu1ew5K5g7vI
wBjkD3bn9zaXcbF++C+aNXxjrYUO4SY9hqxihNlAwdn6eHEYWyU1Ynq3aWIs2RRt
UCeSSJrgkhkIyxwD+Bdc5KWpJw6NqWfvr8e8fPaTjb0i8Y3vXodottgsWR2sx09A
VpI0+CL0jj6wKkzftTWwP139Z38SOcZg3RuCP0SQy//BCIyW4rcSA6ud58wywsgr
MhQtOALLzlDGPOKzL3f4zCEWr9on/o/sVGA8Ffp3bwx6bOjf8ytKO8vnYyA522R0
bXVOg8MHUsVyqsoZbqvou43jWUfd3fCuJml8PNuGYFEWVtWJEJXKtIUL/Z3huNyU
Zhcvs8I0pFdpgwVFgJdovwbJToXT/P/sqWc+EJlY8Jo8E1cUajOF4+Qe8oxQE7ji
Sq5otvcg0gxUkaERjwJsxYzUBCQVZbmcs9wSPa1MeMjnCspc6mkC7JVU49bcdcNK
ZPPahcF7TbdSWZdmKoPxquR1nlsMSi1KIHIB6Ag7TzUgBSE08Juzw7aKFuUNb3w+
MbjokYrrDKikTeVpTMzS1UddaQBVvRlhqq3AMlkwZC9Aqd9sgGRIHFIy3JN1Wh0x
wzkSI9jrWK0YOzKZ5qOL6DsOo7FiFMBTX1MKM95XFZIXn+a71bcXZBrIbvmB1rLB
iRB3AEYKq3FjHl/z8HbfjZvfeJ+BwKtOvIFm40dO7S5s+I6ACXMeRRaspP1+Mn+p
swifKNKXWsoLUQsOjYh5LXMWIEoivYVKZOo1799sQeA7cS9RZH/0Mt3ndhv9UH3s
SnZqRRbuMAwpobaxJTpkCzpw8AuZrsGQTpwoVwynC2i9U9tsuLbPzNmEdZFsiRXi
PTjPSNDGKp7WzQu1+Us6Zj+D/cPaXEV0PedOzpB2Z5iwSSs9judtAU//IOe79Scc
Hf3zsGIM2WNSoCErAq16FL6X78kCpCW/Ycz7hGwFj3Jrufmf2VpyRIszv0SwOkvc
45Uvx4GTpQS5VahbETZ9VYwFcrlQxWOqiU5mJyRm2EuvWHsbmPqhjn7YXKwlpG5/
TNREYKhRA6w9nHL/3xUvausODznqQuuW/vuX+vItj5AYTe7aN7oZ9xkh6rULjNJX
IaKZpZWYaIHcqwX94fz8FK9hcIs9AplBTTiVChBk+eCHVwh2k7j5DY6R7IxLUre7
YGbrbc966UaXPpVh7lQvIYs7yEzcUNrFBkm/OU/qB6HFAqGpFcgFXWZJOmV95QPG
FjVycG/kcTRf1TTO3mD87vzAICPPdN8aTaBTHhryOeKU73UfJ/le4ei6neGWzpbo
Ayop4qwnEQR2CdCxwayYYAs0thWIw5sf9pu+xA0wjJngYcmK3R9ufRmynB+alhPQ
uvBYbp5hyGIF7gxP1XCjVR9hyxYWaBMNwH9BPz9qOr3WvmA5owKfjumZel2OQW4U
7DtcbqWFkQUmtrol/JDCuiNVzP7vpo4tWQRnXDy3YeS75byhfTDHUIMe1YjvreOI
AVpF/dD8rT7HAVTkvuxaV4cWk4rz286WeF/+bUEpt08FyVGaBEsxc7/uGdWLwzPq
iAJDk/eW+Uqpi6UV6lX7ZfiM79kzQ31XAeBDyMMcSXiCJbYrySIDnv3HP2TJrs6f
xGVxyyozlIVCJCtCOdP/AfiI1R65hbGgvSp7t/MFOv/T0PKKIaqMa9iDqHZclg1N
VcybOOuVUI7cw8QezVVtIsepqWmXXuIxgYNAT7f1sbL++uiKnS6TCmMafuRfgSXG
FbB989lyoGdkVSdZoABsC9pZvUUXAHfr+X1aFOWY2Vadn1BeicTqEkGoKd+oofou
Rm3EnnwrQJuBdFR0g9vQ/U+48QpJzjRRB0D58eEmTAwblwPjGSlN1bDfX7/2+UMP
msh+C3dgrgI1NPXoQoKNHmT/HI4LD6daS8QapNiPRiiC67DaQNN38h9MqsEKSNMb
dpO1aE2GCbZnsNnN0yh4gUdUfz4Om7mDPgqrvdhNNgZA6BmOhdWqRz0dEZHqz6u+
Or/r7dJdisTjB9I/eSCbNmgjOQee/LuYRl5eisP4S007CVZP7H47HG9tTuUXKuCq
WdLFP6M8Ua/SvOwwR+dBaIJUGWbH4eeSSujckb1djJNe/drtMUSWnC/NCnBsi/qP
aebPJk3lOEufiKPwRjtvaBcIyW0Clqc5zO3vB1i3lOHtPa6rN6vO+tQcG482/fIT
U83ybJA307SaMwF3vHsRaQes6iKPjQ6Mw7mguYHgzj6wwAsM3ld6pnWrxMOVlIhs
8R4agFBfo0yJSyh5l2+tDMNbBYo3viamuZgquUmyWzxKi0gARv+BXHXG1guoaU0y
m3mhQbLFaZWX9z5ulY9R4MNqRuVMYwD96pDD1p3cxhaLG5FlXnaUirSl2KbZf3CA
YoEKO0mR82/6GOXc6JRk9bxoa+ZLvCmfa6hrji5zQAKM1uBYED3Qt7anAF+ac+8P
/7sDKBzHApd+H0Cy520UcNd2STVSdYoZiptJnfk254NcFvUZD10Y9AVxkfpJvxzF
wS5Edd99aHmyqhIrKX1GyuBQ3rXac7P+IrTBd2Fdb33ymz+7Ute5dxTaDT0+5HZI
WNjiWGQdQ4efvKnSq75sZ1qVrmtP37D+mOl2A6B4HCcO+9byDvPpz3ESqXU92n1g
ycrm7mOdvVUTnOVe9E3dyo5aY+Cn3o4BZy5vfbZpRqdmwXsdJ3xZIn91U7zkrnnO
7Ea+FUYaJ6buH0wnRWMZIagF9inXQnOYSXa0tu4iezTNvY5ZiznQ2Q3dJsHL4sfd
z3lAjdNLhV126qgyYuuy/nAjGFhOCvnhCvV4PgCAQtKlVY/bpeNcldjFqe7UGUKK
McDhk2iglP9gLWapt+T0YNA0AgnmeUpT5eY54tFsQbJO8gmae3cz7dZWtCnpK5lW
1NDTU/7xzuDJ9kB6AuvXnYSMZnODzwB53u8AVhJC2qS6wRfWA2YMzoexOek989TF
0niM8NWuAutTn/LMW7itgalDcGnbif0Bs758X6mNwh+dmr/ffjlmT8nT6wH44dWi
wcYYhgIAM6hEd8RTM+bXHoK2oedkD763ICbnaO/OzINOGiUu20UkV7naQyiFGwHG
njI6WtKd8dN3u8dqDevC+MLjMsaGD0GTxag1ksocu7WkwJCbd4gTEDNk+L313AkQ
Qy6Amf3RGLQHFRmIeZhEpVEceRVJm4xXRX0X3emUsv3yi52+zmPI5ibDQtArIp6J
K3XpPU2dQulknPYL8yYCcqDm7b/lOd4v4ZdwsqOgW9+nvNz+z39Q8juYac4v7BiI
1s2N1mgwTMW06UqbxtMFTfrC7ltFuNf1gUlRhtetDvR0PDx4TLI759k3Q/skf+Id
apsNLmtSDDNFTZIXAGJ39IheVHG9kODV1Mpe6Bw5Ad78/qpxyZQ17B4ggwMtUGrP
T5DxjZJ34O+PI+fz9seyW9Q540xv5eaOeR6FB4aACmKZ35VGJwHXTFmFMJXDxY0v
wJOQ68IUsS5vxdL/JdmhTyV9VtB2AnJfSVaHq+TW5KRjfdB176fsRc9IrLwWCHqK
qrsBqIAG8DCU6ZPY0j46RvaCp1vVpUeI23GWD8UO/AzZQmEdznQPexeyLOJNL+7p
UG0TP7/D6nHyD/6dAXmHuIpW9kA/tleF3cLL6qq6wep5/DQZCQmH7n339IKjU7xm
cMBy2wfYfB88Hg0gOO604W9nJf1VBukX0PKoqZElyyuRAiUEQnQRSoOXwhSjKxC7
s60TSQX/zc+7vK/cZ00XtBSajr292PJ3xLCwD+4623v0B5cJENSHIiLJW9QxPHw6
7wC+P/V6xU3vp8sw2DcJbdhXMf4gelXt+fpkgqs0jeJwC7KlK6RONPNn2XVcul63
ca6bxvH0IS8JtnYkxmdwQARP5AHJlwe+Khy1m1OK0MObSJVUhY4hr3QmJnobFPVl
rIFndUNs3p/pRYJHSsnCm3c2Xxv8JUfnCOqSorjozquEeMN6EYjIeDru2SYccmpZ
ykV0C4Lj0Cil0MX/uulUIVUeHf8AXTGXG7A1smfaBjpTwhIael3HwvDZ3fzNzt/y
/VES41qkEC/DKDF+t/SOAsd0k2o50AbEAHn3ITql+i55w+j8EYDXLOWtgD4TQHSL
sjJ0G65V695h3CRz8q64GeSOVwmZ5E74tpvcotEhdVX5rd9mhfEfra3bqpifcxjL
75gwMT+GbpzmIzSiAX60F+kIq740xS6FU5VHDkxa0kd3VCTGUIUv8zXL7d2fsEse
GnzgRYpY80taLyJ2MgRk9DUFGshD/D9Z6uyukLtOMK28qGT5gj+/kejCKu85QlpM
OrF+DufZdu6l4F2bLHLhI/W/kiNv20GIRhXXzXSDdikTIFucXrJ3Gp4AbI6l0aUO
1dFOT5H0URXCMA8czVLRU57a2paTtjO2mVNbMxBaLGINie4XUza69aZ6eeH1R4lO
vzpdJclBV9Rb6xkJs3GVb+lGyVYjJf4bHA6EsYNNDhlX9vFync3fY/2p1RuJQAeA
xct3QlozQCI0w57g0LV10S20NHD0Lpm5J+WLKba7x5OqRFjVeZuoK7r29Pmeftrg
qauI72WTEbWK7dZXma5I3pgf+a1LjPjubcECZGc/yxbP0VE7O0Oxu24XN8Lf0eTt
WU3zfr2OxwrlvQ9NmKlovLMlzCq+1rkLneWaRHNwQPrZoY4F8IMST4WmJ4Ej64xu
P+BVL0nrry5CACVOfefLPRne6SolyxzE/0FbP8XCNSa/5nbUCiMpovfHKfqCzgD0
t73jtlyeEHrq3nm/Er4Ebsg/cbjY7fLgECvLz2jYI+G9DChDBcmAVcFpSOQF6pLr
nNuBGlFHCbHwI31gJEtVdsQezU+2svWUZrugb/NnYpTcF3ZcF6G8scwzqsKMRt0d
+24WhHutc0HntSDek1b9rgNr1ACbaqKu6Rm0FqLFRjPaAuhXDr3XwmQqXULchbEF
PHrk835V9mNrleR2EMvnb8MVirO/FhsM+Kc+hrWOKbhCJc4kia1DIiU932FlOnHg
ZHD/31n37lw63vIw3l+Q8+HZNQkb9GFAnxFHvLvjAt+WuvJV9gEDD+E54I3rJLK7
8DA2/RFHSHV4XospEVSdv3kHP5l00cOQSiCYTgbLANAFBAIu9Y19Zes9zZgfWCeD
TYTuXXRkZU4yKTcvViXIR0iKtssSpHLD6Lch5ckIa7pEOtkWQ6A63DTyGwj5VBZb
0PVXfQlg1ZITGLR7jdWWJ0DHWOLtdYi8UT+sRVFRZ8T4jO/4Wxb9JBfIE5AvQOCH
Uc9Hrw+r4lMTVS5KqJ5OwCIS8Cq7lL/uynXE7xl8WDwAEy9mWk5KzKZmctTaxDbF
o7LiG0xeKpREKK4Mb/ozToFbqoBf262afM83oF9RYxIhIVcyM5np2WZa3fCKauMa
EEsogpiaGcZSb+wBvHsmdFQSwidzy/uN7ezu/surEXiHEJ8Ilqihl40DmTBHgvJA
Ie3zc9+wUaWZ+oVBhi728sbZFECIE5EoXfp6aT9pW0Gy/2to5AiyuPg1hIftLlqf
f937nuLYW86Ak19VVdu+6X+5J7vS29FpGGhHA0SsQ9Zx9CkVHaVN2awdA4C0EvmU
BD4X2GEwEDyosQ6HKisv7P4s9J7DbTOTa5eJQNrn5WWi5TMPj0wSHts3GBWQpbEH
wwh11S/gaoR5scAQ0D2YhbKEkM0wI2AD4xJAbaPRnLnDlw3JPfromRtemPgWyCnN
KiM3HZiJwxbOrk+owXDbPaP4UC0UaXxMB1lCtogTXxGjhWDaZhMzhYKldFsf+O4L
ZvPJtC6SsTyXsUiJqwlwsdZhpLvfKg9T6sWdteXNkeSxHPmJxMfFcq1fQkKKx3vg
MIhoUDCYeaMusgiuj9QDS41Pqcu4d2RBf04pw3l5Th3H4ZUIpUXAKUN4KHB2Ni3h
q0OloAxAl0fM++cWS2njqqE+C6oS7dF8nU4XUVIY8SkUx/L/UN2rLSFQ8obpy4UN
+ik+8lneSmrVvGk1trbtjY+wjl6SzdBNPP9LOFcKT5WRgw1CooY8hsL07S5DZZcn
rrRGxdItOeIEbmfbFSnnMpPZr5l2zyquSYU/+GJesMIrh14ugRQxnGxdeshRAO2C
756JhQJuG/5jCTLHcgE53+ArO+E5OHwB5HpxFQ6dupk62tU36iEgDFhppY02y1cW
Ll1Gu5WysZJF2kX9UkQaiTDaMdIljECrpDGPzQP8HnI0Fwm3yjalBsRCKbTkLvEA
+hvpvK/SjkL8H92WNhbmSfULjk1bqktSHE/ixYKf6XzSBMMqwLJ6JyP+9oN9GhEp
tuAmKQPI/foyRH51xnptghcxigwF6iDdGH1zE3tCdhj3WKauqIlzPz3Jf+yVTLP6
JLUWr0nBuYp9ewnXEMwYWL3yfrNKkldFHL9tl4O6Kw0x/CrMf6SjfCjO9jHtu7if
Zz8j3eiCZv8ii53K0e8ghCqVwiwr2ilRhGzZ5vIGWM/kmdiVQFgXH1wFaYQRptvy
ODgfvGc1yy6qu2kqbbx10CJxwOLaXi2FCyMGdQf5nK8HbYAwnYm3fyW72SzjwT0V
NlmnatHoe78e+8KxWIS+Rhd7lCOFe/M9X69Pvbn4n2slFSQ2s/vX46fN19GU4ifG
qJndICTd8xWPI4h5x96UOeQRZunQW+I75q5HiozLkWswk/HZC22ynbH7ZqO7la37
xXBYSwPZvjk9Tx09o45e1xSUVMo2l9k1Rmgql8RmCxk/C2bGhbzgqcmTLm0k78YM
1fNCihr3IaWrx5U+PnlDmxtp+Te78U5H4b787YCrRizJeXTL+Ku2oA3LrrvlGUHp
oVg4LAxj7KvZlFrR41reo1By/j4P8pkDTtOcdc6sak0fA8BqbgvRM4Hur77gKpeK
g3kOA8NGBX90kQzoPMIkcfiWBvachjgAyKAMgLn+hUlFK44MoiWwjl6j3Z2zD7ts
lgxjXh19CIXCZUbpQQ5k4cAzavWt3RON1OVBWkr9xXkNLjxyK2i0NFOFnvwHh2ve
ipA1rYoXwXt0K4MR+Rba+AMaruQcz0/XbgeM6MfNvo+Ush2m5kWLq7k0hNHSRupx
7dC7O4OOKQqrGeEd1hSOcgufxzE1NJvpnmVpND/Ts083vv5YWKsTDU7lA1Khzc5z
MsEYTVRSXL2qBBQzRKcwB1YFEW4ohk4LDudCegXJ9DV4NAFd3I3ne3s0I44w+Uw3
vADfJi5XIb4CZVSQtDD5pLCLsV6JTDmgSOCvLLyMD18NevM3vaJZddiVIoTqC7nA
QTd+EVY/HkTcjBInEDzrvfvyz+dZMEg+RFm1OXPqhS/53Bh7IRWrT9zZuuG9QXn8
KJ0+LoeoLV3ofcRwPtREmDI3NPqyJOmzjG+YYf2i2K+H/ZQE8EHV1N/4GX4buh+B
RYDDem/VtoLgWGQE+IJPsaM9Fn/zQmJk9515gP7QCbQVjj+AMkB8Viq+ZsyYbOko
OPVuMAA6sOv2PUqeWiOxh7HT8GQL6lGCLfefQXgmvDWW9JGf2mLYNaOC8IWTfWfx
HssOR+q9TYbb+O9iNEL6vhuRdsCoeMCuecpa5X7FcGsXhJIcTMUiQJ6Dunb0FuSw
929U7UmF/0+I8pWJPaTb638haYiKzZp99h8yCPJrp+YMK+3o1AE/GYosB094Bnr5
3ANe61PrOI2Z8lRAkxs1DMkq7DqgxfB5+tBOhc4SGz1EzSxJ3aICS9tU6lEHHQMH
siSLRDLDhGDooHSTGhUghB/P49VwRwTOLYp9mqnBXTROsMlMumb4MtYE22teNcZz
Ql9tGn+u5OS1GGnBLMObQ+F7bNhHRNTzjgJsrlEFE/WDbDoF4daYYn7K0zevGYpw
XXcfIaEI/M7vT0/yd2UEs6hthFqzs2a1cREJYP2pv8TjmA0VlAyFD0NbthSDjG3J
0GQR6Tx42YWd31Pdsav3ves7J8G3QecRXX+mueuKrev9oX3RCp30RmV6REXHA475
blOJNGXd8HLv1Diblv32Ncj6I/dcyoZAXc9y4G3J8bLrQd49u5J2lSrhF2kBqtNe
SwA4GnFRUxRU0Aswe2EYwdmvEh4qP1zSOBDxWFKyX7Zy536JPOEswrREFNnSdKuq
HSI0IpfkE7AdiyzfyeH0pdgpGZMIVxVP+zKGzelCHAYzwA1Q2wYGgjfFjVZ/E5ag
nM0e8pFDVcw21vLd09J3cmcJXmum864hkaz41PDWDur6kuDv/Ok519IXfpGwi76p
eZgjzDoZDalQ38keLnMTnPEArm15Dl7wFpRfBG8LT/pp020jVVzhHbNgiNGsMw30
cvKCZpb8n7eWHP24/LuZSU1zWeVGb1xZQZied5NDqIIqOz3WpwE+ofYg15RnV+gx
cpp92ppCLK3mk0IQ5BlXaeK16vOW609ZFv4Q5lfbu7GKETYLkxfJ7EqfIZeVYdqm
P0cGCboe4i/VtVcdtBUBaYzJ9VI7vuJeoB62s9ukChNIZ6w0f7TNmgKRiqInKWKS
sBRwUh90HMwcvozvMy9A0drkkMl59q3M0JUtYIV3Wg3/yZ434g0BSM5lGcyDg4wi
J9hlQJOd4Xd2bLdtQsDvaCdUvFjR5FyaVQzNv7Mr08kjTgiKfsIXsr+TvMWnWCwb
23QON2KFrgCI97PV0ySok3CrIDBcxupU6SoD284waZdjAYdLxb4TdwWDjGHNJx/V
SCjiwY3fSHnWo88foplPqaMSZyk1U4Rp0LMMvJll444F/IOr1guyRABm37Mjgoyd
RuNljirclCSxx5C4pxzCENq50tdpFYEog2yrfcbZEtbS6Bzf5KgcTZRRNniV6jLI
3zteQ+xkgQ2p6fbNWoGuV0f7jAbeYsjWQP1b2w6Fk9JLRspfbWnm4Xryt/ataqqp
dFCDQw5EfqChd4wOEtoEN8SiYfQvanTq37reDuPQ9l5Fxu5/dQ3dd5wnAJ7bV0Er
BNDPppZjW2e2pwOVJw4KC/3E2vpHw+ayPPzIZEqEFCJFyCH8oMZlhGzdyOrNWfRa
CnNT1qvTBXSsXmw6j6WLffwiuasnYnx0UDfXYpyVqUuSPolx4twR3AaO3w6rmLnl
vZKF4TjDj6SjH4LZw5nyYPs6N5sfq/vQbC6ITiHlFjRV6PRtuN2lmEToXY8k/jco
KcMY8ZmvsRvm4+Lk1olUZyL6As38KAOvPv2qGX1H6SplGAgFrWd6aU6qCIn6BM7r
tA+2kQ5MFDV4Yw68oww9Fng7l9asqpTvE2OupcQPboaNw+5pNwRFw6wgo93ipV36
BcZflNtJDyIwgk/MXpkQp7psgeJw+wEY343Dg4e1/Rogap66ryYbQAKBmn6Bx8hS
7KbihPnCDMIe3V4FjywYUkLK3o65A1GNlJDdXznaxZmxKGcnbp6MEBE7LST78Tin
7rA8gm5t7FUGmB4JSjm+9XJAVhJHxWMiajzFy0d6PwBe+QmulVmlFyPo2C39Z9P/
/6sqsXHN0WeRYsQGqTGIbFK+6bICpwSoKJkBg/EHM3G1rghEeMn9WIm5JSjMnZqt
kQJazNxgc3xZF921dFlohekOfXHTc+R/CTUnAv7xemeSI8qZml+ZHkx9z/KjmWDp
zWXB+hEI93hHdVs0xDa5wUr9LVC/ikuTYBXtEssJ4WVSrO5I0nGC81s+/JdnjkUv
i2ODPfH5ypwzgdurLUTfIlUFhQ20zIe1l/g/z63hV+kArTVdqg883OAoRTy+vNSC
z+AEmaxKMgH3vuRJ1s13lxsGDf/VOGsgYr/f9c4PuQiRH0qyUzQak60UpJVSbIz8
Vh3GXh58oe4AhUqI0+pYODaOSqYGrOHxuoXpFs7ybra8MdMB7D6WU0YOODhmq3mx
LyKRPTespRaXUvnzq4FZfUAZEQDlypbdfoVmkEXt+mn+9wR1J7gIQZK5DQGwZMXi
Hlg3Qo6rwpgwy1gdH5DgPSi40VNZvv2b+EX2z3LwIKc28Ut8ciZVHKhloQe7PuIK
iBcCfJLCbgW+NPQu7U57Wco5+0enr68u6ESCWtCBu1c17Rsn1EJGvUd+oCr7BQYp
D5EKEigEOa6Ls1uCG5ty2isS/syA7fU5FUMrTt1fy9B4q4AJOFAt0mLVIvF+R+e+
Z6aUTXYmXIl5qExdeEJG33xupwuURkvENLEP3DNwnGSxhVUh2WXHOhBeCE1nNgJb
y0St1vxkDBxvYXLUIDlN98whNMtJhT/NcYrCpIOljm0iyK8CaBOcVt1687Sivo/Y
sD7C9mnkWhIKR1gSuLr+X43YvVuCjZB7eisl/1lzLS+60oOPAFlkdxFAhwVU60hs
9Ogi6DuL2rLArIni+u/dtiyh9juKyJy9BZAI/dVwDGbP0Myiy+U6bS+HsgV7Qymg
6dX8kBaxE+gVxn+nD5hz6cZUsqUGtVX1/yWTBur52BW3RLsXgcTncQbL6frN66BK
VhTrrW7BdJVsdOFBehMsyAU3+0ElOlRXaMMxcs1YFW2oZxhNotXAzY7itAmrO7+V
uR4GH64QxNiWBp3AlJczgTt1omkYjCj0EGjFKpmbgjojET/Edf2AN0kx8R9g3PNJ
+qBQfzPyKtx7VDvkRi1yAGHrAV8L1gqZK6+DTAyr140NPaFkjvLexTttYjrTeGEB
8kpvlWl7noPBg/e8625KlRZ92rNYPH4xlbHNcFPs7JYZQyUbfNNwugf/R7DmaBIW
NgJ0YPdyYTHVr8g8uQps6PfpooYcPszhSTfQUl3TlrVXN2/G/9JU/Z2dKZRVJOjH
ZeAObNo1adJWEoh5G+mxv04xFzLULkOzFHChyGP9c+57z4smjwsqtC1846ILW6Ee
SCmQmyD0KmcuIGjk9LF0wKCwqDXNfEE9vERmbopyPGnCXY4nMJyoqg0NpmLJmmji
NGhhDL45F++4weyqsbTK8Kxn2vN7jH7orvINhIML9iboeoAx/Jn0sFfWfPT4lKGD
QH/Oaaw5cdq6sBeS/ByrSFCrI6fxrcPVPuwc0pdoQUNigoiSxTXQCzf8pIWEg7C/
+QYhM2j1/ZiToiXLjm56/ClmEJBrR8ymFyphuZx8UJ4eepoShf5nBVOEpQ2NxNVe
YBB/vvvNyUv6wepwA9fFFwnrbs1IKRIKdQ+RlotLh7R7rYqp8OJRE9sJjnq0Ans6
BCxUsv+zA0ZD7sU6uaJvOZ43LAiNrmF8T0LX4gYtx4t4w47bqxWlRmNA6O7y+9OB
PaeFIhCqtbgSO3tbcOnviD+O8Bgv4Ssbb6o7K7XQ0F+UxWD871/WvLPi6xOVeS3K
CAA0BnqDjJj1ajnYOLR5ZpbYFGel/KIXiRvQcEcEdnWxLaYFET+VjI7rioD5lgNk
fAyIOdWN08rELxOFGCp6d4bzlbgN3qoH3Ej8X+Q0Ip8fjWiVRa9ZGNSYO9ZhnE4U
NMjbE2x9lODipcmcwbCHAUVC/cJRKn+HJOSE9yk0AADI2e7NldMTaUx7/5cgyGHP
eYlsioEZXEaD2DtL/A21jfgnM6NhMur6ayvqJOSrbXMQf0i99ax1YzMaMVs4ROUm
kFQ+VMi3jnrgGeoAQ/pRWu6tXoIh2xsUssmHbeJoE6Q0RI/ORTGEXfFsxAALrdNi
YDpOVFW4MluxUvvviMr288nFgDfN5cc9bIQWoy0gMi2mOPDLh3gPHXJmj7OKcTO4
tueihFMeVIi9bRmwtYfL9L8OxtGXRiwpeWVdXeAmJKtpgNPydxf9q9dXuakDDAPa
FWj9LdPFjIaCmcBvaCz0lpJQ48B4bG58hiw4pvZin14ddQQ+2fI0dn3uvoESckLm
gEMk2ceQ+1RzDGD++WtgrH1GAE+5uCiXFmXW+NgnDgj98MWQ5dbE4NfxyBrgE3jF
+XFpN7Ud6s2xIUjyv43VOi27KggwmnXLBJbUjPgOQ178/+psYjc0OCwBZdUCFsOx
SbjuNJvr/PvyOIiQ8TykRFyz2lePGLQI7TQZxpKo7IxfUmzQkx+HZSmo4RchU+cW
gaR73RiCXwPtmYUvBaV8m6hXUYUQwpHF4JiDLmTqHoDo7dLIs1AJPY2iGQw/XfF2
QJL108Y54aTCwpoOAO9ZRTmFsxNDutn3cvTzJz4o/YcrNkeUiKIGRpiXJPjIfnat
9FdmRCQbCjNsdmKIxPhG0SFGWWrg1VNw3qvtRueFWmm0eudqRCFjqR0lG8C9LKMd
xaWpAD+A9QGlI2C62N7DJCcEAY9xtdcgTijse1alcZhfHHYFdyfoPRpabG9w6yYl
VmN0ca1KBcEt83/rJ4VEVPV7YNPG5fLZw0otVed6yx3L0BoF4ZzxM8Xsn34IVbw4
oip30q22aHgflfVeNTJJ9DZjKRjk+RRgj8fOd1RjOF/yP3sjwHdHbfIeKtl8DE7C
7U/QN4bXBkHw/J7YY4gCsJ4KmV0ykNFcWH5x+XNpVreWG8l+7ZiC4dvtnRNW0WVv
WxeQafhtFB7i68EhvhxUOobuwXPsOXFx3wub8lVzeiNt9deOzzRLXrBt3ZCIAIL8
OkZEh9sLauVxASQ+RT1XBLLOH99YTEynurxtpvUb+rPUn2JWhYTRNA/SOFkpj8gQ
Z0Ao8N1wOB41hD60ErWrgEw/gKLiN0yzlevjNltsu/KjJ3ZoUdeb84P4nM0PXbRy
6FQYfCe6ExPWHYlySUgcFX0LYRYCS6P7GXwg78EgeJQk2UOeBkew4+GoOw5Fzffr
rGYNppV0F6xUoi/VSQOd53TTbD9nI4FSemx6B4jqVpt9eVLRZZpcbVsujZWlEDU+
3Cvpub+VE0WHDUHN92k9kxVdv2u9B54KiBEcOapJ/xhrdBb2J3fd0ax8hOPHISG6
BYfeb1Oz4U4zrPhvSPi4NP1WIj3+pjn0iL0/EkMKxPIg4NmKTYqHUKaVFQpXQb/e
KE2vDcm0RCmBNKnopRrQ12JEm1eaa04E9Hup8bdOZYjvTcBPUZbXvrL386Avpb9m
cN1fuAbguCks4dYC3jcpXQrMLo5EAjPgryUVBrfDIYT/mjPeaFKOGc/hkskFHW+n
ELz2OdJSap0PloWI2tyl6aMPsGp6l4HLsryQ0/ebKw9c5CVvNfi0UPz1dELD5sKJ
BxAJiAeZ4RJthaXCyarEJdQiiIcGJE66ANN2/4l8a91BmC2gvUaMj1611StyxFbN
3mhM9pLVTn5yPnzJZRo8JvmXjurN2+1uQxVJLR/x7eAGE5oLmd7wHhl9wqACD9yB
9/O/H+LJf1Etn6xS0sE+lTnCyXZYPbhdAZXeMyc2AIgJ9CdICzlMYbJ+xDFb6LZb
/vLXXFqkGJpy6H7Rj+ppehBmuvXuRJsxNm183+jlwwvpCAz+PRyevc/YaAGwAZjr
IQS+kg3jYypDvi0NBn+llkTjE8gY1JouJxNniZ/6XKkZNqiEJPW18dW4FTPBvftP
jUfQ1IoXqJCHclgmcmoApgMHu9BAB7OMNy31gMy5X3RKCPJWQXFhY0bRmYyNGLLN
naR6OwTWocoyRGE1U0hoZqh97QJOYd+Rdyj3GC+9PakujW+UWLp5WgJeJnmBVEgU
i+5P9cJC3jgkVDkvyaumoLtaSLzVD2tG+sTdvMZyq0O/Fm52fKpIzrv2rZdHXYkr
B01O9ZhiXkjOd9stmAHtrKctClnRyS/LPlT9J4wZCCCcHNeqTV6cACvLCYzocA41
I0cRSyOdhJfzRCEIkdzHtafZKFsRyv6nfBX6HTZwP5h1EaGJXHJA/e0rDnj8xxkY
DmXuWaNu55vjjU7fHJg02BkV4ltYwjP5OqRUOGLK06lUN4r1oKyUV/N5c0Q3dUAi
C5DolAoHva5BqJQsllvt7ZziVaoxOeq8nK6ENQIyD0xSFMIT1nikU2ea46wmzliQ
BbbbgSoqfd377KnIuPlQVkujuLiiYJZ4Xu2AuPxuDCHXVZOghhhuTDZ6+7QwGMOz
4glpwxIFnDeWYeh8hq3l5zQEKRDlC9M10uFaTSa3GhKw90NMgnYTlNSPnwCCh8eD
eS1iiLbhpybEpAQhHcs80byrG41dtkGKcmbCuOlK9BuCpXvb+Emdc7zcqjMoOGmE
uJ0KEh4t38UA8uTtJ/mgdg1C0G/f66z4wVlyiXyAbCgSZw+hCxXzYsI6qGdoJQGy
hH/8Js/aNv4DNKHfk5GPYhrJOw2EPacv0LK8+O/+c4FqBwf/P9/v43C6wqKeNzr7
/DGKGVmJCDrkdEzsOcOAId2YOtnmPk3In1ixNlQqCQxX97+OUsEo1Ip0v6iMvxHR
xx1bjs0+Ay/ON+3jyBA23m/g61Jg398D3k+lhHsQ4k0iqqVmb2LDrKo0/nNz8VKy
QKfJWHTr+sgNjiUnweUoLVa4CLFOCjQY80xlsjQKY+MuIWQQNACPFyYA+bouDlu+
Xeg7k60k9a8NUq2KNhc/u2Gq5osPVfCrgHw+hNIR3IbgPpSlwKRF2jP/wd2ppBG6
ZInurJ3LgoyX7XFYu8DSIMYNMTiUmNYMF+cYzsII1IDDndsXNS23/OUDWIKytZLQ
8GKof2buesi634wUZY0W2WUdpcY0ApbMZw3i07tUb3blPVkfgsZhvdXtQNJe6fQG
+5o+jbRCePvLiWBGKn90mmFI8e3hOTUC8XCwDi8dYyoh7Q1vB2fn41XAuuJxeXzk
Ok5rwrAjnBPD9Cag+JOuXWvB/7XSv8n4f6f83qsS3x0cOzkypNtfAqgwmnNOCu2B
w0iXaKLSRhQBSiU6p3SiKF5n7YNIPU4YjyweZCPLoNcPXaQgXRNmj/aDaQcEl9+c
JFY9ESHnrozdJ0n776TyngV9n61NlbD9lrp9xAAwX0xc+L9n2OBrTUjCFCu6RN6x
5qzAPdtf4VLPvmP78DJJcvPNKQPQPfMHTvhPd3ZUUuR3DFjTYgZSQark54AGrm1W
WnjLrjHSOeYTdWymAgZfEbzi7jZ5kwdHjBndCv+bTJmeQ9814qveUlrZCMDx1B1h
luXCycBNCZjhILTNXDvlgl8WR/qneQtJc5yj4v2eg+9ssoneyPKfR61amuEdRMOi
qYYKn1xGynwwobgQQlG76haxWb6oKmrLxTd4HThG72R5Lv8Oug2qZapVyLOqvX05
du978ub0RbxXuttvfOvboZc5XV1BAKBm+W4wZwM8NeEM5aR4ig2osJ5pFVuf2zij
vqbTjw6mgpEL5BFwNAcIHsLmVoNrvx8OILKdco88412AstAIBeqpwuEKRfP3cTqv
+wX0xseT7NVsFJpvHNkWfmitOjqRxqBrXWH9tdYXUvd2ZLdZwK6diUYwmaNpuz8V
8J7RZ+xHSKiCbrWfKm5iRbruuX71RmeiAR1KeNinTlhKXvohlEsjepLsS2G+nX6a
fV3Rllmnc7X0SD/J5no5/5GX4kY1YqE58JRygRTba9cYAvJcVIBkG+oUEZ/ZcuD6
PYGhswTrrqtDUqg9CJ0ARVCiUUOVzGgpzUICgRcUGQlv7mUxOmzd8VlpaMoDXxt7
ks5RFegk1yYMh+Y/m/ePlbp+Mwgz5NQ9bom8N176qCdY9K2vaJ18mqrFHjJAV6BL
msNKYw8l2elOILjdmwVEj/PgY8BsdfBCRFzyNEpQfLhZxfF0kOcP9C9S/SvLGZfb
qXi0xs/NBa83RwH8rMAl12irOVdGk+Z/RydIXymDzxscHA4KPuHKdJtN++wmymoN
VUsmdVGgikjd5kmVnABWfY6hRJYJQbH0CCkKT+zo7cyt6fBHsNiFVtReDCm09QV9
yk7nXnw2+hfjsQkPGlUYKTjGgwadtyyJub76fsKlfb+co+TfFQYMmHth+WOts4xv
h9Mf0kAZUyT8iRwM3Aw+Y3BAUZZd6LYA8mUlkMMYnomAN2LGtYn1JMp8kdxY7ICg
k0YZP8Z5TT6kfpVIa1tRrj2J0Nh/95IL+Wli0Kww12+HhXDDomPv92K8uajlw7AA
zXK6aqzNhWpXe5KIbCXHdyYcrDdPdO5Ce0f3gDMUO6Q8kOH+Vyb8uDqbAmfPUlaK
C5n2rL5wTOgwtZ2Kp7OeY/QQldVAWzAHZfYQhxS+8UIK/03heIzZlabwEfGvpmCc
0+0hKu6cqFofsqAIcmE62JEKzphCiRbKYtMGLKge5hFFo0pK3jfPthZS8lfTDCK8
6INljdfsiMVJeO+sP1rCY3tcpkQQhBspo7P1rZfpE7ZNAEOn667A1d6Cmp2bwDYl
kuSRDSJd/bHi6J3nJ+W0P/S56a4t7U66J1reBYunJ/IITHNae2Ee4Ij+R8BV5tb8
Mq/zJ8ryV7Jp9jAxtBnOBhiDOeUAsFLjPzopP369GZ7lh2YcE+mTlDBmmw/KnMxM
2S5nZWzzRd7VAzcaN3xyYM7CbHC6KO81cGnjE3/Hgi3wkR/jaL2fem9pmWvutzA3
ty+Sa5JJw43RZwiohaqPWDA+sUKjSDU356X+XrYAgXdWVctA0nUw/MkmdlywC8ht
Zd0a68T0MGe6xKylRv9zwcUDMQOQZvd2fVY0m7Dsl51bB5/QRv9rbG1YLX3kw4Mj
ShpKeo7XSNiHVJtSFne9t/OSMDAvCID0K2CxZC+aBnpjWPsj/kD8cWvsKjLpiSeO
HhhskMt6SUB6DD+G4My23YX2PUDeMydz40XKqMorB3D0dthCvbEfnzH9OOuXjM76
U7TLMJqB3p5YQnzhsM1gfhWnVDJlY+TCkcQSf71XF6QevIkYYRvT6aVpuYLsFKOw
c3Dimt9LplRhoNAy1LsmCUFImnZYFn1D1PrIYUWJbn4iqe9MEJprgOCIZjGhOA1H
/zkF8viHjArOhJ5IxyjDG2F7n8144Y49aMgHN690ZXYkYhEcMZbT0ujMQZcdaF8k
NEC3YuUdEQYYY6NPHks8YCv7xMfJza7+NvFJi/9TfzzXcKSt/MUyCxLnQe3xkd7p
iPYCQfDH+D4D3jL/yyWkkZGu6fvBoVaWGegPtu9SnKYJdbyWAinDFVGXzeVkYYRW
dABXtagGhVuza7LQiDsT64ZJ44FMP5695Inos8OvxDOgVRvdSyWfKVbOf95F5fnC
xGPf4xrSP57LelZPIRJ8/eUJqPXY6Hf9QEfz0QuMmVg6+isZwPJvABlPH3MwQ0jX
wln1z2XR5Dq3HTjUCeQ4GDdZKo9VTSR3P4xfSgzKAcXWdGvoBgQt5VWfDl57WKqr
RJGPMgZ327yBx+SXqD+LJw8I+Xh12gCcGJAW/3gH1Yox4pgWETeFbnzZZjgAmPBX
vwFVEupvlVIAYauMtq5nlUGsIWuQbpnw8UOiMUxObmceZfix2Narxd3qOFb3eA1t
AMh/AOtOl7/sQA11KogMi7PqUI888xXLAC/srwACbF67K9brGovu2zMQnIQryoDc
LdwJglM11jqkYec4Uyua7xO6zmvBvAr0apIgxMuz3qg9+1IZcEjng9ZZ2Bb9w+W2
gZlRdHjB+uesxbBDt3KCalp933L93L0yRjSO2cZeoT578mkSLl/Tw6zI5No2Z27e
pljEY4xR/ZTSWSoQm3cfKdqkmUf+dP2D8Y/JikMn128LDmx56mu3R3a1GfMK58bo
LiXAKfze0x3YpmnBZxVrPyQ1nQxMGUbvgUwLwCTdmCDqFFZDyICwb5aCn2bLGB+K
x+RWQE6i1gIorUACRfQab/R19dBeJgJv9JOnj+rV85gQ5I/MS2epHAkyalDgh1j0
LhgrcA8Yphz2DnXC1JuZ22OIpQDEJufFdGIJwJFSVHklpU+0R+QzURfnbKb+aQD0
VEVFsj1y6c66NcjZJMIQ2O8WuW404d1Kqfpx4SwzBXupPm/XDoX+CRREIdOf7DIS
IaQToprkcgihsq9AcfVcgpS3SDkaqsVi/M6ot2+SoqsBP+F0tnYu8F5l+SLePIK5
/rBezxIB2V2905Mw72UJ/y2nh9qexqMXyGmEeonglwrorgyefUdfGGFiVT4eaoaR
RSESe+A7eWx/gaIOp8zxzTflRGmfEcgXZ9z5Rj0m/zmO8waZ5M7Vg4YYxd4tLkdA
XPY38dfsULVnR4QkRbbrGZCvlm/qESZMME10fJsGJ5oB+FXIJNR6BYEkjX+5IKGT
7JaiQDlFGs85z4NTUQzzLUaThhr21ndgCV9i9180briuR7oo/OCiDTbafdJndDit
BwUUfq4+s676QuhvGpyoDLFdMAyMpbj37e9GaJTrzdT9QtEMNu16J0qCOGHewg0p
eI3L8GyY5AApqRMQfimUnsQGXqbdvqp2QtTNLLKtzuEox9XZSpHWBijW6fiLBToT
+lI8lo+VEnmR9+evvJDxv9xOVBojNaFVCBgc0HZZPqV1Y4TtLZS5ipzdui5mfQEW
m2G72cY3YuSxlXruFf1IeELgBkPubmRIlXsq58IJ66DX0Hblf/M7Qv0QIFpK3MKv
YSnY2tmhMF1Wqp5Ah28dOfbZvV2vuJEOqty+dXXC05mHFITzbizZzwJOh76OoLhw
bBDO9NvCfXrViANAw2QknONgqoPOCsAbSnZUT2p7iiuM3Rn54RFvHBd1St8Us1nU
wEHlkyWbFFU8ykBgFVXxvlxVBYZE5WB9Kb0MEnbsIQGopv49YsNuLnL7ASGHGPy/
/vD4wyVPR6hP/PlBXACiKeBUmjQYsbSzfaD+5AE39gn762zvJwWD1PFbV9Tx+C8i
D3KKLGAEyRpzj5z7x8kZTqDSqGo/87it66quXakef7l7umuyiIRPcTnoiZXUTLTd
sP8MgEP5fEBfZWIPD4mktnNa1DX8mRqEa6USJIOL+jky/tpUl0/qJ0lzNMa4mGm7
FEjj8fNzxslkLmY4ZBABhFgh+RXJ0nw2hKaLvC3pAFnw1TX7LEwxypubF1h7IuKS
7rIavEmErNRspigtGb8i+3Bw+k1Zcy2hM9Sq+g+6+K3p/Bg4yXWMQUU7tW/LzLAc
rsKz0MW0kM7rARAkbR60heAaGLvsgWayTGVIjyBxqfmHo5y1l72GkNUN96g28kGu
fFiR9EbRwK3pSPOuR6M/e/TN9eqqe7hrsSuVWHJ4dQW1PBMBirVIA9vFXLTAqTnJ
gNbaSzARaW/6/TXgr5PqS5v9oUeMnIvBQrpb0TXHW7Ji1JrXJps2H0mCm/ZANze3
ZpVEoCgvt0KOBKxrYsTJyqBOniUy3s+BOd9cirYx2fwunxgbRY1KgELdrwTzy3lS
t/Q3HjnFp1fb1ZBK5O44zs3RoKLeFZaLI+GcaXZ9ir5bkgpzusb9G+G7tY8P+HCE
xRy9dlx+VTWhTvjyYlpMOwuOv3mLSq/xXlH6OoPPAZelBAqegMHHkOxguloUsWOB
ai9uqwK1xkgsLeU9kyqXB05waRdB+uwreNWKoVcaVFh6oTS3SaoGJlPecPEAeari
yE8k2KOSAGxwRqfz8R2X95DMTxjui1Z0TqHQZaU0YLFENbz5YwnD7CMlgkhjVLMG
G7+pwEdhYCW6U3Tcqzayj/1CDr3ofjQtXvWnkdu9wbi9E2kBOP2ZN4IMbGajtlEZ
hXePf/LqcalxQQj+BKJHnHA+xdFBSpU3GvpkYqBLOwFOwSQbc1YD6g/P2zZu8DwI
0KzHSBDIrJzJpTlQCRmiqCj6v7rT7vEjwAvWbywwzqhC0rpsvhxrPzn+jEG9QNLS
ZWy99xaHP1BnkWOjbzpGfB4ubJc0ZePYyUNIYqiw+raQSHFztt2aBmTHlvh+rEUP
a78y7mbitxKRL0oe4ItewVDhpL6A3Nu3YGTkDmKPtxVr6YkyjvxEhS0Ze8UmEdNO
rtNPHppiTM+8lrc8f15sbn57NWZVBoO26btihuhWZtS3H+Bi/2fiHpOOJR/JbjXU
FJLT7KUDyV+Htr0m7YL70dSzribmG2z4usa9dDfsuQ5QNxIo8ESz1H5t85YQYAeh
3zF3KuIVUSud+jJQ4ZSsk7W+YN+d7jux+RgZSgzSYwFIm36ciPrMIxLx5H71BQQt
zIH1Msi4PMa8LS1InNvzKFwQaFtPgSs8hE+jHbrsVudymEqqWXowwkHaqhCbv5y8
120NdjWpl0zwiZlsxT+j7G6u6aOGpisnFaAs3pC51TgYTTXy8BRLZriONv+PVAh/
zKO+RZg0BIwCorRNwmifWTAADIAW08Ye4QTYmzh5m/vGBl6OposT8ow90RoFfHV0
1bqNMcvPzX13guGGOH4uUGutcWD0QpZ04JmL1mP7x2zUzIAMkhRENe0ZMkDbIMBK
mDgxf7y02RWdU5PEI3f26KG4/9PvPLmqwc+k716uvMdOZ7INErFmTAGNxzQ1zF8r
2tqkIIYrKEw+/QGmvWBH497ULHKbwxQEhlvc9/ApgqhXboVexbxUQyoLULDv2/1p
hY076Qp4reHvmP/NBmmyrYNlgh/3tgvt7pSk+vBQ8RKLT1z11Oggfl5dbyUHG2Ky
EI/FZPOb4MlMLt3TJeEEdvx5b9el8ZETwQIgshIos1LxBuIVQ01lWvCSxETZZ9Xa
ZuGmBXRYlwA1fyuAr2ZIjPjJdB7gDJvFv+S+ThJvmPnESlA+yeGJIsyPdglHsIru
shO+0DOGen98J4lyoPQ7RgWdCstwWSzgBxs+zZA8MODjLvvBI2Xud+BEDrebDJRY
0FrwowaNCtIO52Mz0PBd9KHA99Z8S+LrtrisHFhVf4H4iAZvWkhPLPwu6BkdHZsI
k3+zyCUrWxflr1mHIl94CI3IRAK8sw0fJhW6Q7g336rzkICVweRiwJej8Drc26Ob
pbydaSzu1rehSomrN8tcUX8Ayk/e39C+v9FC68L2MnpmxKwkSwt1sbErtaiRDbcp
Tc9cekkEuZ4wIbxRt3kj/bqhRblPUtRyKy1xSfu48S3PIivoi2HwehNRsTSvZP1V
ejssYeD/CMhRqFTNgxxcGtJ6mtEmGFexPeZhJ3gDas+o2g6HZfczMF52tFcftQnN
1GAYmbnDTc364BBethJ4dYWmCJbYp3qBHqnZzuvkHZmJhVfgwTSnhYeLJ+YPSFoF
NxfH2vtqxyEMkDvLFq2CjdjElBVyymbMaJqIY2Xb2x9J/yOHjk+WcQUE6h2X/onb
Z9SwV1GDjW/wLF9qjvB0AVECo9xVHtbeQr0lAi7X8ugeLGr0pkEJZICRlytSrYWs
WFe4St7XJmsKZ131zOPWOrIVr2zmpsFq67xDBhXobE+39lMpre+LRnkaLDjcKPau
S4ahx31bAbgfzRXMaIA6ADVp8IHWU+kjL/Ky/45t606GMs623fcYMprNfOcj1Lqe
xBPSI9qxeOyMSOhwgaZchx5cSL7J8rjBt3QdLtaWnxOBRSaIQ1x5Py4Z9tul6hKk
LtEUDYjkCzxPR9OX1TSEv1BC6UFrAt3ESn8dl2RS1EzDwqsTPUO2pKu+QAaRmdDe
oSSimvFCm8aSezVwvVuAlHiqsLmgHsBOqs/ha70u37BZlsS2R6ulGHMG/RnhRSax
FgJX68bMRj68qQCg2OgeCAhTvAc6nKKJMHDfMtcM3waCg4wUCPXAVGyhL+OJvuuD
+EpdGGsaO8/srXcxEvCR4/JMGMgkq46fbBcDjEMPSB4xr3xRHDbsDFzrIIlBWcPz
faZDJzaEI839fn8VVICbXaXlJRi3xc3XBgDDnWHrWodBj/AC8AGQ/xa4OlJJeFto
Hx8FpuMXGfO9BxXIrBcFQmw9vztrlWWPR8FUQyeWqKTCbSqUNBTw4V374DtBauVK
9iKkqzXth83CPDQDYi/sY3m2A/aDWLqVRUCa3AjFhqcELzJfHdpo8bRyUHvTCs6i
ASVlkEm3K6dTRurfEvJqfUs8vMsfkJBtIMgt1x8884nS+dHcyu2mRSfASM9I3W0X
pLhf9ZTJA2iykvNn2QhF9PHeFtImZE4mzpzcXAnxpWAn+1cGU567/BKkIgzWpLGw
EcfV4+N2XKqdca7vDJVUXalNRBmpBRqgqGNtjGfvhYYT4uI7esDcAauBeG5nUJ0U
WAYu2qLF3QG1GTshiVV+T90Az9u3A5eBhOHfOafrNmUECc0keMNwwU6pQAgl1PLT
7hzfXf2as6InVI02BZ6z/+UIzODGKBJl56FZDxGC/JFqSzlfZchvPIf6F6j1TqED
F4AdNqD/Krg1ltKFcnqgdZGyLbshms9+nWShFjowl5vuVta2mM6bV2Si7ksrL8WK
ywBN+ysi4LnDhdlbCjUOWnOs5mzNfLRE0U3KFWhu1WNupEYoytvWWgN7IVuQ5WDt
c/np9AvW1QUqbt4d/rkd68GsaZuJoA4tkj0o9kvbRONbqWI4oLDISy+M2oKx5se4
c15r0kNfeA9o0ATO2BxnyFG3hKl3vtSqzdus8NbfWuSXAC2FdW2OH3yo3A8+UGmm
7MSJNmAt9mkRj3FFbBM2fkMuyz0T0pwY0fsG95v45NDKP4A1hllBPXgpMT0nc+eo
Vg+MU7dklzNd169rg7cMHMhpDl1iWi3QtTYyLpvGls6PmHDTtshqV6jtVyADclqL
T4JUJurvWfvGq6g4RVPIcXBfppfNQW4H4kukiyMAsqWRPpi3QpfEIaCJafNlwVAt
wLj01MRQ7cKDG5d0EYv49b3U2fK70eSsLUcHG6rU9JoqLaUPthd3wjGaaX5peKZ7
ow/4AWsE5gz054ktQxzIL1U+pkh6PWTC4Gn1O8oIf6/OlXv9qHAgC8BB6Ld/6giV
sOmrvUjd1BgoQVaYqou09jRpeRZRXbRq7affwWi5E7kCDNVginjPmGcFvkPskHpo
4zs9SVNe4EmxBK/A/GS9Mvjoz5OM02zA7+tPcd2Gx52HMlgRlhLtFjujqGQUeqw6
frieem/Nnj0u/W8c7MYEWyY78Dg2QBrTFBIePuFqMCH9xOZal9ouAwmlhf7SrzBR
rH6TykKwRq0jum05yx+WLk1a7Z09A2rh6Kp2MXbg4D8LXG3ChMUTNPTu/ZZJU7WS
lCcivx36+oHKxa6qYh4esh7d/fP75NTU9Znjn5gvrc5G7S/ZNlj4a9kb2mdL/2vs
66l1NBLZax930vxw9mK/nq1LwIrGwmvmb006CS1ET7U8e5E107rimMDaQbzNtM3I
PMwQ45KAPL3KwGc5BX32VA1FL9mIssrmgMmqnbeFXMUiPUOQlL6Lyj7DNDfd88gW
Ofuyt525AdwcdgdbqTP5URHxv1G8rTm16yuX4ltN9QPEZgLMpL2BGEeaPDICru1G
tR3hdWbQAVCLcG5PfJWk4hynjcd2/4R0Cj7oBC2RtmhH1st6Z3gApBn72UOB6s5E
pHaxM3Rai1gix4uSB2TJ/YK/aQ8jlyP4u24zM+mZ1ANnNLPZZGbMAT7yVl3JWHxp
umQx6V9OHyy8FslB/Hpu4SW8k5fEVEoKej78rciAGTLykAKzS2loaJ4n/nMFo3zo
ED0jVjWBfnbpz0+hk+jmQELbks+iAb43JXvakuf4Vmo7eJ8sX6MmViMfg8NrvxMo
lx+3oWAERW4E+BdPM0hPGGSCJYOKnTbHWcpOT8Gz59pt1trqEsYUxbRlTC+R2Ob0
CMw0/wwLzC6uuXMapqlFnVClC16U57ESWPTITnPazDqOi/UaBXuBBSrxHZ4dWq95
4SGeeT+/wYBOXFCEIqLWNfsvniXgCSREHugvTrvL/k5L8kQZf3OrZ2hgJOzi1HR3
6Je9LW85NfBMhviHLp9oldbXSA4LVpI6FUAfVZi60gWe26BXhJOTplGUWG6+0Fb2
5+Zm7QisYgXjnd12RmO3/zl0wLwFIjFeJ5s4patOwtgFhm5ky3f42hwcEARYtpMG
Rvlv81ywK8usg/0FyqB6Ksg5dRFBYFjqOes9xNsrwiboztv2AWTyapG2a0/iAC8P
GgrM8u0a6OEuPb/DCrtVu8iQNHkyJKfGqz+6KG9/T04XnJJoceemfk6K3uQ/58jY
tVwNTRatLrWt8/eAacmRw6UY90u7/Qnu8DLlydOjQZxQQQjLXkvb/PcmAlpKG8gz
R5KOtpaxfNSYdCDvVGHkqPHNIzllt6g60u5EVRk5a+uCTxlvtl0z5iIEFYZRHiNt
FSnJQhCPtN+0fxVbvUCeX8ib9Ratf7cetJ2au8pLJYj7VwV0mNUqk4V6x8VbUYZK
XWtvZCVFb84jFZ+Y7E96zqo5/lqqtcwhk1PaCRzrBuShjK7AjVwNEtulAxO6Py3a
hcjt3In1y6z9qAMxN9+Ewuv3T3JsOI91cHosPvn1tSK5E0HOhUtLAi1OL2iOHPe/
RhZ6LctjfxvuhlAJs50wb33nr/JcfFOrqOZfmu9YD64JxkrnWG/W8IyXN8KfV4sj
rWgYboIR4QuTbF9IN5TTFvuozdwuCEFyY20thsxgQJA5acgJrKDP8qT7LxEo02HB
WtE7uLOxTDQ53xUYalgirsB32wYOUONt5JJ0sOrz6eBCohzXKY++XyRUiEJLg37t
JtKjb3rgIAu4cqgDFuT7af4MnlF/IL8lKhw6JeT3H0Sn9YPDInaya4ySNFE++XqS
JoeV19KOO3LRAK+Wec1yMDqNWrbu+VF2TW9Q2xYxD35Y54Y1+jJEsCyEcS/Si7WD
1lv4tETlo/ah3rnvwLjdLVbPqeDo10pD/XXIZyR1x2orFZ0s0kSEFTZnYvBFakbB
F0Xm5SMRQXhDuSY5Nls2+Yy4hrYLFvcxzY5YZewplRItYsshGEJSEX5/JcwZM7S0
IQuCu7iUMpPWf34QNMbv0TfW7KAg8o1dTdK+xsSEFfCSQzrf7m50OdTbpnRrqjvz
yNgYLAndQVC5BlLe0NlGT2GHeh38PijAWfWSIfSN5M9poksrvqCD38+yPRwj7R8m
ODn2ASGoZXe//Cl2db1cnc/DGDH1ZB8gIDNV+PPCaRjMAOqUMVprNYfpkVems7z1
kBJC/w/h4k86yDM/ZuCHZcNOJ93SDM7i0pJX8grXtQFG8uL2PcrxzQrAA0G/df8D
exoWFD9dEpqJ2o82e2N1qeEq9MHdV4kwXWdX1cSH55qgg9n7yJBnIV0zBIEbhrPK
tInEywM8BXKDyHa4TnwtWdJQ7inDv3guVPqgtTwgMhOxG7N8zxm3qxby4rkBNObR
td650O/gT2DqgmPVI4bRjWEayCy8GPITOtoToMigGPqKFAeHSLbdWfIrYd+YYRYY
9X9MKwv8lsKmcezsbHCbpkC8pmARRpdLK3F/9jec8nMSgg/Ursf9wKO4JpQiL4Gn
kLL1e1MRX0hMQD0m9XWCrnHY9iRoYovsO8hpmtWUgInVgY5m14WMSnstLEQrXf0H
06ZO1ixorAKw2jtXYNAEjvAYXkGHqawwGx5kV7VMflNVjt+qkEAOnWx2HF0SOvM5
YTRJL5bGWFYObwaKasFxx/av289evZjrabNGrOO+rIQZP2ETNXEqgcww2BoI37xR
Q6xKq924nddiSGxttEO+jiQk2l96iZvd8FEGR91f+pr2sG+iiaG8j48jqhG1M0Ly
hbcTu5+67y98rsf/mUSMOI9w3cM/PdoJpibaXiKgD2jgXtdRGzuuE7uAWFdROV3N
3Gkff+aQPRWCTjlir25/LHHCN6piCKG5GnRDbpn/SRNPF07UpfxrAc65wkcUjfIH
6LEXTh5m/NgH+OkPtrR8tLNm/nRkaEuEuPvGoqK/e7FHvlvr7t1UGdY9dfACxAB/
sfb/Whl9CMOo2sWjGtVzpJPdc0GbNIX28G+9KqATRghE4654S4+SGPyL+TYHynVz
lrPzfLyK26mDbn6bnnSjaVFcLZtUyyN/rjEr4cQBXubsIR2WPJDsLSCaA2znjQ+X
b/7BQrBMPZKwp7X+dN6drEokf2FK/GNQsCupZLZAa7luca51XtfNno4BzpbpbJXX
3VcZ8jl3rWiJd7VwFiuJuwLiUBi+iv4Y1Dqu1iwc2P9SmCpgwLlyi+cQkobmPz9X
BZ//Y30VmY/f89JqEk2lQ+t1D6w+nFs2Tr4qtZ+CSWW0bktQYfORyv1rVcZWwKH/
xV/qqdWd3WqSNBljF8nknuFQbEgNKXc8wYCVP0o3hqi+VDiwdn335AJn6/H8ajRO
XNjxJyllNvSR7VO/o96bUB/n9tlAXZGFLjkeg8pSKf8o6NxD8l81NCddS/wAzS6o
Lh56ovJOYxV8+MTR7p9s0PO3So6FpI4SJ5n9RFc9qJT91veW3smxy+LI9JUJe+kP
/rzJugcCUO3qlDxkE65ZkhSsXTOZ88LSoEHFGNoYX/829geJwwWoGhN0bTpBE67B
ZPL5M6IrzzI1f5Br7YgFelwo6sSHnCwXr/d8pAJO+J5LfpKseaUpN0kYpbUaegCF
8DEXVzVddrOuaSzi/GnCmaL1dGpxc9LXXkRBQR+EMmiXbzGnJLtLHWAeUwVKqt+/
eS+OfYcLePUhPBMRgZwjth250ZMMuOTgFm6rcwPtU6SiR1aBdwf6c6oaKMDic8nc
M9dCp05KCpRJJFUVzRr9+f4RTBPekLfQsyF1D3GEoD9q9S+RWt0nwESDhvFKFZV8
Ne6M4Xwx8msuV6CoyF1hXGD1+z2jM4k7NEBMROOq4s4F0lZiaiyXfqR8Qmouqj9B
OBPhbhifSXKwqT838WXiuAHLkSAHCyLSeer9fg79IBBsKSs1ErjCNH1lJvAhsxsY
fx9ZJuNJde4M85GOEBHQ4fx6106GuaY7XAlRP2z5y821LdJLX5GBKbmY9VLbijaT
5smScajIcTy/EAfXpJhrfDN4vTVVtIdrKHY2iuvEmOw2gMnSfFylYxL8stkovZK5
7jj359IbXkPT7xJU9s1rNxrD0NRBaRHRYgqGxWef3UmmvGci4yUXX3MTDvPizU78
b0kQnnRn6GXujIbfFgE08+8xbykXaAUuVG9X0jwSUSn2v/xAr/A88HQ77f2IiZG5
sYmNuJuXGrIhwHvq81utjIjE8bILoAGM0CA25aZVtSkUJRsJiJ2nerZhagm8y0tA
wScNobxtPOo9MdQ+RdqYkttsxL08b4Rd5s8utyVYyQDJltQlvK5llo+pdX/T7wJJ
i2gS8dfDsX9eOnRUNCoQMl4BAH0K68SxMqYElrJEHzPEYVXm1HcZjn2ZENylcTjB
B0Bg//Vl32Qz8evijieWCQGCJnrX+jgxjKx1+SliL6ocBSwGovqwtRI9APV2JKMO
G8wnagFp9MYUg6siNQYn2/mXE7QagByGIzHDWaSUkZyfHimZa4lpoO4prrs6CVXM
Buksg7qNpOY2Qnr7IBkBo7Q37Vwx1gpi7DUXRwZa/02k7y0gbLsuhxLWd+UVPbFi
M0DoguNpR9g6TRRjWMQ0tBfioVksaolADZhg4Oc6lstA4hueqsoENE1uwJRqAkMS
WBLC2NdSbJhDuMCgCn3GAX0EV67lYEd8vR5edWC/9z396sZyaLljtkOlQBPCK1KN
dNy+Szbh7Foz9BF7F7CMO1eLJ6V2HNOjkFeUQ2qOgKe5BOj1P4IKFeKVPv6DMiJs
Gk/EoN3mtqSev6uWgEjJdFZuxua+nDPSD3ycuFzIIpcbw9LTUeIoSbHnZXESowiX
06PTlXqwvQrhUyNPfCe/5m7kJQQ5yjSWkNZZgIsXkbLrz4Hm8JWP0k61blktGCbm
3R94KRzWD6/DG9Ku7aXcZhIxEJHax3tso1sE5tAplei7/1EwrBjAhLK9O7QWAoHF
CSDtCffOjmh5JV/fkYlT6szOQCmYZ3zNh+KLTSEn2yT92Fx/W/C4cWeuyD2i1Mvy
da8BXMYcMJ8x1MiGzfGIdxLkm+HlzkSoOqBS4BOQUkVLzJ1wDacTRUK6KLBXCguK
ftbePh8awOPXrcE7fMl3KZ+IVbxSFx7xEtCa6zDc7dNJUVcNkUljTi1n6YnXHXFz
ueYQSbhSJUSzSuqY7YzYI97N2/1QufeuUWpWq4dXNv4VTe0mrh/nP8yDviZHbdBm
jrvY8p03rWTRHKNv0Bm1b1Yjv9bI/eFj2VSACR33iFjswRLde7X16Y5kJQielmBG
VySm33miIaVZDb27w4qi2w/+uxT+TmubgWfGVVjsHjismaDWMSRLZvlixM0j54UV
88gaxnccLO8Xk0JU4Py6nGEhlPVFAK/wW1P6r6n9opKZRaOBvqEq53m5Zl9Y6QVZ
bL37FPSPY0Bo3UzvBskp8N59+v53TVoNPNtCB/9zE00WsJqJLneG8s3/TYtN2pha
ing/q5C1sa1HbgTHnB8SD5zzEt6CH0IHS74nurJOiiSkPrfY++fKVgw2usUw568r
hfcaJqZ12u0jO1M870UIMHqnKMNB3Ne61rC/SStdBSrNG0EP1Q82lC6scvAnGd1X
KeNyQPoFQ9e8ZhsZaFPV7NbWxOEkcNn0c/f5r05TpkHaLpBm6DyYv9lU0oEGWa1J
nuO+AIJPkyB6hWKGdWyimxiOu+UQwJTN8z6Z0oL05jcNO63NDMQC83Vn2oM6iFGZ
m1Fo80KXspx6DDFwSoYLF5Qcwk0Yim5ZT9Dn1BOcome5L5t4LW+eSQ3NZAwQhvwv
NsQIo5j1xJXD1bo/UHjwabw8oyqgFBextx5XSdpJ7anBRANYKnpWpdB7obGeNaH2
S9NLOpIJiGyrbTlSEmukbKHnyQgTLwF53A7Ap2lGi4QrzCbAYOkecaCCl5ocNKJY
8wxeXwHU1efjZszTCaAQFGTEgtnQP6langn9VzKkYE4xIh6XO+DAvHPcoycvNxyZ
ewFiliyWwFNUm2oPggTNYrUxXblEbgsFZW7evPrp3bIgR1sGw+pRwapRzP20ZSTI
z1uqOD1o2hQprMyDCUavnxgZYZevoPGxi4s1DkSS0wUEnAQCAKcEhr1uagiszEXz
LKmrUGiLIsbmwevNHAZJjFPVL1q6PKWhBf42KVQYcVYC6Trmak3zf4ZvwAJDOb7N
QzBtENOv+EF23Z0Y6dhZH77X8TnRGxBgDbHJFvwXIw6ya5OBp3cyFhq3uzEeOrj6
XlT27WEKC60XtpLDN+RWHjorTwayPWRgae69xCHgcjKF+txMUgQI6DoJHRivVFV/
lDYumKBvSzegFtzmBbf9fKB99OZyVcrM7WABj3aYa19xEOITQ3WMT9sp1wmoed9g
l80ZV1dSPGrHSayG+SmPPy74cMjf979B5nx0mV3YCg6A1FVGecOcoNdSgFZ0JlX4
fvnjNt1/d5jEIHyyYtmGh1PbNjX4tfeAcIRbtkQsGG6BzvnwLXrt89K76VqIMgyo
+We9JKM4D+4Y+lriEvSBrv5RAvNWCnajl+iiAMuuWOefg8Zmc5cTvBI1tLzOBt1E
/LYe85ySYp+vEWcpPDCVYMLUWVy2toNKVmtrHC1YI9D0IMYkefaAicLzDPjjQXzB
7ZADMpTtAjozXnMPKgPNBLMFo3/wsInoESbk4GfWZSycyjHZJte21jSyAE6BtitU
c6IDdui74crDRmm73u0nd7mKY6l1+tPL/FgqKvjAtU0c/KqfKpbidYMjUzCGbhyD
g4zLe8KhvPRnOxyr6T/DgVz8QsWT/wttCqy3wOf1Jfmf8XpQBXjkNjWVu7eIRMvr
dd9r4zpQFS/2mpcoRPmaTI7oG2P1OWtjidOkk+x2G8Wtp91kPjcP2NtbzBSgVohI
fn2DM5eKq6xG8/hmp/25eLmJCpcIOKRAKagdplONr7K1e6GK1n7TgRRqoKUC7uI/
35hOGiQg7k5pIBR+RuOKzNZPf/QV8PuC9Z9jCQnWam9MpmBc/1e4hy/xdulD6oEf
A2gDHlQWTIZmMgJ3sa7PSr/96rApaT91RoeQd4AxBrRVy0gDoJMRrWuetrX7W7dN
wBKqEb7/UqATkvV5Vru4XYvmcw1jDOP35OzeRkkjGhqEcU9tWzVNBjBelQA3ZCix
rf8NXIdswyw/ydAgciKYDPrh4ej7rQCDf0P8CNrWAaeszgHJ3mtt/goMk6KXl7pA
Wsl6P4jSqov1xMEA9UdAjWHOdf6CBp9xO3wtx2b9kKIoCVD3o0oDr9kFMV38qw0b
dLSYoMajfK6AWefJJYdmpSI+asWF5IwmcOZCgHC89W4CFO1ZHBuAdqMBLFF5RVdL
ea8sRt2CUXDb+itfEID8Mv4W3ckIbTwRMOBrxfckuPuaf3KEWnrUNLJLxPdFST1Y
AoZyjX8FOhuVo06G7RMSUuyQelr2QZpJ9NCULJemM7pgPSurlicRjHK/T3lskTwp
oBzcefbfESFkr8wwRNbmXOSOrHYBFZSIKRtHQXOyvWyNyV7FF33Sp/lMTMlY10KJ
FnoIhWXVnqDZufvocbWK+EAJx31ZgOSiHSVcEL7QJb15csIU/obS5y/nDda/Df/8
2TyscJL0I4QgS4by6erTs1YuSMxFx8ROFwBeZc3h1eWKlfDlnSQPOV0XwamMcMB8
HACN4pV9AeQi63NrGOwGnK/JejvyLVL0gG8b2zyvfRIUPQaQvOw9e1undjR5YAPM
dWYit3oqDjGDL7Yb37wavCmClH4UGfseHkyy+Rkcu5uTEfat5+TRlji+sCkA0Cgs
vOS1zBH1QhJETrQaTpHIkVV4p1By3D+4hT5dy1GK//vYeBeUYR3uI9RF3NWrbGnJ
WNwJOPjtX+wMGMsppn5LmaNHqKuCtwEJfrBQrEpve4twolZ/E+qyeL5462TTX1Xd
QTN+rCNhnoS5qwYb84vKRyIwGEJ5pKVUwVNwT8F/jP8ouQq/dRHl1QKiHzazQQ+V
l4u5CTAs7bGFmQx1PgSx05khMpVF/BZP/qivibOfvzyhghBsdIukxwvq23bNsP1O
rigKQ5GXxFl7mCAABrRM+UB9EAeIxGYFVoyeyoaQ/tzKL5/87udZALXKusKdrd05
XSoqVdZEC6keUi2GWxedzPzSYkxFqVSPRR2HHBf1MkunJoBF0rcCgHOlSFPhnd+P
9kT9kw/lNBgkSOmPhFAhsfiZyIMQbE+5iBGLFwqPIzoCrvtMNncWUus+gGAL6CAL
Gik3spKswMvvx/SCGi9RpOCiG0AYSryCQLQ4plRV6GBIyDYLkPqKzzw9rzrCvC1+
WFa2jqZXttinPKfLP2sIkw6YffX6mmcyKRcolUnv97AnjVMpRjNB98YsYWdSRSN9
3YqBFZ/OcV+X1g48pZA8J435hSJUaWOLtjOI/lYdGepPDvGT0p9kKYiD6WEYRCqf
yFvo0fBpynQhEESl6OWsE2SBIg65h50oeNRi3hTHRlcN10c+RwvpJyhYIqgFfGVE
2yXQjMDlPLIS7HmR/lms9HmergWZ0uq7DR5dJkJxUm6sfS1cU6B7o12zJmMKxUiK
9DGTn8gDQcshz7MV9/JjPIxqnhZUAwpGqPgCcgT+PB7uEHZ2mDyaZsBnwb7GcXrF
zSfX5z4RiFDRUbYGDygXDlc4VJY0C+An9CuIzguQXSCd22rmWIG/3vnmnXRyqiR2
zcarPz4HoKBQ1PvJ9lWBrDz0nLY3+WT/XN1paBp1H8yAKZHOErfpAgsKWq/1oiev
Ke9Yh3VPTrLCGe+ub/N5SrUxtSfg2Q+5MGRcPY93MB0QdkqJyoDtc/sL3znq7uaT
/KasjbazSQXstvYXEc1gPLDICJuM4U1S13ZUaWoTAdkpnEcEm2YeG7cMyrwopigp
XqVVmCQ3Gds+4LGMIjiFbrxbd4LI+ZuYUZm+fDSc21x1PYUBcxPwMXTuKa3E28O4
WMEGzRlQb6rnibtpQS0u7oS1K4C1ssqB+YqnToJi0tslpj00Y5AyRXiTsHsIhVk1
kp6ja8yZP1SoV8GgBh6IqDwvIzeS3AFQEjki4GbYw3Rnb5EPmobUMQ/AQVN0bEvW
1hqNvyM1mab6TU9JTMTRBFG7011lWzjDAra2ZUmV0J1UGNELSCmCPoHnrzUHcNpB
MfV9nC5t0XXwtnItmoDBlhm3+amqtrEVFbVKf75mFNKLbFybosj2msJxyNvxoDRr
vRvCK2RoaBxusrFS13bzkLBMD3uzdsxmm9Lrcvr2hNDec8CnA1bmkrYMRLaWDrfh
bQZTVqH73/q7wWp6gaBPpC1heQ3WmlB9zW710cGWy9S5qh6z7iGxDAf2bvW6K6uc
hngjSm+TGTp+wJQQyqfxFM7nifjQ19b7qwj16SDtAGUWPlL8qRdN37lvr2niEOJC
TmFCwcE521mp5sE03NqBBS3yRSlsPx3Ml56mFMumhIRRj3GW6ry4FhIfyVwe5V5C
KkeLnmqAla9zHoSa1ZXUTtt2KOOK9MSqGKqHYbTMNxpjhM9i82wLLbv4ZBa3U3ik
teTPB2gQCwd7MsrT07c+rAPQltZFBm1NC1W2t0CNyieQXxfMT49k/E7iQQym79Nr
j/vYRLuNcL0wXWd1U0o+Nj8YE6F9pos5xrc8viyPzrQ8gHyF1NJTlFFEaqml/wLq
381HKaJnvmtbGosvK7Dn3mxax4PbE7hT6nieCvO6B0Y0yOZmPSvu09LyuE+p2YU3
1fHQ7e+Rk3koEAbASgs6coHnozI6vgKQ0c+2ygxUdcEPnwk9+kaehzo53+9CvU0e
7XJD1oMwOE0YNMtCJt7BUFomuM6Ipsbat5EoLLZnsLDnGrzPpsgIAwMPIgZDj57/
dffgjYKnls9Gq9flJFQRnmxE1fFq9KxFoeW++0225b4mPwwZNDoTG8I4qzG3Z4zr
zGJ/WsJo78/u0qvq1/tdgA8TIiZOsPmpDcwgjDm8wLEnHnhH/n+4mKb+YsUg+CrO
c6o25gKENKDqbJ7/QJ5eTSZIinKkIVfFqkzp67s5WtcJfqBy9/jzLcPiZyxLTg2P
VY0nsc9S5SL9I2JB99een5UCykjt6a7UxvIL+MrXGl0g8oMXOM6w3SrhkYFVLVhj
oG2RGnxIjJxpym88l6O2GPZaEum3GTUncxZcjNOTdPMmQlYyuiZRnrEkxS1VrJI6
VacuoJg5EZ2FjzNsZLit0UX8fxfA7F0xvAgXpKYugPQSoSmg6Njg/yGTLf5o4UTM
eN/Vqrhg1wwZt9urEUqavHkLSkvI4B3+YiZatPK+aP2APHftoAK3PBNqe10eU+ll
xrkMIvDlDnbRlwKPp3HBXJabLhELxVe0QJ79LdEE7BW8zTRmRbp5Anc8HAMIRtKe
FdLC+Neo4HCxaaNX0OaEBL3cRPCC8nkNLZXYiv+vffWnj3hbyCAXXicCXh5xNVP9
UjQbxf3jP31c2gVQDpVn/firJp/u0Y8Ce9hp6ipoH+N7AjZl5qfut7dibmzq7o6x
cJTDwVldwgWRwKHfLGA2A5ORTManOA+/TY0o7qbIP8ZpB8qFajfX/wI7Mzw84kFR
ITtmI5iQsUW1eB6GZtcu8C/++/NGBDJgCXiy9A0HkuqnyXrK3TgSu5DF9HY5hZ4m
U0YYBviisiNBLLaJTFGjrchegS0p2RnMbTve4UB1236w/EfXxwavUEpKkMFSh3na
E3Jyu1JM+1B8ip32oGlF5QzfgTQ0BVoUC8ysMr4kNyR76hwiXJa9xXc2Gv2wYgBY
ysQztWbvEocuSElaIXqgBab6B+PWAtZm4nLrGRts5j4lSq7p4Kk3OXctVXzrh2yE
KRHNAQ8YhA3vlpJXx6KikvCc/fatHK1wtoZPYlk1JPS+QpbjpM2d/zmuDCAUbW3q
9p6vsZQuQjXkTDOaGH6E2JfBvzesH/yKKEsyJBD1ZEx5sts2/KUHa1f49CqOmHSY
CLwngNPzKYNXPZzdgC48lT8zqCmFs2KH2pyHo9zss+dQAxr/UyQtRxrr8i8mMcs/
NpeLUgwfQbTAzFcCDjYCjPnd/BLDJwPp0/2C69iMDvpnDwPGl2CmUXG2x2MDP3Fx
duRkzAShmNpRsV9xgOvZUw2jAXv3AJ96l8ZzUQf16gMBPT5a+gY3xS8H5H5inzv0
KQA1Vorr2kxOksUSaZdVt1HqScXxHFqi9yAC1QGsWWnMBRabKRA9MQKRQgnarSx/
yniZX+MP5SaY0RhMHtqPP4hZwN0SgFqvNUdF5oD20VGO/t3WrKhwwzvx9a5K8COD
pvlhHFLa+AqwiJdudSbwOSMiSiIz3j/T2auTCSXlmpJcR+GW0kNsHgB+2k3qmvY9
eGgDiukszI6AtbqbGvrv/aNt1Qn4c4GklWIsI4zZqLZXBVqnj24edQgJjFjSbB+I
E3+fmkXhT3pGzIqAxGXbu8pvZaa1HzuXGXA8cTzOs6js5Lr9pPPrDcL2Uah6zaTt
7+wEhcYxPixoTD4yP0bPSKRq5Cp0FxDUeDBjcSYC77ecBzYlQD1ssD4o2Xw0chya
ghE2uxKcs/N9P3pa7vzGHj0RbU7+aHSm84rtWxp6E1KpmgWVd/m8LwgUA2FAZ9QH
xfIYnRHGvVjcoEPz7zrHYPCPQmFychqqLQZMyfYX6np2Sv2WByVDESMtl+5pzpS0
kbPyXHn/eyl/XfazvONQ3ZJGQdAQK+fY5SMb2T3hxs6/BgMm8oAz3JXxFHYhoeQ+
SjEXvK+KhIWTzqBHgvJcZkjkGUvXV54kl2kBRau5qwZNINR1JQ/sEPBAvcSGcjX0
VluD7z1FgXmc+ZjAdoyMAoogryD8148EHuI1PTRhWu7X7Uec1WTaoe1Ufz5gDNXS
cUsaY4IU+N5yBKTG+qfVcqtF2bfzwjf4vLhAU1FbHIvNDY2/YGl3gkDzcgCClqfK
SLvKuvy7mp94rFyTXy+17dV2yiJZyoXXDdRI+gWUMOTjo/AYUvwkNrNNqHCSqRq0
v4VEbTquWXjfFfgQTKqjTnudaiUhuAxA44aKWFMwZab9pH9SML8Bj4SkyJobJ9kR
6+/vR2ebNySCLr+aEe/WpA/fYxoJvCN7TBQH0VEekgjf7eJ493LXRcrjjNJFEDHA
8bh27D1vcq1acoqtolMhNT1KlM07Hp0T1kaupmfskKfFiO/30vTVYx65t1vxYdsu
c/5H4Y2voiQFGztMwfYfQ1T/LTrvifPJbZRbWbqE8SAv6SdgYyuzotb9KZqNNkS6
FSCu3zlzUA8PiW2ubZUL0sOzY0vpyp5+9f78mQ486VrpS9R3WiAJtUHjdmHbLh1f
53fO1+N0mc4uX9UTtoLLUkLogYP+ZCxZuYxru3pZbGFUFRrrPDqCYOfMAK0OHduo
NB31yIVDoiIZCVhKzboJURuqIburx3TITAvnaM8g0pSLSYQ1ES9Cv5NI7EpnmnGH
cUl9bRR7oR7AXp/hhJhDMktERnrxsAJsg5LWm+2YZ74TIv7YbeJPuIicwebavkoS
kpzn1fGbXJ0GaI9Jf+2PfczARWw4Q7VM26PER9aD+zpz8Gb704RwBpp3cWBYh8t4
lXNxVbHA9T+B0TvA2h3p2yEMK21amTkI3GQ2/sNXqFHr1O/jpBwMUjVtsUcHsLu7
jqb4N+pDDuFseNtz4V97O77k72LyJMPDlD0i7Xlt+ShvJBJpQq/j19Lk7Ui5p0Bd
PEjjdLRVA+l1KXownowRXJUpMdK02vtSdfN4lHN7/CyVCP6vK3w4SCNyBOS63WDB
l193JsfUQRhZOckOxjumcTHkl6yIrLvtsteH4kS7g0zJX9kX2AVLGZS7Uk9dJohK
qFeJCIRnBr8lRsJyrXQ7WFCY3wgYOa3j2YLGKb1eU2ZP9nsD1FBi+9BkIZ1KYMTI
6RzfqqpTBzYElQPuICzBMEt6jyguEbqMsvAP7uHYjkqUvuhQMdPej9QRhobAoIsR
sITYgbjwIwMImtC1X3OY53riqU1pDcq4F4BCiho7aZS5VWsohaWgearhRNJ2VRO7
pr5n+PTrqG3lyrv5psQdwFhmvoiO1n/f8qnG6abaZ/a1x/Y8M4B/2X0h8qA9DsF+
iePqXbk+daTQMP7ScVuiEI14PDMMcTIgn6BAdAko/o/a9QbKQDYqi2qFtRgWT/v+
uAVv6HWVe0E4midFy9JuxTK4ULNf3HbB/8NeC//zVRQ55g4hM6TbxHGYG59D4xWE
aSuP9E8FGpPpvECWHKxsbavPWw4GlABwuEkw1kA+SBIY7t3slDmdSRRCURV3NhQN
8agaw1Vc+P0y9CfL5Yy5A8/7ZhwPm61WcoSHuuQwtmumTFKZxISYfRQ5FGRnbnsR
3AIzOmNLimI4xx5SWJHqOUHD1BRLyGvhzXU6WGuCXthB4nV4ZFWEjaE3BrlXAyYD
JjPEAYwSUFV7Czsdm/+q5qUbFsGqArFWoW1OHcY6HtwenpoxSJylHcxdblgo9yez
1XreSybtAuRfEi4TQ2KRJklpyBCv4dqDkkpJSPK6jWV45ad9ldlNLAio8/xP3QZ8
R7A1k08a5J+s9G3FfglvHcbSjVf+LL+sokOMEoulPXNuk8xkg2+7mikHxji2zYfH
7I7j4p4fA2ID0+gTsfNtgo2Jan3JmqJXDWBhvTn12nkH6XhRreRlCVZQ7UpdmXl3
Vnf2XVG09JOCW8K+eqLrgMBbIgCS2gUm3ehg5h3yo2sG7nvwgE6eq6/lvRWF2ZXO
OTdqwheMCdpU3vPgIauC9yM83rowjF2QlQb6ti4eBmAmsu+rNpS+silu/k7z0CW6
sYEE55V80yuDnF+d1YCn/G8K6UaiyQ2S9I9NvZQjUUhwbZkimnGfkhtblLSASIQb
RRiA6X9NCyTrUpHq/2fQVSr86zTxBC5iCrta19g8m4mhfTafCzBYh5SG7iuC9265
1cM7plXLGMRskcj+cdZgiH5VT32jxLXXFhJYrvd35LBTvzN1LjZSTG1oeMutsdf/
3lB2sBrC1FwuMbX7hZKEK/vEaaEBplKxjd89o488ts9Sq9QsqEH6bTiCG/Q6MkDB
Y8+xBhSuKeEo6VqZdDZsudP70+Qa86i490r+ZTv407CnrKyf3sfq2I7ZRd8A6EzF
oHCGvMEQk5WwwZ0liYz/DLvOg/DnY87TxIkdNZ2X4IE7h2K6IRAxHJGXYk0BEVvi
MNETM1ztiMiFnR+jFBsVoXv7J/fLnSMPQiq+y/DACVIuOgSd29v4JQ87hYvZzFG1
qSAb5tP722mDatVkiLg53/dOKqldRkHAvQzXqGZa2TZBXL11rjj7oFqKFgj8T7YL
SJ79Nj6iuDkGBlL96bvYwOpnBrLN07r7L4BXI1JejnkAji//HfzPEB4AKi2oyYs8
6cCGoUTKkJ+0DfqY5uU5lar8cwMqcLpMSCGkBGXGYF+v1SyMPzQtKP8G/ePzCCV6
RVFPnrbPjhcI5QdKDIHLpNInFooKHrDoHiQycqFMLeSKkJBXdHew8KgYkTl8L/en
+i0vojvKRnqBdghytX4Nuj0b4qYJ89/TMSLHhuWBSEVXuoT55H9zTDLekcrTnOjl
uJgaOukwmTm1ySM4HNTeBeJHCa6up15F4avjJ9PUD4QkyucHROdObKVqfTOIgovo
P8Dn9JwutWSpZSUL+/MrAiVnxbO9BPq4kUWEyJwuDJDW2h7oqWSfIF47cTEKf4CH
F6vNUcmGqWED/vF8vhoJIi+feFPaQ6Tl5Of+7wc41BhPLxQHdEVuHsdYX3aaS2nT
I291vQJm08Vns3U5da/y+zMw9h2VIHEqBtJjY3H9SWywkan6XPQGGYRammNT37Ac
ScErk4YQexuP+oW+xeenwKJ1TGD6bxqTSZRBIWbVZb1c01ieUZ/oKSWHN7yj8gJY
3ibO5uHUqzhIOzZeCuw+HKKtsJrEZyJMQPGnb77ubgtGj/UTPgZ61NwNNztS9TfG
h7iFu1tjwJnVwmOxd8UPmgvx6TqgaGU4iV+er0kkQaBGMAApIiN54aLU3yyjkyNk
oy2WXSNWGrKPQtBWeQVCawZc4akzUDivsrMjtLOqx9LB/XT+47DoPeFGwsDJsX4a
7ASYVUuaKJ8P0MnbVz9GvyYOuYEFHfiOmAt0fnRk1MeuwmwoN9jOSbUoQTCNU6s6
34f5l7WPDR+ywnSfEKe8275yWyajMhvzTux1H5L+NUEuwHRbD5u7k/pAFrq09jAu
pI/7GS5hD8g94fuzzr+VNBxDcSduUYV7UFTSzx3kEX2XPMEvnQ0kEqxGqgeShZv7
clYgmkwW77mCMwrcapVWs/GjlMn2LzjPqmRmVC0/xKBi0srsIOKHh8nLPVH+2nfg
Sl+YyM5PYF6SRDN1SUwHzq9wxZP3URpPHuq7hHY6UdPD90yjDM32wdkBS9Mp9YsD
cy7on73kWTm9uqhjZ3PIMByhm0n9l7X1S7p/EMvOipx4LuG1PYGjj3TBMS885SHt
RSvJgYdPgmm/8g/DfyMUyC3fuPLLwwCuduoKpvPd06T16rhPOOLAY6lp7eU5r9r5
njydpMmI1LWQAf9pHu0GG7Wcz5nwfcEH/DQXOxZv8nsUPulKtc84QvuISpP8tXSD
OknLMph3t1ohshpzSGCdnaKKJR/qF717mbBO76zZy2vpegn6X6TFuQf62lIkMwxg
w7bATzg5IKlhBN/VT9PpawCd7oZU7mb3k7w6LxkP8o/axm95F4drRHFgy/QcDPm9
lBd8/nvOmzTbK7Rymn5Q+OVC4V92XaAz68r66of//oaRCzMXaTHp6tPn9OUbyeoq
/GV597VnZdUTfwFtQ42e+TRJzR/p3h+Jb9ikKOa8GnWFgCm4+6z4YC+Auy+7Tlee
QVBBjdD4stbSYtK5jWqJFKwxPqx1PmAiTY+z8lDSR+ny2TGmreKgrMiPeZxje/T2
OKzqLPNabHpflPWnnneG5PU66VGkQGxnO3t6mzGzB4kULWUcdq2vtxwHyRnh/fwI
SInUx56PYRSyYqffeLazeyBSU0rCg5XCYsWIFC4MiaEsQ8mIxR0uV1PlDBxBfyNx
hjJpgfTCULnMU/jtugjg795LNA1dPzR8+tpSUME/w6uuf4leb2X7R/Qh7YneVlNl
mL8F+M7WoL/v9tue7/bXKnYYvYYiRcrxW9qo26WsjaoUaKfhl3RF7slb/Ny32ibX
vjBmgvvW9LR1qvLMW0ictORjpwgm9uvWuvratG8a1hiBwJClPifLdfbILjnh07SN
ycleR6AEHO+qX8If30u7OMuFKnofBS3eo6oSubFEhOQg15Zxm8Ti6kq+UB3ffeYR
z6+7x26awge/1XPgjD2DXnClerQRypEGku4uBXuXVewsh0vOKPayX7rWq2jx5AoD
nAcW8xczqxLnIl7u9ZdntwMirf6Z3pgkC2ylHZjoI6T02IIVuLijBH0+9H58fLZ9
C6/yoRMlR9obPRyFSwLO8AhqMKF5xegU/HR3TP5QYJBylDw48AVUN3jUKIzXyhmS
KDHtgbdr6onQR7gGWSJW2rh+YIBXDloM7u0xqigub0R96DZ7CYf6TMVIRFDA7vZv
uHoV33uTS7YpSSjge99hxVjsQT2sZVHrBQbkUv4fTaBH6jwMXGICePbyFl8cY4lP
Qrs99d6YY2eSWtK0FyIibQEJ1xNoulG6CqAQsPencOJvJak5sc9gbqzcb+TeRubk
xA8KRReSKAgbTU6BNQ85b/j4GRUxRLQFbTsKN7C8gzjUK8Rg0H7ZGbOCWoQd3mb1
rBAYditaOrvi+vuwdZh0Ccrw6HTiQj/NHTkkHriIdfXNl5oahH8J9dA2VC4RHp4Z
N+H9mQwxpTHPo49VFEPHiUoeeFDCKaEPVTkN537fER3nCq1yME5xhJGZ010M0sOo
6HOvBS3E3LwnSTkZ+j8wfoKMfvXO+rBfc63dbk/X094uBeEPBL/eQZjbr75GGVgy
jjFg19qBAkKkIwhE3rMxakrsJ35545enM3c4nhqeq2wiD2vDOwVw6qqwx6ppXc3F
oSvzeUdbyTJt212LvnUhjDTt2Nmf1vs4qCyURjqkS1//Sl6SIZOFJXGAOEZlFkVR
TBvpGTYLkl+Ldxbm08O/SbJ5So8I5g9n/SdIef95nicAnZ9Tc7lwUgRpMwuAZiZo
zziZ+SgBfChrXOXnY2+nhi2aH6ro/aF9+JhI2OdnBx2qxpXTCuZ04j+WJTbc1lRn
6tuSiNYhqDSoryCoT2AGcE8YXMXl7EMS0Lg/onbNu6IU7W/lH2w2PA9LwG/Ozc4z
4do0DHN7zDc13KKnzD4kbdYQsXYc0rJVKH9XvrilayFKYHneud9esc08xEA4kYq3
kxrmoRbtswYujPMRZwV1QcKlSvM4eiGP/RF7QRGE2DY8BrmW2apwctvRdn9ICAC8
V6gpDa2hS3yTrvMS4papgtLviH2JlT7aXvNAV0JnQ2k4Lel4Ez21FdVYuuF44r+5
0RSiJlYrSuCPFxdOcpMDCJLU9EPGiWUFxMDbSHBI18CA9lWp91s0cxIFVyQZxb5t
vsx+WV7CcENaqyPpK33Kfu88bBZdVahA1Lo5SUmvSbBGNyH+h/D3ucLCXl9jpSTj
ub1iI5x9AyWTFxC5vlYlYmMjpzl32bMR8JAh18dHVETfbIek+i+wclmMonc9Ew34
hNkLKoScnQsGxMWmjaZ2Qv/YGhzhxt7RW4M1nS6hAaF+rULRJIoK/uE8IeAOAuzb
LZWf/rV6U8mZ+nf3MIWWh4bubv0NwcHlTGCRZGWAko4xce9mAO6HCmHjxcGpB5yu
VUZ7QmZ/v1sMDlFubLrbUEj+VVqWJZ+JRTGkvk0ait++nh4aexRvBT+BpXmObil6
Nwpmg2YIV2mEkns89ZGrH2zLJ7VNyc//0qUX4VSPeJKqa5pRYvJIPW40me4Xe/zu
3wBLr/hSGWKaWqaeUcx1kqMVRO2p93BWh9LFicr28HZugpKgiS0BS4PPhIPnjW4O
vxPmI4JhuTRZWYcj6v2IT6EV2cdpKr1w/W9EO0+lCKvxkoYkXLAO8PoQ63v0HSEp
N1snVENCrY8r4JMO4fv1RvEoRhW6gBFQR4AHmQzjy6jPdr3aadvkljSQV5h6b0xH
iHgPovMfzLuaaiEx5iBQ8Of2f8UrcVGgXdlqO7nM6QmHjtMQ3E5Cq5zJJ2/BM2S9
E4xLeGvL9gwzvpMkYQtmEilU9cCPzeQDkXHO94HaZu3B1EThuJ5UfL6WzsvA5cqh
sqe0Ac+xdop4sC4LIAJt04Q1g32nf0UgbTEwNxJjqDVR/zsvli03J22jx5K+nfa3
eCAi+C2tb6hvAbqxVbYgE9rnwBeTqhdpWw2tLWzaS5SpWkmGjn6rVGjub4LbHOH9
Z1nmsTFg8zNzRJCOUd+scvUXTMyZnajquTI3h+0ErSfnVpbYZ+ygGkpx5rpA70Y0
zJGa3jvuccehVDIIJf0K25Ql4UxmBrn2N0dEFIpSNTSMePjMD9kNTbwbMgZ9PN6W
oE3tPbGFWwWMCtvzhPWUh9exucbZJz+ZXSWUXXKu8DZeXzcBogDJzq/eL3Zlx9MH
ngoXnggPb9IOseQoVgaVws7coIa4BdIURy6AFYZVrCpv1boAZ/aDCZmQO4Hloc7w
QGICpOjofJZJbsqNq3ZKz0AUHWXQbFE/NVlRFlMPRuCYrPXR5VUrS/hCtiGyHF05
Gs8egNegtqJUhVumQ3PwbLskTZprwWkHFPKAI91umvDn20oeoKiLCdzNnGjo/c5o
v+NYzTOT4KjktiVp0TBWxB1hHklKBaILTssAErSNkP7uOuQdYzRLJXkmtROETQ9h
GDuTlPtMz5MosAVMseyBgJyHOr2wy0/wj6gv8pVfgkiRXVuRCCRzGKDqL6xFNHi4
c7xgD5zCvJjCsVnDHXuJs2YD27c+1efYpVnyPMG4PuDjcqR8ktdxja1tv5Yn+Vei
ZJ9yprAiilX15p4Jb4m9XS7wxfo9tTTRSsMir0nK2YFUBmCZf1Cxv3a+BWiPuHxU
ORJEBODSDU0lNrERBAHD6DU7TssfmnJe+1cqcXVt1dvvW9CZTfLuoEsZoS3uDQdQ
szKfZgj58pkP2GO/FFcpI1fIh5iOyqXsHVCZJ4HvDDJRayPVUMtFSWT8cWMdwfgo
o414OzZliVQS/2gQkdO+ucONQzbAgraNtItPeJf6sRBoMZDtmw2fyfWwBJgSWZgu
AxXGOTzJeTdFERYuFDUjd3vJCnVv5rmmTzJnWS2/7MkmVZElm4wmT0JlxiNkz4n+
5WqWd5SKM9qicv91dlUoxz1YcVOBEbihTV/41SMKIWP9FYuop8um4oleiBgkclWO
PrYE5nrpLa8LyajHotAeRbpQB9ea9HznTO1lkQGUcn+IdkCQaaepArvlNgJftGq3
oTrhKMJEYFwCxvu4xxupygCUwtP6LDgfW2NCwl2OnSAxgh6Ky7x/YybeYOPkfRr2
+TiPTjxCWNji5K5abCZdEkAJEnLiOsro3IPtfiMSBLGGkXa6ZqE9Z3EIdDG4xS1L
TUVmsEc7Q1cyON61wSp5ILAdhAAwoVcmSZDThxyxgdXI7dATRfGxq6PDpnoyAl4n
u/uDlkun76IShj50DaCPsHJUFJGXW3KgIcx187BVt2ZGi3DMcSxPugNwSF+x3uM6
kcrv3vruJyh9o9XMKYH85aOz7OwSrRrHC3Pyt35giaoqd2MJkqQykE0bcKk7Hymt
gXJQeYnAY/9zxfoCdmIhCy35VTNA3IUMCp7gj93NkpJ+Vf6I2AWnp/2hDPKWqaLv
ObFZCkWyjaVEXr7ryCTkDHqU2t+J5tflYBPXJZRTwOnETSYmMSdZF005KPyBHNaj
Tn8F+3l4DugfqHm5gw3VwzasKwAm8FoxrEyZvoMSVG5GiTcP23b7A1dwdIMZqLCb
K5WYnGq/jTob2nIKEI9bGymoQvgfbeBQiwHiv73bydeXVVqA5opWBbd30ofyVSGd
crQSk9imrn/KkjbkB79HM5ifQullIfJkqa22O+VxTpX5VhAGt5cdkl69U5mXF+0R
t413VLziPOyq4Cb2YTyptKiIhrFnllL1gOtdDLulmysXXDlYsjpUPTVXeR/hLvQS
foznk4g4du6vC9HQxSGzailPzQA8O3misjdPbQyyYAAo8dhdrY/i99GfOXIy5IUX
crHgprsXFG1+mH8aRbZLqGZ3o0K8H+zPG3noVNEAp0wWCnvXif7nkLPxT1hA0KxC
Ay3tVSXLYgFw96IlNBM388zRcrKhjC/eIavyyPHAdUFzNWqFNdmSCxxjiEEZ9JGR
WA2hAKodOnhXChvwkiszwk2KbbsGgnsSePAsD4Wc3I+2BWuUsI5K8/htDmfRzdXP
8BdEKdDTwVRVo89cmc9gx+JH6S5+yi5MYxwMHzuhdF/FearxWFpvK5zlM6qz0LPQ
rz52ex8P0HvcRaG0tubNjX9GdYHjX34RIbxWcTnXN7yW0fIixhMFEYAeCuFLoH47
wuzARE8/tQ5NYsSanpNEa2mnOcg+UAm65DUNEK4lYF5RKjSzuthM/WAkfMz6HYxt
9nSB0g/5sVvV4ndyKlhkuWF5Wbo6dwwg30B5O/b6iagdLSoZreOqtb9OcfU9Gokv
L2mt/dzURje5DRrewx8hX8mf//6k3vVv7qG98CU19bBTcrSdjDmhT+JPTPSrjwAu
OGYbI0wd9tyxqAmsLi7GojWl2EjXKCpP2e90OtDfX5dSD9JBgUN6OfhHehQdXYht
qunHNRZjiZUe3UovefqSoxZ7Nh1puYRaz54TXQqFnPgPECUxfReStZo4K2jrCdNi
NW3JST+3LJ0pFrmRVGOHIpgTFAK5VqVuWKjDOdOEdsDdIeIesZsjTYgoKtimykLZ
lDZg4jvNy9iQUGpeC7BBS8HU1grCeRnapsofYTafDNd+qidZ2WeyiuzkEHupAH1g
4E0EoTqZD7SCAm8kjjgN2PtLV2h+RYj8j8duSRAIm7kjHOrBPHu9RcqFo7+jUfBL
fvaSzlb9p4GkhyYfNyl86sDhto1LQc7Sx9VU1R8kTqy2Rtuk8Kv05WxpCrHB5ooq
b7+uZq1cofd6LpeehUmGA5AfhaHMTZLAwTq4ibz2YfWz1VihdbkoeAuW0ORrMxT3
TbAe6NT/sBjUQerOOB7gUJujS4lHYHHyHoCR71dQl7jEdf8lKJE9W8N46twuC3aR
w5H1WhbepRk4m+wNPYgDqqgUT8ievDLxijfNMJLfl5wfMrDhKvfyta+3eZ4RI5Zo
TBoHmIIe0F9mY53p1P3hG7nHm4vMHsHDxhodTejjZ6Ky0fOyou2f3ubCcnHEq+vM
dmEerN+vkoY4YHVdEtc+obT9WKUMjTLZRsDJSQ1m8g2M6fvK4PO3PIDwAR3uOiUQ
sojVaieYvy3IJZStNgreA0JLykE0p06VkeKeXqPAme5yKsHuZzDAe/aVabxZxEV9
Qo8WM7vr4sg4VJgQ5SXj6zhe1DRXMehD/LmHRGsJCzsC0eQEsetED1BFrk2L1T6T
PrTpB1Qaar3SFZfZHkpleaSVX+xsdFuA6GyIj+kZykazttqdzpK8koeuhSuEYLvR
+lqFwcmnKFbJEji7r4BBqhtjH7ntmcJ8Z90flq2SfIcBlX8Wk0eXnDoHj9KPH/Ol
FSUiMC8mTTyRvjKOMEQvI3hYaaSzYLMh4whEndo/vNfnR59pchV8ZUL1LIyDcniA
3UUg4f/MVt4V1dOl2a2voNb4/UC1nenOe7bSkqFfW22i5VC2fLvB3djWlVZhHpRg
Y5VxXpglk1jiPgypXRbkac4z28QLuUC8fn2g5eCptDihQcgO5uTLF8DhPhGBaCq6
MQ4ZLOPbWKlZeMkapHx/fMnx08fyhZgWr6GAY+NcJwOklYxhx25Yj68IV7IakMfD
3dSs3bPJjoaz3bySB64v4brHt3xhyBP6Q4UQsKnMwXL6zz2YXlmMVi8wBm39I3VQ
CWG9EcVAXtfTxdZc/UyeN3ydl9gWTSWle7Cwz+zJkaush52su6X1ew42OjpGpjvj
A48ZIwDYGEqUVs31SO4KtxG4HMSLgFxu6R36NhM4dIvOZyQM3djfDKql0bjgu/dz
S/YX5GSjg9Vtd5yqgfHy3Wm01FTgICAHEoPzVfGDYIYQbKGwAl3TZAE66UXubSIp
B+xNtVIfjar2B18hPR8wEVwVO2EEbbYArL11ppQFhHJrQeuRb2TC/S0bluUJDA+6
ZMdhScTD5e9J4wrWMVzDAmolOE12HKy1xu3xVThWrkDGR2eYOQy+XDuKXLHwSBs6
71wcW28fTiPIZdZysDeAEAdV1Q+iz99DaxKzmHZRW3Pmams9xVI4Wxh2OjwtpK8l
tESYURUOda58CJ+kKNSTVGHEIpkw02HVWSBrGjSKCNwLViKKtadMkUReC7fnWOY3
J5jvflhJ6QxxfLOr6Te6aFp0PqiSGtxUvwh3duwCTVSrijsiV6qBdIsB3wagYwNg
SbVbSH2EtZnGii21w17zHlleEmw4VyRuVmdfDfLDqqRAazC1fwrEfbF9PSGQqnNe
G58Au1VfQeznmVIRWj7BPEKdLtPx5EZ8rZSxhgBZNcl3nYNVkqa3TEE1djzEbkwP
abJOSK2n4xiIGWgGL1u67MqkDIpsVOBda0CZ0h+A1xUoMyKEQX1TxztfvXfccBC4
pLUaZjJi58zNWBUFJy9Q4Hf+P7cyH5+nx85aEu8/D+ZhY3k6e+fkCOkJ0aRpDb9n
9oPzN6ndLFQ1fWnu5qVXT6vKLrybQoHInYzmo6m1xNuRqx00EZOu7r6gnaFyRtUF
KeD71l78fi2VS0gsHANwnEuMP8Jr815xYGd1SDBWoOHfCPCEhhuKmlkjN8qTchGa
n+FWLwpvhTxyMTpbsu1zhAchYotVTwoeuLC69vjOtMpRI4125QUTciLw9ynCFvAy
czBuyVhIGQ31OqPQEmFBYqRYmS+Ly/ZupfFhyj2gTVnz5B3hbcPi+dELoTI7hjHj
SqR1WUCVXWCphEOLCuznsR6xCENghYyMzCXtft9EDlohWmPzrKDqlnQeiohFbsdM
Rpz8vX7lG3+zYiNXwurKlpJxb/28Q/BqMAQYZ7Fl/TbbDtigT45AeVnEmVmzPEXT
KF/uhx2W7lo+TJbxTXTuQe3CUjIGi7gHyLi/23R4nFDPdLanrPtQ1jPfc85CIp9+
B4D4T2hT5TQ10SmavF+qYAj8HvsDPmJ2ivSxtRcs68CSTeWB3RH23KISRdHYZJwo
WRW8bpxLXvQsIZXzHx0W+Z9D3LZ0o/3M5PXWBI7IHEUGe5m3h8Wux7VM1JQ0X5b7
ZL3tjUHjiY95OTkZpXIFl5ZgZ8p63+6miBG7NwTjyDRQ6tdpKn5lQmMf5APBgYCz
82KWWxHfaSOYQDD8kzmM+H6/6fMlFBWoNTvCSEYZTdukVqljOggijdI1ZYfJURW4
CMIewGVqE1IOrPWWyUGZz5lM2+pIqWVJcNzbhYEXMrNaFtq6zxaj40xhE3/Q/BAL
vs12Z0p695vt0u7MvVvFhACbMo4olyIUpfjgdms+oDHOHjl/hmcQtgbKkVIoqg99
UIFDJgWad6ogfivbdzKc+S6IA6eNmAgDwnxTbvkK/waf7MbA4Ffyp3M87tuxC09j
v0lNJi0BiE+tfpu5j7p0FFkNmDF8Wh7c/6byCZa06K5jUPrqOjdt75AC0nmDpOY0
fwzjRVRMkmXPpTt3+0imewx5Cft3o0GJ3VtSeLgFHUmFECyTi0s+WEIMVkDl2xOC
/LupWIaglu+91T8Ct/NW7ToTbUhfS9UIeCVvQXfXGaFPsTVq6XTq1YGhWhnSMnTl
IybRZOjmYWucmHqc18OzfJ7G1xXVpdHTF2qORzAUYggkCcZ6/tYu1k6Ml49jcd7A
6NiyRx7X/BjHzW+UgwjWAEvgr+hkLoBD7Jr/Kh9wCop221ngRnGklvV/JszZGNjK
E2vTIYH0WF4pFGoX6RU4YDlBtJplj/9GxMzX7IgId/5/zK2DRBfKxfcy1tpnYDgM
p5wpLsSHYv8Vfb/HqWl54xG0dckS38plO0GCseBgEdB339gCJXi45YlCt57DgEdI
8H7VUV1D/FNpH/Yaxa6QFRf2DH6a/zf5we0S38fUknuAief4bMtAJJ8eqRhJTsD4
dY1CH/36lVBOBa9JtY9QsvZ25bBK+cPn9rT+W4yiGMlIROiOtrgWnIKTGmJD3u2n
vltDctmlWfp2AF83/D/p/Wza/x2nLGg0BO1dExZuStDl8X/ooGYpvJapKkoP2V2I
Ug1F29aC3iPnQyXuR4RB3g/rpOgndbb0DDnBtNeCvwM0Z7RKdlmiU/BhBNO9pDCf
tNXl3BwkXOMhhuAgDiTCyRHc822lh2n+QjEblVKH8QA5spw5hzSzI3/7mpe929IH
4fEH/EIdS87B5PzCIfuK2BLdypdGCTGPjFOpiMO2PyuWuf/+JVqazDvNNQYnEuZ9
Do7mMXUztBitGXw82mnFlnN0CPqPxhw7SMSqf4uoretB/RACZzkt7xoglLm9taIO
7G9R4CeDt0QOSulZA1vTRDyND+rKzSv6Z8SZrPCFJK4xu9RceTVMN+bkVPvGozAN
2VrpJZoaUP6tIT4xjv4x1BP+JInMR6jK/OVjd09iM+UGYrWe11AQw0DHCMujhsQt
WFpToWjsv62ok8s2C1j+IquNagmdV0bahM3B/StN7JHtpeNkynKUF9ibwwJiM/kv
+SYjZ3iu9vYOnZG3OwIVVvlrEPYgOkbs3NFZc/Y9EuDIKZNNI+Ys5GnTarWd/SGL
7klDSVvGv7AaL9htXRQ+kJkwd7evnaNgAmiTTAgC1aGTSLTsY9sdSBsDimZ7p48n
sAy3c7GzWRHJ15l4qt1LO2JqF/O06r/zWMrArEgUn0wIA9Sc0woMGWIfZiM1EBTc
4aN1VLB8GIhfPWaPMhmvhmQcEbnnuIdk5+kEZ1wEKmH0VHGQUCLHPH7mChBNXjol
EcLggyfQATMuoHIP05tVZJiGNLTcX4NecrvoYZuEI1sC7DUcAYwXhUopAIuwTNyR
wKkgetzewTVVILLiZSwA2PZrdkmv9L8vbN7Dg5KTCbRFihtncUhn1cDlNoOSJrGJ
27HJkaG9y2O1JfyG7GzTLCxQTLO1DRCh/5EKVm3Ez/v85/o7R5c5PRbP0eZ/Mnr8
LMkKrMHRyyUE7MjtUS1pchctMTxuB7ecFjw4z31FWLKeNYm3GrIaqMb9Dn58qDQ3
La71p1KzEi3I6zXMhQrjAwJ/W23E1AtI4CVVguqTnL4HblK0joLxGuJ57dIJUOuN
TQ+wqrftwVcH8pPKwH3RiGEI8wkFtEYu3HCkT8C19q5EZciuQ8tFTx4/Kaa5FypD
bk2KOYDvzm+IArSbPUobJtrZx5i5HPvrCNM8oN8qilww9ymjg6xRw7DWuGE4pV4Q
Gzu8JF33qOyUhb+C/uQ5V5gz7bX7gr92YcIRhCBC9cqtpt7o57h7s+K51q5ticuG
IFNnsJgVzHtv+j1df/PWQN2Y8+A49/Xt3cZoChDi0EU08/acRlLuj8hFOr79dK/S
L0kzUm7mgC5hi6RnUvZU6i9wFOfzN81vwLZ/x+i2L/DIrzWOEeUWevlpoKY1dwRQ
NctSZfTtYPcoHTKyjER3vuh5vjKiymD7ReyEK6LQXdV48KaxWVMIaXdqxfIBiAhl
X0kk+PpQWodR6MmQmiCo+VxhVZOfcMkvOG9LU/S1tSL+ZlZ2pBOBlHih+OGWLJqD
FNMRochjO0LuiY3CXeYiaRhug/F9Tywqlx4rd/HrHeNKQpxjcHphqB/0QMx/Bdyo
Zh9+QHII2x8Jz70W0Zmp6jrSoqivxqEUDS3oBwD4FjUBP8JDsTJGd0hgl3G5JZxe
S5F7c3uAkDIcowE3QcCv83ljOxOvCRjhJVObaoe0QUYaGckcIdbh6lis9Qjwhpd6
8HWq741Tberf+J/OreTNl+AyoZNrQWju2ueHelQfbPGFlFI7ZdGVz1YHPQoAYnEE
c7yIhnbR4E3Vdeh5pkPLWEKVW/w3/7vDri+HBCbVarUiidzNXpYTv9dg7ZE7/DP1
vZct+ldUic8TrnbmEMePyTx2ZlRhyHt/P0Ui1lqx9RvP6/uyd3omZKu6W47+kVT5
SxPoYth7o2no4PKuezos3sF2wHLTyMEX/waGp48LcYy7QNM6MFzWOqzkW9iGKrFE
btrwYK7pOBNdoHpceYJe5lw952NZQ1RVs9xUfgltvddfRm6ZgdLMas4Ow3whjU2p
3Ou9GopRHbXjY488V+2xS3pbvxiAfZViX7168cPh2Uf77Go1gItspNaWIV2p1SdB
Y6noNFpPWhjs+WlQyCWHvS0UJb/bhLR6xY1WxQCjdL8GCI4KxkuN8mVplkOeUZxk
NcavXR1nzeeueBz5sn4AVlWLIvFVhaoefS60vyyCQ2dSajSJfU9JFLK/ELzm2tkl
AF6WPZMXTWMPvi9ZnaGrp3JP5zvteJX+Qn1nTgO/xJ8NT/s3UorvUBEJJMkKT0O9
WsR1IkrzD/7FyZAsOH13VhfLl+i8VV4nZWg3nq3gVdnuG2MVuKoUvBqqflrHRqkA
Uw30mulxJMk3p7WAy+kb2/1MZlvWruT+bH6f/8dKH9JuFvBvy/VNzzt3Q0fD7qzD
e80Y588pm4Lj3Jp2yZz3rKoppIoF01sjKbNzurDv+KZpa5EX6Noc9+zbv1lYEDnG
7wJZtltRrUGbNiVLnEthomlkScu+wh6KQ6im33fCf97FyOLnpAUPq83Zla9it+u+
dXmaDOYGJVzNwwnk+4Q1iBGms/rfb384I2e3GWeS3uLg0UdPkVADlCLU2vkvY0Ye
lyZ5HkQlJanSs+EHh5l6/5TznjfnaMrPmY6PTr6hkLOthk4Ynp66cgo5pFIg75WT
kjiFlEAYjEzVd+ji5JscMCqMAtKP7DXVx7FF9+4CynVbpRDa8nayZOdzhY1qX3fE
moIFhCxcPP7738DBhs1jCiiRRRX1sM7WIRGNtoSS8rZPmDHLzMFWMcFSNDf9aMCL
+1jrtAzAB290ENYMsZIs3uvxDDZoUD2K6EVEABFSBWJRl/kaIMwzzAW9xvHXmWC+
UeeBEUJWncDQyWRWl0xRP7DA7qLjiSaS5O70EzGfmL+j5Xs+LIWqwjXpe1Am9yHm
quItuO2ArMgURg1itkxhEFLJE7YNJjOtYkOh1bBJd+3TKa7JkuRivgXRxbPxjCW7
IsBeqHkOV/zobJV6SxN40IM4GO3ABVfOLzJmm7YNyy+lB4ROcvwLgpkM/qo4QlsU
1sAGXF019cVvgCk5Ky5U5SPQwJBdC7fjaP5y82QPUlbs9Uh4wK9bI3GD3Wcb8GOE
UBSMPEJq+Ff5UxOCH2CcR9NAq0g5C4KT5sozMOs5Ww1Nfe4wmUMkVtIcQPH/Mypt
7HStLRClwps+CBeiFAGCUC0iZCHUBhaEgG9tguDAsa8EpoJ+XwaUibdw/FuglqBo
7Ss3Mc3Y78bwrkP3q4RXXok19OV16RlEuenKuu4KFO/9BQxQg3Wm3Ic+kawUDxhm
jepw5IOFDEqKgqJn2vLlUbL8Sykrzvm3S7mlIPg17ZTjr5f1vqyD6RvUs+S4Z7a5
8XdvNaXMx5MC+Jk36hzvV2XW3tNYX0tUcaYwoN2SBJtQc8uCunOOUgWFvOTevWPQ
/LrHAmbf6eiVhrLg2ayje4xhOqI7zs0PNY2BEQO2I4vHyey5GFzhyyv+pAshSDRz
y7HhA+R9ShLi6NXvgMayO0OgWINMWTVpgjvnq6IQu8D/0I90fXb9s321K3L1PvoP
Emg79GN/+I1cWU++VvS2+v0durgDrOP/9BSRSAnxKrIAJextmUNG0v6bH3EiKg7O
GcJ1i7tZ9Ex2RjeOQa6GuvGcerTG1J5B9VGC+jlhmpqthWziKU+vBxIEwpbby7jl
2E/pTCtD3e3lQVGcDwAygzkfFrrPX7Vcg5NH4iiBo7hmhYwSDi1lGlk60DCCT5dO
rVjZK3ODZ94bdxmDJPx/wNeZzputpN9A6k2VWk9h169/3onhJ1FQDmbuCFfcU1VL
/k/58GNFO6zAf4ar/8oVurYz9LkotSyHtAKZs6TOPYq+rjde8Io1REVSk/oCE06f
BKm+fc7bPNBTfq9GyCboBegGtSO18Uc037Ee5VIVI+gX72StMcHOstsNdQKJv6t8
Rcg2BACRXu0jz3Dmh5t2v1+JN+LUA6tGP6S9N8QXN12iH2ul7RfTf3me9MCB4wlT
xPY1C2b2rhLSJzVfdoaoPfcon3HC2DKZCSND0acofZ3jUR1FoNkKEp63MNWMS9kk
7FdYtpF3IeEaHaGVE2+sgtYr4PK8z7K6tlMBLJE02iL2w22nriwUX+obSG9/cq14
4dmFo0L50SB2F1/7uR7v1MWnnQ+cInvZo+vyNtca1xIZ5Y1YdUZurnvNSKIb8FAU
xsa2gW+h3/Agzcmc2zeVf7MdyDHaaokcwvaOmsEd4woWL/1ScLYoOOYb0OrqK7eM
YWun0vtLypjyoEnILuxlM8IMqgXr3/eWuiRVb258mLrn+K9cSO8GXmaMDqNAsXbv
s+GRtNAb+8Uz1U5q2GiBsbli5EqSa5gNI41wvxQgM3QfvslWWBzIsK5/M4n7c0a1
l9AuWmuDn34x5c404z2zwlbV+ZJISwW/d0voLCaiYKH4GCGwX1Z9HHzFk3Hh2qLJ
M2z5fMTnM0zuwEEU3NNzi3suVPeg5Q9qPJToeNKVBGi5kiM8dlQzJSK1LLp2aY9j
L68yz9TYDV4cDt4Xse7nFw3Gcu6apSYoMLAHDs2sUUFRqcHOkBDvlAzljCKbN6Bt
M5kgdQjxoZSR0TPgeizBDcBVVhmYdcAn/n3YsFE/EnYGXS4HTULGfEZjttgIttsF
ZHVQJNgGX2AeqFjxR2eJktqCX4wgmDHgFCnHkbxv4fCaD6pjKG6bQmnDXv6iqQe/
5BOqXaIdDr4/2zHg8UF7Jir3vZAGO5jD3e8qyHotKZp4pjPjJQIX1xIjVwzUJ7Mu
qt7/wJdfjg46e8S6Mp8RDM4wvEVMQ2fUWetBWAmMcWwTBW1nTNowu2mUMrM2q5XQ
GjBLRaokX7L7BJktS0w6ef2UlcLHpyH4NWsxCRoy096Wb4GcDwLxp/LVfOUB2ybL
NA7bqqY9saLoDext2R55+qEDp2sL0+ynpbIjzGB2euZoW1HmzTwn0xRkWOs3LKib
YAS7l0wKnRb1Alcb6WKI3h1SPjJzOv6fii+eBspROB3b3LoaX88NXiRKNKnFiBiA
wDfEsogYipbJ9RZgJudSHmegGYBOZomOOY3C2HgWGxGKAx4FXcrjeRhmLy5PKYhE
a0qJZND9LUQVchqJm/cypo01m/twB0cZgiTmRkFE4/CbxwKwH2LHuDUjRhN7sNhh
fG47fxEzLlH3fyysCoSno956FYNfrZxoFLZ/wATaBVH5IVyClg2kduUw6pcCGo0u
V0ST8GOnUAgVFTCFqlGcik6HEgYQHyUjeP9KhRG3YA7zUF0c5ihrZuHpUY+P8vIn
DzxNA9KsB2++8aVJuaf5IErbXmGbB0NJv7bL65zgEcx9f9TXb/xiE4tKR38dw6Q3
N7U5T3JT64bWq8pAi7bSplebaRXIwCzLiCrm4hY+vsoqmJal9kzp5EXWa7KtAPvo
E5qB0OtsoAkooIgDlqxrxA4JUuGhllghLVkOZ5+FyqOWiU06khGrMNGpRPsg8LzK
Ry+rHHsJ79CJbS+wTSDXajjrnd8ycRzxSs2ldylK2MuujTMD0+3FHyISMMxaB3Nb
7isrpvr4hJs3yW/t9viLKZ9tNS9HhdZx2Mzw/wgUH8EwCTyP2wacygQtEsp8ndWo
IboFQsrU/KZqyjBtKJfgmdJam3EYfbCTKIS/ozdoz9tQwTtzTpqqFXiXcqqq6c9L
LmebNLrEhb2p6RiNtCu+5QGX7xftBYxHlHQKUUdGg1raV0sRKoTEssbhGWgtSAcY
ujjww+gJsBOEqRVf22QpMHiALinUcmzl8z1ZyYLijF+fKGWdyO4YwEhr40A5KTnd
zmrGywvy97kLj0V9bC8anRUNm5ulg/avQmGtAZgLRXnUrUH1JpHiMsb4Cf4NkQ7b
yWllBlO1B12qcqqzK8fK6hK/bajdUUV4ey1iLUS5szvhI6jZ+eGfgjby+h/McNiQ
tjqiAhk/ACrwtUPpN9FS2nrJjsl+zqxtXlVhQtD8TSgezpairfw1E3tGE3zmUa6F
rkxrgRh2jNIYCyZFX9r31lZfhmhOpJnjHVOUHatfb9DIpDpjNGwCgQo1OYOnJwI/
xD31q1xBVsB+FasvYP9Tf/dGeHh+NSCf8hnU45+FfxlFPE0RWfZ/3V0nnYZ/5Nk9
+sx3hON2y8+O93bj6KDw9gZUZDEeV6JfKgvz60xR2ORTo0JWy/eNB+EYnwtWbZEL
Fsg6pQnsQ7Cw5ZEgzruYYGarft0jXvUlEnVcY667r1ncYebaMPQgt6oUaw7gQZgt
nv+94guX/4qykAjYYsfRIxDTn/Aj7A9zUbaffNC1XQyvEsGh6VrNqs38Y/m0qjRi
6pshdrAwcV0e541EjWeAjGB13NC649mgajg5f2roe7cw9vyWtX/IsuY7IPYJajY2
QpMS1qfJoC2ter03E4y14C3Ja3WNt9RSbicbUsF2iHcaMHBwyH5mt0Yxdi2Tivwx
0KPSQFM0KmUcX2JzSsPfzXlhVSojzgusMQI27Gyvu3MnUvLdoju0ZcXndJOYhNfS
MxS1RikF5XrXi5c/P0MrzLbrfj8Gsmd3ofhjEqDCfMa5to51z9KqrNj20ULvsvTu
D7dgZvqv1PaqkjutzsZGiqSpteRiDBKzJjlWkDTpI5l0AEPNhly2fjNh7BFqbIVi
CzUJHw6XqFZZ8uNwkJStuArAtwa9xvA7xL+8BcZ81igHZ0ruAotmIkHo/3kfVCNU
fcUUqErO1Sq//pegpMvuOFn7m/vBATVKApOPP/16lvg0Q2gcDpu5mTf0qKuTioF4
hz7nwWUVoSBp4aIVcYZNhoCtKT+utsXg3+PpXDhKfIbVMMzXmkj1lcots4rQTBVz
l4fagk3dWPA9MuQykBDZyJj7eEIy8awsTj/zBYqwfJ1JYZORUkvfUymbz74eEnwX
KRrdeebCJk0u9ZvViylOYnbMY7Ieozzd5AuAJYDglmcwpgoL7OnjjtQmF+ykPBoU
ZAguzTF/Yk/roGDOHgqLDBJ2TCRzxG3jtLHcNwP3t80aHAIlA2hGYKI8qCugHGl7
e+fZNeR2KKcCVuXHdfslsnlxGZ3RfyWVw6SeBv3ov4DvIntH2UDlnz3r7gh1zxOy
vojAwWlwImtVF8ICo6upgySiUPFayP8uraxGSvimgCv0Cu/nob4taY5FJPmlMGls
2KXp4OakbnY/BHDk8zP52Bd8iUmJ44JB6//1h4rfn2z/Yih4CXRE2zwuwVhNPgtB
a5YRim5fn+m/wdKmcC5VdBb1TrDFJ7kBZkExMFrhk9BEU6q7rcv7GRvyhtbLLOSW
8lCoe+CNy5URwD91UN+eZUBGe+oohobSNi2h4AKgv7CSPNlWvLqjWBUh9jFMf+Xv
cf5IkgiVRSTDnkZjE12p6IUE7OfS357p2DAmeqtJOLj9TVTcJJAp86GWV8tiw9uw
gW+N3IwklPPHAT7dZnNbHjYsY7BpWo7HvochWes5Bwj+rYFC2zTpZHY/vzUbqhhx
ucgY9PzyBYEaUKGRmpHo9QukPkoj46pHe19K2hiNDK5CGYpjzEEz8D8E1x/BORGR
nKxVZ7oEluDpK21VJNMV1gPxef2xTlhk8CCHtYfwwzx/wBT2rPQw68ugI4vwTc44
+W8VrSsrG9LTHEZIA4rj8SRuLU668LK5M8OVrHr6JIMFxYSt5BMn/4gYPO//G2iE
tRL0W+zd76VoUBlFN0j9GSPFry4sxeDQ/8/hzG9NMgO9EdUp+9qADasoYAS95cb8
zRERKa6KiSiQvbHC0XbaicJrb50QsGBhUAc0ib2NXeFA3h3Jx3jsPdxgcNljIXda
lQoy72EeWQMANXDb9pVPcvsF9lAsSBE+R7aUxTlkI0eXMGy3JogiRbCo4tKmMN1z
NopPaFTirqbHdmcH4QRwPtnM7Gr07+BBSqSCy/i0gmAXJjpJ3EoyT5oFr/BB0bbL
60VyZtc5S80EW94TUQHZPSGaGbZFq1qP/zrGbq4G5QyG48k91+IogKkqjHDd4HXl
yuXgmglkzTwBmdPPXnE7B6FHxpCb6DEZFhLRphQI8JSKsg//g8V9jT26LmuZWi3C
sDPfXH9UKPJi4uyqcWAZ5WUsId0F+yZlPvXKGxj2oGG/tND5tYNYjV2ii+MUwTu1
7hJx6AoYIzuPqLQ+ldJQKttyl5curGgC+23/UcnLOFkP8NgYEnquexmrX5RU2xIQ
4sU3dMz5qNc9rHRHJ2G6+KLg+Dr9OyY6sHrjuRo7/dzwJKh/wkTcCjUOK9aZ+yHc
CybTzkv+uN2G0bShHsP4kTn87/ST4TgJmvRp4Ur2wPD2jsUtYyhMs8/RFZARQshn
b7lq4tG9hrD2lpTPXc+MaEVzL8IGkjxslYpIK9smQnibFUsWelCoqn6HZEpowb3G
bT7tfiYOJecD/ppQfcbKAEMFV+O5r0ofY/VrSfGewQcVINGVssdTAOsmQC+A2Z7h
I9++5LL0UwOVzZ6nsJOioZdcVZQaytfWQhD7bibkS0EY2feD6jD1VcsEIC/rfWsZ
ZjrAfQNc7xRlaROyhpxPXoXs32FFQ0p8VRzdeE4t+9wqpvigB7l8c8dL/nAnWeTS
ByIfXbGLs0pSykdVI4lcI5PLugugC6Ud2J4JPUuAyIzsnS8PV3m2+hATwFsU+5yG
6PvazkAMSSqUUnh5wu6A0rAOA60aCb/sTM/XHdy5PMRiMT7+5Tn8GuGkqA4B2NoG
YHXUAxxCuhxKwXk3i0zdBozBhS+dW1N8BxNp73aSK9DRThdibzVOs4ynt49phR9/
qEBeZY4exaRzz5hYZqlS4gp4zhzP92jdyl+5mmm4LOL4dP9MlCMktn7ZRrmkAOXP
3FiLuKOv0ndJIidylaiP1kdFyOwRQte1S+mKFgHAq8P/AOazDyBl/pyujIQ+kJUk
MiW/VQChuXq1axEGht3FWDTLgbsSBH/PiCWJ4xUV3WVHyJRuQWPQI3LTwWYxiNBk
FtqvTxd9SEfQ/BL1hZaMLeyrWne8i3rzWe7tM6xoZznAczZqsNTiOrqbt+upgWtT
635FaGXLlUl0GNRFnvb178AG712fdc1ydcK6oRZf2Nd1R/NQQ3bngTqoEw8zkrwX
itPZBAGDVr03H4q+R5d44x83kXWPkvYS4zQHxDF7U+5oQtZ7bVyOSm33bhGBTsuc
kxKe23R6+4TIUuZ+3U7km0nJxmGELgsK9/MWBMI/VbwHGJdcUJiivwti+zteg8+k
xIw4S8h39mKOFgBWbji0kzS6tHm2UIHV/rb1z0bpt5v8dDj1SVkMQlMR2mXxriNF
Rml8vagClLsukRo6ye+Kj2tTSamr+rgnBamUPovSeEWu/0hNLBAE9mpn9zXqMYOw
yp+2I67fMvZPOJkIfbb0Zf+hcE6WeKfa4w4YV0QmQtzrBDKVq8eoRl/0dFSkw0QM
6W7u0EKDarqlAyyelLsrdl/navwRVTQwd9X9VpTkuvvwbBc+bAPiUKkpGD16oJii
0bwpP6k8eoYoJcV3DSCCE+paVc12nUGT9gAZLNx048n03HvrPBQpYdbdl8H3quGy
0Iq6kDKanc9kZmmxfvzUBOcLDxqNQcrhP2OFJdirS2H+oUVtMqVdoBzFdCS5uQ+/
dVUeAtBz+Y1tx+fOnqMofxrE5HkfAuftz86ZY9+w/jcYlT+lHtGOoGxNiWYHk7HZ
twHNlrcrld7QvTBawspTViZRR/TpskDezYqf7dFbrkM3a7cREqZmgsiBaTzRDkqE
svDv/MOOxx+9jc3gE1pRlaRIH53X42OahMYcgog6mHICGwJlWs1pxhEqQmmE3vco
7CegMqfOpI3YOaeXesomdIYbCYl+RXeLxU1alsdxw/eiN5VoQ6lF+eByHTwEtAEQ
HDNBByLfSTJ8L+kJHGDFXarUxmP7eZDV2csb+9kaXUMGHMrTz/X1CI7/b/kzYlu3
AkVctrWq1bFRQDdWmqP8Qj6+qiJhQl2HEFAonPKItmeTOwfYv3kpii4VqKku+dJT
QkHmuSvhXQyEwtM0ExlTPvVZRhsQGagXoQqSpQ000Oy0mI9f92nq5rJzzv73NhDY
C2NKEy0MvFgISrG971kM9lqK4OOMST26CdS3jgNkYjalHHbFELOYeAiGK9CXephh
iB+0HU3A6BncKu+YeP+VWwyZdiamRng1396S5ac+tkmOMzjmoVnUQiFFlZSFlRHx
XRgox8CuGF8mwgUM2IyjNSY83RfDYgnx4fKoCKdv/hwmSh49Dcu/s4ovCZRFtMhu
PUq7oZ8BpiOfL1Injjd6q0oKy/DMZG2EVyuCZNGNQ8G4Jf/xtQemf58SO11cIBgx
uk/tMsSUWjtQDUUY6L4cn4drPGAcPrXrGep+sGkEtG3Pu9Lj47PE95/XiG9wsu//
Je9V8iG/t828eht21Q2yaF49g5ETujKrtVtV5NCKNcscIc5tTfGFBqCVbROrl2Tj
QA41s357UUp5r2vumotTjl7sKhN7mh9xTx7w5WBlUOS/LY3Y4GCLqhR4aWu1nNAI
rETu6rcWoEjMEvIxqfSpyL6vuxuXXCaWHi2iLBUomL5V382IQ6wDR+EXV91lbT3Q
pAXRl35sDC17J9PjxXdzxU8AJaLSftfK/Z7mDgjZ4IqwOUG8jPH8jOMWhOJFd/LG
m42H8G5NLmJvUNWiEuMCe62yeXyVHBK0mttqUXWZaepH6i0TBAhq7yf9db1XrjsT
eTWNNme4jNgtNA88KIGa3Sc6EO0cWdiDGuR0s6GPpflI+P3CgNu8obdMQc4en0/X
8tbWXiNmZv7IJArUo9T32WTFSVbEopbTbDtnR3WrS8PdR8cPn8/geALOXNMNT6Sn
UPR6bjS630PRzsgRTi8sRpQSMGqlgom7tvY2zyPgs3W7c3tEkW4cRD+9TU9bl3fh
BQ7Pf0VJlEWy9X/QzKSX6nOwszQXIBy/Nal0N9LLqndyz0H/w+QbBq8NEk8GcU97
7krfKKErUh35LJGrsVUfoZiah4YR1xL2MBQskRvWLh8QCPUHrN/xWUemcaixuOyp
g/8y7HSXpP0LiIzfUCklRq3CZZSLjVOhlwSII2rzSori2gw3gY8wlUlAcEB/VwYv
Ttg8vgTuVoX3rXQjYX0WvTCiGJLgEGiSicrMKOyMdq4Ds+FO98GRI66n0sB40D00
wiYjw0qFe9PyX9g9L6bLm6EgB4KGeIzVE46f1IsUrmMpr0uRLlu/mMMjzhHgIdFt
eVoxG4Gu5+9zrJOoMjrIe7SavSxaK4kxEuz+oBIbcD5T+loTQN7Ule4ZRMj/rImh
x4riIs4ImyghfP4gT83+b0UEYuN64GsMatqePHEIB6LqH/CoOkOz/YgurVwS59y5
wBBIJ1MEg6DuTwn0kmCLfhyxHTfrsFAl3M3QBDhanUmzTYHZ+PAMVkTh2vPTrlYi
dlOT1vJcpraRdc8/GEkVr+O3V5Hpn0y1UDRIi/Fs66UJ+UvARx+A1GFL0R6UGff3
rsdQFcGrkWG1PtGnQYHvt3D6i9f3NlxGWPEwhD3BXsrLTOyxmuEGVqBg3q0myxG7
2lXXaFNAOVkwHq71KqBRSaBcNk4nFt4rQPfVdge22juZvrVw8l7mn4tTLVrwwMcV
ELrEd6ZxJWaX7paxZmm3qmKY4gjmV8Qa7XHs0/Hsl1ZzPbgMi7samVXo/6DsZhsy
h816azw1OPQqZNCP2ht4klHMXQzlZlmhMkq0SPxZaA4tTcd4Tf9mdiV7lUiDgSs/
rxPm8xl8SQk/bVXhTL7YF1Naj4xBmaEaVEt40meT179hWUQ3pc6C+T5it8RS1AVY
+AK42laN0wF4Nb4DuGtoC9G2rf0oljp5uDQnJerAkp8fuQFsITFopwFSDJ+7bLUd
AUmX4kb+LycCEyhY/M0uYqk7sMZi4Ae3KYIStwKWiOOdtKNMKuKe93aEqL/E1jGE
kGiahUjihwKwUmgqH8wOcUFBjSygo97wZXCa5VPXDotaTrL+0XxdBjZgdwKCiHMz
LOI/wNJBWpvrop0qxKHNTGPqzscEnHUmU3VWGCUYeZbR0iuTeA4LuCppBNpv2gPJ
ieHo0OzNQFgOwINAlw5LaO0OYShlfOQNh/ZnZ5/FJco0zL7bIz4l44mdhtNVJd/y
nsZElAL3yVwnLAFFA3xv4HG5dJ7SYF/KpUVgQgNAuhi/rtncAS5hHklF1h9LvYqV
/r2YH6kO6HqtO9RKCC8b8Di66MzzAI8MfeNZi9i/LSMRq5PugE7AR+UAo3WTGibM
JEQfdnuxoCei8mReH4F/MmkeYxN1lmIDGVTHV5z1CNfSuI1LEN8H/MgjW542ya1n
D5lio+hLD80M/h2aW7Hzv2wcWNfVnAOMn6BvTHNHuvm5aajgnXbYPl+AgGgHxGk4
1y97cj+5bjllh9ALaCxCUf3FKzWixEz3B3Blxh+PRMK74cfzQBPN7Jsh1iGUf1vZ
2x3vro2Q8XNZzEp48xIwhYXlgTSZTStBAmLqMmiwvica6STSK9h7Cjy/Hy/giWcV
92RIRX2pWGDq9qedfPiwamMi6YEOvp8+TsADjpfs8KzQf1NiG4FUtF0L0+PwAWLt
vCYMZ7bWnxLb51T43AA2I5OftnUZ4snwq1UgflOBTjCLHUjQRIfYDPwv7IJejKSF
I+tPXVJ4A7EYP6ad8qX1R3NXkbaBius5Jyuy/GFIW6dKvHST/fdxDT1ybNqrYr+U
IsMBzGWTKT2C9IGqwi6jQRiihWClr7BcL8aMSH0CKYJLdv0ehVPQ7snYn9zqC4tT
Ebpqgay6Fm9VN+cMlB5qdAod4ug+pZ4aNy0m3HX2cE/B9xeNqLM0f9Qt44O/yvpA
JYKB1BXsrzb+n1Fl54WLf5OE0576ixrq7faCMGJV/342wzZBdZM+2x8ixI9rh5lQ
a4abgXbUF0JC+nrvaitIfxec2ht78jUGO9E4He6iR4D+VCd1t+cD3vnow2cNyjfD
zqCM44LDewWQxXyvHYUX8wd8GzZW4HVmh6k008H/20DazL5T4j7Y9rSeELmGDE1z
/bVqRs/mdcB11TZ7bmuU8gqFUaQzA1EtYJyKwbqKtY1D5YDciNlgO8RxtRBhF0xI
TqvyeplWrqT4jlFugppsODhR45QRsz1WR1Ar77lNgcizRfnEQE3ELY5putoRqsTH
q+JLEGZKrslaV79ufyAdLmtUEr/apMsLLU6CpE5YDQ6SZNoX8RZEfGNFe7H3t6xU
/FiEOLPCgcPLoeUXzaTF8TS1Qle9kjG+hh7xtn64X4uXBgMcmJX0FbUyr4PxPjJO
EKQq7l8EqY+ZWrmLTR7EvuWBlOEytzlsBUkRnKJ86dQqnUi6BE2z/nElxXBPGZu3
hqnFb6xwLxITuwHFloioO98eX/jbShvMhnlBeKj+C6ZT4XIoeGhV5K1pndKybNCR
GxIRAXtsWeJ+8ziWliv6yUaXsP0x4R77A6M9pC9Tv4T2/xJdZIU7QBFy2BnytQdn
PVHUxGVQvWPiHgI8NC3W5sHwd0/7RCax118MVFBqWT2hU3tJ7+1SmRqa5ffjaVSZ
LDbwPAC4w08YUThvQ0NsNipMi6sqloaGqZfScovLYwN/U+qn5dyiBiBR9++7B311
MTRIuv3J2evnwQIjkP2zeNEdNy+6LjYKLlX207UELz9oopOP7nnbzOwvVC4z8byy
LkVQP7qSqSF2kRXIGHuAlX37ItnuP/0PkO6K+sEnXBYXIgGoEbhC+zppDM9ixpaR
ugahcHVNQBMn9S+dtrPBwgew8kgHPv1bmAQAQ3xWE/AtFQeIvQkPk9Arim5H+z0z
c9Z91CeENX07zuSKIShF6YAugip2l9nVildCddEuz7jqKwMHaLtG5BVlOGM0RKhy
S6hYtEZif/SB8JNoSxflpCK2eNzQ67dsFmn1ypv+KrX1WyraSSfgDbiLgEwG/Yys
lrptjVpIfyvKgupZA1p7YID10R+GCcPfUiU9syH2nJUh1NGfwh0o/dbswWUzm51u
h87uPtCKgv5LSitSPVP4gW27pYeJvdN/PN6cdjfjixSKQqMEokV4qetEpEM88VhI
vEfVgxRx/Q8KXD7eqbzhWFOHkN152jS/SUsDXuR5wVPOJJPU9WKYlQt+b5EULzDM
I3hR+c0fPZpot/uv5yfbkgrVOtF129IIAw/hZ17ayyjAsBf53GtOyudeb4hXvIkz
IGy6vcFlrF2f0o+a5tYzzJpS1uZRKho02D2FTmaZiD71X/sS23hM1ziJaHh5Uzwn
yTGDUUiC7OxQlq79HAEBFXxrFXRnfmbKuVfoMAvjzIw/r3hl+9DtfIDUBjivpldk
rWNviao6t5fUHG85EpVkKidTmWP03BSUSL3yzpa8ZbWCeOExwo66WatVt6xajKYD
jdHlwGGhdnpF1zIxq/cxZ2D/wMai2rxuj8vEzb4Tr1S45coUqcZb1pT5cfchyWKp
2IVT+JQbDVEKA7GfyT9q7wxC5TZQbSSsRjd2YVhBhtdwanbHPNxNr2noCSpozyZj
s0hframsu1PHFL0OTp+92YWoqqXF1ktBsBrpSL35wCWwHEb5MphFfPQbONQcr0SN
1FLrc8DmsP/fpFSZ+b3nxiOC0IV7kV5Ry9sqF5RCQYpDPUql3oh+XIr+bYKb4NBn
Qc0l6uR3yipftJiIgJMm4tiO/Y80fwbxyVkr6nd0Zg4+/Wk+khPTqidlGyIG5me/
Nsv2CgRdjDcijqquuJsq5jr+IbqGaLJOTk51AMiaKuV7duK7sxnPwS0FqGu40bM1
VU0Ydgea4OqCi8FlenkL48ythLWuIPAeE1lATyl6qRA5s2CMsY7rCQiL/1wigGNC
Sp1kc1cISxBH82XjlSycMiDbNwFYXGNRcYjdvHBS33Wc5QKObmYGSMZbFuRZdPCB
zAjj8CsPuPGWbviai24tnhtiaamSAlaRolmlz9DTHHnaT6VFCChtsLsndK/DM3vv
+C6pVZ3WT6UxbEoxb4CmpOJV/MoaXVar26YaaqMzk9tHS3yy58a8eBnR5uwp3u7w
57PaPhP/BRApgyUdj8sT2/MTbTxcd+rWAvuZqPtb0GootsdhUZjA+3OpTCZTWAAl
QS8MwICTAmjoQrqRFUGPrGnJmcZBdBqoLw+y0/vunHV4HDqyb++DrCLVQ+502jP2
cCB+mb1UO9e5mASRWnEYqdaSgUJRgv/+W8VvVQSt8TLRqEfqN2ru+OlcpXvshoxt
EkBowpCdVXwRzq4C1OkEYOp4rUoP6hR3ZzjhIjFki/qew48OPlsI99fORQlsknwx
JmQpA+i2tz5gOcnNbf/bv8QbK4+w+tnD96ehEulincTn98H3cbfIzGvaWgtB0EES
kw7p2I6I5lLleIL8bGoWqO7/DW8afhCxn/W7gqAuIlXk3F7sYYxfVz36My0/sMQx
t1bXK3WB8KisjZ7RnQHuku4vhLXodh2HuhU7fxpoliaw/JlHVZ5cBHpETYl6njH4
CD+JQ7takKcBg5PBCUbRtyQgdCFHG3tW3W1CG+p4iG4AupV0hbxtsEP/Sb4KzXvF
uaowE8aK3pRV+Q1iTmyXSpBaL9HxCDIlLBKv/CBLGZE6/O3pUH5fwp/GV2t8Kb4v
1Kqyu3jet+lydEX/XLMK2OJlC2tDGoAx5dXcVNcYv/8eDAxkIZDtHoAtVy8fm3SU
0sYhZrlpciSd/0Ee8upyy/b3dpLQ17FDhfmj/mpAp/szlhLhlU7wbVdHNO61WgEO
yLj0lF/dGoHK0tmYsLWVEbebVVthvK+XvQT5nqTdm9WvNoxAWZ6mbs1unEAtnnJ1
QRejskHlEzOggnL8sucQFCl2pO1NwZePrFi/NFoz+bh20dttnxG/RKgjfq0d08Bb
OQ3ElEnSulIpLtC9qzNog4NtndjpNeAM6xciF20jDsBqJJzkl9pURQFnEA9fLt7V
mcAnqHSadatn77WWqEB0jL4Xn2RptGFYjjB3lPi8MKcsueoDECbnVE7/NOl4PhYF
s8Ik3rUJHSRm+sGW6t/2vQsxi1JhY3o5uT5lDVtIxVkktGfv1oMVqoL0Fi7N1oM+
63xrSLnJhUYC5vAZlIICMBi1Qy2rzL2uqWas0Ss0dFtHTHOOOWdUaxrkCRHbZk0e
ORrglToApKhZmCuQI4lGRioRoQ5uEqNHZ4hXnDY3acNiYpj3qI0cZZT8/B7czlL6
EgIsg7cg4jiMNxRShOIBKNDIzdYCT/nZ+FwjyBSSlIdfJjuDcA3CdQ2d7UJw4KVZ
4I7BUxOFxpVGsel2EtYoZuzeji4JYMzLMOpGrtGAlP2AYMUJwI7VpyBY7bAb+KBa
abd10AbtAaWSS58BdHLZdIROjncE/aQCNcMGgabwHTe9Z55pyOwFjE+JwujyPVyX
mSsbV1TKqyJ/pQfmPI0HuRNJwiQKfuC47lBmzqM9i4oxKyVvuzfqP3SOeg/lUyd4
/0XZTcv7zwrlTm6+3xdpbZ5JOYNLvGYeelJb6TOAXOIKx7vgee6tv5iTHk44ZMcf
uwemPrU/dbzYMMQddiuU8gLfT1C68CZ1hEBu5D1hCUVSZcytK7PhfR2jmvh0kyzS
HVApOBQxI70DHMneiHNyOdslITi5eNRmlauM0OfEBW4CzN2JYsOvWpmxKB0+l/xl
am8URK5lzPJNpvMupu1XGnKRHwR6Eb+j8B1S1st57FfJYF7NF3lgj7zGWyOOhh0m
PwV2ea6M7SotC0CXgTUvGM22kCo7nrqLpzBDgTQaVttdJ5AtrqticBcuPelFSwVy
3n8TWGldy8qWTDW7Bw05XYJhSR4sOW77Pu38cW7IH4o79HTFHmu3SVBDgvjFyYZ9
xW/6w1wZRobY141BEaD4ksTH0GH5cpvc9Rb+3r2r8idVSZxzbWEL2KcMkSqGQKHR
2bU3MjI2QFm5cWJZwERkm6AGkP7veG14eph5E7n7kSVdyTF2sz8ZcPBXCQE9Ofv8
uPKrT7lGLOepCknQyzqb/iOwSwfWnCX+9sctf0lHUlkXKubFppb2oWK+1LVTWqRb
rGGE/AvqAGBXwUEFF4AlXCUx5LW3GDKS/p2RxsEwf4R5kDMYgGv1sqxAQ/a9XyK+
w7oes+oDXlvhWIGMURJlgzoPzqBhj2LsPc3g6tnCKojrt8OooD28PBh8kzK/wlIb
7ZAvqmOQRSxWUw55ZLnNEN1KMa7KGY6jnAiz7Gl/6E5hwrChPdcgn2bgl2J6JoHV
hAIrHVQhNwhBhuYOCPja91rJEij/OHPKabIpp5rXgWjW5HC5WzDqxYf3eEQXX6cv
eWYKxW2wM09CibtXNx/DLCPJI7RCUZMiDbiBZyhXPLB3fmmlNouk13rcoDmTHPnt
tnO9lwRDZzjp/WT4Iw0hR9/4ZRO2Jo59QjNqD6MtVk/lFQtO0Opz04xfBwnCXPza
SbWhfsBPAGwXMiCVqvrLcs2+cGZ7Zt+08SnHDObqMsOJ0XPI4VG8CrfzsI3qNrSv
HPJbOFUcXnLt54pFUJPMbgtslkkVGmz3tdZbxGnzwGcg/bWf+B7hIYA1euqxm+gZ
WIMzy9CT1LHFRTOfOuOaa/7XE657muDYtoJjbPaMAmarNPOap01D/noDIesY7+2k
x/rWd5mq9FxpdMKA0SdfNQY9eIefKKDVUNGlmW0fbWOnNKnaQXeIyOd1G74PsB1H
IN5XE3RE4HuxdJ4PWHBDOPP3RmJcCGicZgjTxg4pi3gXEZYT3qVq+EYeUFyol6ez
oYKHo0ErwFRVS08lX40mgKrlBg3srZ7l09HJPVXDJy9OGMGO6J6wQuuSgyvC1R+C
ek46t8YhGtojS6oz13wM9J8dhQkN4+092tQn+6vXYgpC5cZ+ofNGb5j/ThPOxYBh
teF596T4lGD03BY6l0gM8ZBHZtuncnhT0F6d2WdpBxU4hDpAqy3EP20JSjYWdZit
3uuJONq0AgfWmhhuYeLbiN91WSkT+0fLgWr8MwMW8BrfXhu9lb8ZNqd7W/Boa444
wbu60gFKF8Gv340bScNFi+TfDRBs4OC+S5+q/rI8oCY6abuCmK0cFmo+FiJAEUaX
uCrHSIfUP9Kb9X+NmkUH/YjjtSoJ7uHgPyDS6j/d+BMa+0i/CcQRMlDg28pYKhHm
gRooVbTNRMqxYpChtg7dk9MU7QHrtTVDBGsvZxRlxUZmMbJjZK4PU9SK0OFsVzqN
ALiUjmW8EFfhw87OrHaeSJc9QlWUoSpIgL/0jJLaQK9eTsZZYug3xAP5T2xEtI8C
5ZTwCn2eiDYaDRnMN5KUhFz5QMqvNMFuQ7FZi0859CWW5oG82v2Al1SdEYyoZMfR
xIsZ2qSnALtbSahn+yAXTpIZJQcdEOB9RfL+ftgzgAhKC16PVXG7w2XyhL+oVr7z
EKV5xz8ZTq10BmgZRKdYvCqm8fnnRHnh1CydlMlfncwOZQDPAmxLanWyu06X5kwh
No2Qo8oLTJmbBBiPtF0pEI4m229uev8GQO2spWP6zINViJ+2PeiSeaCo//KKq8o+
k7fPcPUf1vY5DsbLwDRM3em2fQYNYDJkD5WWoqL+NdfeR81+n8wLrMu7sUCyXnRn
XyRngnHm5XEiOvPf96VdgyEziLs05LEDX2JPDdwWQ2U7N3wjFANnJ7pBzYdswQwn
UW+NeIuJFS3cDXykaUeNWWMts0zb+/zl83g0Dt0wJqCHFsfhtvoMGMT1NOTP4mzE
2jY0HLZEf5dQT5qLzYrW/GSYRURV5gLfPiqen7JJ7f442DqlNLpsm9VGfHnnw22X
Ehb4my9nrC6JSWzngseUFaVoytdLRcbHKd4pESnF95rzYVG7Zm0smUsYy/XgZvu8
7vaktf++Nmmi7XgbQPLfenNrCP3aSIgGg0/4p3DmE6OtX6cxrt95ZdDPs9KiAPob
MQPw3aBmBAB8wgxz+ZuImA+zwyT5JeKvK6CYDJjTwsQHAsmUQf8JukFL0NKctsWz
p4hWWHIRgyb5EgzukhuiAhaHSrFUKI3RREK/De0xXDPlTB1mUuAzbLtMhnhL8GtW
ymRVkQ1C0ymtMe8H4WKoNCngVXW2nSQyNiBAKhb/EGoyKdD6cn9iOgL6O7OzVliR
AhiexMZpTY45PKuhfhf9I+2vZpMCU4vrTqFPoFFXbwKRB4tptcEhAqbGuGQjx+ZS
6tXavdTB3Fmp9BW5BNh314StL9UsxFhv6n/haGg3qqfKYWFDDGNjfPurAEuTsa0c
KTjyZe0KUBFbjIHpbTGYRIjS+GLrARlXGY7CF/Yxc1aIUgy/lSdAf5EqhffIPYSU
8Y04lLKiFG5aWt6aSodtShW5FaMTt+GQ42UXIhNK7Vy7rCtrHdF2eepU3NS5rOoa
cYJkSvJ9uvQxaPCZeKWcaEFnlPzFYY2jvPjUj0Dgpxy/22nV1LQz8TG+B+QaBBsm
SWQLQUnckLj9yBXZT413RfBQ50n3UlUZ/WkwNzUTTnO8ZhIpXna9VMk5xiwsKS3N
XOFUx8ygXuRPucU8BEijDE/jCOwmCrzBx35DRsKLpI3HlRJVaFLudM7RLQlXBaSX
tiMo2Yw0gkDJetOYSHjtlr1bwhC2myEFd0GOQkd6rHuDcsHKV44zvGP+72uoBVY7
3QtxdYBxC+F4+5ZG6I5jysFQTh9UCtEPNPNYl2N4sUk2uA3gnGyyt3hvXbboZn6C
uZu3W+9XUaLK6Zd2WcmTrQOcKByzr0OpeqkqccYObn22w3qQ3POSI9DjNVxnMoOr
8FG0oN9IBsxNXXVC6krhpooVfKoHgd7Zl5dtq9Ikdsa/dPRGinlLzPQRtVaAl+r6
Ydt8Do6C5fW78etacAfLLPip6JfGrihRje0vXv0SM127/EnjaKeDf3ySEgQjm5oq
eCLEK6H9mX7h5q7vSfrFk+Sv+yRlktQ8++C/U/FezWIf4iqNoA7lSiBXzpjDSvM/
YF2vI9S0+IGLkG0FwZPBpcXy0mXgDmztqeOdHVCHjXZq2Emlm2FLhUuVvoM+yIIu
FEsvm5E/M0Rwtl5BCDpqcBn7+8r56aD2T/3I2A3J5VEAGnwpYx8+XGkMSsqk0393
dyGzfqaWQ41779C+Av2Q4WXcdaDuS1YYvSByYZ+K1jS+FaITQhiD2jKzbW7js/8Y
5nMq2dLJ9T7GsTId4vCOpKox6dc/YaKf6JxvR+qRCTLBbZVSVkikMoHDi+r2KZT2
sgxE5+M8go/iW8afa5sIKUMqQR4m6j/QV2PKdCWDxdWm1dZliduIQIMWTZsIdmbW
3IxKDrDiAXmFW0bn+eLjsUaa0bY5NwP7YZkwXQa7hiRJHMBDj9Viz+J6uOP3NYki
aHC1biHXB7HUqjxBGhQ/j75h4bSaP79S6lxP2FIxjYrGwqjV+CX07un6k74y7Q9r
KEDKD6oRTYDVMXa/uXpg1/BZOnRfUHhVf+webDaIHHC2NdL7gWs7ElVx8MO7GEGl
2Q7mQDRW6821CLS/fcdD7dLuCiTghPVG7GcpfdrRZQzFC7NQF7TEaHYij73AsSyT
Z8ZiwhbEL+Q2cwMRkXQhdgatOiU7VCCkVGxWoNDmNiKpj5aveT9YJWaonfdcOi/7
S6avW8RxSoyxZgNcjqi+V1JdlqWZhGtE+1Jqw1WAhw+9CVNhSreA7oFdb5JjeQ2v
R0iGcVr8zvSHhioP3WVcrSJWLDp/aMX2w+dHIwdISUzqS5gTGWo2LWr2671DkL35
dj1WWZw35zgMgMx/hLQNfEUcXEXaVb3yVPTbLXjrGSt3LZp5p0CxkQqdhn0buR92
NWSIZlmzfHbflofbHf8eTrugI8my5JVrTcPZCXOdYOUCGAYSkNxF28vxqJfLz+f7
PxkeT3SVNnAoEsR0p6vhzNBZI7FiDKv/lcXDDX59m8G1Cu7PJKRai70J+BN/HvoN
45CsWtd8TcAQdgZp8m0cQRdzXxE5R2RunZd9NMPo8nPtlnvAwY6StN628qLykD19
sUwLMpSyZraeu2G+mG6HL+y5furKkBpxCp825Au9U5DU/Qpgdj8LZMtrLVZwsdyd
+5o0YuV5VXk73EqpmAPf/Ui11r73IAW2rvHPcUKHOMChQ1tgQmiIucmNyRDwERGi
goUwC+CoZ9n5nMHMlgMujzaBBxLracX/k47QuTLLZ61sOWH1xXxyIzehVg4bhgqw
TV/AEmAnYonX/GlqXyukLD3Q3XkyOED6fmu6t4LaePYbX1SUipiDHFPvJW5TyW5U
2CS6NT5neT/qqU6zUCB/lnEbJm8R8XlLwEY+sc3qUep8Yr+vk+7bO77G96u1N52K
c0KlLEJtWho2A2fDTTjYzt2YpqpNQnsrthduTHg1Lse88++I5ItEyRAiMF2mIGKL
oiKTaTPWCT+p3g8LrmQRefKtFq9ozkYZ3EBvNX+gthHKjpIQBFaMwRsYp3SSvyK9
dZxNmyQ5vuMQYhSaYE2gXZOJI5GelHfjE0Eh63Gwb3CdCGWFcGM2J+Hg3cPQQCBs
hGo2yex2jI8elzNcm88HL/XwO4k4qoll7UDMeZrs+WOXfSNh/G1mRf31eZFTwWVV
kuKP0dR6IP63v7o7rEI55X990fe84oZVTmvE7fIiOg4mjmeRLfRVvPgvc+eiUGog
7yFYPH2R06OUaoE80snkj0x+Wh3l49+mxHeJ21jamC25JRf1/00KhVGUTTfXJEoX
lpJZANh/OH30wN54OIfhS7YidSOxVDkn91orESrDU1Pk0EQT0qUWQ0NViJ/fZZn1
33CmV+b3w4TmdDbNzJQ7UrE4lL687gJYJs3/lnU/3XJCQq1xw0hm+Ft2cTyaFrdF
2yyl2a2yOX+fZvj8kjoa5DOuV7whwKUNcIkGtf+05weU86O3HjLo1wpiU57ayybr
2tsoipu4AykeRMCUnv+gVGHZ24xaVvOwnaBpJSDWHihqaUIfSZ/Jcs9x3kSemnSy
grlg06Jl96PeGKsMOlUteqsfGkK0wSsVbBELiTx/POW+dEfJwm3tVHpu3tx6OQ0g
KCIiI1g0nuPRmrOoMI/xVNf7bc+pFKTyEBQECjh625AxqmzVpK/l8hGoRocrqv77
/7edKMFXq7ZSdzlOkL4nBBofCv0pmwIrgchQw9z7GQLc/OaI9sERoy6K6VmrT9Nh
NWgOiNCZsBs2D6o+X4SteM8YT8eKFYHEBvP+BszbSDdjZ7Jig23ZIFUCMLry3U4j
InyK9XoEu1e9ocdPNoLfekDW5AQXOv4pAHyCACY1d6cKa2oyOgIeGPrQbiWhu4xB
kXLWW6nquHt8sCZyjvCeA2xNm4E1M/QavdwcNOAQUhXl4+XtwOSAWBcOrni5M25R
GOtJPRzPwe8rn2AurTOzn2vxgk7NlON8U0XaSlVFsYB+K3WkMYDbOuSxdIWs6UZT
l1U4OvRYWO6D08+AbDfGQTkq9nintldOp+usX4mhp9jmtGuCoOjYECRtjBz4o/dz
M2CBatTAafF4irC4gyGMMcIjx5hIIhPEvZWGt2lo0H30EUi1XdV8aAJG5HeUfAkZ
WbaBeF0k3jqOwOBUOAH1yRAgDNfKEESIJbHtMgHzJbGMAvz7LI7pFo1xk2pUuPLr
s1mxYTGXt1wc0ZZYoOh0HU+smVDiCsPQcBim2Af+m59S9KPOEMaZlzcMLCdrFxgD
b4ZNDPIZXAMC4KGFqElw7ku+nLjaIUtKzO0UNFTjkW5+98xi70/Ja/aWLKEhzlsZ
ih8cW1eszR7lcgev31YxfIcNsq1m9VWrWZ3Ao84L01ybkKMwetuGCbePUjQ9AOtC
Ej0ZqfAX6SjX5+VM6mZdSD5amjf8y43lGdKBRKAlqhLPKhlBOY23EMCdHFHVXE7t
wdl2K5IkCF0nX5bth6sTFy7X8eTwVTIqs6ERDj0VC/fqNfCIpeH0mUPjQkZgisvj
JlXdO2GrQQW6+CzYxTj9MD4gcnZmpsSuuYEWF6wu8vm3mBl5Q6boS+aTD1VdpcqL
luCjBDztlMl8I0qdqhI+F9U+OWy17EvMd0PTtIFFzHglTA/fYnE+z/t0XDW1dtAC
ed6eYI1RjKbYlD58nf2LHKzofs6c4gbn0lrQSoryKrH7RaSN4uytWdeGeIuswwUh
SBhIDFfwhB8VyL6ZlUcmQejuLbdDgXGPb8lqvApLPwyqAoS8bkHsovnI4J0g6Nte
xDBqhBgjM0DPex+KikEqb8UISfxE+gFqzGfKgc7K4xR+1besa93NGO5xz3G24Q69
VXOzI7KuHr7kBChuwUWwhf5ATUu2C9Q/zUScHMct9vwJxCH9awu9g46Bw1aUAANF
BDSDBu1eJoFc5uClE9wcQsNA4Ss2ixBLktLHwmlwiMNe9ZZyuY5nkl2KyQcbNYdf
ML8rxBwODSnX6mYaq4CjXyEUU5vtHYcR6Nz5U1VXAceY9f3O0qGyKsGIhfo+DGY6
eecxIfA+ig+Bg3usryDjic+SD8g6Hfjx2SZYJT8BLrW0Mf/Ly1WWHVIe4I8iQUZk
IGHDKVw5uNSKs6wQArdjny5A1H7XqlC4+66iq3lz50iL20vTMAr/SwWdRELZ/Jn3
bAY7rYUF6NtgE/q04/azjzLXBptuLuGvRliKmiKH3i4oK8HVBHwCJtry/fLQmM1R
mGxEPUOBUIVBS6g8AULxM9WF9ZoEVAVzjYVSu07SV+r3/GxLYfo+AarhxgQLfgRZ
lXRWzn2FUDDwU5Wp/ashu8V/XmAS5F/SVzb8/EJJlyCQuUG/g0c86oFNnfe7QUuv
dESQsPZltMoYnSRP2cTV3JFD3MODuxBXYSA8I+yMSFvbobdDdX2qN0yCLhtalJEH
bdLUyeOqxlfH3zpufdnrpvJnev2iDgJ0zbzEGoHh8hAJXcDiPV44me1QElgIFRL9
PF7e1X42ZGw6FxO9m6S4Xz8BvBkXmAvF42UIwdiQgJ4gn1hammVTXtAZdXWHJUo5
kkb3KtlBmYYPMUDXJTfitYQs9+Qn/gzD7xyY/vox1a6GrmbVqvZQbLEmEZ1RDEss
DsVGPLGUoopLXNN6dsKJQy2PnkPFfjq+lhLHoMoNxnb4JUYay5SfKl3/7SoiVENs
dg7hNgDsuDgrNW2lBve5gFnI9fen/cP4Dqqi2Pnm9v409xgmHvmpRU5MFeGL/YE0
J5wiy1T//CIALFrmfSa9Y7gbc6ncefNRrkFmLFYtGdSxQQGjSBAsZTKMMJFbEApi
HdBQTDQ6I75QMg28UwmRcaamOKw8wmFkKwtfh4hboU8Y4/7DwqozstX/pfK4JwAI
XS4AB4OWEIGAenG0jG+T/4j1UeNHp0demYvDvgezyFrmMkc+EuCZJcPqnvcWq7GZ
dXGtsY8c37aFkFFRA63xQNTpjlSjyt8I/NlbPoPcKOgFj34t0lATX1qDc2yDGlgm
gung8BDY41uCLlX12erO1ReXtmyaJT79+pnTup7P2l+pNBzM5G9C1zDhG5/WHhfJ
KHoZ2v0biaeEdUXO1fGHviBPu3wSpT2mcH5Nd4Rq6B3r4J53kfXBizFMBOv5eTq6
8CvMu2W6tEM/IHvmWusYQ0l7C2BaIcdvrRUkC8CWHhqwc66bnOG+8drFqSVyMQzj
J9fAM2LGm/GartS7DkssaoBpN0wpCCP+Cp52qr/zPEw5f8tRjaSW/QuQGZT+C1KR
auVzCX54Ier0DokFQRkxtVIMSpBKWzX8hLpnyqUi6+R6CzG5f/EHFVHZRAaDV1XM
UwUxdemQpt7hBKo7RTolC8D2GpnGAiFVQ90L1mb0bMo0PyEh61OAiJSbRfJzwX0f
Kva5Lt5+KNEsq+Wx2sFEMafGrmDRLDDN8q7vHJZACJpSdWeTPBFI/udxsaW+h6ge
IY3b7xieIO6GJmjLbvC4qp0wJQMdRr/xubxl0xhwVMDZRLVogDC1lduuV4juDJtR
zRFsblsjxVtcCE+OPK9fE7pHjueiWnLTdO4ksajYxk49A8PiaaffHutoNfFVh1HA
wUOW6JILFLniGc8IpC8ECnVOewcRRZyhqvmGvGBJTE8ipXj56FmNcSzJ7xKxsB7m
/mwXyW0YqHXmMrY9SiGkZO88fLYOjiPBjvp9QOxAzWpXp2CXl+1MYdiJRlF3byhO
oNhVqnOJV2p1wUi/rxcmHYBgtIb99myRDdJtdHyQhaNKTCBaQFTe1MydsITtIIxu
sI4t70XD1+nkgu3o69CWcHDzOoH35ysQw314CFQqEpwbJYDIQES3gnLifa1ciawt
+IIDZoXuorDuFLKCb8v96UvWT+r4K/lsYbe6WNH18cJMZpxFcQ1S3LSuaR6N90rQ
xZd/0SWv7rp3PwC7ex8eqE0x3PHe7WNLWWDyVAEKCM0Lrxss4XaBtu3iT1d89l8k
CVrMYkXxFAATPEnCK/TNAviIxh3qghvDu1RE5OMvlAq4Jj40W2/7d6kCT5vGzLA+
MQZHohojoX9BG+M/zYHcmYVm+GndcGhg1J91/wxM3mktGfG76yGULEeAoBCZz/mN
m3uWJ0ox7/jLX0KE9pdWFS5VJfA9Pzps/ipqXnnzHCjBp8ZgQeCuH0snMHxJxu1a
CGmeCDhuzg89PgBnzNv8FkyVZGFNFGbXW6mJ4cRPsUE=
`protect END_PROTECTED
