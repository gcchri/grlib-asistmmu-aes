`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O8dbCSXIUJx854ZTTVbQ1iqyU+SEwEsaaSufA+DH8LlVva9QTwrcw9hEpo9xPNu4
8XuJ2hhOIMK9Ovyys/tlNxgado+Ny6DljlmQIk9uMjBk3DblUV1ThWELGF4cyuN6
AjHJnlroRjciehp3dFK9tacJbkE40/kenXOJmdoefSU0w9dtRfSOozI2gvITRl5H
aUvIWt8v61SsFb7KjFmLJUXFN8q/rbrYemsHpBGlKe0iAvR2m+w12BdjPJdKqn2k
f8aKHigBVBDPCXarTtDYUKEBZHa1vbD6O5nxpYbucnza92mHG51VUqYuzIKvNcX3
AFNfh36LRbVfYQPE/a/u4w==
`protect END_PROTECTED
