`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5GAXzPm9dCJcGerHMg7hdRw6p011qmlLiUpo7hue4Ng2VLDInDnU9ygRrr3QLv69
fWOEooU6fIBm4l6ZwcNnRt+/VTV5UKxq2qpQbY+TwflBoj2o1meF0rMjxbdYfY18
h1uUGABayQWYQVAWwLnPl+egR9j4LBKg0JNkhHSRZLxW2wwnW+4uW4nnjJGnrNbi
MPOx57PFHH4NQib8TbKUFVYzTR8Wct0IgfaAX3L0Ud9U24dnWL33IEeHPw0iauoe
Byx8t6LiKJS7jVWoQTUqsAE1gxO0ikD/fw7nwhJnuTqo63w8lssEf9Aq9trxDJSL
hfS5qhvRd3A8xk1iIQc7bbKD2vi1kEyJpj8T2DDGyJOY3X4P3Mr++cuddwDTlb+Y
u6mvoh71o09K8IOP7zRm/jjAdC/s4gWc7+QL7lw0WgCuJ7SIR2998Ljy7Uwr+lXX
27q91BglcLMtdQqUigTVVheE9YkBCQUwAUJOOorF7l6KEq6xeHPrPAnzeq5hE1NN
1eNdQR9t0F32og2cRwYvB1Ypvb6KXDIhArbW7TmC3S7Dp1Yz3CamYdr8Y4o24mfG
KtFw5McyiXB8Qr3ElUH+zBv1ZvbX3ZnGeSEr9KhlX9mXo5YSuNxcla3bl7piTl4K
0TKuXGjmfzaPiwFycPGcHC4z9+2EP6J/5E9it84ujgtz9yWTG5qh+1+iVk7AfZox
HbEKL1JdMe0JhmC5Nv5nrhOEmKQFCzNczG9M4Iu5NG/+cQuX6fpZKbS/K3K3/ImF
63Fj2NUtfYZcHs/cLDQOOw==
`protect END_PROTECTED
