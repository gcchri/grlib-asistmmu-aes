`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y0s2RAgY2Ngm5axPq9KK0dvWNOHr8an9Cu4ZiNTjKZf/B1bCqYANxzITwpmXvDIi
4XzK8lA2ESXVgNvOfx7J9ubmXLEGlm/JKjgY2sbqQh/0DdiJjSJnxVTYM9X2GJtL
GZVEpx2ZJBAJjF21IPb/PT3HVUOBh5zM7ec+a99bmRMClnPwJJcSHfzZwOehGGc4
/5uY8LiwaiI2lsNN/T2W89t1ojJa3LjSTu5ckXMbRCbLag/+jCleNWhtUKWm0VKe
g7biV34tcKPzHyry+B8vEYQgsJKw3AFcdmCSzobNATHoqc4+DpDz8h9CnIKMLIBo
uN+JccPhUEFwF2XY8Y/tMQflWuFHOenx9mqdZ0GuuOoVPt2eDeQ+im7pHhIETIi2
jH/DaRpXG3HLhNdG50kHIhq8zQJM+RjjnSeydBYvfgMSG55CW9/j7So7y6lGPrgn
zlDGZJOGxmiRnBHjcKwk/WGes1EUFQht0GmGMxtBPE4=
`protect END_PROTECTED
