`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yCr9XjPHMsY/JWTU1q+RadUG5JxggL+feIzrzUQjoOfJ5Y98jkNDHklMGHo1LPWv
1ZUjTKpgJx6HczRvoSllfcQaVo37Cd9iHJW4ho4Md7Y5c41tXxnL4FevLNl+vD3g
NmBXRBAD9h9jUm7GURVO8RsFUPj3yxtJ5M4QQNalzHGDMgZyoTW/7nmhN9cHNpPo
oRiosI+XSD8d/rpg03Ew3HE9wbF0CwPnjqxil1W4vLix9pbGAkvGtwxaJVAMTYXM
Zm1WM/zghHPH8TSCxcptq+ib+RJ3T6xMaLLcMUFBDpKgr/+30hj+HI9AsM5ZXhFJ
c0BenXh7AMzblfVayYE2FQg8NM0GvylFNW2xDehIRP+CyF7Z/E2jPhNvH70OzS1m
0C/5sAEPnQswjnqJst0WIRRUfwlilLUozXNXFjRR5VZ5n+VAojXuc9t7BDhMCXso
kMaEj5ShdLWL2OmfD+iicGkDo78RR+6kV16jpvI+M18cEg7N7B7wNg7Esvf/+S4y
l96Z5i0fHRYVCyrOFCgXFhidRkHt+gaBh53sS7XP9QzXErZ6SPVTS/Mvm3heyoeQ
WDdmvnFxQh+FhVUgkkPRFWVLWArECfoY9MyOVoelIcntuNcB6TgshgIkQuhtVyX+
22qA8gjhimrLmGe+3aG0dgXriJHr/m6aEijZ0r8dNuiosqq1oijbdlmJ/ujBeT7B
fXYZTJ5mgPaK+TadKptadXx7p+ixhddQc068yEaHXo1T9OAturd1zFeCgMyAGOdf
Now5qZB19r3p/NOLtbg1aVhDyTs9Bft6dIrOoeEb55zQEsevixatIwe+fqxvY/73
Dz/RS9Uf6u8H6XQzUulMQIkCVdFnXh+8e0UDLZsJ/ClFnyKZH1Hn8hovohH1RzVM
zjtRFBZHhvudwXdKFi9WfvuCWWiGw+3k4UTh05R8V3fRvoSRqB6vOm7RtQB1nRnO
JORrRV5XRLEWV4v4ET2XyTzC/cap+B2UjhIz3tBfm70M9kzxz9Y9+ZkNMM3KrIUM
46zc2o1vcrWGkQSQAMMUc3fCKVbJL3CeIhmcimK004tzMJf5mfe3VovB4bJ8eHWX
T2DrW+nOx0XlmQ1B1DFsdGUUkyvPTzUty2srlRcUimlJag57Gq8H49XhwaxFZx6G
WK0FlvXyMDr5sosTzLRrrl7MrD0v/2Jp2JDNlopc7JtM8EO0+EBX4pS9RRPJbj+u
XhdLZNEeYYGAB4gA//bYW9n1PA4z+Jwfn99atDq9PxweVolLyPZrsKLbKCnyQek9
jJRypgI1REIsQTA1tDvS9J5p/++g8eTdm3jvBmZO9X++wkvQIZowjNh12nOmU7Gy
KZHUWL0z7yisGdYug11+8u2pFBxErNuON4v0SH2ZXEY/9Pn6ZTyoscpOYr7O+UTN
kJW3GM0tzq2tjk0mSv5rdOnww28Q8L6b+QVPb9FsukaZMGkp6ce62cfrbikFS4H4
DJ0gDvwMftLkJDMdjOzQ2QfnpHDZxaRUFBgzCHE19KUEsP5yfsm4Src5yfZAULRk
GMeNht1gT5OGo+L0Zb+mm5mrU7GRIXyuM1j30b5TSrY6K1KGpi/oe1WYFGpX05fN
ZANnFp5jHwgTYiyuAgJvylGgX8GSguyEk9HHLFOPDQYAQnDFfbN8YR9qbTbix8/l
0Rc36nrufRGhHu3OXenIRfnU95rCCyMiSOHH9Z80GBPK3leIzNafv7nUeYWSG742
SoVK2GrCD68oLAcjJB++KOCLDY3P1gcpi11vNfCAaHGPkzM+4I7qUuPTbM5LQ7f+
rEBT77ZJwb2/pFHEzY1F/Ho1RLtVnfr5rMJiGVRt55wwVX/NUoU93HT/FsoZh8I0
YVWIdG/LkAB/ir2Nw4sWtXpehOkRnrEToxySMiZVlSoQ/0pAcIe98wuCBtJfa92h
ciXJUX+eOLo4dQEvQ9Q6E+OlLo9fR4sPoT0pTHMCv55p+ectN/nZucuik2YmDpGg
xrWIZwv9q4me3okIHC9AbyFs6MXHbOQCDvpQZIb+/DSbN2x6EIFosHod5KRbj392
A7B6OB/ntHEAGsi/IVG3/Ew3boWTZ5tan1RUZAs7EAIWzc5tTRp/ypxyW5Mf0ynZ
3pcR0opO2UVndWInAXug2g==
`protect END_PROTECTED
