`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
07M1Gt/kv6IOKToaGb3NhJ69Ay8A+7xYBxXrxgifCDNIZmrNGNa98y/hZpCfTXLe
z2FtU3zvufIMnNzGq4MawAQ+gVgIvXsJoQ+if+2VjIaziQecpSzsK82GPgJrMXkl
XLbj/P8CGfHF08m7FK+tKwM0haWD++1D36zBAdaPbuZn2pP0Qe7dfc4TOOcEyU9j
8zbNW9vcfoAxtqodlP9RGp2QzefD3AtmblF/rWUeKgBk1vHXZaOcDBqn4aTaaTS5
1QNWvD4sZZRlrSiDDiPRGjeUV9CiUwOu8f8/y7ctQcNQNJUCFKfbZkvMEe9kkkzP
`protect END_PROTECTED
