`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uANOGTbaPGVD16jqtFzlxt+eeqgLeqAXucOTW0bmjtMkU1dgfwDQM2o/Zi7PJVbr
FiWm5OpqEhIJ7X/lx0W5APAzYbYb6YPa2iREvwv03UxiaILP5mRujfdIo4ZL72Lf
LsVNt1jVH0/jcvN+cFC4sf9RnLikTQbSySX2/ha6ql+hKCDE0ZyqcPjtRHxXefcm
Ssgb7L5H6DCY/TScPD8jPO/qhf33+StAyg0S+qI5sWaT3e8L0YIsk5b62STCfnwC
1dps2wuXSOUlu7oYCxFYjw==
`protect END_PROTECTED
