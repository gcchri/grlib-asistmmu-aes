`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JaqRYcajnCrosxPhMdRlVBp9nfGFUS8A+/WwC4esU4aF+vVS27RneNh1BunSrDEC
ppYJF6k7cS1SG1gBwd/87TlwN32ui4dhZebGW82pK6det1imG0547A/MO8fwt3sx
Nl25isxjaxCuBsGAkk21jj6OBJADcMHDPMltLV/FE9povs6gEGZZigzaObW2R6lx
MUtg3+1s+bqzR83bOu1H4vjnCfHBOq0NalZEDtmOtBL7x+yGkrRB4kk3/gGX+Ww/
Cri+Z1wuCgYLwyhJosoYMgV4AxTMlm2VCnflrqS5Hf4=
`protect END_PROTECTED
