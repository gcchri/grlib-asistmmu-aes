`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l78S5oROjIWZ4DksgpuycO1Djghsrxf6RxsIoSoEISncBmeWHzDydv1ZK9M8MQm5
dRNrTUCmJxq/L5w/sLsmPJNVIDzwAAFIzZ2c33kDoVYEUTN/LL3zuLW4aZatfqdI
ekHJ7uj9ZJnX4xyU3qTrAPt0hdwppFZu6nwR6z7MWjbXJG2Ex3MDkXs1a8y8nzSN
WAOrh1zs2qEi4JE8LYdH4nYRUErA5mT48tN/WTI3j+EHFDLVL0NdnVw25zB8CBt1
mBYh7EXwNQYsFkmmEEWXW3VXxA82hwQ3d2fxSPZcHcsGYnHMfrHa2U5xizLMJKUA
o/YI7QyDCyAAb6Bt5WNEK1WQpVuFxXqk/cjaVTi5KVZ4nA9stnaobic5NpPLXn7x
cchYINBae74vMWhs7mjcck1lT6Aoml0IcChVKzvAbFumq3uwGcnNpHAfk5rAsqS8
`protect END_PROTECTED
