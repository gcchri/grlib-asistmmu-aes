`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wuPCkH0ulpFsKUBi+Di8Q5BF0vbM5lVZhASPOBNrOxvtlunERHzPAI8LiFRTMujq
kxf5NavOUhFFpX38ZIJ5OD/lkfzcdjbYAJrhS5sqvSm8vvDvB4E7RJ3tXYXUOciE
yd41QbhuBM+NhyvQk3bAllMdFjgBL/ObaO652VeFgc8CpFtscPAldGcRwrUtxHtL
BHUix607hnAV/EE5AcJlxXUJxsDWcMrG3M0hsBROr0LgkdcQ0217Lr8h1TVo5I2K
IukkKewWd48S2IC0BDjErUElFIR8n35WLLl3GeBf5RolI4JwSVKVI3gWns+A85fQ
1d7JPfzjaMRM7mo5hdWitg==
`protect END_PROTECTED
