`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
teNc5kMY60AH94x0CUgwzKidH3HAxW/GY1QC04pNMWfNfE+Tw4g/wanFxyyKJ7zu
hBehYWpMWnOKfq1gNmV8plakATsZTNyll5WtOlBpHsKcxP40f5JX85HYEdXzjk66
fYJbJjtxRpV5idFeBTb+gTsxfgywef49uT/U8yvy3lEspaUuyt9JKojXA9PVz0UM
Y59lxLrdzY5H8dFaNyehq0hB1oU4rpopr90s3IbqY2W/L7YYD0FxlICwFX6sUAjZ
4HlfZPsdGc3AVTRfEcRJbKv8krB5R2uqrHGjI5A2eAC0nWUPGdcbG8M4Syvb4vqe
93Pr8NJq/q9Zh7oe1vQOibXT0QxEHlsPNFQj1w0SA3ZaI849um0VRTa5KRChyDJK
dihD5iPmCXkjbTrd3fZbOxFvgudwCs3M/HQNpl28biEg6qO8zMGvkbP2wQvWPRa6
dFHnbZWzocRvEIzapEruMSfIiMpvRhygXpBPKtOEg6/odzaMtxIEPi9+OLkOHto9
f1eJN69FLOkVdti8Ul3FHEdegXS5Rf/nD89gmx/ed2wp0PXJc2tGN99Mp7j0eSPj
OTn/wCPNi1LXslzmvD8WarzUu5qOa7Xd+H+sNVKKQwRr9c1YwfnzAHBku0qOcpRQ
tgIsIZ092/gVb+6Wz/4jTIlFrzkygzT7aAeRyVW67ZzNH1JRDHIA6z4P982RTI5N
7DE25HZP4Tya5O3ZWLgCoS5jVksnjTqORlODEw0Yip0h95q+dDmlWSvZ8BGnaOrq
LFb3LAmAaSwIyzMLouPmPldMAK8VrANfyZbvJi++t0oyN0+FsiQY52X27Vr6W7CJ
ozMFwU35rJCEtcOgKVjj3X9lLj9mfRAbLR+cksxplskrTVG2VO1lle5UkrdQsh6m
0Ip/x7r2xoXvVhgG8ghfxMj8Wg8Jv9PF6hIvr/ifW4lD6DW9uEW7OPigGw3qS1N+
cHCKM9JSGMhyTx9rutHaMXGHdsXlAZcI3IdZvW6Fksy92TYit9PAzmCZcd/WjhoD
eM/9T/2uPruv6fsenFMhLj3yqUQB4DWYbBZSvhcUUVtXTjRaDtxexHCgaQuO9Tv4
RT4xLSsODmMv6px9lkqwX++8RhbAejW5cJwJ5q9ji7RxavKCd3mgWzE0WmoemLRF
i2vXs4NK1uPG3WZ+9+cxdcw4yf279LyfBcMuskY1qBoJTFWhpG5u4Qf4cMj4QkO8
HTVaUUp6EFmcMs2/JFCgwR5p9al/zZtPNdZ524EEw7DRgJyLip6CIUBA5fquNCL8
hpRTW+8gGy6yEE7v8I28GXRBZ7U2Qr/Q9IbZibLJvtG4OeyZIWzvgFmDr2VwiJZZ
8sQcKd2tEdRW4tLijUfreNl5DmMIA2urOItoc4qp6QtzXiwZfwbwdDNkrYG4JKjZ
NMDKXPSPy8zIrTH/73QHwFg9PKmjNYxrz712tTBC9l50EDAuxoMlysYVzzq2259h
3/wB33hTTkOgpjrk2APc0Z1538Q6rBO3z2tMQ+vWCjWFkbKF+9z/kgtNyhceB8Ur
l8JtJ8vBah39BrONeb5aDH6Mi96gN+MTz0HzcxOmP5GIKeN4Qsn1UBGMUInLKmcV
0iZlA0N56VHHB5USnoUwSjp3VHalXbjvWpxzSyRR4uFcmWBR/PPw13uFme6aMGcV
geYk/PnLP/hCj9RSfwsy9NTH3LGRnUVuR2s1kQ2n4p/uFe53G07cqx7cDZ4OpZrd
1HmHirbUG4Y+lWdtXfW6cK6kCTedFT44GoDXgDlezF3btE2BQDJjfrwp0DQ7GXiJ
dXCIS9Yg3fgG1R84/URfGGkCkorm+RD5q+fqHdurdhJNe+1wn0WWfimowZsGYzcw
sY7XDZjGY0zTWL9eOWFIZpxeYc2zO8pVq4H7AWii3ZSJY8hlD/2yMdd+pK7WvIQC
hfRDFXg2WQdBiJ+z2+oP9cHt3X/VxQ4EMzagnTFQgl7i1SXo3hk3LG+kzM3Z3nAy
QyT9TasCVqN4aTrqcOi7xeNhOLon5M89GMs2lsQFBMwNewYTjZ7k443Hts/yFjbE
jG5Vp1CUyCMYwdkj1EcgK+WfBBmWzd9xd2DMo5OOpRSWwICOCFsLZccEtgUML1nt
t/GXSI/eReY+yaV1Pjc5UiSo24octrWbueD3um4M2725CHgR2QLs5V0Texu/xyEw
HumY05ePKXrdjPG48Dkutd0w2jS6/6t7XovwvCFcvESt3Uit8bv1misBCfqnBy2n
Ze4Jz4t9V1Afz+25uBs1+4cMgXrwN10Si9VHmJrs26VXex7UUQM/x9UVVGrGD52y
OPQF1CJDf5xTUA1jdCYkfiAr4rXQU2uM27Guh9lJYNSJuc8k1JeuGtZ/Uc5kQtIl
ROEbamUyeMnOz0Ob/8IVqk3+x1WxWtCkxFAfO6MgKH7nRe6rBLuYm13pZTc2HXNw
HsphZUH9mX89uZ66lU0VJhFNo2SIOvP/w2pJdmVA/tuS0Xg7/61/hd9eNdGXjQXW
tBBIwxBGNWR7LuC0NnGX90+s3dDLedvjzpPsap60c7XFwBmDnGHc9dU3gNbTnxUI
lmvdKbiwDpFspWqGESkzrgRst76Zf/cmjq8EdFnWQu1R9xixmE7FRNjZrvCarL+e
wy5i4zXkgGw7cI+OEWpIKE30xom8j7Uf1G3EQahW4fTyXAXYviAygD7RishVYrFB
2aYmFDLQbZS7q8ypT78eil1Tlt7bRG/LreaoomeRJFntBFwXyJVB6vnelhC0IDUR
VN4oQOLo3AFNR+Rg2t8xjTi1kO8HzI+UxD1xkyk7x+Ojj4xhvt3gvA9yioPQGheX
K4lS1tW+gN7MWMEZgpeZXzpMBXjyuN6Z67vVaV3eNTEL1iBjeSO4GqmSmH3GziBu
BkSL7/FTT4AQRjUHWE0i4trWu423H70IU3mZlfAKMrv14lJznnS8mZe0hGp2DzhQ
jzndn4bnvbJ8ArYJXkHRu95JWECz3OSa2UVK0lIFCPep9BDpDzgdHRYl2R43Gk/R
L9bA5eDWDWSwUIVG00I86AFU9HjV+BASkgeWsLCr4A17u6SGjeWqa5mQ2S2ikBYo
Kr47dusG3eXS8Ztdb6KRXyiBlMkpIGlN1GyehHPrJh7OGEpzfgURsSNS81HvL6sj
1ZaEkAE1AQLAch5bLWrIp73dG+RS4mFDvi3IdSFgyUtn5j6KWZ7ld8VLt36MsAlZ
7oSH+30mHwUUKSCGXJn57/OUIGLr93BsZt5Vjc3tdjdCmHe6k1hoJQf4NI2T7/Pc
0pyjW7JTT56r+T0L2yTdGvXTQ5p40gByDIEKB6VayPG3PY11xV6tNnp6CZC07/t1
9FCaXJhGdQDT7HKW9soPpdZN6fMI0GfuWdOAf69lqoETCvWZ82fB6GNtkP085tUi
Rl296qv5DyfbnfQVI38LZ5/sZ2kj+WlMzuMWISpikJx1jCLzzJYc4I67F6Wl5qOF
PckAmG78WKUKKIFSuNdMIV7xE6y60zJIAhcSD2rG7rmtjQN2jdoWgTrODRRrkbt3
HJD7x0Zt+R+BgOh2+/3M2hYc2eRyfDLQmtodR00diD57oPKBqE65RK42Q6kWGFZA
GVuGzYOoJPMVRS/MGyh+X+ZTNtGk6PctqwF7572ELjXsx2eahjgICflbynFZuVnM
Ee6CmS/w6sNqF96uC35DgVRVyREz7t1GUIlvB4NDBQJRfbDfCBytNQbSj1eZf8S3
f7MYWcGQ41wY1gbDTPYIJLCrQ0qcqYX6tdsikJMxQufnGE/HKKWDhMKROGWF4CjZ
Gi0iaK7z+/wh7KoDOHFjnU8N1p95ZEp5n2BQ/pkd2eT9k5RQ3cbMtqltlMIju9Ev
3ZizFEy5n3jCx/L0AUZMBCqo8sQqwDUc+Tnl/Psl+nd8lwCuWuOcing0R0i63NaM
ZbzFwZVb+f/5zRNF3RxeNnkjLN3WsyzgtICfcFepcn+4Wa87gPDVUaJk/iYjKaOR
kT0kft1K9TTOR67tnzXE29Kc9KpRktja5Q+ZpG6YL1fv3l4OmPWJE1JwhvDGUIyy
LB65M0lueHscXvVEyvZfUG1fgj/v9/F9bMz0D8B/x2lY6WncVy/GGEZvNUCU+lQ6
FmLI1MNBN38et7PjmwV0kRgr2wOiOWUFeTzno33bywJYZNXO0apOOzXi/uDUc0Za
zH1p8H1NBRr01c1HolwGW2VB/Jl+lvI55vK89QQ47S7W7r4zrfPJyVB4YfQ5eB9a
acro6iG4ur/JK8zs8rdiwcZxU/Vr27bfePQ0vLp9GU5VbOk1/CtdUMGUT4fE0uaX
8lI6FEsdm9RKwAyI/yd5q2MrVatNnkV2pyXdK5qQ9mUb87L22AHaQGRAH43p2GDF
Og7zk8Qz30h1TtbUJc+KpY7DGwtP4nGtgPFTTPy1YHXQ/ceYngIuP5MRDTNbc+AK
eQgGP8xr1LtO2L2M0Mz5yZ+wgt3lSUMilJLIKvQNNAmPr5/JlmKFCNE221cFyrAc
016N9pVnsSzB26iLhsg36Ei1IE3babXdJ4aTcX9hhOX9lvxjPgxMg2TuMT8VyDj+
Vt0PLTKXC+puAJqLDSg5ocL56U9WvEzGdxbmHoaR0dOt5lkzP1vsAJa2hb3b+p8f
zA2cOoiK1u7iuNsklP6lmnmVKOo1ZZzYPTm1Fm0L0jtGk1/Uef8i98EeQABU7CtC
jWFJWTS73uhmdJ/K9lNCgKX9sSe/4p8WvPj7nIkbdDQqiqMoFm3SPGv5UBm/f79G
z1WQ2g3lL9gCmz91AZGnpv1Y0HWBM4extFVzb6wNAjfOUd70q92EByPmRmgGlc7s
tgdOsay5vqqqkZPRHueQWrK/PC8XII4QHDEYtnLirym401wSJH8qt9oZgxbJihjT
xnFCij72TIGUOn1vq4G0byqaIgPRyDeN4UIuBx6i1xgiqHNDzIfzjqb+z9YybpXR
gd0cDegusPJiNLVxm6Makydlptl7oMaojO0K8zBGbCYslea9Ty/wt/gw04iqqyF7
zI+wkmyK4UpAPabK/DgHVZsqRAiItlL2PI31Dg3wZevZy27WsdkeU1Q7ZO5s4cng
CgkV27pj1DnH77LEORBWfzEwSCJjT4R57I+V9YuJ/B+zD5iiyvro4qyHdtFkKZiZ
LZBki2hJjA7JsS6MTWHuRWJ3rGWrBPDMsqn5RbCSRJPnZbxkPGb5XMaHragRWJwZ
Y701kQSI31DhBZv06mUZsfJ1uQEkXVcrAKqgg+YqwGMRg/icfV/XJanG0j8ioUC5
cS9yEJVss1je0ER/PadhejhK48TxdE6a0pB/T04EMrgl/8NAD3kkVWdo59I8uthP
iQitd9qTbcFDVoQ8P4xdl4UeMzgr2rfhNsaU+OnIW8n1obhgIxJGBSFaqOGYqwvv
zNxuFog/ikovmGnax2/x74JCYWeklNCH06C1R/8LzUaysvK+nTQI+7sGN/YBNWi9
mVtBjDGjHfumI8JIdmFouatJYDUSQ4ZIVpC6Hm0bixLyuNHiMRGnCcPfVfiABL7f
DO7s2svuBTa+fKFxmoZpk94AJ0LKVpd4SIlIlW1sbmanJ0oIRpFzjtRhh5S27HLS
/4BMqm0NBA3iqGNciMlszepBTYlbce04tFwAq4/soi/PgYT8dSJd8SdOpmvduXRI
KfZYkCaYzP7Yzf9dYwawG2gF840UeJ0Z8f5w0gNwFb79OQF1B4I49MPwkPTM9emq
j76WXIo8dXy46Z922mMZqSFnIBumrTEG/YFsZYpY6fVyrkwvw08Z4Zue9g9QzlbV
heOXZNVABYF5/UPv6/CzZ4h0CmbHFxFtq0VDQ3h3F40gYqn7rpb4paW3mDjLQXgn
O9tCKdl0sWqDAl4KE0zc4r8lEFd2y4r+2cW0+HKJ+9jigC5SKvj9FyFlfUs9uiMC
+gKqG4nqvWJ9EnFrYHgkIXtPu0MPwAXSOtfJvq6kWADWvt+rGSku9Kw5vnhgzoYY
efmesh08yWI4+MLcbqCciCIJmrkmKSS28/UeuyQZBhRvizJYcvyCFZcrxY4l3iqT
yx46yeHtR2wZDpY9Up5RXpTIORqtYL+tOofDppfWf1WAovdVNEGzYpi3ufE62N1a
AyPTM5uBNoA9CNO+dCp7xFXOjj82y4wUIrnpJkRwmhaEhP2z1pOS88YAOEmJj6Rz
NVLzNWrX/DmnPXytjBDwP9oMXTzR2BxZYrRkBAYV3zknPvg5dcxJeTwfKQfVWDbU
nzegxB4gZjnDsP8WV6ZDPPNwlzFfvZw/UP4gydOMzLflH/YUXO+vjXwkGFOeY30S
J7SWO3kCSWvOfarD4J9yAEDpSrGUxr6ao1d9NH6MpPe+hQMehjYtQ975kaz2KOVI
I8ZhJ3oY0xXvewhov50Px5BxesgvcnsbZZJZ3CdvZEbYmRMrT2jkzfydhv1uGPjp
QQFhQZtu9ol6TdTtwbhO23lifHeUqnEpfCWKGcZjQzligJKCY99as1brVM8vusxA
K+VMXgi6o0K/bARUgS0GvEEY/IHSqPaAMVMeLjPzXprxynOB8ZKHcc9kTZPZsRzx
M+GVleMFCGAwh6E7I8jVAyr4LO5DhisO7/+lOAmrXnCCgMoGRWOe2f7TTvZgH3uI
Mp/tBiVmVXWBn7hk17B3oVpEphHbJ+EjLvhsIaOb6zaPAuJXqCV2E1Zg6t23xXIq
woMgfF9H0KEvcyg/U9BD7EckIta8HBqH++E3Tb+Z4LTQFBoSmgFEx8dEHtXwG0qD
Yf01g3xG/sf/w0aJF8O3wMnYg2dIZJRZm6MRSjS0nmqn5E4S9s+gUnrNmLwghRue
BSNflijzFo6Q2F9fUEV1/0c8OJKEJVdnIp76ibB25nZ/Yj6/eUCSOzEbwr/xSDU2
aoIKMFGZ7mJjWs/L1jrxnDFFiuAmEtKgElBO8FAA7MMjRV2LrZLOCySmGRYSOKu2
8rFtP6vW8Cmigp/6c+w58c5IaGxpsXsheAaMUqIAn0eFCIwjZbZrri298SrUpaLZ
Gjt5tpYBO09hSWn0q3yYes16mLr7W7i/j2T8DzTnnZtOojuMoE0/FvhxFLQxvzvP
qW/Arf7IyuOpbvzMoMWJRmSye2EBoNZ0eEWiyIp8ttPT1VQFX8yY28RHZJ1W56pg
QEK8PrG6jAma1S172V/Hpg==
`protect END_PROTECTED
