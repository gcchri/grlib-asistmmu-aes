`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+9IiKqkvpM7voFOqfbtYFvEuLIoUi/R5DuNyKCjwDq7qA1CbpvryNZZslW9lvnef
raQhPItvaX8YDStKXBeFGpKwxv33SCTOcUXDHXQBi+134wWrcrLaBm5EYxeyd9Mq
Kn2S0fXYskFobqEGbUYx4bspEsHIV3lBQqKuI5KomwyUbbwntGJK0ItodLihW0Ez
PRjhncOyN/NQhvzBATbl7QeTEVsco0QNEbkKkr2gg4Zwsx6tHv5l6RPO47zibC6q
4aFNwMJVYQ7rag0JmqiV8w==
`protect END_PROTECTED
