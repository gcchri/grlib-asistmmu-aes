`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
32e5jWewd3U+eSU3/zDBVhrvERDVZWvFo4kMlPacRqz7TD2Ax6yCHHos+NqVBAa2
RIAye/bM823FLK9gzGopfz8Wb5Ewn1/E6KSPAy7tHAX+UUKWBOU6lv2y6cW4zH0I
2w0ouEEFXe3YXN+wFL9cys22aFvHkIlyAJSIsvFWR0QDjKByaev1zAM+TzP4MhHI
KTUtAPGF4zP45zGvTtacmhYCWAH+BXU0cm02V+Po4N1wFFFjNXC7I5zrm4xo+A0N
HPY1eWgHT35lbEIrhPD2s5K39ndy8RqCVgM8k9ll5vFkG4PfYfbnGOj3FIGYWQ7x
BfvY6smTF84yU+LFdhedDHxw2A56ccmRnpDurOVD4NbtYgxRcGcVU4Mb2mQW5NTJ
qn1w7vqqyJJk3DYZ796HJx7oevR0shMPeOAa3gz8qsbQ+0kOoSyWG6C6LB7SqTHe
Pm69W2icdptkjbWTA9OsFladzs3Om2Uz8CZejfuGhxI=
`protect END_PROTECTED
