`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XW2e4WKm6YSeesFU6c59gp7JkGNRRY1J9vWRNX36sUs5r2ejzbAkrWPzRq7ydsFz
RXod0KC1ZZSHNXMUP1wbvPWUBuS6YUts+5mjs+aE6DPbULZ41/n/QZaevEvWvrZS
UJYltklxv7fLMvUWXWrVI8dxYiL6o56u0ibxAStdox6AeyTbj6Dq8Uzm3ZzMLTbq
Bd8e0zUSH5pjPt0T3hq8DW4amiZeoMuKSHlzHDBLv599Pk2ArxYpv6/pBhTZO+M8
Ahnbnklr/385iUuo8+z2kQ==
`protect END_PROTECTED
