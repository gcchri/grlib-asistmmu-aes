`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NRoFzEExmEPxweEd/4g33sqlb9Wrs5k3Sg9uKdPGAyITuofBxDlVV9QTwHkq9TAg
QcHlNy9NW9GrV5/xmhtKmvLqHLRT6d73MPqmfMZyNml2pTpQJmS/DkFi7qHOfD2Z
j9q+nyAnnh8UdPOR+rGNnEjFjYeaahpOM6hgHk+Q0ljSUNdDQxiBNY2Zt+W2U4SW
1TpJdGeT4kB8L/eha3B+bFyA7jopx6hYczi7Xi3c4vUeuiEr6D/Cf2VPt9uKPRkW
uV+f7p/H02lVJdX4fa3uHP511de6CdqZtdPjKLQdAmSiZb/Mmw8bUXX3RZiKUuow
W79Arwn8NIYeoyA+ZciIQPgJ48esYZbvuCS00KgYyPxgriyg/bFCw+eVGQwJ9to8
ds+Bt+N7EPgHeSa4eSHIew==
`protect END_PROTECTED
