`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0q28ckrZBIwiWgGQ3u/jt/ZK277dRI9qtErVJWMPP/P0hh2As1tCbvtgg/XGDeRm
cXd/vGFwkelx/BQSVIPITJIoq599OeqaPUGiS3gvs/YFWFov10nnC59/gTRoKEUe
Jy3NDcbyaujYTwd75Zj1rMlztHBIlhf194KAUFF0ERHIgwuUYzQmlWejLWV3eDm+
z8wDqSBRiwOgkvBmLOLczIc+S2SQdhfVtqpJfTuuUlbt1qkAdz09yInnU9zDw58j
86slZ78rq8UsFRknHaDIH1SoUVk/QX7Vy9Uh9UCXVwrnot8poIPce6wE2fvC5L0u
hqc7Odws+4tJfHrZS8cyeL1Y8FLK13wuyGgC0nMUdDNdIWuVkIqgWXvCm8BqKLoS
ZH69HT3DXWCOKbOoQC8FcEuiOxkTib+SepOzpMFCklxr888G1VY9zd9ywkp59X1U
QTeX61SroQV5TmfgE40IUhtnEZARexvBzkk2d2qb8DkN+2gNcgroCJ3vSTREv0v2
UcskZmvdu2me+wuuZDCZFthWibFF5oN+QHyVWkTLDRFCR7QlLHZcHh6DkUpg1qqB
1y9/JeyjkczwaeA3IQ1RNDASZWoAPh/gyjtDBuQHFvGsrTMv4n0uZgiJcLenqSNG
lD53N4fE96aZ7ccRz26FR4PUm8CE77oWezgWDA1emWBnHy9n+MF1dqIdLkWg35/f
zECxMnav43P9YV/qx5nZNg==
`protect END_PROTECTED
