`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EDSG09OodaBWD+XnkhXz7YC83VNWGdzsqI1VxfaUEqVy0vi8KXfVVaDDQLvqx7fW
upM20TzIJFKCb9XJ1H8gaQlQjPJMJj8P8zmtUofEoph1ZghADhqNntmwGgwjtn9x
yhdceQZVqc7dovH8AR/LjA==
`protect END_PROTECTED
