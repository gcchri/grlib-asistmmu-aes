`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4XeJOfMZikSSWPobXaAxsfF0rvX7mu8qPUowbvbn5e8gQAvAAC9KbH35RDM/FjKg
uw6x0keNbiYSuKwYuSsPVFKrmZCsbQEh/CplQ5Ab5KvCUM6rXkjtCErFFitRliyf
QaFMbBMXs6IEO9hOrgfQGbntkXALZ1Bn4Ft+WvTQwBg5pXEWCUfWx1SnN8/GPFMr
ivEHI1awclbNs4URaaDiDQqBKS/nvyoyKVyzFgHhQiZkco7ksohOKBwQkyG79xuV
1uyl8b5droWTyggbufdOHzmIk5IOgpi1cji/GlC+ZcdZte5yJATp6za2B094HZoe
z59N02nDK5wIzQTV9R4r2N98QjAej4oZGSlw8jb4/qQc5Z02hsSEVFFGl4JRtDIC
5dzD//UGPLxoktpnFTn153K3fvKrNRPeg58+bGBg4wz9L2xhuEjgj4zIB/HlKvEX
V8YgHyw+7l+6Tp/Sts03txqhiMlxWwcijMA4AF1f85HiLZqgTha4kpcrXiC06lqJ
ubQkYPQTmZe7JaAKW/IfXYjzB+Iqk3ymDN0O16zJZSEJ3PulG/tX9aq6eoWAYJ7Q
QQqh+S1QbsZsrFevFf0lG44DMvMYKZFbLIx7yv6BgBZsnWFEygLCC+AEWWMHEsdx
+kiYGyoy9Ufm90HGC6Y5YZvnk/yNgyerEMfB0Fy3D9HEcjl+YLwDtKMvak371ihb
6y25tplGJl7g5wPJiYxmKw==
`protect END_PROTECTED
