`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
njxACd+QqSzr8T+C7wFqMPOHSBkN6FnEt8qtZaREE2PD58iJP9p6+Uq6o7tVCni4
kMnF3/lDtDRQaNmEaBeO9bSW7hsY4LRfNrBtXzRk8kRB1T/dENVryinE3MhO0jue
4FOsS08+8YgJ7Sc1HCx7mdLcb3K1xKmukVSBb88CesERq0GWguJQecUxeI+AELdy
v9a88+/wGZmMYdmBTSXzNSO49ys93bi+ivLJ7lgYOQtDBLDUpCp/dA5TrGfky8y6
r2+Utd3VqfYduHrPsILnPTQP1BixGOhb7ji2+yAeOvuLEQVclUmp6gjPsI2eRHDS
X6bc23wN3ymdY+hgyYyb2+0RMh+1oecDwExL4/AbHzUiXWuMSNcKLszVd9wGyOQb
LWexKNjNLfGi73T7+A8tye6FkMoiFd7o3HsjXdRW4ZmAKR4phZjYSIyWsBbk4Yna
J5OflREMKhry3ONuFhsse8OiCjyAJ+EZeDwBIUVMP+EyHY6vcxpduFu1ROHJbasf
jjvlbloCizPIY3Dhg+wPsuzCFGd1C0/p9c7zLoGNd5wNoAq22LNHDfyCBIkrWNkt
9IzopoG7u2O6vPiPcs4uSaKTeXYcYU2hYItC0So4q/MDnLM4uOW0HRiDcPrbkJKN
/Lx2NM0y/KhsWYaeUzTRmXmaa+1tKA3aWEs9koUUXkLhzFkAhKxU4RUKs7VpUmOI
Vic3MKUeYqikTJ2Kw6U8qEOpyMm2pfP0LWiiy/Fo4WyUPXcVl50faB+k572VvAwF
HkvrnWo8z5P15FPuQeuUjP4UGjb7LCw7doR8tmYHYLL5VhkDdF+++P62z0q0oG+f
hcRNyGr0ud09XKncjQMLsw==
`protect END_PROTECTED
