`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JyDql+/esFSTHn5AtLIWGbC+0vwptZNv8/RWUo65b9x9MzmWAqyrd5HNEWMKxGS1
LJ4mdmcr7b4C55e0F2reJDD6z5Zfdt8eaPrk+i6pvak0JTO0a8cSgn3GGZQ1s2FP
HFqhJvjUZkcuno6c0hLvwioHmKntC2OJcXhSh/91Q6D5g4AjqOYKeOwZFC40HuBg
gWfZjD+UvlP87ZIJxXJcLz6QS4Eec3N3V3+400Ej9jykKDsW/M10x05OiDP/YYxU
8FuGB3knzMviPbxJOF9OCrDgSg7Qdk5IGHI4x5VEEoPTjPsJn8y0pFNHQJKJopk0
q8LRU66Df7zQg5jUKAzgvPkt/bz1jxSVwu1sOj7fDzm1EPMi777CPzDIWy8gU2ZQ
K2Lsdquoc3r42pIYkyWaiFYWpEJ6KWWLADUPZnsuQ5Nw+3rgwPqedELddxuyxGsU
NMrqnv52+7AfXuB/Zf4cQu32QyrmVj760ihiwIaRAo7+E9lxjrY6Wq3ejkc1pUOT
GhEBdnEaSk6Oz5S6E4i+y8O8C0W8yFE2C7dp2b4sShs4+jooSv3jOnR8P2SAEUwX
SC/3toPLDMqr2TFS/xCuZsQBYGo4PJZOTmgLkn+s02Q0kDVYtr6I+6JHzpFy2ta0
4Uisze9GdPiOt4IQzyoC0pAz8ZDlHaJqbkjYlg8ZZ1zHiCu6LhyM8YFvet1hrKLw
KB3eLkIc1a9mK5TY9MVXqXyxFLEEZkSFJK14WYkidKXuZcXfVajgf3vuYGFYOwC5
mClMjWEDe06GUI85wLww3v+R+1uyvWNrF/EPQBBGLecsSSXSMS7juGZPnSmfnufT
imPjtibVVJ1SjqAka+p3i14EKgerzdWJoBDvdxIo52mdmm7LFBCGZLKf5kMMj+Ru
1qaRkpvBHDhhyWQGPFrJ9AqnPzcuQbxCbX3OF7o62tlmP8VcO09KB8cO5BfMveNg
/UCclLRPyvhM8ZASuiFk+Gg55hM34jmueed/ToC+kpIJl/YmSwPAxnJfG8hHy26G
IF1svuRZz/m37rUF7O0IbsIR+8NwuK+9XSGz59DBoBYICbYrTNpI4naF4R4g69rv
f8qsKzsRrl0GpWgy9nEGAi1a3VXa6KKn3c4aw4HdX51MAYU7Gk+2Ju+NYsYxaArr
caL4oQxn7wBu84scg+yLBg==
`protect END_PROTECTED
