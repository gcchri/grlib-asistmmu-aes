`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T3JDjMOihqB/A1l++d24QHFKm5Rx28UUE4oMSX1+XGnaOD4K5yVfkMQqyBpjokOw
OBxswMgnjds4LC/727mHPxubq4fdxx0wBojkPvzSPQgkNlIp82xk3UILBIsJqisV
eAMAP1cXtSqOP6zTqg2GVhtv3a9/4x+WGbn9GFP2zAQzP5HpPeqPDwhHzzXTXVu0
C0/dwEE466qK4a1tqB3byPeS0/TGjfoFzLmMZ+6RvtJ0vZMcepKVjh7vAAwDU6GS
y/cHIEHKiURi4T7qEL3Qxg==
`protect END_PROTECTED
