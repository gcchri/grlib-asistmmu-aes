`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3EcP9g50xSORv0ZEViW93QVHlEOTcOYnIyseZiWQJZrRDqN0xQ+qIBpWhRelH1UB
iV3Cc9qkFJ7/8N3rsAEzAQOOzGy6HnZJX9BR4jK2v12d5STDN0i6KpOIvRZ1e0AL
+aGH9QflcGtFfgaSlZ1e5I+pMAYSjqfOb6xEjXGz2s+7zE7QzpxEFeYlonsCj0S/
R4HeH4kDIB9cktCPooqV67BAoO5ZdM5gmPNMVCujll85EsC/aXzlvz/+jQn8raIS
3M9746UOxy5P9MfbVVePd8eyEFbFaCIK/8/FohMdwdV8E2IUWwyd0HaIGk6Rtd9b
PqjwyhYimh310d0tpGv5YGG37YhqV9TVzdI9Btty0QsjipOO7LQExoItTTO8c0W2
6krYSCMz4r+yB55Ae8XzLryj1kroZDZrcg/Llr2R31E=
`protect END_PROTECTED
