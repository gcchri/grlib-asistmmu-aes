`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uWAT5XiH3hrd5bgUILfZaLKUUQyjdRTvs8vxmIqZcZFAUsE6LIFJLHuxO7hbrk74
hUA1DZSlapTLIKVLaP47ShcxpNeBPirzJrvzASovEALHack3RNr7QvIBQ4U989Fm
ZCxYPZDCgZ967oHRh+9KC+KUXo51PFZmKGuZVwPvxK7LCjyeQW3hD9WJHspPvHF0
aROnNe/t5rHe9EoRjPgS1qiQv06LZfvjc1C9HRANdWeFuX0uOVFiK8A5fz3c6REx
cbB0KD2qlW4TSdhEaJs2XRbvzR0extzdeEAMn0xeMLS/T0+uufUPYsSeUOZm63qf
y0j5k29ROyJka3w+8kGOaPatgXe7OgTyf2Ou6wt3bs3p3kyPVqq4WM49lkEiIcMO
4wXMcPbF5VsvqDJTN9d5+rnQADXeK1HB4zk0uaAzSeVuhGuTjyojZwaocYI+98qO
Wo5qytRcLmjCNn7BgWxkB+orwgYzplR01I+q+v1gCLE=
`protect END_PROTECTED
