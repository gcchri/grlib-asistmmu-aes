`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eS9jRxx0C+xML9w3/S5BWRE99XFjcVLwP5FuaYwgnN3xUL0JHAtoOhR5nHMAmdIt
jr8j8sHWsJSyQYWM2KUs7ienpDsPezgKyBpzTRvDcKafjfBwf8DeNAWnr3fPRx23
xhAOXeSmIMPSpVcLA5n5LeDx6lyECk8yi/OQAH7AMBfISAy29CTwEaVoBMw8xrYH
kjTyg9VEVCNWwnAz0xMnGRrD34QNwRokC2RgdPQ7OSa9gwvTx/AR5u9aCLCOwuFs
LnAA+d9DAy2Wt8SBMjdi6CiKqK31ZMueB6+bMvGVVggSxaOdCqkf19fXFW/SqJnG
hEyFqC2ZuUgdviOgdKqBvFw12abC7efynR2vu88phR4HfDkLlgH1ZbornkacCuwd
pb71evAigXujf/PJOwH6IuJ0N9I/5y5qLEpzNbMU5kCu0w6qVk4PqM32qCFrEc7Z
80FmI0VJbiekFAuDIau32AE0+VgVuxnUDS4U2bZjG32iBc9d6t8wuq5zg7XuD4G7
57LQJrZIFvo9fOGY/akGUe7e2WuJIAXCGJmouhoipdF9yke8YWB+lpeT2SNnxJFG
EjIIudAVwV+7MUYQtjTOayHGlzvLShLaxdjYqERYGgSDmRwGy4qCkV26EGNAbJfA
NyGjRg+CZv8mcbwsGPZhVSSz20WfYAFZP2PKGMdok+vJOKFmteYydr57BHcvQgeB
zXZb9Ei4ybuI0tE99mfY0V7pI4tSyGwxAskMbUZEq4Tf1ylKDp7eAj30sNgFz3yE
sslJ2Uia33eWf0kUEG2J8z8x4lA8l9sJPoD1wH5nTMj+uXUsxC9+8Zg/ROYb93sO
0sSHuJhJd3EIZ6nDVxDFuUjaM/belB4ZDzpQFOrlkR8z3kMGtH9EZTqMr6cCBXtY
hd8RavlMXuQJWUsEC/QGZsdg6EXPjXYyND44zm7L3e8M0y8u0H3p6AfXDs5jthqN
ZJd/smqRQMPbBGono+TwWqW2ILGmUextz265VbRCjpR96wDC+rYRp7D+0QfMQXv7
3rjCr88uumKBBiiVI7iM1MSDR06GD79/U/z7pKs/F3LliU76qg+SESZIK9T1FFfW
Lt9XcM1ubopM4BrECtYimnOSnE/9OSZ3Cn9YyI6FXtWf2lBZyQheKziMuJDashBo
OGC5KOL77o6hHe97H1x550rXGD6h7Amabh1Gb+pPhe9nPAXSalv1zh51iqZsT4K7
D7pRc64Ho2hywoShm0c1actInq+B7I7xvcj0PEaUjV105jAiuM2wVOejCnE2uX3L
hYA2bcEXzvz6l3Fihzf2iyg2Hz26PC/yUrmRWalEW1R+oNWSTgQKWcGXHX8L1G0j
4vmkcU2dzPWHVDxIFvGKu77g5Fi1VfbUAqHn9zr5JJ0UQuQtbYXCbtyxtMD67v+b
9iBIT9ziyy/mXFoaUOn+4zbSuZrTY5Y1qS6NyavosC2SggZbhGkdcpi4z8pJwKhe
W3y33LE9m4nEMXeQA8Efm6exN/8h0hf7Nir01mqEamDHy2x7n1djekOIREQ5q8Pc
eLt2U2rU4rY0G4fwXtLW8pJ+ZiFPv+rTZbxAqA0t2GMFuqXpNIU3yLOQcveHFrLM
C4lOLDEHmJMZ5ZTwUsVX30BpeoKRuqjI8BxW9HoxWb1QgcLpxJdpEbxyt3/R/EuX
P/TRQ9iyyTpNOKllVRtDrD0RI5n3xTNI4v8EfRc612dyPWW0q360wn9DEZzEiAiw
tDCDC3wrI3kKPqSZ1ZAklmtycpkefJAuS8QFt7J5MT9h2vOfygyiJunFtXTPtdiu
vemYDahoVPihaRCxqisrUfPP2bt+NGPOOm76ebhowdieCI2lnL7l0pUOdpfF3HyK
sk/rCuUQWUqi6wWqLrn2O5J5qmBcqprlnrdgvMzDItspUqcCWTou4ydM9dDdLr0a
7FgFZOQGijr8MkK80aq0SijX6m+x0unwq0HgI3biLohJvuPxsqVjXkqQFt94n+35
xArCBZwFOWyov8tEjfydS/b164yz5dfFwaglvX+i06vkliKyTnTMPkkR2ust1T/I
DiKIk1Zi0wJLDumghnf6ytpdMhnIWAHVxoZA6jCScn2219gRnNTAayo6gM0afT0z
ja52KcT1AhigrdYJ+IuKw+ORk19yc0WUVlwX1mAfPA/uN/HmyJctna1V3rxwg2rT
AltQh4XxrmvqaIzJjz8FRN+yBMlBQpYtdTHEyuLLC5bkB17/9YKG032keocyEC7G
1ArW27KUaluUO6oNaJ9SEMpC8nGpvTnujCW5/7Ot5wO+5IN4OInnhdWdkFf81zEt
0vdDnqbHSTlhRMbGjkHPYY2YJDYobqjdlJ6o2r9HKW+1GwEY1pC14jQsWVDsIvZs
TymGx6IOt8L2PDCrshf77TJZ8bZdeQx0azKrvkvqKt8LjsYuEFJzP69wm7yynr2s
ZB+eOPe9mDRxkPVeoEGhj6ySdIKD+3/GRYxKmLQSO771GUb13yYYwOurHlzj4tFc
lPpBC5QWClB8gUDHQqeyfqvmMAd9fSOg+RflUe3S+azUO0cEwogsE4eOQn8T2Vvk
mNgD+xmS+bYuiVoLPvsSmsH1m5ht5GpDKqDq9/UhJJKPKyq7QRPT6dK3HMeJIjll
NMvydsvDsEVWE5JnZANxMg==
`protect END_PROTECTED
