`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qUgNuBk/xcA1p2drTnYZR+9Zeiy0m/f5vmvtzm0z8TIV/1m+mBlGJAE9mif9hsWQ
DOtK8OrmG3cvEXT4g9itrNeprAy55ehzAi6WQckgyh8cr+PgMhGgwSIVEDn37qrP
nyCjYQFoXnzZszvEqPil+76v/dx0mlgR+kiuVnXMGd8PzjzNU803ZBG5YCnZcle4
j9PJKEyXb3Zb6s3XpGP4eIqeFe+tqvtlVFQbftAnfrLUGpGUzcuSKUZ+hYbOyB0T
gEaKaOFvAf2OBJDE2x0DvLsQyJHBRgUCGjkbwqKgfm6b2ae+mf5ysWq1Wmg7Z0l8
AYoDm1B5Vg0FEVwZ1uM9jFPGU1cwqPhFbOs8AaEJVc3KCz6wBlV50hl/fQBCQeNp
NmjeL5zBLqmEku0V/Kh4cSL2Cg45GasMgbgi+G6ibI+sHG3UtZWESUhDKLD6ED97
tUg+NrMXUjVRfxlEb6J5CjFec2czOnudRThjTjywk6IaFO74pxryhDNB7ySENiAR
NXI61Xhw2xGBPsk1RQqtHMTeC7irEoN7MpHdXHbY256UJpO8YzukI7Ru6cdj8m9u
9jRtJpjlGEfB5FV2pjiUMb7ahbfrBgRBfnSQsNHhqADtyyGM8cCvSQmyS6FAfizH
LtEOoq0effJNKz1YduTzFrtUk4aUNkuAg8Rwruq4uuhftoqRzAtezMcQHKR/buyn
O/FSbPxYCllg3wO/PwdmUV7Xy+ulYJ+BbOi3vmTQoiIhYuWdWTKSRBWlSkijiYGP
S0n+UHoBWPpYyadLKSc3rDwbFWGIEOg5o5PDOicBRrDFwgsmJ6lHCpBGm3OFrwpI
sJgAJ9W/aqTNM/YTXCQl/uhb3LCFqc2vjlDxxHqEnndvgu9PfnoMVFn5YwqN87jY
915yEsoCqWlsb3E1Wm1gHZ+uyE0tYmuQ9iqs4cTZhbU2Ja0S3P1U5J4CftgDJxW/
`protect END_PROTECTED
