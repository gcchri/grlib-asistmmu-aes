`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mlzvARpLxIXqjDLV7hCYyTsoHxdNVj6MxcUsTlWLjZgm+YTfkXW7TbzM6v6lKsyq
rVLqf9Iq0PG1FJyfZrx5OACxQI8P73YNNmp3MqmaFXZbOv9Knldyh7z/wlUKn/HM
pgMAJXWG9CLYK1fcJzL4chKeNy7L7OJrgjuajeVkpKzSBwXjIdelX03AsGM3qaza
T68jbb8gjZa9ZcwouBDG2DltmHcsD+/C7d03fz/E9qN1fHuBY0Bk7G3xmMuJuFCV
PnH0MQ3Tccx++F40pAbl+m8CCjC256THj8D8l9y026s=
`protect END_PROTECTED
