`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6gQdbB/GkiGLhca7mg58PVFLboZFgFuD0ybiCcNIu2YieDWPBXf7/bkk7ffVNrP+
RVkQy3PbaD+9i7TX9U8JiU+Wes76XHE4FoyY8sjDIYjtSGnwLYrFTkSkS0K8+M2H
mdJUXsAKP1RHPeFqK6LU7aaB2ZhHAvqgdnbT1euUW77GAdrQVRwPU6Q6RzVaMtQH
lsZjN5iKv11wSONLSfubVYz4Jj/vlQJJ55jHKbAXKLhtdje04mavjU4nNgHErI4k
GQXIiyRMjilOKui8cpPC7gtyExnT+JSn8FhPnaKnBZVzIfEVIQECpQW7l5SFzHJP
Qc4LfMU079xHo2Yu3Jg4dQm0TCDsl29GzqAEbjqdyBLuvNi8c5P+DKQRtTEIPaF8
8fn0DIUQrqX+qPaiZsApVya+KloJ/ii0Q9y0swZDjqu7dJTQk8TR67tnn4BWRlnl
PkF+CGGI2FvLJbtIn7zAX50ecxUsOKV0W1oy9xk9fmZ7soeDjrPSCv7ksyr61SHV
GE+kC0Rh9cqf5To14tCBC+5ti8QIK9414fw8c7poWHeeOru5Fyp6mIEG8rPcem0M
IiCvPtK9Na5/DU0vHeEF8R8aA+cQRGv0xJxzzwJa+769v2fTv5+jIGSFRWkqSnTm
F6VX29PwkiT2IgkPq3klVbEuv9ZBOkaynYxJjt0lViUqutJ9kwW0MwCOtRO+C0LK
6MA5psNoCQVC4ZCfnGL98yC40pg0YMzEckA8/Nur5AclAO1iHP0Eqzu6e4DuMl6W
eyUyIamn0Vp58pEmA+Kaw/FCVWEP7ou1icYb1j+/aR2haQCY5aPSH21u2AZaDdNh
o1QrLvF4qIc0CV+pVD1TTb5BU5146731Ja5CTTkAtvw8nVUMIBnS0KJUfnXa/dt0
0rw3MpjPBCYh4FidW4x9VpTTkyBHBdh9MrBlSCW6u1voJ//ZC4yxnbFhvKd9hTIy
`protect END_PROTECTED
