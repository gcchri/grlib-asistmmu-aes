`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F2FPlXoZ9WbcCBrBMpXG12dkFhdQ54kMhoV7NDoZ24OyCpUxVNnBk4RsqfFwLJL/
BiAnwYa5v0y8UdmUkLS060g+tcA+kob0voVIiJ4Z30y3qnoLx5xW8CTKdFL3mhP+
dn7PRi6CpwIm2a9LjL6Gjxt7hS5nKg7D0B/q09nTkbsSFMaX/gwAd0MLXr6+atzV
laJBueen20yH+yTI3jEec1NDKiTwT7p+mMD1bCkujxSm6+Iaq7SEdEUZyWEdWQgt
VdgGhKWDMlVpVZdYeLJscVVaQou4PlpeOY5+Qtrz9U+wz61Hm9m+xWoA9Lff800s
7MZoqo6/fsJsdc5uzENcY3l4PG0yk5mCbLeIjkj/2Sxvvsk8165DnJ/w60e6lDsZ
FL8s6fCk39QQYL5KUmpICIhzf7IM4tVWbOOTDnHvh5wkim3SOADgaFSWdBrT/Lp7
r2H3k+8Q9qB64vhc/57jh9G6FuL6P86NHu/2FHtNemagm0eWS25LDcq/47xHPBQb
Ey1pjQnZ+zi3alWmZdTjLgE9SyWtBdzHVR/6oe8qmGdArHvsWujT4NqxvBW90U/H
6YTVXdBn/ArjYhMdbP0EP4dlOkR0CjpibAU/hf3aeFEIcMJ4EFFFCtEhrI9v7XMq
qEuKGM6gx2xcUJPv0grq8+KiRz7wRCvoUw/1DBu+ZkCCcuh9/D076PHib+9aznbz
WIiMpyvhtmkP5Cxk8EJq7WvA2uWYi+WGASDuw/UU+5a2jRjxLIr2B+uTF8SvEP3B
Q/KCD3cenaA0sBTboCnIBLx6bq8QI53Y/i+KrgMXh7ud6Nj9scCS8KpJtvnFN6Q2
`protect END_PROTECTED
