`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PKMchb6OMdpPRPMb8jAesM6NJYuSBMQ4ojW6+Dvu8/x3L5z5cRvD2jcCPaWheqxu
dn4jp27f2TYvSImqhFc0VfPHrrIMWLYn9laFtR3YU8DEaAHY+R1FHSYvSIPe1wiH
pXOsXT8i/Nc7CFQJWuKw4H9FdhxewXovuebiWqGuiRgGRSFohJj71z1ZywvH6OMF
DVmAmgzm6weSilWPX4M0bdh5uMyBQnGIU+e6nX5IFy/heZOUsj9wqQ3YLbN7NbqH
CwLcPcFC0U1BfisjSzs34Sy3D6BvUQkjjP9M8Diy0eEIbLm4aSjevlye/utUI7Mf
`protect END_PROTECTED
