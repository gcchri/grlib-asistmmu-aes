`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3TXpeGHTGLIE+G1/x+eh/5Iv8astlLIjZEVHhhjC/AAttG1A17lMwwsDvubTbv7U
BWXx9ixOkd82oNd266JrLCOkm41Fr+BNMtqcQBMBquJwXIv4JOeYb6YtYqTYC37X
h2bLJWFHf9yTUX/FYZWVzMtNOLXkcaeMNESlNh+sq82rAQcHSRkKexma8e2SJvw2
bLOn1R6Kjbz/qp/8sL+zkMuTwW+iFwNPdTfTBrnKgZ/IXL2NSVYX4SNNj78cddt7
02nJdwV1k4IGzVZFC0ccXE3yt1/iY9H11Wxd9a7Nf2/uSi/DpOimPvAn5A4VFEGE
QB8TLhJaNteQfjdVn3frwqYKHv6yuxw7At6YtDfDVCkk7EaMUYyqN0Q2tNrLSAZL
kZs1NT1vy+YYvifZtP9D5WENiAA+WCy3UffQw8WvrNE=
`protect END_PROTECTED
