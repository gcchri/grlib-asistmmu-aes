`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2EIBSUOdooVnylC6vRmUCn6iIqEtwd7qBuF/QUBARKp5gebwZnNuD46yzLieC8eJ
5uXmb5F3EFT9sMgYjYrmqeS0wbTlgVk3NXt7o42Lz1n8kmBNkFz0AaTk2rydhqX4
8uBeKFrruo56BmbpvE6+e0064g94G1CtrCuE+Iuq1gbkntcn573cEsS7wUhUGhud
5j1tm5jDlWYCTMWYTYz9yq/p9iWRLAB1WjdZdpiHEstciyvb/DstoZ1GZhjfG8C5
zDfSIcpUl4jpk+Fn/2vlEUcVNU6RKnGamQOmHAp+wi8RZdNV9jpXt5PO3BwkAWaT
JcGsO//QgB37YT9kTbltdX62si9szlW8R0EbWzWZ4DkavS17dovIBau8vzx/RqL7
qn1jEamtvq98krA1EYGBy//I5npwKTO0o3IgPuTnJppz2uDKCCDOLRbQdFRw2bOw
DLNybpfd6Tx0K0lLhv9AeOvoE9nTLsaCEImMeJia5UfhSHM6EXmX3mkmekzaXH8o
zo6cxq45m1mmdj2KHi1JEvpx8ItgPNNKyeyYabZvhXxiEd5uTYzR2neaAPpPIwoh
`protect END_PROTECTED
