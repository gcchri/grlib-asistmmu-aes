`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sN0adtsdZsJOM5mAVIzd+BPAk9d4h03OXBlzU7QT1DTbXELzPKlSjALc1U6HosAT
rkEVhpL3C0M8ABGEMMvhwZ/JsGObsKRcKyheTxWajRdtCU5Ld3OeMLjvZ4SITqpz
9XKRLfDfAmgbseLSrGAR36MgLBlKlnU7++zLejuyEuc43VXdheiPIygaTBLqaCBR
ko/CUsYTXwHlChnwPao3bDwJXSo/WtF8U/F6SAOnR18/AOgIDmvyLol6tqyQZaHF
NDR6v/2GcfiJHOIOKtQVYjMaJaSbRiAgbzfmOAEN9TPMAcPpTNH11gH55E41ijGu
M5C9wAhBKen0xdzbtdn0fd4m7M+ugRx2DUeYcJKgk+1k/SyXwvJ6cm7zScu2hWBt
+mun0577Yu6OzRrgICYCgR8tErpkEyFE5P0eIZLVmtz9GDTU4aRU+87xSkXSwykj
`protect END_PROTECTED
