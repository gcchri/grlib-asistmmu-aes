`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1+nIvKhCXPGzVBu/DNW3lebHhBjUkPX7eGzp8QJcerC48VZR6oUysMphldJDvsTQ
RVq+Tx9eYThkLf07DgwNZAUxz3hDHfxWl+WU/t3Voc/Z+toca6fjnG8WvOhUceHv
ZaqSZXpdJ++rVUaEXVRsiy3tUY8I/Mimx97txJvj3/8/IbrTt68KAq9A4+VXzXIW
cIwoIcKtuYEbOdaSK9BHYr3C7ThuOdfxcGjOBAhbB5qaT6lnFq5a1VwZsaNQH+MO
9EzvGCgUYl0eSQvjHrQY+g==
`protect END_PROTECTED
