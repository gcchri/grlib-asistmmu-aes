`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tmy2NdKkbLHNX5OUceUj6NFqm7ugc38bs7Lz7wPkuX/omoDMS3vtLv+pbwLCQtzV
3gK0XiZIqejQB34DNs/01gxfwFMuqYDB2ZLJGx0AexumEmfvy6901fkXCNMppZ4Q
IeHHgNNI4CKHiLlrp1c1vv4sDoJQN2laihPFyutHv1ObxOqzXFMC/XDnVR3tHJ0x
TLLypm1CQa343d9xIZ8Kn4MU0gfVrB2D+wp2Ksb8e/0ueXXtoLt2jTNWuFtFMVY1
twmU8fuG/B6MazHAfRBFd8qtmVFgdLKlhA5cAECjXvs=
`protect END_PROTECTED
