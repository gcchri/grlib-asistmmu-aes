`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GqYdlLXwU4Wtqv///5PgcieOLZIxmzBE1+7N9ABILjqTJY2bkStehHeTY/TSa57r
n1pFvM2AvmHUm3s+lQ/Rx9Nk7gegTU3CIRm7vPDXSF6RWzAyD/WH+t9F/Yc4Z0EL
GTF/F5ltSqgQp4hDXqaKaOgd9VbLoE58McaO95iJckD5BFvBgdOct9rDET0uC1hi
N8VzSXcoAavwIvsFwCLDT1FQdaykQ+xbU6ehiRg+A3Y9ZjszCNRL+kUCI/ihmmfK
JPQS44xn2ERcwqFjgan9Xjwm689LDjNn1Cv8Vu7rXlLWxo1Hz+w8bXw6hs7ci2l1
HmErIEzEoF1wmND4MvyCT8RAq8egPyU0AQr5jAFSN4JyoDM0eXOrBI+VMJ+Q7Zjd
e8OPw/U+0W0EYThrtqpqLSV+od/kPoPfvuCWmPOBbcL291vssXM6Y9WFPXm73lgR
FxODDigK/qWPCeLAhVYxY6KfCn22gYOJrnQ5wbPyvpaSGpjgXTl/d6M96uSDbsU1
oFcAhpEtbE1o7hi+e2vkvEb/Ua0EODwFzqNQJxypKktpKgwDOWA4wRrf3BE7SJs2
hQHvhbUNopG2ER1AIq85wwOn9pATVPOtQhrzDcsphs6a6bfvX6xapkao92ABBbfY
XKRxVuZCztgbGP+k0uFTgUWfRLYILQ3MOJTO+bmD+IyOt+nCjZb5frjXUn8Zquow
PmoUHqYwxUdjM5LimSp1EJn8FDuF48HpLJ5TEhPEnqMJfC0XzTxwTbBUllj6pNG/
8kAAJOpmeGFqweEgt3TUcmlcHmJnPWhu+ROFcB9RgionMTcQm7CJEknSQgP7HSF8
KcUMBasofdcaYtcPoGDDZg==
`protect END_PROTECTED
