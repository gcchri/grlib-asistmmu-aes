`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mIpC82qu6cXCh/s0XKLTxcbddVePpbDyF3Q7NndLh3R6bwMDdFsBnh8/NL8d6ogG
w2zm9NZvMRUF28P1KTMB8UOU2xJkydLvSwXDtrPqu/zqHdXJdR1z2glVRHMEukRz
QRNQDhXuKvaFCQzih2I5mwNdXF2VFv3QbffWTE8JeoX7A5SgpdrFa7L1Gd4phgT6
xCGHhoypT1oQc6NIHbtaZCgF97jcRJRkqWFQ7orEYEMBu/KQCHQ8ZZTIhuIQ1PxG
xHr4IFuOw+YZQo7f6PceL4luI3Rn1PVUeHoDgR+eekMpqsTFE7sllUL9VliBh2o5
NHO42lwVAW3QmdaTXBcVZTFYPkUoFDqhjj0zPiHK9IQ2YhikMGEy9CP3MKBcjEK2
3OM+Op2XlLP6MucMaDhN2DB4kJHljg5Yd8UJRhbRK9/DIhhhYM68jG8lyXmGF378
JMEzBeFfuw1k2aUYFOqsshis0D87NFknj9s+L4GoY3PFTOZlPEpExvdnG6wiy+eX
QT4S5eh9eRbUqpOMLio1xgbIJSSR/s3PVssKZzCxnZRNcD+45jvHOIzL0PPzKqmn
U7/WHwufL++UW7QY8d05cgYEjcLtQzwvwqqvxybYZ/vu/JnlIzwRD6d+wu6C4zgg
BpMQaeMRuCUEJNn74aeKfh9/sIOISl3x1FT9+Z2tc/ej56TqorUl2bh3/w4z5BIM
LfPRXbampqfoUy333zZi4GoAtpHFwgsk3kN2PJVSfYefkebWB5K9PBnJLyazSkWr
0o8TnKwzSwgdoydmvU4EUk+E1Y9eZfkMUrVp0PNp0HOPFz7xMCPMdhC9Mm2bwp54
7s5T+h/dMymhucXZgN3hulIeGaMNZnpGxklwc6nFXjts5RwO3tbDuJGe4YtxYDYC
ptrMxXt5qC6irCLMGowl2dvgmp0GiRUYsTmDgNnG6fxuPxDUX/X3KEioSnWfqXum
pZox4piizHEvuF3qCh4uNXrtaHg/UktdllT/VNjfrzXykXIqgg19Ou7dZsCuF2y3
ZQ2TCsAyqzkX8BCo//LkMtgZ42acpboYt0G9gyDBoVGJ8Xlq29rEEW8fUBlMAdtP
7q6pYOqwhry3ylRg9ScZspvLFB+f1fKbhxz2QrR1PkVI5mnZZ/8r8ZM+GgpD2Z4w
RwY9J1QSsaYIgttHAQeexIC5emOuviAJsXiWxMPTfsELrGgbbSzEktlaXx7no/Ru
rlsNDdSNLuELYCTtJavwN1Q8qBd2E5PnzyENNk2wWSOQsQtCUY4PvfiUpYnQzt5z
eACruyAKU9F6SKT0qrExVTENqIvgDeovIPTxm/OCZemPrJNhOTeLhl6DemXRCW0/
nNsp7ix5+Kjs7AdLoe28h4drcDRyJaw8qCgCdHYk7mNWs0Yge8Mf2BYViw8FrcxH
vY2AJ9jvn0CHSwbbpbRUO0M9hTfwiyVabcJC6z7ZKsKcp7LeQK1sNQMMYRLTFrhI
btzpe2g2TmoWlRKBcad+EsMsQXmxnLhZMVzm1Zq127DJ0tUsE3kg2OUv4fzhChXt
BxHT9R4QeO7uNuIn+SiFV9nGW+qL4BBXv2lXhsQuvQRtqeawF65eNrMsbFOR3Cet
Rf2dtvwSB8Jbc7irl+5FTlkHFL1kM1mN0Zp7B6edB9Y9zdSvoIsqYdpfQZcMR2SS
TMffVWh/fIKKXgEL2rumEDt3QLVJjAm7jcgapJby/p9KIdd4gy/hr0vzZfeP8iOj
iKGzuiNqsxl4q4hyzcDYJ39ljMNabKiqMjATtttc5pzsaSaoTEiG0Wmb3u1NveKw
nsNN+OaydxDAUJ+0F60NsxDBRvbz7bcLj91Bt3KqkVZEVJkaiwfb2Ezn3wp7gTaC
Z+wTivgN3G6Ei9qVwwstQly5PFXPWbMHWKD5EOH/i6rjnLspgq1vIn5B5Xnj7BFM
UJB5nzlTtmM1U6O/lZCrTGtvzgCTahVHrEYOJdfbytKxG3iSufw4gFOUqzYmUZa8
o5zZFzXXRyx4Ug76KGDYonmK7X2koE8b7LVGd3Z82QpcFng//5/a1rSVYTXQ65Pj
yODnFl1Dd/hCr68/zc6URJn7w9OUGUWy4wqIyNCHVvhkenwCpGvhgo18cNFRoJGe
yDMqtyDJLfOhryk0vVrp1jk437UgInMJ0B4usxzIVJWbjM8w5YFZ8qts3KTl11ZJ
4o7T0SCpAz5dCKKXG47MMo1QJB8JaG4KPpD8OdcWVOT+aJGGHfG19qE32ri6N/mn
lLUJh3k9XCCoP6KJY80MCw2UdqmJd6S78xU7RBK2l1luKxdVPwR5D2QH+4VcbEQ5
KqNsK+CMMs3y0x33ZDyCjg==
`protect END_PROTECTED
