`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TTKfFq8BbeR20srvESfaG9Zjn3Q9OSJri4faQ2n948J1Jl/gol1PPtwizWVsQylW
w4J71FLop17Xoy/Nfwq4a2t/JH6qaUM5MXE5jtwJuk/P3vcJja4By3KmspB/lirA
G89QP4CctMM2fDSvjfTJWv3w2WtKQoZJkfPEgO+1sa+9A4pkde6C7pYZqhnSxxMm
OVpaav3P9r+MU9s80e8D61sZmBADyYZuynYR26XqEjv7lBBAHsOzk3oHvyUamMG9
2rHXU119lZVEuwzB4xGsU51ypGhwLhbRwG3zzEw0MTrdZHrG5hw9HR0XtngvGZdu
+Q6DjR+/92W/XpGPjr9N81Wu0YCvvkO2UcKYIBoWZmCSTY2kbLUttIyLrKZlloke
2ufu0iLEW9fvFWjJYehFJROmPiZRx0pL1konCPE/Gz116J3bBI0eC1Haj/sybnhO
`protect END_PROTECTED
