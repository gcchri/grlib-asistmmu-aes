`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bioZZkL5ksTEf7M35t9HLEGbj4HgiZKtnUyvKH3Ei7rrG00onQc2VOiSCVip9Y5R
D+11rAwXnxh5T3xa6YQra7P/92M6sWBOK4k4nq/sS9pnP/3Jk+sO2lw1qWxlyxNz
Vg7NlE3p47nwVqNwFRvbs2gKc98vJrBhROEDrXqaqgUaZzsTBT5wGhLmp/lrQv0j
2Xrh8r+rnQAm9x0rnFfgldVwGyTbhtAxpmlu/LmtnD2IamTE2mEKdaohrk34z3si
`protect END_PROTECTED
