`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TEsj9wU8W/hupfT1PtLI7QRZ4WmQdQt2rnHEiDrqoBpgdYWBEmvTmiLx8HglnTzu
yDKj2Qjy8Jb3/R664imP9JYgrDCgPJHenI8sYipoD7uqmNVYFOlzPt/oKYD8PaBJ
iGep+p65V1shzigWszViacZd0GyVP0ALAE/MfeQnDiX1hFvQuvFAG5Pbss1Xs5zp
tyDzGxYSgViENjq8k9xe855KxpxEQPMupTI7CvgWHUUrSBwzKtiYwoxWlEPvO7Pt
6ep6PrtWnyP+SYXS9ZTj+XMVyaNVE609lqYSTzAOEhzcuMH9G0hqZWS/7PeI/KF5
CqXs2dhfhWxCkmT8jTmPoiToSMcv9MUs5q+KFmJDoq4aE7TtYKuX9uefooVqsJdn
C62BOlc8XeVE17BEbSjPHhgT90B8eke7nse11eaS1HlI2wR/1+wfYTjaUJwszdpL
S64rS57jOZ3FCcoZQq/bsKHsby0+5mWlrE+lcAhk94QUzJTjSvNC++GxmwF+/dcl
HrCQbkTNLbRuMPQFBGZ0I1tMSotfMmBpI5LJKalVCcvjrttO+VDszN+ELqbPxUSm
7HyiYhS9H0qFycPdcYU91238l0JFq7oZotGIjBK6foSkwzwTyl5H5vYBQsRS/YVA
0AUabfa9k7NzMFzy1yOpz+UOlgzU7lSDP5mKgQrN3V9ZVSNN9U3+m+zZtgTzCfLe
6I/hkE2fH1TKeXSgVBvUfUv8hBIvpCbxkX0eehHTiW/G9H5L398f8qTcROJzMZRY
xKw7cOp17QrXfqfwkhXBdkhMBmZI9/pibgF7u6KWZxgZv7S37hwGjC9poviNklWy
bzhY18nYheTPd55rcaGBg7NecL4DxMUOGuxitMOXisdi224hA4Osvjzr6F4MX7Mm
K8PcVdx7kfKgycME096t5EMJkqBvkW6XGrELQ1x8MvZrRw3wlDU0T4mvDSOBqPmP
2rMJfMEBq1UcNNGBHQPs0acVMaok7V3Q8MfltgyMw2lZLepdMvGG6RBUuiej+9Tl
H+2ad/Dx7Rdlah3HbyGu+lwjQ9d9ZIE0OMmbtdsIddSdAfHILn13VKwCClEZJMUB
9HAixNlKQrtrDv4ecgq65w==
`protect END_PROTECTED
