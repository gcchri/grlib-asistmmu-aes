`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qhBsOSb3lnKXluJviFJrsKq2cOS9WFXXDsERDpwQmQFsetVlpbWldhGVfiW2fTLO
Z2WEHU55Xoz7n3Gtw71Pe0kwDfO3atJGuVhwOCBjINtElBO08PvW8W493IKCnqwZ
/bz/3vPHlRmwcUMZNY3B1h2+bGz6+ViSJOkAygD67JYYxHl68SCVCI5c/X27f0Mt
YOyRaqmOUnwWaH0latDzvTrKWgA7WEHgSphXtt/GjdKTphlOs3Ana9Sn5PMv15mJ
/fW6m4Js7MD4/un/Prq1mD2PjeV4opX6fdWDHxbtqL6EX8SH9l8t2qvswzf0BzTG
DYWe8E15WOiOGynmgVI5GUH5PM2VjWcKPlI3kkD+5lGwTR/gV8FV50Fu6pP6xXAA
DVzHhX8hcK884yUY7/Ms85Y/uLHkbtlRqENM8K6QUjqjxTItKUqWjOFjNxA2BSik
MBoJwWX7lLzi5eZaIafWp031JGDJSnJyuyKII3nsJ+U=
`protect END_PROTECTED
