`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YPyWf9Vf08KJnW9zr4jyIa4VSpd4lxecu13z6rfamo0GVGD/hWgG4Ul4hod/V/go
XyiENqh4lML0Lw34rOBH2PucbwS6BCM4EnG5RcMNw9gZLIzW+Hnf/jE48sR/2f0m
G1BZ9W/rYhDQMx36VdLdkQjYmH6nsUSqEZpm3bapqwkLP5246PJc0eaHMlZzUQ/S
6GPOYsJ4OZaM8JPcR6a9JoSnPiOO/BD5zqPNDcqSd3k66HQbntSUkW70NkmWt2Np
nX6hHekTdCREnZbUHoqhyHKXDG+tsD2H0k6EUCIN3+1nc6CgspydrEVvzfKqATaj
zO0aHQUnNRvzxsPOF5dH+0Y/y7aZwmVuRBPzt9Gnoec9OSAvUi612VaW1eQ4ozh3
QGdx9zXwpEvgYT+Z6Nlemhk8mNLwCrTiLICdn2HFJ+nFQgd3fHGbyLqbri6YpzXz
j8UWMBHUyf1ujIAEq3BzRC43lKGDMT3YVNuJYR8Vfx37Y3wTyPMDSPvdfooBytDO
dKTX9SGr9v8Lx+L4HNB3hP/eFGXJO3P09PSuxk7McWJTMdanUZNcVfKy9Vhe121J
CvQEKL9SDAdVRgsrUSJKEP0s4bb3rHOnmloZ9LpHl5n2HZOJJ73zpDUyvz9i+ugt
xrwW5+uziEMkBItb0dliLOeiWAqZULuFVjATbiaIFlITPAGTCYKTN07Yy5JMfvT3
BdN0sXJ7OW1+fAmZWq9H1GM1kUf7iPb+xmCia2kmctv/Vc5Py9WRsuRTslSN0ePm
A/dILrqj1bkgSZYrMWEpJlTVVt17EJRcWYJIhfowYhrCwbKml9iM+tKMbO/Yymbd
+50MjfVUmcuTOtPiyyzDAyuwguh4x7cq+zWK+76X+aX5iIbHkZ9QU/zNdgGaigFc
7FsDbSEKUTEK0+d+zv1mI/K7OcMtL9ABsJqLtCtEcpTpY6T3uH0XA72vDNi6h3oH
pdCOpes21pNeSGLMnalWlloqdwD4HcOblt3xxWAfSIfk/o7HDGePmujyza7h4El5
BGxZbkU46obA7f5FT9zjYePqrgTOUjcnIgWl0pGSqBIeLB+8vbYqhbtAm3WpvclP
6fO7Aj16vYAx2I+xb9akPO1yKrYdH56e1rAtrEjZm4tXYBL7jRQMCrLRkScgvvTL
sy0pU4H4pcCZumtq8NukQ9Ya5Th8b5M3voPbFET7/VJdN9xJ1MGJlR1jHjE+urMW
Dv68ELb8MsijqDWYXggIezpFJvdakCtXdaUY62mn+YKylvDyjgWBtkJTz7ugSEKF
SYZlhXU66x1MQuhDOy8sayDfI0GpeXEdp256z2EvDFlR7jMwbu+p9brhzpd6DuiU
IkR6WTIZV+24t+m73p8vel0mccdji+vIWqUTRUJIq5MQGq+APM/GKpTTywqP40/A
mgqRHXwIiF7x6Y0G7ET+qHvZghbFGXEYgPaln2LBKFx9D9+dNz4kBcYKzI8V3dOE
6fib00105ATZYcRf+Wyk34bub+Ku7wZeSOIH8h+KLBcwMT2kBEX9Xsnbswr2EyvL
sMtbklq84KgDTcc2d34rkDuTJ5BrMoVzeP5bk6nnxMhyCTgyxFWlCmRjt+ppBHqc
3RpWBu9kdn+/P4hU/JAvNhEU4io+VWPafqdIDV9z7n0xfZLYaLiIbRgAxzW9NfTh
nPOaHSiPanZFFIFthQIlMungtGoRVGs9F1+eaHAMWISxhAssY2r0ubVPIdXErRDY
2emDXsbvEjNLp8VLxVgjA1oNUjd+G9wL5BnIANOhhSJ95aORxvZcsE8dtda4VvXx
DGgjvLn6GaOyEvAMIUFgoPjkVXm7Wk6xRrUERtH3BlSwIvgMt9UqaGegVvPpM2A4
DwEkEB41qPR4O0IRBnjqi5rwEDZW5ZIXu+0D5uzUgFWBsxK9l20Kv8WjS0MpvKDf
CRi6HP5iyHBBZ3EPXgFXD0r+cyFDHyfliexWsGXkFocwzOcUqlHwJho6B8LbDr0q
8TiS0WNDK75rkqcJY6KgxXj2XhNuNUuxSsp+VQZKJfASjBAOth+rpafKK+ebSu4I
2mdzZ7xEL1HmvQKkqL49jgjPNH6n00hTv2p048MGeP+g+FuULXqclh60EFreZjyz
LxymGMS552jl79xoPbLG883RtN71JOZxs0Wf7pEDxahnl/jDuLvgsLsqSWQgex+a
eYwWM+zF8njG8cTCphZ+XK42Oi0QrjdzxlB1nQ2AIUJfIEVKXXDnqsP5T2X/aLuw
CIlNSVIgUxNvfupSJZCZ6ThRcZHsFs5kEBR+uqGeSUU=
`protect END_PROTECTED
