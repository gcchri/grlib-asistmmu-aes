`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rb5ppTjO+mmnFMSjgy5NznUadWocr+ZeVvBTKMxU0T3gPDTOFcD+UCvJbNrlgw0U
64+NXDpHtOm3LFhueVxJEaWMA8MfmviS1NW7Z5WRjDkjBGT7uGfnreOYFhantDql
vENbi6xeNbGkxPGyLhC+yaVBCqw3GrdP5xYtkQ2aYHqkQsh4KyeME7NGEo7xKACD
fG3/d0UeLRvYT0tXpOlfUlrLbLT6rIF1XEopTK+XjDV0tpQRa6PBKPuye7reNFUJ
yTlf5U+Xq39v4Z2dHUOIcv0OCPqBP8IglrCdmqyF1MG+OgGzFrMTo7MWYIGXTXl3
V5WDgjfo3C9cS5jaQUsBFWg95mzGpNH664sFoHcj5ulDTG24J0MichqWCuxietq9
pG+9ky4EijZKTLA9z6gcMZ1+mcDs9o4/kY8ikq+9dhYvccgC83n+b5ZpqVQLNSPE
xrvOruF4Cc1ONOnPXQh3sVZep1rum/j4RWHKNMRldMFPdkGGHNrxZq+b6ky+2Gqq
hG+xOUK6eOKg/1FDvaRrGy1XvZLnj5c48iOOLZ290XIyzVW6yPFpaDLNN1U2odaG
VX36KKTc51lZbaZ1QaeDbkvymxbk1f1v2Ir6SMsJ7PVKiwoipxjbvPQg7PBTwlID
khbkD5n/Mf8gq+VZyFmvdlYRYeQGW5BvTeKTlvyo88E/pXzSK8fOGrm6yyRAwdwe
ol24smdJGtMONWgIhkcGEs/me6Z9DFbPaDpFZ81MuP8h3NaRHuNF3wRc7MzyWkCT
F6apjfpgpEJF+b4GL6mfIQ==
`protect END_PROTECTED
