`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1rzQpE8qaQj/DJbdISuSqCK5OkZjG8PpxHe0O1zAszRPvXNUg0JjshRo5FlDijcT
pItcUWYr53l+LucmAxp4xOHBGA9Z8eVzC7llpWm4jXV/bFvYxgFX3GK1farnh6u3
3hjFzcsbFSZTh1tbefcYpqnM9hE+EMN6k2Hhyi3RPL4KFG0epfXz+az8b4xn9F22
2GVG2J3Nka7GFHEB+QPANErelXn+W/M/JSMgZh+YgzgKL/2oDBv3S1k58qoz+a1w
dCCXmu6OHf2J1pqWd0hTj9VTZtDaw4rZguNRWCbsQaPd/W3fRMuef5FnPFcBCYt+
3km0n9qCyg7aN9yVXK8QsEGTl7fzKerQTtfOq9X0K40+OvNu1n2S/RVWVh0qBwGo
`protect END_PROTECTED
