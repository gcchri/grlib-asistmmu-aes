`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s4FZuZefmPSaTeY+duXIAaLePVAIs1rg3d9RZoxCdQ5THJ1kaPv25gFfdYMJecKa
6g5siTVGeNMv2cgmGWSwpu5FcCyS3CvIRuHzuwFDmXeigNjxPz144HEQQg1q06Vp
n4TuV/YlMCRpemZx/a6n9wct8mQJtqHL27ZB10qQrxy+H596V8wRT2JE6JyudBt8
HrumYAMMBJbPppNqr3z9DGqlPw5h/EzPzRBjl7QBqaOOfJEvaASJ9ua6RueEemH2
1k1YzLjO6uIa/ecyBTcxOtRNxg0QVXN5VyDGFrbUQF5QuPJqFIAYkkbXp5pAaFX0
DEhHnU8+kGh3rhQPvqCMq2TFkpbw6GidvpPalOSBYm4ZwgxfR4JHLTc3ZIzWlGGC
OjlebXZa8dBjEEIjidBe6PkTC3aLYkrdzB2JCCTHOyVhRW5/7BxkQGKlwdqHt6Wd
8awM+8HAweSMkVPAA66zKRbBp97xGt+kVwNVLHZc8acu1u1cHoGrjPgKrkrX+fjv
blMGeu+/Zj/d41I/ldP2WqW5O7KGzgFzfNmQAiE/MRkCmhcVpYry16aoyeUhSOO4
UAVqrRPEhOIe314ydu8T7S5l1YMKsysawuS3D4gLLPyPh80cSra9fsTcDXCzABoI
GKYYd6tg2agCLMmjYt7PQrGjr4HbgTbQGK7WhzUFEqQsYAsAALkMC4VH3lD/G8O2
iCEhT2ZZIqf+q9qAQIyZWw==
`protect END_PROTECTED
