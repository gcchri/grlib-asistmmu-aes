`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
otImluxQY9BEGktgS+tjVrWY7bh98T2xeNTAMIS6eZS1CmBLpdst1hR+2to8x/i0
z8t4l3V0KPU/sFTJdM0mg+bn5OZmg6MQtqPEUv7Db3Q6f1A86isRRPPBw43+R14P
dOK29e1RK3dO+KKP1xOSmAfByj2D8944gze1gVprBTXRYK9wRJxOEU4yWn1RQdq1
rUvMEPY3Vcd1YmNrpqxdowhQ1kIs1NJTWFhVK1RONiOaxPcGIosNlKWiyt1zgZ0e
kQpLOd33a62+BofTisVxtnRt+Q6hXbTIXi+BkQzsmEJJSJkEu6OG+zmp3MSTxmww
Rz8Yy50+mzde2emj0v8aGHACXJ7x0J76t9UyQxJffiNAc3UQE6y0XblWFibQIh/G
9iDZq2OREhoGJk88qk63Mn8KgFatOmqBtOPOAJjJLUQdp2/kmIF99xHMTgIJND2n
005ANI2uEcALQbyju9SC1wcszhpBlrYJtNzf/cgtCGxxkTdGZYY82g+/uCf5zpZ1
2cJi0EZpU0XkG9PzVC6/7qRaolR5yDPQPmcUFQuxLkG2GoSA17f4WtU/CZXrhbsG
VKGZDmO5lvlKXKgJOk8N+QX/VtX25uY0olUa5x0s6kHNQAOMz8394RisBrSwRBSr
ohTZRKYYktje31IHs/NSOsQdFAgQI+/f87zgvXNXvTDLn7jB4ha0iCXGyQgbDybD
/0FrjUM6+mtH3FsLQ44/oAldEylDFXgSeD41K5+ONpGo/aYgkzoj2FtyRKVTj+nO
iMVCfLI2aVTCYhCpStRg8C77ALPkLgmlTvz06mb63UVbH1D/seS6FZBVVZjJfqp1
z6tDYwciA56cYqdL2QfQaEu7ODCpKIlS9SuJoaGt+y/syjIco4xwFevJjU/v+Y9b
ud394LJGV90VO6PpvV6i6ewZyjCIAOBLIndpG167T4ikIVWAz19nkWhc/5p9GEJe
yKsm2UhEo/Vtne3wTCkY0FmF+Vu4q9IZntEJlI3ov80ugGHs2p8e0UX2YGB/pw0g
nIIwX09JLt6mgY4FGEn5GBZgW4XLLa6zO7MQCV76IKWAZdxWWeP9XccuSlzhjF7R
RyS7VRsy76TUYTnlrtS0xQ==
`protect END_PROTECTED
