`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LgbFxb6kuV4zerKZ2a/M3SbCk443yl1NLI7uXW3mqP1ZBw27SG2h6T+4k9P2HM4L
O6nSyfuY7V7LUfHF++d7iGSLivaKjhZb+wXSPTbPAs4yLOq0dQiYEYnnD11Q7VV4
8aSKAbhF0C8yYd3ZxtI24vDZydWmTgoY42VvtquNjkCzzBpk2LRzXmyuZOAjO8qB
Td1N+ViHjOMEUGieg1KS054wYoUosvfBi77oWK3uI3zlmCdvrWu+HBoIlrUvWJwM
mwD8ERzDOJgf3w98lUa5sOE9lB6+T9JjVbB9idIM94tochs/TQ1DgjBsjXsYzSa0
tUp4n0XheAs89a4bVp4tD67CmP0SjiD0eo3b9I4aDWGua7urJBjll2zNyN2Xlkpp
QeuUzVNgsg+jWyha1gsmIgQgCigInrCVD7yJkZQ6RgIfeopP6v7rOCO17jv+7/f3
mTukJXFEolTbZz5VjaM5c4O/6dyIfozQUPTN/CcdJ1vTPpZ8w7l0VeRF9XoeyjSA
P6VT3v1SJ05kGQ1FJmkNZQZQKbAnWEg9pPdGad7fnbNWD1Ou7NvSN6kR6Vg6tw/2
4OdY/aasTSvncSsVv7GiKZYfP6/vfMYv77Dt9fH0ParD/U+eeQzCJmBGV6c1GxtY
7ELei/eM+elihF1pfnNWlg==
`protect END_PROTECTED
