`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DeDr5XdEPXHgDS8nEhDjrHuDy2MTctiVoCxfJuvvr7MQHR+f/uQLOk5/XWHuDVX3
63pDPIsNNd7FRLVw1qfNIostta+pTqoMFv/bbte63RCQKL8TYvzspGFz6ziZ5716
LFefFZrALwqS8aMvGFcwVP3nHxswsljKM7iYew1rj8wWaHIXXnyrdcZQnrl8wqIa
qdlkvIjyrt09BRnLSrhJVsMJJCvHnbmhO6i0HrRvwfOUMTT5xNX2WINHK8ZFkI/1
ifXNPP7CBe7s/ns0lRHKNg4GifLLCYt07R5/lKSOTCYJmjYhsiELpwu/rXV3huDR
pPdgv2WLk86izh8aChQMzG63skBe2EMhQbNx1pOjdPsuKMH8gASAJa+MQ/a3L9Iz
8V/0fxmWI18JnJaGJ1wR9RgFuDRKL3VXzSWgUoZJO8xobdirNz+co+kvbRV2xh9g
Tno373MJMBEqyxUTP/+9X4oX67qlHaO8R4DLXocABniMI/mb5BWZ/Y7lWm425xmS
aW5bhnkaeKE4EHbU/4gSsfIOVBnLeM02LoV68n3rrq/S3jmJppms6thLUWCc1mLx
`protect END_PROTECTED
