`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c5IVVOlnDr7SfeS62MK94mD3wCqKcOFmuoY7xYBwR2tBl4xa/PBosyoykEz6oms6
c8HwE9EOl8BJkbIpKrMYE7oGPRrPyHY35Lpr/9THg7Ev1jT7PKstr08/LQj2fDw9
Jc7s/ob8c5wuFgeg0iqf4L9jVHt6+RlTjl+wI4v09lP0UJhTUeecTLODP8CE2W81
n6mNRwfNvirYKgMfOLU7D3koAn0z+cDEovnIiV2jDwP4HmeGkY4a+S/4qLclalb6
qwU45S6I1kZYcxxiz/agNDtlIYlKVh3F67d3/H+rpfXhqhYNZcfgtW/RYElfHwDZ
Mgkri14Ug+JsDucFItdSCGivz8YUG5lmXf4mqyiiD+zN5TF9EOL6JfIRCScA+OaD
L437z4+ITFBarTy0m1ZeltKgg9EgMlJk37qM6+5mA2Tq0uX9cqKboKo1HJKpiD6W
NnHZ0Ng8Krxc/T19qK8Sy4+ufZL29G5McbbDSW+rgF9inxK+xF+trDgo00rB+JaS
`protect END_PROTECTED
