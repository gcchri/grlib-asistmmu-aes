`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5vpGRaDQ6j0qvQ6SMJGr79dKYD6HWVqU2Eg1ZzrwA72SPZTvyHNGNk75SA7KSOjd
K3rvKU8bypvR8mP59N/rbdN/H7v/fOUIfy3Xms51sSysaWR0j1TDGPcOXuHprCzD
rgFvGKqG4PnZXmQMoqCGRqTcoHYTBeYLysRjanARV4OqpOvanizMWM0W5FQTzAKB
QiNTWcxp2hZuH1K81vANi9C3IUV+ukdhn4Wuru0bAKMXvhYE6aarkubwzrFUK6Wy
yvcmKFbXzIQVIepjnW++ydkES6EFgVifCHWcDdy99lDzNB/41Hcl025Zf2n0mE/r
BY6pPC6gWAdfZFcEX7M7WXCviZFJow8jDwZ5dY6th5+XBjwyIYyijaYjJIBIkRZZ
s70c+dlfhgDmKLqq0T/guW1+0dc8KS+P8ahuMIMt/Foni6/5Qd62Nx0Yg+S23afM
zVYSb1h6uq1gAYYeeI1FcNI/AObZYmITqi1UHPbSWdhUJkBqFtnG1LbqVoU+LeTs
5rSmJBS6kmkiI4dAppqITaQMOFnbExF01lk2Pydot3Ye0bB0MBH4qaM60VuRjzAI
ET4dB9DCfpw9OxOZnKHJHXqblegBOS3Avo3KqelJzq8uWGZMab+3NbP+9u5r/1ub
MeulxO0AMx8JHE2dViVzwRV6KZExKPXdjJU8veAQT7tesDikM+eF5VsynkT821AG
LoUfZDv5H3JKoRDaLXOfJ8OjnwHVvpplZhawbVnWYPIIToZgNPPMP5zKV9KRVKRZ
O++Cb1nhKHtG6Uhx2jBBBV0ZrJ3d+4n92x/8t5kQZBX95lRGAytrwkf9RHSQyxma
sAlkYnVEQOSWwR5eJicYksasITl2Ubj391KbV9Hl9QCFzGlUXCDrvDapzelia8wp
BbiIeMhmGQq/XSrRcE0RkbSqkIxvwO9ShgF7e25v9KH2RLRBXBUZzAldKYNu8+Mu
86UjmJ6WVEvOpIS1DxWmSJ0HGDzjGQ+wins/AfDRUiAZgiQ4qAfF3Kn9GaHmH6va
jBUJVDXCQR8MiQSOV9uglhE1293d78L1HyVie5+ggV7BifXCniAGSfKqNdgHInMl
eraFtQgjKAXp4fZBwnmHHf/HgeGHLkFbuHSPUbbxwNc+GowMCAoX5S7QijOGspfQ
ue4EdkRF49FVo3ZoKM8UuwoHkgkwZNy8RGzdN/B99BqhuiRqPprvyg44t6eUVZ4i
omxHzZMUi4hTGt9g4C6uTmDLQ69hblgyYAIFejstVehQkVcOCPn9XIqX4JtxdfQo
6FFMnD+MF2mv56uFRjHyLXNnmO02TkvphlebW1PqLV7AwaTMqr119UaRXtDQkf7l
6wroppM0FRgkJbAetHP1LWFg9O2eK1kyLGH7HtrCf4GpVUFnIolnE/83MmiRC9Is
jCJMxGSum2qtaRg1fm9Ug3sEG39zX+iv6u01lADZvelo7DR0oncUNCyILmIRVkAP
CnF2w6vrBq5M62qYXCBQmnSe8kbNzNG93BMTwHESt2MboNl8ElvEA5knk0uFP+Ht
bhGNkgeqN81VucI80Zl3bTa8+7/3nYwMwEMhHl6pb7zayzpdlSHG2OigSegBBt6C
Al4gJ52ekCIoIqW9StAhYfOEBtrRYLNc49B04LxbOem/rAkZl7WmLiB23R/vvVNW
5g9t6qPsuCTJtzLzgQuOimyfNNT4SOzYhkUDIs8+rSGycCPNUpMg+uwgijam4F0q
CDzLMKivZjXQoK1v63TVHht0Lhf+QBjos84VgudxUnGnHSv1jw3l4NNa1Ov76TOA
3oVIoXfmnbZMoP9BWj9lkmQhtoM/AciKEr3wkSW7DefLovG3O54YQiqxp1pi5YCO
vCXvZTIK+dgcRAUH6Ta1IKR3A133g83iamsw7DHfcruKBt73NRmdE06U0hJhInkn
yROQUnBw4hFOxkxZGhKumVTJ+Ac0MYysIXyB1fiq2fcfq04AYjKkWqr2YKbg6wuN
p6GFDAY1R7hTIPuuF/RAkjA8Q6WHApk9cBk4Hm+Znh+nHkHp+GMoyb7k52/JcsRY
gRPv5OLTziKMeaZzYhqy62oXi2Wiopu9B5MDp/3lYb/kx2I9Sehqd/qkXtNY1bfz
o0bMASq4a8JjYlGm8D6Vc0ZrXBlxbY0IrVwfCVaUkx8Uky/CKThgfhJeijxvJj4+
VZBkVcLb1b/Ot9VFIsWb3GqNdWHaNXSxchkk30KP6/M47uX3Q3q1AfO89McYyGSc
DvjuoiHw3z7YseocBjRawxtM4Y2XXyZPDAhTiHJm8GbNEyU7p5PsGbCADGzVy8bJ
pGehhY/Ppa2IYMyGGSfL06hWzBYNBBzKeDt6h15KBdgRhAYJpfO6VFQK5u49Nfxm
OVQG3g2386nmcc1NfC+ttOigoQ0zhFwMfcW880EK2YTwqd+sPlOpWodKc0O7dOtU
`protect END_PROTECTED
