`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q20F49mWXusdXbLD+rWZwDZKXdSohTJMT2A6ZK9qYsupWFOTGJCCX9RnmU62RA0U
RZB7bOiUxptrt81PdhGAIdBtiGTxteR18T181PmotmXgbAVlnNoTvC/p/vkcGLL+
M5N0rUnJVHFK2CnYu7yc1xgV1A5Fq5Q/UVWf1kDDyTHdC4UJDoMgRck9k/sNnPQu
Qz9X9DgMDMmaa/uWC0M0QkKGYSpRTz77rt5feH+MIV4OrNjJHFEcvLE2tEg+KWHy
f2LxkCBBkF6X3nE4R0ffIhuliHscCekV7AsKu22h1wKfFfY/29ogyoatt0tNE9Ln
`protect END_PROTECTED
