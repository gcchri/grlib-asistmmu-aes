`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G5XlaD2uayDH/1iXKe7Z6QcoHWKOCKqyxoz+iEZO1Q8KALZUG28IeMvuDAD4d7Ng
zw7QLbX1SblNThzwhv0zDIrVYW0dhW5nWcgzm48Oc8xvSztl9y3RQ09CamVjp/Qe
iToWAEBA3sgUdtJdB1nLcttEfWVL0XjdvClKIlDxcnhtoIisOSILIAtnPozwIfPD
EHazo5NOK6A6sBUeJp1IxRlk4CvEvF8m18v0/lW6xz7zEbkqEoxyHXJ4yYjMySJb
NreSknZSwpDTXkCBv+uG7O00kON2zPX07PX2naN8xRZ7ovm5qmbrNpIDe0yDA/iX
cUKxuZbPfCvGmM/tPeUrZSJ3sgwaFNzqqxisWpwrbI/goiF/GM9rmF+JlkyFPH34
y+7CXIjRqWUNtmw5c7s6obS7kXkHNkhZozcl3L4kR2J9NgHESyWGCLAYielZFhrh
nh72+cGbxHSzsVOy9UjwFv52qA4aF/CkrXRExQ/c/0XM8x520NhfKJghutGGbzbc
dr2j88zJhP0Q0oPw6o3yR5KuJtY8p1I6pYSiDVW/0Q6vJpXTsLeOhdUzvJvgE5mN
BvL7lCkB3ds6licMAAKtt2IcLSnUTxKdzTwjKtIihRsnNqxwRbGoeBXU3JeHggvF
5pZrFaCqg60p1I55wwqSVQzN1LGAC8Mq3ADCv2C0bq7FkyX96UDP1YwywKFzTgG1
PAZwurSP0omS8TqbyNdXBSFYzedBN8WmzBbSKFKyDR2fE2KKDprTAZw51vkEMFoR
hVY6KN95Q2Nl6EClsMV6ZDcslpcceiXZ0PICCqlR7ZjMdUPlXJ+9VZRV59vjDmUh
r5qO3hjNI/4YpPv8Si9nBOf1gIKlIotK617qwB+crA4MNn1JlXp6TjmvvSoeJv9i
egXcOC0IAlE2UEOd8BW5986awdvZK6KgL7VD1qfbSvWvv93Y6ml8P5vQVndcpeX+
FmAgPKHKYODCx5mGsBerQtl5mU7wc2aeJlkr+u0aeLDNtblBSOS9EBf6GwZUXIru
95a9/UFcnCv5zg+X6lUoTW1/9kTVyC21eOkGx+CG5cNZ9SR6Von8MESPX3XI/1M5
m7C65vVsx2UfecSRbcQd/jx+zxuuEt/yjWedgUf3e0iK1+moBTsmjmZawsyJUNF+
HZjsrH7z8PbA9g7SQH10FZTE3bWGJQPtgvBlwmnwnY/dDTOnX+l+8BU4eBHgvqDh
RMPxlwkOcaJtu5FxopcoUBYAmK6n4HAqQmqY69wHRgp5FcuWmSTjYAbCEGq/6AVz
/LfymPi9/+50cGIbOvBcG1IA5wwH3oj7U/6fzwtTGTathpOB+0lZ6oKa0llHCzW7
C0BuAuk6dep6mD5JvHFW7ktVIYt8kXQEPkN3ACUEnzj+jfNXq4fX8Vnv+b4Gb/tQ
W1rmHV2i1dU7aAkhvSwhNda7AKYM039qX5pDTg1Wo2JSYje1Xhtl5uU/PjIRRMce
ZVzUCfBYGvgAmPECcndrCsK3IABKFzmpvWWB9UZ6/AvU6/NjteM62RsmiHJY7Aay
vblwXf8ZWm7nmA3GgQrj6zcV7rGqQW/RZCRMQjnBXCd9ckA0pN4J0sH9i2rhZTf1
/lAbSjDhMYUb8hxgD6KUmcXR+YHmAIsXnnCWCd/AUYSPkvPa6/9yE4I2y1dE5Xhn
yEZqrRGownTvI/1he6x6xLf4FA+cdptzIKKoso6nHVffSs2wlqcLR7o+OFOp7d2K
nihOEyKbBYttOqUjLLye+d7zpVnOfbcDOGCdAOn4Uz+MxlBEjG4SFobrHpno3H7m
nGtLqm9nPPYXwpjqOF7gl0p+6q1XgZcFD0SQyNx7qMJMGHLB7ih3mppc4wZzOmK9
l1G4MNYnYIH6OSzBlz/4jn5/rFZwz/05s8dEWdD/VBpTimdZ8pTiYZuZj0vXLZyi
ZHAWMmtPQyKgbCQaISYA+9MYEkNRpry2KTvDS4lSHw61wj2o5xVsAvO++RfPtYg4
2KuASjyj6jvsQ5GDYGYXaYohSIyuikc6Zf/TGkySFtAgKLRsX9QZ6LCUjH6iGbBX
tuLlAS0o5wzP8+RXqD+0jxGkNylZcWYlXfutzQZRX6h2MEq+OpmFC/0+uozJLl6s
GyTFNEnAkw7XUWF2sUPGC7Egi6XjLylIrMnXQPhEsW3DMlkYACOj8OcfUxplwh3e
fhPGzqqiMNGyofxYi3z1Nb9uaXJ0sxDZZnN9yHdXxz/toVJHq2QcJ9WIW555OWwY
YuLNe9Cqn+/xYq4FJF4D2olN7jp2l8zqroo7oKVWl/YiT+wqSbQ+JzZhsIbquV0n
BeaCesJwJYAup4gu32CUbkDz6pE7Zw5sdEbQgjQrFAPbOBahW+MzDaVf0OPgSZOd
yBOcOuPKVFf6XB9B2EcuKxqgbPUsCjEG3+cjgsvzNyp8AD+2m3zT38iEmCd4S+Vi
L4mfW+HRysXPFri/q9Bn09/7mMeLCtH4OQhu2tPoUOzPn6fRpEnavswTsC7yHbrN
/fFaH5OAJa1e4jzyQ7B9FyZgxR7rOfMLVpG6rD65D6RoESID+cvmW6bvEqWqUWpV
WjWwr0jro6XuYFb4RM+qMA6kJJb/pTUfOGzhfHDEhmRupwJ8n4aVqBPzd0WClnC4
WgkOV6ZJ/cCKrCpFM8YaXHDd0XfpuOORyQWL5tcFexpYBx8xCc0Ob2gfJ0UbSAdK
HLFk8Ni0lCeu5km8OWCfsVvGaoTydousqDo2vByPI1yyGsgHHHo/eOy8jYLR1wMw
uEodf2pvslUi2fEl04j+aNGWwICu7Zn8qk5c54dFGdAsnbqx0BKpA2FJMTRj+o5l
e0qeihwzZl1P8I9K1+SAv3qWYh+SEgsg105R+EVKGoItxectL7LilNLMHM/f9uw0
Mv3LWOjFXuhaYrV1QEHGSHI/3qwoOMOrtVySt5bCkOF2Cn8nbApXmXmwF8ng6/WR
bFIZG+MoxcIJjtsd5/a3ZAw3HGIeJWxZXqMf6wJXnMIPR1JkFrGFSG0ZY9jKsyeY
XXrl08F28XPeQ4PaUixine88Z+jSw4+DSnDBgDcn3CuzRGy1osCFziF3+wh9lItl
GkFlV3CdtnWDizttj3wvHfJczDfVVObZhlueqCzwSYL1GpBzdkWO3AXTh21+yIqO
V10Qa/TeuFinWtSkssbPltCryQkZKsvrAOP8ooWR1miQx1tnmIAL2sw+8OftMI6P
xr3KknnSfMoMdUZh5b9BgULSgICf1L0WnaOM8PD8NzevE6oME1hLPVRpHEhPrkJw
8o335CBBftrKDg2ZcS2UJL+ymyAUh+sFrqkjrk7XJpZGrgb1QqNkj10dcV3iXJTS
tXTMhU31NcChsQ0SCwRVwBRrc7J5fdFqWIw4DpZNeqFWRtdqZqVv7bAN5GQqQjsL
/c/dxfiOg2MMXap9zEOGnR2YHET/fzHzUJcOwDbkTyhbgPxRZJRvgtxu4N4TDMkU
gVETKIw/NXkpa7yOG7/q6ZJ3fjcX6nFyr0XRS5NqcmgjZn1vNUEDxus9vHG53LcA
q18M7bz91qt/VzYM66eHA8FFq+sE4HLJgYfVtWm8W0tkyoyp6LeH6oR5YoQdsJ7Z
5pEVr+GeRT6D2t6vM9RpF16dDDE/OVa/secv2afLxlupJsdbozEeq0JpsMKdnhEI
qD9FYR7IOkdW1yAivGT2jxyAQ919MLEtR5DAOQGBzsSPoZsup0cna0WsbZDF0253
D+GGVS2LwmBz5P4tel2uO6dowuVPD0khRaB/Sd0H6P3DkJO8Gpnxq9Pu5TMxdRNm
OV1pOdFItR5N0WRPV366RrgW2o+XnglvTuLGtF5QXNKF2mzOPkeHBvqjI1U4j+iR
YV78Xdy27KTDBIVucuHBUymCdBt6lzzmx6Q2TkcS/kHBcrmZjUPzRmw2mT1YHRlw
bVrfuoQXYHx+f9dnkoLN2KtE1EawJx9DeR4Rk2FhrcSKy1H2sN5fJjjPhiP9DB6r
Zy+ew5+U89gx6iOVwc9Tffnu5eho/fWY09QdWqcawKA=
`protect END_PROTECTED
