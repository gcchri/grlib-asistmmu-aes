`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lXOYtKYt1X/aZNZqpOv0gqaw23twT0Ca61udvaAB+/P9bs8f0n1n5BmZYBOk3x/9
pHXwlm8yIUpQIKpd1w3TWJeWoKyHv/dMAbHoSUplFXcAUl4JFdKAW3Cml01/3rvb
N7Ac014LcTr9PqhbEMXRlvgLYyk18si86E9nz6YnLdBD2/WjpHjo/5vw7g0wRusl
trk6W9lYA17wQnoTAbL+hsGITfn8fgdhgsbnsB/np1KfIBJbA4qc/9NoE/BK+S4Z
I0EUFd++L7/alFsG9XLomJhzFi8y4u6yoGyOmKDI2mb/Ddvdc8m7zfDeWJLS/qeo
/nGHg3v3m2y97TapkgEgLU0eSnrKYfPm/7wmpHHzBbY9yNtrrmXMPZYjsNqd1BCR
6L3H3/hxRofD3tBDHuHjh+/0+vqei0CZE6luOXSA7M+yvMvqpzicy8YjbkHbji2I
HrIh2kClkwhOv500oCvZK3vZL5mszpEM3O/NNURy42ECIxz/nPFXo59o22mF19Sa
RMzXGTsFObkhn5CNk0Esv/U13r0hDMWOR77oqfwEhJtSmPXTlNFUcpZVVSQO6ziL
O59qNmx39GjsYORifJNqaAC0Do4SDc48WwjHNi5u6MIlvHHynefWDVKcIFOlj/7L
X5DFbNJvWacdriO47Uyee88AogkgbYHP0BWGWrOes9SApgOQV/nxroULtsD5LzxJ
KQdL8njbb7kSdFWr4IhI8oNaTEcvoC+wz4CYgDXZP5UknoYnU4MG3u2RIOCxL2aF
vvkktC/sRjx1WSNbgveau9VICmWO/xxCJJy4634aMsvStkWYwme7+YVqcpcnLzmQ
SlKLKT2eY68qW2SMOPvLzw==
`protect END_PROTECTED
