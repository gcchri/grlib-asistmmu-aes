`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z6y3WXlhrQQoONAHXNc2mgUJppyOSM3c1/Nu07EjJfee62byKmg/RnykgKk8o9+z
KsR2fCSUOAACPCXAXL9ilqOwQHkov1aolYZCgq0XpygonO9TMSrE32J3Igi/jEMf
Xw2rt4IIpCfrdT8HM5EWhpAd9esGEGYMabXqpIB67b9AvRfAIcmaVu1iqbFE8M2V
wv2b9Ni3paJJ488Bo/tPFiczRPuP5vNPErOpORiLZaTcqi5wYJztnfWUI9wvwS9F
ztskpfg0eBkSJjWMtBuH7JkNCACZzXYi2UavGpWLN5ZLwqeqo2vj7Ku1AmJTVejw
6LXYnSBNly4QBOoq2sICFsYqXodY8/29qJwh39/OECRcirOTJsvkWnUAmjJw2GzR
dgvQxklTcQC8hEC2WHb28w==
`protect END_PROTECTED
