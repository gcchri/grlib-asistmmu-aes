`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AKB2661zI4f1cU2l8KZmiyOxOEa+qd6HVHdwq34porzt+2p6NjuYI8AFYcgfYm82
eRzOs5VcqqzhPS9zLxGn/4BMOe3TGO4D/8WotMA1Ozdm/kecrIxvKcacijf/vb3n
wTw09QOdZWsuIs/qPk5O7Iaq7+zhCng8Qp2mWigWjeM95lnCJe8DTjXWo5TXx86R
ZoJLa1JzZzfSPpVkWHVKl5BVVPmKRTdHnHQLOdQHLiiB3GNIpYUCvjpVBozc7j+f
5262obsjROwUccOZ6YoE+tmCMppGzSKSo1b5NVgcN3F6fbd6J4eHLzlQ669QK4Vu
XGxemmqgNPAknRPNBRpRuhcjqDcBCwiWlGU6xOTf7ax2QFFCNRWne4aYN1dk6Lo2
NN3gR083AdOGL4xjageRIeWzGqy4VvpxtVapzujtj+Dchvj7TEsXrAIdXuYHHXzZ
CQUSbbtAYrmKhvUmbg3K6LPSwTbgScrJuazK+HaDuj6X8BXk/O264+m49UdpxvDb
ilCRO+uk9j5lfbKcuCfHgvRm2b7pq6iYyd9iGtqKVCwkyw4noWQRmVrQB5MjWQ6L
44INNwhLwk5YzLZn3m3WPk3+dtorH2C8caoGswlm71K3m9G1WtJc+rHivMyyEGQB
kRKCej+rlsiE2kmslDHuq82WwrrE5uHvwqEN2zNSjEel+2h4JxdTVC0D4oaX0Z+9
0JnOkgCBnwQUauNWrJeB/g2+S6mcZCk3dFGhEI7ukBTKPrHNKQqi9HGUW1RBGUJK
ioR8Za7Br83aRcADcOSZfgpZHypIjHkycZMfHybAHyDNZGeOgNhES+9ea0+d5Gb7
xMdAj7VANaGUU9Gn0ckRV58AzsEmMprbww/TgL48H6M/v3BqhzC+oDxWIshMu1nK
sNHVQzkXa7rZnBuxyzGugLiqrz4fffkwNm/kVnTnTjbMZvZRSsOspC9i3bvs3C12
4KChFILPLd++0rFsKgiA4qh7HMMiwt7qxIvdyu3OmYg=
`protect END_PROTECTED
