`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
epi0EhyKGZXmLEPeXORyafDk3pbFm2V3VUCmrK4jtspqvTRb7p7GFOAIOorRBTtk
U64I8KZF2OvbvRSEe9yWuiwcWlcMR8ahi+CtBO1S3Dqdyrl3/4RnUoMhfQamntW5
uUJWK7LddZSiMuzxOcRbSnfuXEo2c2fmrTsqrJv6Q3WG8Qwp8QkbVT71o9RJh4WG
DLNxWObVXidcW0GTqe0pJkTKpt639rer0100N7KZ4fWbRiCDN3endcLuPwnktNEC
f+iGev768IS4ClAXNOTN+vo+Lxf8I5K2W//991XsRrDeyA8UMJMSdh1CeYJ1S/On
vvv8dmD9pRcEJp8G52BQMJZZrKLvdSLROqgXS65CHwyXoTNtC99tI/ZU6BmoPMuE
b691JZS56ryl+WKZ5Z/TYeVFaWIuucEjnQH5X/7Qr1vTFeBtkpMht/F3yPFGaegM
mTsX+PntTDajl0/4zGsAbQlL5SdIGSPMZqFpbfbGh98+Xy7mw32t3qPGRY2pPsYO
yA32m4iUWXxfwb01SAj50Uujf1J4zuJgmbJPzBJpdQUJNbHsZJN+BnrVKLN/UpVT
VqfjLKO3duSFUkBvOqV0UWqU5CXYK9EGW6JBr/xx2YfoIr48g37JGjYIHe6TQBE5
/O8D8tum0fDP6+PSdsuGXu8AwSXFFGbPiXKuRKF7yPMrfiCVi/EoKfD1dV6LjHEJ
wSsKrzQr1gqEKu+/MqGMQak8hQzoA/6WO/WGDcY4+JavL9aoBNCNNDtl9enO2zZ3
eydi3JfjgFpemsYFbmy+ToxUTgSL1E/KUzYooETKd+WZcyQVwgKjK/FR1j08Zckk
nh2kOnEkMXKh8BlAV4tidHHpkD0hFA/yPnjdKmPcZwrEKhqSZx1cU4EbAwi3EXoP
6eaG2Lf59dDTSy8AFy+2JamYgZR2PyLkL0qD+Ih9hbQ+J06O+j1PnPMyypG7sMxh
BHZtr6gMzQFaaigUytkb3TxS7JVzIdHC1A5YTasIQtzDoEHGogWumuuc/+urjtk6
rZDrQ+5ObFQFGdJniCmqbWk1rBkli+VKT49mjcPgun/++uejuDoPg/T7Jsl6mAFm
CD6X0BOc2i2jJ8jd6Y3Xxw==
`protect END_PROTECTED
