`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pY6+CCG4nvIjYksKdPPzamzV7nwePjWOpP4SQeokwvTno+vs/U1G4q8wRaPYsZpv
0EjZ8DgJrXr52jEKDkEE1T0G07F8NHw4X00wfdtxwix39I4VGLKMa1uqr4FtPcyl
as3SAlxcVYDsqMQtt3HqfvL0NjeA21vl1o+0zGDlMOkeRcfeL0V/7L09SGcJb3a3
CpahQ/W8bgph6JBtBxYpiKmSNM2lIo2l8k6KRGwcFR1sk+0kRpBgYY6mvwHR9jer
z66uq9JN4aPuOZjNacKCrwziXkN6d9Wp6KneNHsJI8Yz9JukS+k166B2qeCvDH7d
DT2KiNFMqfzgF1Js4u4nWQJ8cI0/5m0afI+jGepP9kLyi57f+z/rLLZX3Qi3k3zW
5jCFqhfM7aOf52X8YVrsGPeWCamZKo5FE+lc3H3ffcTcco+j0mh0BGmOd6BnVzUV
GGR12DDg0JfNMPxF1a8iAjmJxC5ZGCEl8QteWh7p0XSWF6yMEN+OJ5PoYi/p/Grz
3xf4qNDSQMrJDzPj84lXEG8P7MpgzYOzp+g5kI+h4l3x01qm6GZDE1XEPZPTiuJj
FDn/iLb3sCg6eaXfDWUipB8Eg4CLbdvbDrJ6CkyTLDLu8vpLpknRnmr97vC617EG
/Tp5gmWCQUDc1Z4lKZoXzMSLRP84apnnHnaGa0sGyHePD8cZ9PTxXUA8D/Pd1T+y
D6qYvAkx+W+P9HjGcZhUGDZcgRcTDwoUHnkvRfH9DI8=
`protect END_PROTECTED
