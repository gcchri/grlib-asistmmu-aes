`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+0cm9sflH6ibijb+sjakUwBJOpSu6BZ0zifhWTvQch/EO4WefY25jorj7YVV7xMX
bF2X/1PnaYNW7XvxEnvgODJmKTvYdaZkjsD/6lgnQTZaYW+4O5yQ7js7/yqZfHQV
EjnrR3BwcwkEHALnIQ6rB/yONIglXTKYWaT08dv3rlu9QZDVpt1Y2hUbsL4F0yjV
SeTu7ffWNGBgwIUoCHmd6poq72T0OEhANQertQC+Y9is+K06LDpiC3rgwtasqrW2
VfgfYKvYyuKEuzJxfQrgllJ+0piHMv86HyBsWmmZmIFGdQsX8fStdqB14d+j3X+w
QVRixCrnXGZPMDdomYCoYgmJQfP4QX1xI09tayYq3mhDRvDetGoTrQWnxgzHmtKE
Ry8mBRkXd/iot+hcWFK4KnniQ4rZl5rF60hRljyF0DKQXcmFaTMPquy8pKp6yoja
PhMT4ny1wQC3C/ySsUFh29t6UwPfe5rjsx1aMg6BFx+3tnFUURBDCmmzHSslH+x+
rPzy8mGCvbQ5tdmkhhMT8YbQDNG36h91QdA46qcB0i/Dv6D7Bd+9FkoKML6vVWte
G9o6EP1Apu/knQDv0DgAEOmwHP1McZdCzsmxJ4cwiwVNSsd/15+Vlyxj1NgxPrUM
U9nJrHqz8NBWnvDJ5dtpaoiEUgNQJmKZf4IJHu9qjAN1GLa215Vr+ldy58Fjw2QB
7YWDUhLE5dZGsGzu0JMhf0Rx6wyQqiD3ytgeXgJfRqgOPfzLXmiV6+CqND0enf5J
hZEJ2E+mn6NZ9XvVSDXbVzbA/sb2BmtH43wH9H7WY7AwgLFfFslifslvD8gG/Y7T
jDRzggTsb0V5R8QCe4wEbq4czjTWtn52wQZs0fv6NBzc25en0ZtxdDakjOEHnLPY
iSfvxVf58w0nzkSAbnFXeT7ZJz0SSvjziC6a8UQnseMn3iALEXb5SaVjrT0bpz1K
99e9icy8JxptpJ0fIOEByXu+7TdB+U3qlhHMeHM9OrX9zjVCPIzxNkCICYMif/lX
/jZKG1wBt1ufM1Mop7woHgypNZqw8zkR6FR7nv+dYuUtXSxoVmhuNMMY/xAtn2Vx
IMUKzvwFH2xXYKtMpivm4sWAMP0kJk9M1AziqDWvMxmCYCXCmfciBF/cHbOGsl1f
/pwuOY+LwY4nAxCntul24JnQE+aV7k0bYBhN3Tf2pSnwdaI+eyhlZo+KlaEi7yxu
`protect END_PROTECTED
