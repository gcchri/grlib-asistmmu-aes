`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1i6rkD335Hr8v4QWtdp4XYvxYAP4T/Wv6BX3WU3JgJWuMPGiGrkxkdDx/5qbtNAD
GoSr4pVUKzqm+5Obdfv/OwOPhp9n2CVRnk9Ny727KwSLx5oT6itDtXjWCaCa/d+w
0qTpeq2xo73XO4dcJpSAP5ZTCOg1HQFCSJjcdke+g/vRuIDzPGeYRG7683mq4Llm
5eqsaxda+3UU/9s1KLjiN7IHiqA5U/ypu17XB+yJYJwi3V+07zF0hHBVFwx8NPd/
xdosXDNe2YnefoA3EX2Prorr3Z0fyvJJEqaNkbYozXr7UlhZOZai8nY06/dacRuG
2UCGGpmbFCt0Qy6Gs0fIr3UDF96eCbN7PxVEDJmAzhHICNFGCIkufhedMUmA67y2
szM0ap7xDPGpuyNXTLZ9NPg0lCawoho7V8GoaMEOyzk=
`protect END_PROTECTED
