`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Cr5DvU+6igTQSKeODlkYwX97vNtoOPjrRjJX+mIuNVxZtNqTvFi4qAsDsli7LsU
YanBLh2iWcN/mp/V2Y2c5qNV18Hokj6yeTUNzQNU8woBvekn7BGXHKOGmkhhtdQ+
b787Pb+Fs63q8ouRRIIRiRPwnvuYLqz3Lxm0SW7edLHtlwtOsri1Dg7yQ/dbWsEY
jCmOv2g1UI90CC1zBvQDSYI6xI5aOOgmCsIhxfdNQYx4vG8HCDMJIOa1JICLzMsK
7zvOOSPUEhUvhdMOuhqYDjqhFxXqdI1WWCpcxO2uvg4=
`protect END_PROTECTED
