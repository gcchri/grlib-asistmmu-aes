`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zs4abs+sBQwKkYu01uZsUSJ5Ar/ZlcdUq4/sxVESn+6alelWptsiwY2HZ0Bf/Wtg
SVie9zGK15hjrZ8rDg5c6yCAbOB40Y6Gw3UZqZW4GEAuJ07TrE8dZemGkSlEJFvR
Or3k11p9wPTqubVOsC/sQ2uc6JiOvDylBfnHfIBpt8sTWBlFrBcXkxw0DPkf8TjQ
NDsuqwCaVv9NaWs4xryA5fnS/8XM6DTwKLPvRttDnsBmVqK6uc8/Ef9b1oS0hgOF
9bNlFhMmUkwmVzU7XRDg23/y4dS5tDV6mr6oLvptEmeGid8d3sscsynG2ePTLJhi
btKNwAayTZSpUtKMLUJrvG+mzcHWdioGiav1kZDrP3kEHtHUCSVYaM0Zvg1tefXh
oYGkuoji/Pw6gqv0tqAYql+GnSbF9/Zb+B3tU4x/sCs=
`protect END_PROTECTED
