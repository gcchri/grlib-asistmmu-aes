`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vzrSfFyNxdUC3uB7v+lQQMQY26bY6IxxqWL0WdqGRua4X4JxERoLHqsbRztanY9/
73Hkll3PEXTWKeCjhsFUgE6brHJgJkpEiq775vY6w1WlbnUWMrJdNxpfr9QTC+lS
cfp21Ji81VwFOAVG/Tu8/RiTpCYMnlx5PNRGeyuLfXtPeKbjhUajLWUCbPvF39yb
RigNUZsUOoN2Ur2Tbj4zjhpV8F+B5nD1APjexB1hwKsXCSWGepNG795Kpcee8VUi
QXQZnTwDMLjWGJTdC1lvBZsTAkYlvRKb7X/kVXgvErau2ih7E9nz/GOoR+URED4S
QN83vC60oIf7S+OlN8ac0wzO23qjJaEkZ1eFrAIi42kmQgAzD+k5K1sQO4g0vIMs
zG9zLcXGxT5NLYsuTYjYWkl7jJaFGmtjZtCQJQTU6YPDjGJPAKBbihGJfFTxhzsl
DhSir7u4bLrcAJ6x8S2vxJLJq/xNGw3F1vDnLk1oVy/rSJtjl1WMdw3/gGGy+Wh2
QzlxMPhh0KMadRyilM+hIChs6iyDxjMHtgZyraT4nRfpgRRi00ozKy1FeVPHymZw
Tk2hRhj9ULtFnqf+JxP6l+LXtmxcSuSE2nZzYztMdpgepEUKFg3GtfOMzNWfP0pW
rqz5QwlMTUQZxE5J6HAvdg==
`protect END_PROTECTED
