`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cXTeYvhyxQWBIyqOAh9VLg+mXzM6ACl4fVn2TgPJVglRsbThO++VV5+Y9KoEPUwq
flgmjtvoQA+yM8YO2dhI/tiSEotRJ4/YYvEMcaiW3XGKUKvHSiHzaNSCI4j81QG/
LXx/wOR4bMtFkw0640JzpMDz5uB5DkGzY08d2ppF+MBIlwyVsHuNBYrS2Ke3/CbV
P8yzNGgFa7HRF6akJisdjSQdt7+vQKBIre4doBCeQaOy0/I2/CwlgCUdrZZIJJP4
jxAzg3VGz3jmGZSjvn7r0FAfnCXajINqFRNdhz5kcN6ydyIvIoEjuAZmxnGT4/Km
7jXRGtBd02p5q8gSG/LP3Q414a1WCjI1qyEa7ny0o7eqHDzGV4dQe5zPlxfhiqfd
6lJSUBeZyutG3ooPaDXfRTcB3Ha5pc4rCP6XdoIWJ7S26ELmCMX3LOx3DeSCJ2SZ
BaPv0GYbk5zoV3Cg7JkdNo+F+jojyKm3fqkecl+BV+Axgp4UZu1fIUSrJ/QM/r3R
4R98cnEnOE3X7CuLqoTC3QpXu+9/SHNaxBeiBKuBc+Ty+GjZLBmC1LmejECFN480
PMsBMjniWpqeds7lK2m7COeYAFeZX1+mjMnfAMfg3dc=
`protect END_PROTECTED
