`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aIILptYJrWm/YmPSxfHFH7qpSpKt3i5qG7EbQloM/jqQ3Fkf5v3ipBDijiYB7T8U
ic24QR3RxFoqsd17HkR/pz/Har0z98MSJlAZF7WNaxETbsdQ7f/KAAZuNltYgKf7
HG6JXAT11nCNyTWqnzwoWlG+y0twVORHYVWZT3oMSUryisojEs2MdMdGNoNyctdD
JjRVwBnbv/lLq/nMPkVZxSxwjlajXBKDl7zzCdYz2Q7VBhlL97eW044quh8XDJ+4
EJroUW55K9QadDDA4Iy3Q9zi88ReuLWqdEY1Nc+vKE8JrekjE0fSB0NgulWAtZSO
eUa1tGNslwrCVbhBMyv3NSi6RLBYl1DVD/+WRNX4Ir9umdeL6wVGLgA2yZxffEZp
lJYEh4riiuMiXOwR9fTcFYSYrxp1yMjHQEXfhCHXd4rIS7lfSGtg4NdKLBj0R0lc
FQ4JQalDfoJmGE9qpAnnEsZq6ELIlBGt9uM/KHnmXkZVDftxoL6px3G1VNTNPKKW
339IkKTe8K6ApZLpnBgWauBxS9KiQWMIE/XArVId0m6extnCyHpTW1ri4aSOnwqc
jpVsX0PsZENvFjLEE2Jyxb8/b8t+IxZuBFHsV7SObg77Bb+Mu3/NLa7/zPjmmeQz
Ib+l8gUa3kFFicswJ5Rx2D2ztjkgvMEJ1THKMmc091bavmWwnkV2Yx1Tt2YTWF5k
W0gu3HC7qi2Ze/+WsAqFa+rZwjz1WR994updkRywl3ht8+9DskRLK3wuJQSGKcCP
6cNHXAULPHtadw+8mH8eXQ==
`protect END_PROTECTED
