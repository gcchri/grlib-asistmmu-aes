`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NjrtDs/R1m/IeoZQnPvwO5o3hgfyz10Ij2r3PtRRikvmzm873bmC09aRr/v79Nfm
3lY1p0IVrLJIiAZlQQ4EXpKVXReXzBGGWcgNyJ0f8lDWNlH0skDG8iIGkOTCgg8p
lJn/R0mnYTgjMW0RFtxQtSmZernsqmf2BGx/Uow/yNW1ESXmg62EUaoFn05nSL/j
o36AaxxcMb2A1D3AQRB3Q2nhSV6SsLhlE/4BZdtCQjlk7XVDp9aH5ni8c7gOj6Fp
K+h3erMRXwUkx2aCk7E8WDhU27uufIB6OQbqGa/vbo+wzakstqlOc7708qIqDEIm
f1kVij1Q4lStX1judYhhvKxePzRvcNPobNvIvJnMsB7zLcZ/lAp6TqQa4Wit3GSI
ZF0lXXI8zXcJiNa9nXSOBV3NTMRWpCIdSbYs5tdXX1MXqiG9lYUWRCitTkAX82oV
rLpByVe6wO95JL2FQSGFfUtLExBIu7+rcGFlE4Umz32XB6OtSA1XevMbT2H55HwA
ylrvncZNrA0xZGqkvo2RFgHW4ze7oswfEiZ8uA9P2WwfZguKrUBvgy7oRf/4Jd+v
U0IS7gTAe+0upDlEned6cg==
`protect END_PROTECTED
