`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SAqC0yqVY1e9Cq7THxNDkQMNG/ZXrBujR9wGFuPTCUcwdr8ySxboWvFAMDBNBegy
paruSS+QoHSTOnqKxbHrtMH367QnWmjfC7w05KJ67PxS7/He7QaMeqpsGX8XMbKC
Fz45EMPceH3Lvny4Rc/317xhqGqP9GDOV9FsKGrUeCWLXREXkylX6p6ppIVrEHTc
nwbhv4LlzA6lxKXgU3l2Dy6kZ0HoAbooEwVQrUEFEtymTTBzvEObZoD2yq6w6H1n
oRQbmWgHKEumqv/tifV53qWUTzGdtv4rA8pqtwhsNKLDZMWR42ecg8u8XfAEjK7F
zmT6HpqcsSw++K+qY/m77OVlWa0gS7Jjz7qEf235/ey2Ez6VOiJLPxxFl/fLDj8h
i5bueon7LZcue7iKEiZuHyZTpdPWa/D6bAId784AseQ/XTKFD/gBrhHnlcHf9VB+
F4wWJWs2C0tG0DFFCZ38CzF3ghP1WMlGVlDfnubsPtqfZibbCgcqFncxPOWQtHf0
IjRP4E7RtL7nWJ8TMGeomipTRnRS25z9ZLjt1V7ZzUeXyNiH40A4oyvV4hPlMmDl
Izk7rnD2kBzEtIf8XjEGj6yWIoGJke0gPCmB7KJ+L8psW0m1xqWb0Vz+kGHzVWtZ
ByOsv4UbwtXfOc5iTzg2ExLiXbooPES8fSsYDyVdMgO4u2FoamZKep6RiUNZ/VPb
Nu+B0hZvZdgC43ReRvQ//8HL2nU847WB8uvxbgthCzwoJAY1m8QZiWN4KnowCeAs
9qgjOERoTe74KgNZII15j8PGJjGzgg6uwUNNlAynKWP99p6S5KUl9zASqd+tL92p
EmMAgVMJX1WuREQ4PCSlN0LI40PfvrTTdvjHWCopXfZJrLPe2PnWZE4O8m+QSiiF
a94/e9joM36a4pv7WF6TboAPRkZGz8TozbGHaGEKRiY4qSn0B8DuKFMzY0k0CkIi
kuL6K7wTQW1CAwE4o9N4YEup6pEPO5wOCCCvEEspCkyh9q2biSVft3bDkFd2S8iQ
PmuyeebiTDIetSQN/7M208NbigrEXDvs7f1+WGlqSLRHbtrhkZoe/HS1h11IAaa0
SEGirKNjF8XTBoGACEq183lgeLRvOmlPDVebLej09Qi9Ebmp2rf//QCGEoyok3OA
/IyVUC2UpaHgB+rrZgH7SFyrHAPV8P8CKgTTjjhl+cdKHgmSaI2nrinKEzJJO7ch
giKYq3EhY4nDIUGinynHaXmWEsqnDypopf9AFCkuY1uAYNHu+2KuEQUtKEQnFfH9
aZfITT5jI3Jy1E0PwYhn1uAthLXQVFHmZV8vewSHVeYvLp8QLGoII6yDaQ9fcFcM
7O7Yl+mrWZ1JnsrFA9x+5//T5a0SRTE3cDCJJvtleyFMbMVzI7GU8gJpEqPkYgAz
`protect END_PROTECTED
