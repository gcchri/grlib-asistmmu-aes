`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YtdIInckHCUVzKIbqohEGg3MGgSBixarSd65sQ0IYnCWMBSsuIAg2jjXgD6yJm9u
PM9j28y8YZYfjQF60CKsWkfgo4sOCZSivHOsR1tQuHiYn7u0zEWc8+dIEpz0Z958
tnRI4TlpxC05LtA4L2CyM0WD6PiaR0n9If0vm/DMGRb7zPHkygeBJGZLsjt8+iqR
Yswr/NK4GeOQ5kKpGmRgPfhGlw0cP7uRS2obn1ggj8Q/yxCZ4y9qybNDYq6PKH24
HMIdALfDXq/tWI2pAuIXbf/OUVMIiSsDcAp/k7bdwHc/UrnjTd0ZOhcDaT/4V24r
lXFAq76p8LlWMBo91In4lwA7mA4ToqKcXtgQ2NHOWf70BTrsrgBEl6sqmjG/DOcr
HO6pykXPbEDuOGKujiEMGg==
`protect END_PROTECTED
