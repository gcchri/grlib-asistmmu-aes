`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YNTRhbhSnlyPgROyI/waKneY8rc3ruN22YTcicuoEMJncVXqomagBiBD1b7JW7hm
wIn6gi1la2FZP3T7pnQjmLGsIrLhVbBykEXMcRZqaIjZ7KGNkisGLRPw9AijgXA+
idOucbkoN5jjTgRBJFO2z3nIyJYbUR/5LtgARqFXXDCqYPnkm9xPnYNBuWt+Z7IY
67QMXUvm0XE9RDjHuys6KWfgJVW8gVGcaE+qdPzaLz7OEgPAcHJRHva4emVgC96z
gd5BXMK24dgbaczdJiVd08jOZx89Hj08+bvGs13gu5Vxli01l7vIknx0BN3Gloci
BFuBS4XR7QobiikCti2fdx8HIqk1ZTtB2QjG6BpWM1UfuLTAv27RmO13V6xgbj+Z
HdB1qtrwpe+JdHINw7HdeX+l5IoIY3MtNhP7HMw2xuGhmwSd44aMYMI9yqJGODDl
AAc3FE4x8jMLZ5x5HL1/m2bxLz9D9LCxTRpw/JOmsNSJsYppdm7m+2jOEzEXxsK6
VcT8XpbH1blMi5tQVcNI5YViBA36nLQoD1UuHzvJuN4MfZ8Qsuxg/2NyjrTNBhLl
2KLOwjjbPlSgu1qKIrzmgsymme4zh7dyS5Son9HtHe1bH1za1d7xJRDQCDuurqRA
KC2sFF1VKJ4zDrm7LDIX4yoEEbGhHQ1lYHmK3ec6eMo=
`protect END_PROTECTED
