`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aGM41TqPdbYuZJHFAsrOdNhAyzb+qKyHIn6Jg/tbLH+kHFSbkskzJBftBMCjCmw+
K2KqLe86kytLX54xRYW+ZbySlgYBHL5FXFjnOVgriEpy4PAXKtGPOpvrjaGgcq4B
9AQNJfyHae6QuHVA9QywWix0hBxpM2B7y1sv5JfY7QibMImOCekQGlZchApM6mUI
k//Zl14qszq0vzQcpyvRPWkC9OfAptIR6LPbINAIgKoFUCC6i3jntE55Q52Eo4B2
R0FdFrGRkMWxTAbURJCGhGCT3l9WeLu0E3t7ZuhXc2K95+JXmTSW60RT0WFygsZY
4/80gjUMaxPTo9jIJLNeqy41nnWmtPqPYYenIAg6pQmweeuFszS3C92HKNte/dyI
N7Ja/KF6dzSF+ZMU4293HULrK7lZSczMA6HY4L59mT/4uA209QXSGAPYTWL7t4u4
idyR2gNG+POi8/2iPR1j8ElQcdXw8gJ9NHMMhChz9ogMFCLqoHiAKCgdjfas5lbY
nqd/M4PQ6T0u4rJPTQR9fZyYrPYUERsoxL79spgeFvfRCjhR4I+x5L/6jK7A0xg0
kTwuB5egr9WhWXRe2fDRxh/U0n68LxQNr3ZkooHk+qcIv8n9yqeVxQlIsQZcjB/y
qlVubKURXdE6DdPeOdESzfcW3nfk7q2xDy6TpRVeRgG8aAznI8TxRNBifd4h+GEu
+JD8hm7hULVRGXcbitxvRgZLedtx5giW+GDyx9JGWawxszAaJHkkAOJlc4DuLsxw
dYY4YfvZxcW295LO926XmoM3AJ8tMYeqLEdMBtNC8M4XErbjRbrh+dgUaSUUHiDZ
fTqkPe2z0rLtsj5CKT0jUyHuksC4L70+BnUcmdpnl36cSgCANLxLZHLfRN8tD6i7
C46SL9EYoBRzO93acfq5VkDN7bhv1vwVfoFbWVF8W4sFjpGZy3NbbZvHDwECW6jD
w8AOL+2Gg5uqtGVO3A9V0r7ccCnQ/ZCxdYcpd1VPyGKCEf6DlWQP6xOPPnBxIxqN
atxhMrshYrt0jxlWGpbToA==
`protect END_PROTECTED
