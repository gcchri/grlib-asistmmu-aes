`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LO2nDHgfRkIw4rJLxnGBcGizsvJCNoHokFfXrax/r7kl4t647qoFflfI4qgl59Ow
49sGltNpItC6IwDLFtkqChEX5bPOpmnAbJaD8QfrqBI8B5iV/PbEB+OCZTFWMDOb
J+VZoLa1Cp8+xi/XW1uHXkNwJ4y0RfOQm9t6s/jae/oxQE4EuLuWftphVxyOJx3y
4ITTpQ7aagCFs05xFzC1ET9XuYT8MBjqzPq73XH0zGtcvwIMSDG/nHsoikEqDGED
wtWDAovq4qSchSXQT6MQWZtBoQe6xqTzIoX8lCKINnK728UuWSIR0zjqc4BlW4OU
1drecgnUk/yrTCGiznXyEQ==
`protect END_PROTECTED
