`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5fOyh5lWTVTmTi/ZTjj3zBfvbaJzgZZLscTcnmRpvzJ2IdsQHhT9tHYlMgVeOC3A
F6w1TfTVzo9k+3s2+ES01yT1sDWncJrSOaucrNS1LwIJGQ6SQVWnugOn6FMzGtpF
6EM+G+Uz05BJXSFZgd+WYltaMRurZjr7GyuYf+8djhpn+8DDQHEXQ6FHPuxk56Nr
JNacOVrtQJq+mp6/UuUMi9wfG4LOF8FbXrmdYKiYVCNkppwkJaXlKHWl/q7icLlG
JWB4vHQVgwqDQM6gi4bcD9KXhWyQKwpYa/cnrYl60ppj0EnjLxFf6tYHWKdCds5V
uDufKHsl+OtLjLQ8vzx5NFB+WAQYadysfxhzDHv+aBBXh5uQIjIM52addH+PBnkJ
RSpsC0isdQp9TlONVf4MbuxA7C5xqgbRwAoVtAcox4wIaBcfNpxLbg8s+lYoXX/E
`protect END_PROTECTED
