`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TDS4wf+ebY+u0UeJ6d0MaIFFIJx7HGOn7wIugtqM7OLoNNJAIJd8xUP/LbydOZnm
QemfOA5PnIAh1eGhHq0x6K6yP6k0fPylgZqK8YhoCVo0jVYMjbbUJSHyDhQmWDwi
su3LJTH06MVy3i5YEkcbeI3nd/UtEcr8Q0xkltl43YEb1yweN/2rEKkriYSOcv+c
kVVVNDqxSQhCC+LcLp+z+yqHttbK5AHmgolWeRCNyLBsVgzueDds77iLyuUInUgR
OIUPDBecckBYkpwoNH5Dnk9oFI9Xqij5PaSfWEfQcnE+6Ss3bY1XKUfctLGnlvAd
CQqCCYFq1yXcdk+IERnEBzs0y5bM+/x493aYnrHRa/tZKqaUqNAcrazjmk24nECc
R1nlhW6X/AeBRVcH/qOAGHbleJPYAbrGhoOU9/HEl5l9uk0sdfaNgzVmd4Fiaai6
UmZ1QxZtwgFqVIGuUfHWuIXxQ1xpbU6WVwfaYLO61AHPHOEzq52P9H37CRfX0erZ
QVLJEkY60ITqk05mRrMB3gfffLOjuXAqOeMf7Un+e75QcKQ6KR8xdxecn8wbRZX3
IQgxCbvyE98kj2Kkt7/uRDarZiqhnntwG5U69tPCbBoFhtW4DlNmnPNNwplWwANd
/gNsAgkG+Wk5zuPf6qkvodRiNzur4OKG0txKVeMPHZOXHIXe/ZgLtwmYUfnVMfE0
SJPSFYW5Sf7OAmGtTj1H2ay4zjzbMDlFcdihYByAnujMIp9N2rL0Bx1ALehXrvTN
CwkWn7n9jOjxlGpBmZ1Sw8s8DeaIgCYNMlPfbEa5H4yCejBkep6Go1C3vYSEzF90
a4bSDUwpvJmxuBeJyuMUPtzQq9bjnxkODe5QH2BMpxHk8hSLQ+Od+y7soFQk6qk2
8QgpgJH2ZTNDNlcNRQ7WyGqGu02e1YTuhUiWHgwxD/V2/MP8Mym44P/X/PujEWv+
`protect END_PROTECTED
