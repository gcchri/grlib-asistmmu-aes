`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TIUQoqHAZ2i46vfd435hBbbWsDbgQrQ+008B81sB9fgz4iyMxDYPZzS+HdE7GOcZ
119/YQ/k4N0v+Ml9cfNN5lHFr8XQpfdweBHlUzdSg/VuCuLGj1KZbymImVKFm+9W
qqPYsFq8eaDFmaPIwVO1cfasp3wpZv5qMsVjInFP/J43+4rng2QuuWNj8xelJ6St
2i7pXyiv3rh6itwv+46qM2vK4Sgz/VOODxzD02JJASU/RC4na6/eEsA++3xBO/mT
1MfTA30lwgV4AlARoCEof7us3hRFUvbUZGSOpL/bYHHfl1i6dXK6/mgwzO7yadch
xc0zFDvb6vwZXF/gC0jtT+nlMs538wSHm5MQek7pnZ/8221HBVSxaA9GIFNjN8q4
U0sLWvsZNpahfnX/6TSyNiLZsj7d7y97yAgF6hliH09WGdZJAzbscEaeixeco0hm
oEECTD0EohjG+9wNUsZGLlLlk2hAsxhRCZ4HUf0vP3lg2dmipKRvfbcAUu5OWc1N
Iz47d9td0wEY8pWOKfN4pUs6HcdyXQ1/np3zXQWj9WbdBhNVNlWJvV63Dkherboa
JGzZhtLIY+cKx0Pd3/Oi0n3eT2vyJmPdgJdYY3u5ziuicrVyCLTQFum+HriyisvE
MDE3lp3yhjYS587W9kI876iM+J5kjpWrmx0RGxOZnNy314kpzPnD8mpSKASyMMYl
`protect END_PROTECTED
