`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xA6WADCeIRSfWx3DeqtCrLCCy7oHh6dlxziKburBPODmeV7sItZB6gmL+71UYNsJ
J8mU9XY6JUCegdWe40dUMv8rB4cWfb1OI4y5tWZToFQLpJGTMyi8Yse4cI9NmHnv
6ZpOqN25N4jDr4anq6ykHld3bcPXhRdall1WJORWfMHiY0LqKLZna98U/Ai5I9b8
zocAAVEm6MdsqTF2S1sj4+2BEbF4DDd2g8gU7v60QQaDycFiGcQ8NISIvuXOLPT1
qkjNef2DnItPCWzu43TCShoZak6VUWgHioIFH8vlXjTQXniU74UIR8XfB29xP8mW
uvR3W1Xlez0n6vzkkun/OyDmWwaGhElGsd02gybNFGWQ//teiQoyjIYA+Hp9Bgdh
VH+NvkBIeaKeVelD9Q8pjQ==
`protect END_PROTECTED
