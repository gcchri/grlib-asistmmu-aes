`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sOKMHArErm6XtXgyQiqi56hvhx6iepU7XrpyPNTdGlwlGqi0M1d2z9SIPIeP/1Kd
EmKIWMMRvKDWXg3DtntPKHC3XVWalmqi6mpXYKbb+uzdQcibdaRCn/6ZHTtpZhhW
QnpkZj9h+IOg1YVcdcpDKBOSSkAOmIj0icoWZ7dzZLtRZyQJHq84FKss5f6W9FZ8
brdSaVxgDeBvsFGNILPfBOVefn3ABQfhBDaCXR90XcEodMBU3R24KvBA+1X6pym7
kGyLJKvDKkukk2i+IfFJl+uKgYfRMRm7Mi5LHp0hYbcS8GCI4TSa4rXxnVh4WpFB
j39mkWQlFqKVuZZASrwBSEKmMP3+DuNp9UpbLjsc1sEtmuLL35s4NuDNOcIXn6lw
SdSiCtX+Z9wwYr4byfcOJRte/AOORzM5hYHe+LIFCmeUkMt8c1ORLDFIXoy+IEMc
q8v4eZj5EmZwFxsNPUKgRxfBVYMRA73KvqyLypKYVeOJeT4QWgmTKSAPXIySOaR2
/mYvSY2X2EO6qLAbT7AJFSgxjC3xj364uPccY0L4c7z18yV/uLD5CvO20fdfNywQ
cGgHghtbWiRjNKI+jo1fVPPQkci5GY6/GY7p19FBr9eh88kFtbYGszBp0vr1OF+u
ybPj1S605EwunNML9bFAxFDeNLrIwiRaEskxkegMy+6SFH0DTQ2dVLQvQBp+DpB3
RHvFir8xSS6v0Pb3YKrzJcs+Ad5TOsPAzlOSSeq/BOlxG+GWbNTQiinF6ebnA9Og
DChARTunnHZ43r/+3bC9OphUEkTC5XXm+Zcuzzjb264dQFJvZMANCCwcj1K1kaHn
5oHow/yR8XnfSTAVh7P+i0EO9Rf0fzWsqr+P7o91EbMC+XsISpjgXpw8Agzg/86j
bDc09MtV8/tZ/dyhVysgyYVpJOZdTaB+qKG9s2xqrGtiitQmTPXRCAUGIlvUYjZx
yfJBeQdiBo3VF8URVtyqGlljqnyKPd0ZHARb/AXKPIszN6UOnWnBoabgZ3YACiZX
D15iokU28a4AKPGbWdkGWtQAP1RI7RUKreLEEaLoyCk3rJRnCl6MgLDoJ5Gc7UgE
KVZC1ibQsounqWcJ70SZVFIxv+sv1l0JUFBBvNoeKfRYpNRAK+oLsMxgH96060pz
UGMq+NYG7Wc2vElUutXp+9vPWPGAdGH+gTMaXLCGHaqLyvcAIRfvD6lM4pcV9QAb
ROf4CGs+5U/HLx7aPtR4Gg/xMVyz4LYdPOr1f6FxuS72edhamZpmDJOWo8HxY3bl
CnoB+am6/TgyAbCl+rJGYFW0BXtT+83QXTP7dWirkpSy+uJR6whaPCmE23mLzOJ5
w7LDIsP/i2aEkHk6utxml5fDIqfGS6u2djfQY214WH+Iyz/TRZ+v9IVxA38ipHpe
deNdATBzjYpD3Azi9XsQGhaUu2T+hi+/9/mxWTvIzxBErChjlWKL47uzAh4EsKiz
bWDffHqmzH/ASDx5R/e6W5Mza8kXvQ6o0zFA4tkOkgEcTLCy+6p9GNE3In8y5iiu
Qk+zDKsWItewIoAzTCJnSuVBXDkXYQ89qdgZA/TV+HtjPhYBoSntQAWEQX33FO4s
pFW+f7vJ6rMAebttDhWgLplb0MQW1BBiqW1yB7xVNqshlSIryKq+x1QTXwGaqcnX
RG/xN0ylvxHb8yUxseYIxXCsTCFpMJn3o5jcb3M9R+U5cvd6slw5seKOevFvF2o+
oRHlPo+okAMhdObGOfR1N23p4FmfuLw9nWydO2Icbh6nt+mCU/MwXF2aFNmOlKwo
Aw/48RaF6luPVi5/sssfDjjwfYgMOWQHFOfUjyOoGBlT5PaPI4OYX58Rv7JSy8Wv
ZgYE+/kItLX1IQ6bGjs2LxEhRIwBdK9m50aAstHRIwcvnAVANaEksxCnifikIimD
JYKXd+Rnd2zt+GoLqeko+AA5WJQR2zfTM1aJMRF8O8Z9KwZ+J5PQ8A7PjUMAgs+J
ZPGTCmbweIn8b9FsjNd+YOJHxQqD2crnLzGe34PE6tzglecgYWBQ0gFL3aW7r50E
2LlQPmzuAIMe7oQkdyhAhN+1PbVlQDdMEWHDNE3DGSnyL+0tmt2PRAuOERmv8IrL
cUgagLsAfb6LLiOIQ8qB/Mifa5vJxjjQmesoWIMN2vsQJNmVWw726lEspcZj2Pth
psIB7X95tALEASWafSnAAL0TWfsAVfF1OVWQAKp8yQM+6lOx3r3ffMM+DHEgxR+D
w+ZeCD8NovMN3JI5xcWd8rB3hb0sIFKcT1TWtlBVPplfzYNKZYk7qqTohFhrALtz
VKALw0Eg79GkLAOToGxMYuk2E/V6tOtsoc6EEvb6YGyFf3WYMEhblx2AH6S8Chlx
u2mhS0CdCG3UXA4cXvDLeUY/AP2RhcAe0SRWIbmcbx6FY8PPtoa/KmW+Rk4W9YL6
CO0aYugu5a9chX/SWngY+xZXXFFb7mBx9kDgZ6zz8S65hSPRqLI360tfm0gvnJbv
dyqzSg5LWw63s9YbrO8DzzvMJDoz8Fd2G+S1YcFUsK+1jp54ugVaQIH0UtPclN/e
67igydwQDWJVfI0zGyM2Sl/h4Adpa9qkkxAXqfjuzW9XsHvTkzlexjYhn3Jbcul7
rWCNGbrTME+1qRvFQ7ehPoTLkkrltOVskQg5tioYhUVo6PL0EkKkWBaWBUOTFQsB
KT5gHiN8dhh27Oh44D9JvBaJds4sVLORlcc7/0BQcg20fxC0IrxMrZDkXFsSVIvD
QHoUVym58rHstm6GF7CLE2KUVywNSOcPSAlVptatNQHuBE2W1EDMg0I6VNgi0ZRD
tUNT8f1JtFX8019vbl1yz6x97ZvOwT8sRJsTH0Bqcs6Mv2FGMG5dHQBDfzw95Mbn
fmzO/59dM7woqA74uezFfT3bEKO3pAwFOooiEuqNPRS+yE8zYxA46+td+IKSCJfa
AsqqALs1NvhVYHAeVi5b05FvKyPSH4pBQdTUpsziO2Hv7tMYFpp78JcQhYfeVwHN
wr9Mmt8QSEMfLBm03dQFCX1C0xUMBKzNc4H9HB5aFILDSmOrY1Z073IFBDTfXp8P
CXZEI5znlif4DVr8DxPrpJFrwfU/QcF4UvpYDbC8osFRIfnZiOR+hqIcq4pu1FTz
3iZY7cVct6PCG+UfjffOAyS7jhJbWSMeYEcYMUwAJcGO/xe8oJONXb4T4Dw4axk9
0am5lQVixQNnnOmS7PZi08juyCPdzVl1Ka1HmnoZwwQuOamH/EvuY7Xb2HSNGNAH
ZeSYIYjKV2DjmD0oCDYauRH+7DwG+QHvDoY3ddQEslGlKvOhtDCycRiHynYu9XYn
dFbLyBE1/Xh1uUVZyL44qzaFzyjWJX1bot0/R2pH7hgVBDxdfyBR5PKWtKpW1ae7
fWgXH9saRJTQl7O8CTyhlBgmzLBWQzlSxg0vMGCmx6oe0DYd0/p9VBGGAUpPmTyB
HSrJS0gez4/7dgz3Ljm2/aN8yJL7WWCM+4rLbqLNwW0vj8j7DJ7IFvErrNgoM/8p
OnuYMH1vHup0dbPPLPobMuiNIr3NgsuWCEOH5i3yKDpvFE9bZliCJHEV4Jv9GaNV
L0zYTwIRq/KWl9mbMdRAxrdsrUVVwKoKDME806Du39og3DZvkVSp0bIUnHMsuLnD
ugqYw1u3FPid8vtiMsg/ToC01yZ63JCNyAoF3+6f96VWOA7rZq43FZ8o7trROzfk
cUItYLe5GmRgqTYSUBWRbB4kgwyurHqclbY6chTP5/2/2Wp1sm1CosUQ5xtTdPJk
83gPEQpL8wxu7QTcorIaABcV8rI5uiWZcmQH75HzAL3zGGM8oFBi763BP7q3xORA
0IEQRM1xQ/SZZ1f0ub4SwsmIo1m14lGP+jtEXCPLZ6AJODwxT+nJFy5op/6XQ0Zi
Gs2PmDHCq3mv0qeGXTmqom/OkTD39FZIC0A2V2xPKXlOkpxjB0rWOJBi6Lk3p87A
FiRUPx52fudVUPmxJqg/Y5x07EXioZfQ6nmGzw8dVzJKgNiKruBaBPP7NHy4mUW/
hl2jw8YVVJmyqrEI95hAiulX+BKkOuQ1aAIlxv+kK+cqIM0tKQVCPsAPinUZUNtd
yiIRPIctXHR81Zitll3ntoRolg2Z2UZqUqeVkzFE4yfCBb1L6YpLUn9ZDJgjvvBe
0Wk2DaetKFXPssBeIhkmUtWlG/Ft1Txwlep7vPIudNikPFufoPYVWPrBqvyOZCNs
D6hsCNRAiA7k2cQTemZdgW43mkU6hmWfMSCwWpuU8TnDWiETf+a/BSGPkOnU3lzi
MdzgROrumdWwIA69VcKbyQXueCeiFAqkBRpxUXK+YUbFXUYlg8p6Q32BbxW5ruWh
25YPKy/hP2zvQDQtMqCrxY+tLgeXoKqiNecSD3MSF1z75BlSH4dmkExkeRrI9cit
xpmDYvRxqDC62EOzUw6woJaeYXCPA3WRDcx/Ej73EEMfphZd+4OpRs7ySGcvMbCt
c4HOWGoF0BalolAz0zK3iRpBmf2xzwL4TQXI6I3wr54=
`protect END_PROTECTED
