`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
acWf/yOF0RS/m3oPOw+YbOMY6B9CJ9flg1/I2gKeTfh7tb/okfvidaU3MqtEp7ci
ETpQqkUeW6kx+5JiMUCXaL5VKx6BHUDaOAO2R8F/7jhXrkNlSgxlfhORwW0mRoAl
aFGiGNQl64FxRHy28lMDauE028610ZjA0i3NFb/KNwot+G9GOCnAsBKNayAAn+lQ
515D7hwGHHjMnTshx8oS+tzcT4sxIpnCSr2KJ1lGOzKyuvrMhvzHfvP4r6IbYO75
5CaNUjj6cnoEBv11ZyOnlFivlMVwltfdPz/8YKzy2Kkr5YzUBQbNwNK1TdxMo4If
Q05QL3fHC7B9LasvtOC4klr5eQKEmI2GG/XbGqbaZiXD2D9b8o4dYnJtSBIf/VHS
ZjyL+cdbhBKLUreJoaYuj0C1HoEdTflFq/+gdvRhrgaJjZ69tgDeHPb5S+8UAg9f
sCHfUxYt9gPVVxtNcM+aYT5LyARBvcfH9vFXh8OzFSbGpzqfMnKen9rEq8gwOdAX
ZhoS8DOgC/6LMWAJo2figym1URJBATPgSjyJxjUHqNAyz4p9aEWFR64Wp3HM9Vwc
`protect END_PROTECTED
