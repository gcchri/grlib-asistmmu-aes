`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sGsuopKv8mcvy7UcULC1Gb+k8BKTnMCE6yGJb6jhYbuSTxxxSOSUx5NVKjWcZcEi
skeDW/lJkMgf/JdJR5FGDqffEp25zcgzWTtIapdk6fVk5ZgI4klxu6yHgsF8r6KJ
g9yhvsvIfy8x63v6cA49l20KxE0k7rt9b4jAR7Yc56LidHocBgG5yXKz4Iu9eXsJ
LedFt3Bu41Ntht2QaRcRHnEup1Ye0q7IuGKgi/ERmUTIwcB5Eff8pIyBg169Y8Y0
NcD8AUYUzGSBSPxeS54IpRt19cO8XPbO++wlOWl0NAt3tq2lCEb/TndLP5GLz/kR
sfZ2gBjj0Z4NegVEIf3KqATkzTGw+vzgPO26eylFrhB4Li1pc4A7RNJmK1EJds6g
L4dvqgJjxwJDauYdQvZSZSHfOi8LaRPpv8wFcZj7Vk88NgtP4zuW538AywQ43omh
T1bg+D9i8Gy9UeT0Tdo8+l+5KlL9XQN8TNjEnW69iL/yQAh9Oprghw7zEk31DhtK
`protect END_PROTECTED
