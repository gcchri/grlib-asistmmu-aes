`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H8yR/PoR5T0Z9Y9TFRoU6GvtXc08RM3DnyEdoRkqJdRP1BS7rUEo8r3KuU3M9phE
IQkQ+fCO73wSY4fJQhJIusLQsXDU7bkbVwto/Fl1V2D/P2hgdX/r6LY9Fvv2Jbne
YfpKxHuMdRx1aoEbqTlydk+omIyzDPONIcw96otGaZkn1LbKaXMIGRYGXnsSGEvB
Tg2QKRx3e2wOY20xNeDHR+7EVXV1WCrpl2tLcoQ+8fxzkNfVVxo1LirGoWZlSYuV
icNRVQyjcwUXe+UuuKU3tF4KrHOScdf67DxsLoBDGWyFu/VAOcbLfiCE/bh08rbB
HfMuZm67DTNus4lKZ4VfjNhd+Q+eMjomSaFFmFrd3EDUm+xXy6GpHlZeHAhNngpT
mLWsPoYIrbUkInBQTne04GFw3P9j+PdrQj3hX3OmF6ruOGqGZo7xLn5PGlbk5TX9
lCULjgsHXSvwYeeoDCASyg==
`protect END_PROTECTED
