`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1vtMM6kMchB4yFeVbvD6/dLImkgNYWLsYv6YSfqc2q5XWnKKK30N+1eIDrjv/BIN
M68z8CfckjRPtsd1GhFW7+52thN1GE2pZc8iefkP+zc4O7NycC/qNeCN54HJZUoA
0gtYIXHr7nePe8TOpi4xZc7dPLrT0RPiEdbOsoHKyIwNvGgbo8XHBHp151PL8XLT
LW8EeBKKTAhSU72xh96+XixkFy1kJFqy+LXUicTykkpldWApWGcilX5up4nnsUiH
QfpaTc8qnZxi40isGG472w==
`protect END_PROTECTED
