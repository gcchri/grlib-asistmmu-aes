`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rO59ILh3q4qatu8uijRYJFEWCg3InzATeHCxrXU8XbtqWHujvVDNtgEE0vGcRYsI
svgaOto5e+2N0Zuc4agdkQlJ86MlS4R7HDqP5+0n9yNotb642RnkdjTUa3rI0u5E
kb9It5PcEWcuxeEy1JhJdn7h8oJ/rocj8NOSbGW2uUr7qdzLKG/e0oZor376UdUh
bhtixpvFtALxcxoMKu6FW48F2vT9iY1V8gwLF5kqI7ZB2/Ye+zrcP+v15e1CjKGz
Kd2LXZO2kGKPoVOn1p+i5iZHL3k+Ix3OxvMDwzmgREIJis1IkN5wVzwcplgvv5/3
M5YIvn+hDUnO4S78FIbT83W57zYgW8qmaIkUC1kSjNJvqL8GFvfPMAKfvp3dgxkp
TUzspkRziORDnf0xfF+zMg0TtIZl0L9BXYY/hQv+8qslS3mX13Hhyt+HcqpoYsYo
XWB54jB7bwmYSf00h7rawgXSX5xqR5y5x4KkgoJ/kVm5XMqPCyBaAqKOhtlUOtr9
ZDIlksUsTvrjG4WUlNyoWg==
`protect END_PROTECTED
