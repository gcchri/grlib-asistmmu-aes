`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oLz+2Bryp++C+kO7xkZ5jenRvehDjJXnUcA5eMHmJsYpFwp7nqQ1n+z8lnwqXkF0
VcFGJf/wT7wvpDSt/umSDYJBZLD5hJ7Rstq0m32M3lF/hhJkHkW17zUz8HOi2FHS
NagdRQeuDsZkbT7YDAgqwzt0tsqNUJ+JZZ6F8iNBRbcyxMc4EuLwlibvCJ0kinat
imNSxJ9nHvtXWbwfBz2v1uw2Nu3ULg1GY19qWiDEknHV864pG8eusMbRx69+jEYq
jnuYBEXMSXGbzqw87tgm4M1a1fNNYj3s5f49b4Ua7iu7dqKffCjMkB75a5uZuh5F
BTsLb3LiqsY8RlXyUXdu32R+B9lcgSKCwbMGmcVLshsudcwOgw7Rk+MZmJMLRfYp
CbtHucGIWeVZMAdTh5+Z/uc2twHdc6kxInY8IQ15QBGcoQj+7PcKYKLbEq4tRihj
Jg/AQRcFbHE98QMUCMRZeLanQquy7HsXUtiHTzzBA320pP8+OWY+nk+3Wjo9xvzO
LXltWKuHINYOlr7YPD5IIdzlXjS9Jy0h0gq5jPoBrXcrEFJe8hcyZ+uVzxQ6Cqjn
UHtMk5otL8fyUg1CB7zk9M7K2p6o+YvgZ6FADR04T6FwHKNb5ThWk/dM9XqUERwz
eBzttm+kyJGCjjTghoOk7no2RZc+gDGauqQLxC8pBLU09l4dqN5LKTfe0KVIsKPh
qewNDSpH+k0rm1qlwtfa5SYVq44gu/rhBkrfHnvn+NJ6uYxmywsui5ZtDV+6XQK4
jswDm1XDZ0zxJYKw+ab16VeV8JmDK4ZthRPZ2wju7L3q2CKv0cQq7AF4sI1iq6ss
IvDqWKzwn8vgJlcfs/7tr/tCi634e0bBfMJ3hznlZATX0l/qvKqjpYJjKgK88DWT
mHZAjcFeSlTUcYSd5iJDgg==
`protect END_PROTECTED
