`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
seVaI3q32dju1oS4lsrBrlXUmxZ/HsC8JLMvJTwyGVZUwPCmD+x7sIM6ssxPlMYJ
Uwp7bvuK0zKEmD6YeAMpwvNSXHIvy4yIDxLCLZKVCeBLUN/d3ENQ83G6YEN2IfBQ
3YqjUDmg+6ltaG+ZfWiqaTduuxWZmGoLGnnJTMeeE+11uGyqV/5jEYCOZw6T8lOV
FH/V3cZHbwU3DHKTf4NR6WS6A3ATPhel7CHDf6PIR7Oena6AWp184zSgdQ18lg+c
Douf0wctS0AryiOt3vR8oLps/UEcmHvt6BXe1ZH7E7KEmHu5n2+iDYlCxapfau+b
Q3g2R4WmY7zIBLXpw7sxHfW9bpFWvyU6MWH/viyo+FRl7RUO/KQVBp1ZVbdPIWJn
iAVUjn6Nmoo0/16YTjbTFsPgfOInFVywTz+9rmHoaIpS2dhiuFEsiQHInvlOvdby
fbykP8jZRdqQ2+2baNxY8r4IKTdsC0r40Ih/5//+hKK87852XSJhyCDt64tGa91G
`protect END_PROTECTED
