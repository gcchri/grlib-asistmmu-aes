`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sGVVqcgHl/uPb9DzImejr1zaA+uVx21cBoAd4o7Ps4y9rOBLG683rysSpOQI1H4U
si2NgkspvPB77av9WchtaMtCE+EK99kmGp5DXNDUYre9q5v+hlodOcLObndECzas
j5fW+pKADKih2kOE88NQJQ0v7QZHjWAUeYwIbNt8VOYu1+uh+CsdDusm5NP6ZLQ1
AeF1gFXTx4yh5jfVxjeYcpBVe0Z/9RvjzgT1PPLKUrWGbmD8PQdzhN8Hz4IYg56G
u5IUCqRxthG9fEhcq2TNo7+H3nopcqx+ib+qsB2fM7r6HQ9GS/rsin+btFeUFHAS
VA5Luj1FH1mqHhNW+L2kScsb9nvEViUo7M/klZTAybTQOR+a1gTuHhxhYGwwL8o4
rj/D8x+g6XCBaf/+nzkq42mVvq6Pfc36tWHCtCwnbJtfSG0aGmnfoXpQQGvJPqqd
uP78ufbj/h7EcEVYgkm3KsTX77MzYiGedtVQFUBuekx8sDjtwQ60RF4BtLBe5d5U
`protect END_PROTECTED
