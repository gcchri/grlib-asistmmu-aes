`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GFPSRquLLnJWIC+4JH70v8wDHry2TkF3w/+WWPDCZnL5RbC9oAH0RbxC5hNU2rzw
ZWPmPtpJf6F60tZD9iyiKzMnkwrZ4TcnNnvXse8GvMBIUPOwBEiBRlktemTffjL3
rxvtcFRs50r9eF/Ltx1mP+jHz88jC4mBMaO4yFFvxsYsi0AWgjzO9XHir5MjfWzf
by78ST7747lL27/4xVfUbyk9EZOB9iF0V3aoPJfX+70rRoMK/N5snd7LCbbvZb2b
Fc7Uv5G1LCAiTF/sdk+C/gV2o5DumvacbcD1KFGWIHt5BiC2J+p1u/0b/F6o3A2c
FqLZqMMTdLIl/c06FqKXx4ZRyM9c8rP0b4eJICWe43fB09GIEPJu3wy+0jVq7vcX
vC8dXU0MuNYuMZJTOIGIoWIf1s432PtSkuSkDvExRFa/Y+c0QQ8YDncOLmOC+x1X
M945NAlvOyrTF19VVBXprMzn2suh8nVB0auxsmQHHQl+os0X/cJggdasfW7hfU7K
ajuFRR2UIWy1BzTGpVosAsn+Cr/fwmDfH5OR3FLtIZ0rXEWi22h1bWNKohAoXcEu
itISSPzxxaQ+GEDyiwsJTteoB/BQHOHOt8NACSzWJtDh35Vkt4myUAUlHw/euy78
wGzVPLcYvto3zksBdhateYsz85HsUx0yzL4Tim8KmU8kvEQF/Rp0HmqjNEkM9kJw
Ur7xH488zOQDtxt6fwWspbaUvZS8Lq6uexMTtMkCjrLx1HFvyUKZa774hKq/JTy9
fvX7754Ey5WkkG+LCOq6+BlhsuJpHMnnmMFZ8JRq7FD0e5ZXtZa58g1+c0spCtNO
DlZVUnF+e3o7CnCLrA2Rf2eYyK6sBdn2GZyrsLY9wSpBuCKntxKsYp6whh6zl1Wh
1n1tHaWPkmcOsooitY7f8HFUSx52JDPLFnK61o8F46E6S8Eyep/17fRIiB/znDuj
32zmOCbpsUiHVykpnKDclNBmO0NOdDV1Twf+k7P7YaXAcwGdtW7O9vzsvii8JfuB
u0WP4BK12y1w+huS/Wny66qi8JUxO858X7MU2eeLlMPTrcWmg/Pdwy/aKWPgJlLf
xnWb9965LCwJEZ442ByE14U7i+6+M/Iw9DpNsIPtFRXa9NQFKNO2ljkLW8zULpYc
roCDI531LslMoHx6543v+n/TWs/yCZlPdQpCvd4U2AuqinvuQbIS/ouI/CPNkye1
L5d9gf0iGJfC6CgbV11yuieZ9PpeX0BtJFkeVq9+LhquwjEL/xNNvkwBW4+TJlWp
WjXrE4stL/ALN07iIXkwBlo8npJ7gipYbHxDYG9paVjOVKbnVi/KNKKECa6l6IUB
jNoAH+V2y7vUf4p1RIZZyZ8cF2zNxuI3J7YNofdj71tPRRMm3jsv5h/dgjSAnEp9
nOjUzkrtI+YTXfcPoSHiOd7SR+89ILTR5iroiu+saGjAhjmYsLoRzP90HdJc0dg3
KrWDVti1vfFOwOaEAyk/nyaUQMQcIWaeo9aQCqWrPog5vx961fQ3cZWFs960dEXh
JKnNHDgFUUzEZ9ola9UNcfnbRL3NNZfocZ+3/OBXLljQH/r4CgTaoPGFw+23T0z4
`protect END_PROTECTED
