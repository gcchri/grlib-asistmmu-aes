`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uADTO3VAb/D3HdRGyALNdLO70Qhgnogl6ohHhwfYIf0F++NGFrI/qGUkE1LrgabS
tvvjuO4z/fowhpstPNlLnIApCQNAnQY2sdWUTcSw6QpGq0QbxhuqGY4rCRCsqv+9
PRhee65So9v2ibrXikgq+jEeTHMXLFymgd9Sc+x1/rVP9biH2aiRciAP1g6P4RYb
SoZR66VD5hlOQiOlIzJr3wJ0WVL821iKzVqSFXHUe3EWmRJtczm6ZqQ5AnBmz/0a
+yId86nVd6bQWAAyVVb88bES2nRUcCpvDlCvWWHmKxLhNDP+fdOG6AdbMbkcwgjS
HLNtYQVW5llW6Ni9Bd1Gc7nTT2sfBctqGf3Jo/6daVkVuH8jV7f47rFP2OiwzE48
grtmurctBT0A8+emVjwPwyyzFeRshlqRgEHltu7GzQJQ/OCuhebHfCFRswqEU6V2
I6AF6EHnHEJBlJU2ruayyAM5H8y0/KTTk0S9xltZlgqcVRqjzy3xFg32ucw3NP/i
WxUgahD5LVd44PdOaJpU7CzkS8g8Xq7pt3IwrwHyTxITnKYZfhRf0aO5QmAxVB+z
Pcht/CGHISXSk+ORUPbfG3/jmDYszP6TFnfLs7qzhQNY4O9Lk/IrfCzeCjBSn6ks
cr2H/sCYQilnpv2ohE8kUdGc/LlaZQa+58rHRvc9yLWviPslHSnVaL1G3XQU9Cz7
uMFDr1mfWBGY9vIRQS96akIrbxetvirlNnbMkhIsaBTvbstytf+Q6zBp1rc4LFoM
Bbfj1h8hnL3kP78c1hPrdJ9YBuBrc3Og52ZdoibsnakHKTQaVieVJHirCk64Gtev
fhanhdk9wkvQ7jbKoHLQyHBq4wsSh/Tvc9MpDAMlMA+HmNW/hMq5bjHB5qpRYf5J
iZIUoASVeSvihnHtZ2Tj5WTejVxcaeSjIRyn5rf9vwWRszyzuEuEg4ZFPO0WO3aD
LtkjtyJN21ylXLn/4u+hQkNWPBrN3SntNiu8xhpyRKG2JVgpyQDez0YWquAlW493
xawBuCQYauh61fweDYliaQMr4llgOLhZ6OmVF+GI6ulcgD9/zqva87nVEq7d8I10
QIGZgU5edLqsFHLjxNF5t6nr/kIZ2FpNduGv2kDeB7vsN58j78otkQC3sEVjSUC5
9LgD8nWqJoCmelpQ1ME/ApatX/guguWr3OupWywm8qMduL/xZ6mt2d38aGSjl4AX
pztFxyGdOYlyUl/XcsEHT8CxwFvjRO7OdCTEgKWqfFi58LH16ZTN8kxKRAMVuHo9
uMhtjW7WSZuAQaX90pf0rAyr/rafo7SqBEeyB+akIDbgEyt/MZ+gqThbNcQRAmr8
Ga2JXH704Vu7N9pXpbID8v3mazII8jcjQPbjFmOQDMpM6cWjVeOyTgfXh/lSMAAb
/oQsW1JM6Kk0z+UCF4AhiUrkXarhczHVBws/0x9buj7NWEmXYygYvSgnJDcgL7wK
9T0G9yq0CSELsCNx+QIlKamCvTVBt+MoW9joTUCbGmGIbhveJ8n5SagXKQYq4rw7
1++/AZuFVvgjCpikyz2xqPIp8jcM0QMi74BHmYUkRbGq139d6QHr0C1pyaEJooX2
Q2XciMCcmZxeQc9giR3BZpouviOhSRJqgBQjSmzBMVq5SEYJU7wgnh2WLusv1JiQ
g6376N9SJobNPxgMlfvZ+6gzTWESZlCcKc9UYlj9TbAIUKVS9rUL32AKWCbKHXWA
9Cx4A/d1HV5u09oT1O4gknNvPNjsZPcK53iN78FlW6ibMn6+AFPTDTQailQp76Tv
DGl27pMJNZXj8lCMDP1H7VqKZjUmje9oE1k+5hZmbUKwvzduTb2r485VOS4u4DND
cG7UdLR4JNBV1BYN/FTcR8/CGSF2MzD3PgR4Og/b6+oULBt2aiIHWhv0kaJD5XFr
9sMlT2y+9BhYcQC6bxobgnxh8YZOWpeJooTgkjAi3jxG8XcGbKlBicYo/q/z5z9Y
ZDmfa0MqRIJes3fPNKMDU4Ftq8URskLhJKN4hy5topV/m8mZGweuJfzSsOYfHfp5
ay/uvdNwJQJAKhFzr8fp33EDehJxBmmnUrG1E6PEj2d1HbsZSxnDVKN1DOh21TmF
xztirpv4c4GFXCNovmPJ6UpQD0a0Yz7QmSXCH+RBWyNR/9na2MqIzxJjrNLKTWG9
vOimN8OjgYHD7vSykj5TPeZdj4FmTXTtXPpHlR0VV1NIFEutJ5C3ifWJZ8j9QMlN
DfADqB1SZmkUOCJJJqERuA9PnTI5I83bW8nDNbEw0lS5liPeJoKVsjybU39ZMW/x
G9a92kJ6MmDfurXL3aDfxiLyLkbtKFhXr8DUYpzp4gdPQZI2Qhg9Px220OBtHKxH
WPv4Dz5tIZk2IkXt6oa8/qAkNhRYL7JygQcqMizQ3//qZkFLHI/rovWh1dmdHbZj
pqixoaLCiot8WMy86dDFbg8HEHnz2Q3MxPnaOL+XAtNdJk5QETB2Osz60j3p/yAI
/98QDlVOy7HI1tOPJx1Lw7geExMGC+0Xnhx4656NS9DHDecQoECXHQ1R35ULw1Qu
5Dj6sh7iUxkvlKOdrC+sAjoow8Jds9PNLZ4eeAvnqZrL8Jzx5NQlDRazVHlPljK9
H1SyQpLosRgDxZiCCalUDf0k9xegeU1pfS8gmydk8FJZjBlTzW+QBNpYo5cMWgsG
SMjI/76ABMTOFQW86GegKSNAwRz5FJFQQ6Qpyv0AUIaA9npqduRFjzcD1txlLqss
fThbtBRkGCWwvHJ9LQU/wlw2QToeMmMftodlt3p4DuJ9CgW8ni+KznKth+76r7h5
gK+zooK837lLNYo6Zl2B5IKTH4aopU1vfdyzS4CjD2aB7LmxrGAFfB14h17cGBXw
Y+ACewuqGXAil3pDty9jr6b2mjdof98SdroI+awRw07Ufhr/iQz+Durs0Yv3W5vc
NwoT1Us1EMcYCJgOfyDeDFgmiNfro9WmcGsNslO90r6QgNmoMh5Xe0gE4h9Opk/F
A3whhiIm6gt0iSmmLmIuYWY8bQ0xM4Kgz2+LK7VDnHomVfDlS4azD9lpPUnNMWmZ
PHdsI7thXmDjJGYDtiaQveGN3EGst2x5zqAUzLFzIcY+ONTtTKVouwN6CtqiJZbS
LkDW3+YKxSaNw2IhiSHWVpTKX0uQ/sFO80SunQ3YQ1TYCJfTsMpZvwgKCy+5V4lY
LFxZuk0msJHWK7fBPYvu/YdYFYOrK4lnlb0tZe/jj1MUWywQ+qFwm+pBgKTiYpHu
zXOxviijcrUyB1rzN/uLWTVi0m28PERICdxj5ZsJ/GEz/UKWbuNY0WULyYT/hqqg
zdjsXpgHX/K/PSC6iyJVei7zWAA0uYy8VNHXgST1A1LxpNPE72/72ZO7BHEfx7Q0
`protect END_PROTECTED
