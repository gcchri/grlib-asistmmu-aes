`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9EL8X7yifjTjy/iiJD/e1cBflRhASGH9dxlt8LnCEurOQ5FaqPvFeAkm7+yx0f/5
Id80HDTD/StGm3eyaSsRm8v7nwU/nnq174gYYv9ZcrBtM+YoC2x3eOX/08i8Ga5H
Zbz0O6f1M++WFm3FP8N9FkXMM7gEQaV9dGdjmNOAY1/MF3iGo648pa3d7Ow34Y2I
iegVwNt7wpm/EeQqD9TT972TE/B6tZX0dgDNg3e+Bnhi140KvWv46YSgGMPrIm7I
GJCpU0UiwcVDoX93ap+uR8LGgNiMnUu1WKF4opTBK8moxHwKkKc/ihZ/iTWASmfb
+LhBRtzhraDwDnHmdX3XfOgH4c0j7iImbVsxzkG3jWHgUK0pnU8cdnW7Des2I9IP
i1rU0ragDWfJQmKg5rGHUsFgtk7E6eKG2MJiGlH9+9VuTiG8UtC1f6YwyJSV/6Zn
absL9xfXideeKBjf4umv0++Uy07Ea5ZA4j9jtscSj2BM1uLieIhAU8LOnfl8aDPx
kTJo064SxRHzCgpSGKPxMK4xMYl+kR2jfAg2F70hg9lkpkPRlv5zJv2VtL6QS4Z6
n4vL64hzirS4i7Ztmy4UMfnGGux7OHfrTSuh3wdi+3TvwdNWfWjpqKAZmvohQ0pA
9qtFgtEcXzlptvUAh9hf+Q/al6QjxslNXNvuoc3LHDUAoS0X6WUWta6AxYRQ3fy6
5TIt4IOWNxD3uFvQzwFrLA5ZKczNjNI4mYfdpiu2tc8FeBRzHOEYrQOkfzZDGNsk
wL/bDULcW7Jh29NOMnYhdWLYVLA1n0InHEphGjWsYBbEJnXfKOnTbfoH+aUwaTrz
55Z8xp/bHdEcISPOjmu9UxVs1OlM7NhKTYvlL0/VPj+YswbMDrWDxDLpVkz+G/Ml
9pJogku2RHl9dzgT/U6zD/4BWxC4IMdCYruljQuiJjcgQ5ZlH9h99yl55qobU5+X
`protect END_PROTECTED
