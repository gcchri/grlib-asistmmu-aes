`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z/Lp1pEMSWafHDkE2TtKepql9pAvcfnNhI4wAM4wDYEz1k+W1Ah0T9Lw4enBOKgP
DRw7uZIySG5GUgrIXQg68WD2hhtGqftyqp+9eotl4z49863z2h7TNVStk6x8jMqe
qRJL+q1DEaSlpbKH0X5bRwrVfHekjyvvBwH64HDHxdVdEBsgRE4/RFWpzam9dqlz
F/nehKa+MK+XfvOGIApTYDitSM6STIL+8XqcyC0yY8HIpV8IQfswTLswy3IFxohn
+uJZ2vX579ZwpZP1dGrwSDn3/zQZNd2Z+pArsS6dmOWqC3hvlFJknjZ5OkKpmFz1
4vlAa+lenZbdhKR12yDYtEBpu6QJ+3lwegpuuCQHfWfMMd8vKAit3iZqjeuvjjWu
JTMNtORsrGrWTiOtIcdLYvqO4AnLa13oYjWh86m/TuGMQ0xuG9r+inANEZh/N406
s/65LqfHr/JmS5Vv33ce0f2QN3j83zLnYUEXV1bGE7E1fv/bBXhj1INqjOMHhIAd
QpTK1I4P37p+P5nnfoP+49WCyiKNndSHmXEESbE9ghhd7jZJYh+jZWTkBMOyF7zu
rDzhwlSdz2kuG50NQzQkhu5Dt6iVQBPoU4omdJ1qUsttEWSyWkzw937X58L0Ddds
y+PT4CJHfTjIp9iRKhjLO98fe//BgOCzzooda+j7FtCd8ijT2AIGGotS29ZrJLbs
U5AkTkg4HEN8ayETIuJ48H1v07kHogQO5pZ2/mLX0PpRjSc/2yr1D2RsPJ0df5eO
17a30sChe/vBhwD94lzs4qlkYVFwMi1TbcM1Qh/hjpUpWnw8Q9QanPXQEVWng/XW
aM2FnmDKBOyN/HNLkLoheE3WRUdwV813Au+kbRaC/0Yyq3BWuzQaGu3HVHvXq6UO
evvIy7lZYjgOlb9OaziC7pnf6dD5fcHU0X3ZyzaUKhPBag2NRba1uyE4FOI3idiP
QAwc8VVzpLIkgBZIVJSVKLOZkVXV31BtKAdkhlTTqGdJfuxBY/NFMIiP3GQ5hozD
nA/zDxt5sONIX2wJOAAlpZBvq6vvpWZvwgigky4PGIoS5OA8PZ2irJzoqOyAkgJM
9bsyuWFckLw3p2fzUn+r0FdsIKSKcrhoPzFD0a2wK5tYdNOt4bHvzkgzD81+GEob
rwgpDxJg0m9GqALl2CCZg2d4HHgqx5U4nF2DvZEleYs=
`protect END_PROTECTED
