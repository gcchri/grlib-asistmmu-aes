`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
btM2aztnUkqX6cNpTCthrsU/8wnOyH1ThAe8mo3mbu+wRJ5cSQFa8dbFVFREX1kb
cK5BzG0Gqc8gSzTaRzxQLn/TUX4m9eG7kd1zjaiLo0gHvskkev4+72/spd0g8w+4
OSwsvPMGpHCTT+XHW1QlrsQTPAIKHz0uXGmrGy9kOFjhpaHVR4szLk8HhgVCXbM3
qGcUJ3JZW9tLlo86Gb6NohIxmb4hDQcVDbtfurR2VoabPpZtbTrPMYUhSdijaBcG
kSzR2AKCrA4KRY3MShTP8Isly7ffsktvhwss2ZlrGSu8gT5qbiZeD8DfVNdJiMez
67pIehlKfmPgajGbrLWP0OylwgKmmao+HlZs+bq0xAq0UqvLYZL7HOrUg5H0Sfof
O41N4bWN/a5kPW5nzfKG3Fl0p4tPc3dTrpg9+22X3xFKp8A3vXJm8gxQDKveUtK0
YCd2TSlyYXm1MNEmXQWjdPxx4enECsNruB/+DBUtwLqyc2iX/rMrPu1ueMJa9n50
tIU5Kw9Xk+bhwmzWuGFEP6pjgCZw3P/WtGWBkBzkuvo=
`protect END_PROTECTED
