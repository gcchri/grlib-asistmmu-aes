`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VeTnJaAsGdeY1WhBLdurON8tWlYDhibRfquCMoUiyPJ7GUxVYnt2du2RorK/mX6g
ZAboCJLWegknRjwZg5UvVgCUlR6/RK69KO4GXKRPA4um++60eGG9/x/D0NM4GUAI
wYwoBx6wPdp7NjWOsSPt3DMmtD8qSv2y7FiW3ZPOVx54VWqD0Cx5QhQiOFLIqpzq
lykwHUr2CB8mvh1UGStlawgNrC/Se/FPYSF3s/Dc1iKMB/7pLwePIsJyqNrPlKDB
hfoPapPeXEIyzO5dGDBMR48pFMunckrU12xmt2rKDkLvsZKyI1a3U/Q18qgllU9d
rtW2KarfuYGQfMTsaLk2I9HYrf5uPPe9i1HIIhX5CtFXqussm1BAukV3sAWyz8QE
86D1oqLGVndjCxzBrcYJlnKFQEnl1ajI4D6N8hoEq9Zlx8Z99IbN8RHJztEVIMgT
sl2rJQCCoyGjbcl6SopdqNqQkCvizYK6lSa4FUotpV7ahjOOhwt3gQYNQgY5XVhk
Pg0PeCNA0jlaFOvkW59bsyCNcm9J0gLAIdOtz3XaCKI=
`protect END_PROTECTED
