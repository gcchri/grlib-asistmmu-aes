`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FYO6K4fHrp1X21rTChCeFCrbUXhNcaIjXCuFIa2bAgMgoy+4pdy9LNsJzeZEWsTl
kSPirfWI4wc37QmmeXDDQONb8XC6o+D+CMrpHxPUCC3F336pvOlIUsmPeyaGkd1O
qZa/OXmMNoBlcycKg0hmfgNVRS7WMzHEw42fHqOdK5ga06dqrQN7KUGnVpUrSSAq
HcgGwocKOJDBpp1wbv8j82uF7vk1sXsji0lL9VK10PXiuAtCfzmCoCrEUIRVcTv5
z8Zitp5bTYOHp/WqBk1gHfBssFk5otOlfRqM4irC3LCWDnzRzrY4LJHf2PorOJbl
ZxuozqFQYALw4VDah+A61g==
`protect END_PROTECTED
