`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MK+ws1eT8dIuGRPSNRob3V4DBbD2yyWOd/LSvpbc1RukcM8tXc4sJVGMqwcF9/ud
eolBUS+IAx3Qt19u5T+6Fhuw5uzXUKokIjTx5eirhid1E7DsDAPjaobvGAGTg6+1
y7q0EhTr8uke0MeG1Ewhz53dvXLZcro0GwIsFF+Qm+zN6SarwfKP5QHXZ1lOAIFZ
waU13rLTXD8WQHiO63dT8zTaUOPQhJSRPtl15gsvVywCrk0ShhWkvU6sKjyMsjC4
UXgiH7SPIN9FofDZawC+HMG544OErIqa6e9g+PClI2XTKCgDx92YS/dks0g2FNFx
zSzwgb9Xp9G6Amxh/903fW9buvB0is76Fqqd7/256gMr8n7Xpfg3h7Ln+zNz2Lec
`protect END_PROTECTED
