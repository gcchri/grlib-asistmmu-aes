`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o5hj4ssVxe1YrCwKkmYpGBtwL/A1vK/zkvnkJ+/K1SFHqMP9kEw3ThsQzF7SKU37
hrTraKUT6Ct5hHB03COc/+4fslCEWj2iChBvXm6eIcQffBYttrDOFT3d/7kSqmu0
oqPqlJaFBY/dhe8vJrjnlrZHp3epA9PueY7CkAT+bos5Al6usg9LDtdzd1TgjpFj
NBTg+ATM+DBF9K1RPZsQvs5EudNnrcoU3CYJPX5YVv2T3cbOL0qeJ0GFhPf7RBPb
nKk3l0901SICW0YcajIzCQi0yrA5ANNhoOWLKVhUWFoA/VOAhyxyC1GvnZLYmNHs
9GEp0BOQLGPyrDwJCF9v6hMNicgNHFd955Hi9z/z+sGZvbP6bGvvJlc0bXlRmSig
Dm8fZXk+7E+ls0zouR63JniUPZQad822Zo9ABN1YGQUOoa7QDj5L+RwlZOtxSp9t
KZZ0ghAUT+OEukmyt/9gp+6Wn3la87+WnunKOoxM+KTFTR/HuJILwpULml9iIcNI
HFMQO7oBJSSB2ag1eQi1RYyXD6ga/lGWnSEO3Qnr7HoMHatsZnlZOPH/goxoXq9B
XQKq9846Px2IGH2lmV0G/pL47+P5wE0Y5m5+VNT304muaS0MWav5rB4Rm84XG1a0
ziAHeUMMMazD0v18U51SxkGTFsODUmBX3VUi2ycYfxOH7Z/h7GFmuNsJpcvt6dCS
zxVX0CwUzxXdEsEbXo77Iu61I6KVeLaqCK0S1NQ3ZQTXgYHgjo3xANwPGMX/Jnbe
p+bzaeE48AWO+toEL2k8q/puwKFUszwk6GjQKEXhv54287xlrCOY8fn4hnvtnfZf
PEUH2czPWvmN2ocIgvh6Mz+VS/2V3xR58UOl7qQViwUJ2B20bhaDw52+wIvbiyIG
ECy4WZHBO2nohSscCrl7wM4kT6fEllQm6sDykgvEu24DzsBxunOojmAdpSUwnKLz
abbdz2EIClol+XZghOCbH1l1gTu20xpcGwp53fZArUkdyeGJ3kO6JTJrjro+KPHS
eIJNIWwkGwlJ/nEdfCfFNWe+Oz9PQdrWJTnhpdhGij7tbXKswI7EATMyLawGUx8K
cKqC/sZkGp4ycdAeVByaVJnxufSKguPI2XfF7GLpxwK/NwM9cQYKeBApw1wb0Zcu
O5zbVmDYlEsOoJBYFzSNLyU4AErOWYcxfqmwSSeKycR9mYFKe9q23w9TyQLlE9Im
1EsPYjzZCEw92swqEEQcgJIANggN66Y7XSYVrmT7whfZJ6KyPqmlIF+iI7YNVVK6
t0Mow/MD1Hl7pliuq7n4EzkbwtvFRgjqNi4zPy4o/9VPh6keEjV1I5dwWpm7rMF7
CheihnbBYWuLa1edDJG+ybHGIUPYWyY5F7/jDgNp02pkcR4C2GMRNXS3bpsX9kTu
giQJHRmUFdK8XNITqsm2uZSitrFhzf6vBfsgnJJOM9oWBfsQ23DkI6p0iOkv2x6Q
ssTX9k0dKzsfqSakhU7dyqZEvjVdjrtV3ovzvCPFEgNz1iNNYQ73F1L/0ar/C4xT
QXiXIw9qkQJOpjtIMdI62Q7Ffo3BbMB++1P3/pxJaT5127ZkUPvGocNCFGr/1lBN
vxbnZHEislJ+WmpC70ESvbIkx6ZE8MEU8pgxByXEUP3F/ztSMfM4K7FwlaOnLt2x
QU9rdyagtdfMiir2VQqUZKJiFzI/YG5dBkPbeC42aUWK+LcHbtuSBMdataOpX+Zh
t1uRF4dETHkA+2ZP4BlUvEJO6reBvicwQDe96udhtnDQpF1y4yW/27iGM/nuY63/
udo3uf1ti8OktomMaFnnDpqrpU2f2/VzTAIOPKPexqKzvtedJm8grRX+nPd7O3mh
2/HqeDAGcEUFfVmkMVnLmqW3Ts6o9nZtPNhB+zOQVNwkILJYQOp5ABvVZu5wFrUO
7YZxc5cbGKt18vCPtvQ9SW7doe8jsUDg7jmT/zcbHPXw3RAsqbMMNIw/6KnjmNC/
`protect END_PROTECTED
