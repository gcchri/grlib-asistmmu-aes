`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CqOdBruoXkD07hwSXn+2O6z1A/mflpTHQxuubrHwZEMJRQhQVJQ5VKYs09XdsA4L
LkVAny/0SSguFK5W2nkOUNpcaL9ASHwI6qWjKGs/FRtxDBkjDVW2zr96sHhCUeVC
JhemqiP3LVwpwvpReGNeiWP7MAha7pUs2LS2vDYmJZx085S/tYQ0O9ekzTlttOGu
sWkUfPMEicrCTvnXBo1M0UXnqU5POWU19lPABw9/BF7SgEsVNV60pC9ZknR9TCBM
auFQEAZfhE/w46sASHx+zPNlhI1o+M32fZ4vbfl3BITJv699xrk54oca3aUr47bq
ARKYwIy73Crv/bHlobHoe0Wk7NZz5TXZ3EaC1RvOZtEYyNwXDAUbxmvdo/y3fOho
`protect END_PROTECTED
