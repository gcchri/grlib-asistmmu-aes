`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1eo7orrYQCD+s7BdIsLZ5mi6qjiMGnZqzQnR9yNItES9P39c/yB3gbAfN+tLVtHE
f4O1sVG8/uJ9it8i/7BAn6aCcFhmUjuUQlAFH7p7sde25kC8/MGMC3C4q9mYZux9
59NKKdZq/RGPKtX9lyFnTENxVX7ljsLPddSMQVISUCKlq/ubmlOzDsZeyh5gU1Zu
AWU934Ztt+q39RiWATj/4Px1YRJMv2PdL2BsLxmqHnRbGD/Ysh8kFq63BkFQZdH2
`protect END_PROTECTED
