`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZcgPkXLkCzp6oaAuVIn/Uv9HNo9OtG4gwak0ESTXH7w3QXx40F4hkzeItEfEF3Tk
lv+hnWIhi7/zDujg0WDUy86qo0NHrsS6AEX8syfxg+5QxHyxOFNax7dlCjvoL8AI
XAXDohaM3mu0CLl/qD/T3e7Y1DtDQ+LMwxcuoCXiMrhzmSdQZMNVHLz37lJgAB/v
rjmZz+n17eHvTb/3PcZnfPEiqEhEgs1Wrzzb3zDvivOun0IbBlLobocrYH8nCvOV
SOCiMpLbzNT6kHzfXzl9seJa5c7wm9UvVXSgY0p4e8CdaHVpThTU/rL9FZ4CsLgg
4pULmU04pVPijFy/kv9DKA==
`protect END_PROTECTED
