`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XRLPxVUG6Yx1oaNo0Wvzth833XaJSy3yE55m9TkF5B0jzA7Oyxx81bVk7sQO5DpG
ZPkYkUymthbc+opPPnzDh77Uxn6+gu56x4B5s6XbpKbhktv+ex4vmGaN4Ii3u5eh
kNHPqIYenrVsqzLdrXijxVZw4lebr9ksjFcNFAd8rKp9Yy6IFNd88riLEEd59eRU
L8d4B8KB5GhGBZRKZwyRB5irdQPmqTVgMY0NGFthnnxn8RaBGJnqeskBCksiYRtU
+dswLjzcOCNa+iNI9XsHD+fZFH5q/kHY/luxUiprCPwWfbAa8XU/5fJELUCk+Efr
1iQ0aWMDef+IU4xZiWdVWfWaABaiS24Q7Fr4xJfj/xPSGvP0HN0uhu8cOMJF86kV
osErbR/zaG/1Vc39KmLkJhca+YPKs4MKDT8ZXrNVB0syu8CZN1kSSzULPF+tm0v5
mNUXtzBfQ57n/O1rgMVON7lYBHQL7zMgWU+ow/tv9fHbu4VzK2J2Tb866c3j3gBL
SKlt9Si82SM7ciP1slviWjCzGbDi1GaiHkW8Hv91tdVOUVseS50DsCH3fdWByI/z
`protect END_PROTECTED
