`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rzzOFwMB8LUekSrIm8jdHRf33QOaK6jcsbCm5u3tZKj+WgLXdOcAjuSbgEdCQ0A+
9WfbD7+X/qeJplf1PGZ1QSsUvRPI1P2WTyMExVGpuKYJdQTSRSGKKQFp50LhdmaA
vo4PaWf3XYkAERKhUCxtSfBslAcfV3hVN2fHSwIN4EdG8PA9o070g5UJOBPku5kP
WFUAVVNXD5ROs9xliPCA55QgdFOG1oDwZvkjWmo/D8VRK+rZ6KSSLMrHtG+BaeFl
SY696iDTCInFcI41Wj4q2zPCHjV42baVsfeJRZ6ot2Oa/fefMlGsDuR7w+DosdHr
DIrKzCQFO99+KmMu2zmYckz2odaCUJrfI26SZLwzE77O8RdPMojwgGCHepseiVSb
F3Y+1D6p5RCxRwUi4P92fCO4yiF0uppYSx89lZHy/AH6C1o5kp8GDis6ex8+YGDg
lPFv1A8Iy3uOGg9BS0TgUFV7hDY/Z3/sf4UooxM/Uhw=
`protect END_PROTECTED
