`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g6v0Vgdfi0OME0VX5nd1DXG5EIMoJ1EE+VFGkcaCszgNM/ESkA8oPTJ+h82eXuls
ja9nPy8BRfO54HOssK5CqI7PZDxsEA0YBqtCyxBEUtItaunZ9yty+2yL4Vqzukm9
qHOXPWYPIaLCQ+Pe8QEUZ0Nf57Kh7mYMU5irQuJ2mZu6cxwPuSUbs6athA5CERPa
uNjjXyCM2j2EfCqpvY+yO75bP1zoug7rJgxXJeDh0lCT8DY5he8x082hWtrlYzyv
qh8e1noAn5gQrMYJn1oI0tyZdO1KwL9ebhWSaf9NvL+wYyHGFi5KoNhsAogWSs1J
Gpv/mmiTyE5JDzMT0RFTmZXOzDach1u44sR7/pXi3WVEL8J/h2Uz5Sr70sjvA/61
J/oQ3vXcvQmVQ1he+pIapOSgmtcn2ePacV3dFg0UzlL3Pq/R6w8rPmnBpvwbiA3i
5/DN4YQxVUEvyeZpX3oOzLe6+nu/EYoL7RTgv+OBwo3lEiqTTHwZbOnCnEuar6RG
NRUn/EXHMDhEdgVGmBwYOukMh+ru/2tns5RH3BR6m6pGv7EJVTR/KXhnYMy1dCZt
7ivooOlotWGetpnDbz2p28822a6x2UypxU/I3kZIbTnadV5jgN1GlkwRIl6ZdCk1
VT1oUl2ZUcfIPM2GP7d9cKHGyCcuxGE4mskru/BdYLYhN80W7ipvmCcuR+a6B9sc
C9u81CDF16MW+vXGImt6m816HO3g63ZlX4C7ZMmytbHvkSxsKahJ7tBTM1RFsrIc
2eTMxooK1Tj6sQhAcQOrsi7zxvFQ0WJxd9QBon9c8ajQg/Q9zMDlZdYl5GS4fHGp
JHHpQHIydcRQHFMTN8XABmIAE4frx/LCmX//EGHJinN7SQGiz8E9EIf/PNHDqTho
vZlr5x87VpMycJwoFOZTCoe5jUcouq+ykHuqiqYnyAqVcGds6Qlk0S9j7e9osMZs
g2TvQoF9Tiq4dNOJYioNZ0T4KutQDdjPTNo6Ob55F53z4GqRG6k6S4gtZt3NhBp/
OvYmhiHOXnVd7QP3YwQlIMXvo/Wq56Y4LvV6e1LZX7b5dkL1btgUef2iGmxLD3o+
f6txmVhIePZTcd7tEf353+TtRUmMHYAajhuNpSNZJN9ZlQ2JeQTRmP9CBjM+bYJ4
4xoMX/3PeTh3McBKnjYxYSZ4Orq4m1M/WcgEw7koBUD8SiS377hgVKXONHwKS3lo
+U5Z4PK3vJaSbaU3xnNkiIdIY32h2GZpdQsnAw3WEINtQfYiC/LO1BlIBSqfikMF
+1GjOdVOnWwUfCzpzXQ6pS4rBXq3oUEI5SVLLlunskMTcU3AqIO+kxAS1Rm2TXr9
awroQfFOEsha7FnvtvcW+jBhKZaFKAM7s6EqJpoP65FifhaG+kIHlcve3I+PbQle
skOeswAy2TQrfI02rCi8e8TxwkvFwXIIvqPZSy8tQCXnSSIZbAyQsj4HRfxQV20D
DxG5rlgjcvD/qDKlx6uEOJ9pHCTjgVsPelv6/BJgmDcpPo5Iku8aBixHy6gcG469
YdfSKROD/kT7pjuh9PVdqCddeyatK1oS3G/aH1dz1KYBM/FMVURHnpl6N7w+PuUg
5nRs9hF92sVcy0/MvB8dhyh4I2QRR0NOpW9y4nxf+R/dn6tcl9wUqkySOWAj5Q6F
ae7gX+0xzdYtBDfmgzyn38Tl3U/Okxo6h6VXK/trhGzp4wArkyAqsdOwFjalwHEv
o6+oMQetYhJvMHrqUjDQsG2qoBlLvp+fBtY/ppc8FtF/2AfrUQmLheTnxDAizhrP
ZhIiVYkxSPvb5Rio6D6fPMhxwhyadJPSFq1Hdc3d8CZlPiCgSmr7fKPAMuXEi5h9
ijzOoFBHl6Tdctwt6LHWER95lOm2UrO0e97esNf83XEX5HW+QsR1TQy5Z/VHp+Ia
QAOsXCYoIGsAvDPeBcTuFkvZEn0AAu+OPhrVTGcLufZwZ/SR9ZavOVzNAbW4MV+w
4TMerbCHTsWPCD3rRtuPpzxtb0UfvH4CEltmywcPZZXFFySze6MG968q+sTWRXe3
Ibn4w28BEI343YD6jb8W81kl5YBHK/GJ+ZrcAq0JtpPIf1UErEq+036lVjZPIdct
3Qc0HYJQdl1uMOpQItolXtwyq5bHhYaeP/I0aaMvY60OQq3GtYYHMQkDyjZIVAzC
IDpEh9YuLxLUJNl7HXGpJ41OFeIrkbaDo453ku5KThobecumipuXyGtCM8tFvcxJ
8roVtJtamc5zgZ7IxVpFOa+d+9ORDUgIqbEuxcryOGhCX85SKqqSxjnlLvWc0xQW
xDvv8F3AnB4ru73Z/81Q76BzRxbvr76c4awROiqpTJMwf8t4/qLARcTD5y66jU4L
ckR3EPoT9qZ7lcUjLWsOLFtihIjeXmrKPjWqULEad4WGFBPa7dO1hlRMk2z2NsD/
ycPe12l374bSpa69Izj/D9vZGRTarODeb7kE9hO509kTl1ya0Sl3J20k+nYjbKdy
rdjncu8BOPbFPYTpaTcy4Im9PHQplAFhvEwVr2h5U9x+OCcAe3sCTCH0NgTpgiFr
0BaAMwPw+9CeonVz9GctLXp0+Bxo7BoZApu5Ay7qgZSb1KlToD32md0FzbHGo/MX
qSnTZDZPOKIFC3x+TLfvG31vKFsw0aoIieT0T3B++86LGhdT8/3xxovuuz7Gq1Vj
renFJwBjBIjuh2AN7ehOAzKsQBHHzrwMpwazxYXwdQ9mDIc9zrZ81c8bm1/A1syK
92fjBrUyKXJh7GQnHB+lxJp9ywSGT2ph3GtGhHxGmtjkc1BAsJ04Hc423IRycdlX
`protect END_PROTECTED
