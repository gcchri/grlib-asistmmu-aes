`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ZNeNfxk6mpLl5cEKlfSf/mex0SWkAgIn490cZN3UKK31WvjA+6meDvEtnHABa/U
YmX+fJoYPW9DL1va7kU8g7ixmrWt2pKVo5OAhI+Lsl/0S6kMnPrPtH5gPr0kkhqF
mmxikcZlW/NOkR1UszLz9WfS0NMk2ZYoXuGqmZGZrmfLzp1xOL8qBKUNKxm7BOJA
QEgordKAVkeyp+DBf4YxjrqyAWwvR5wkryWPpQaiQwmdtWo+iK0YbCcojBR4VoSD
WpWXWR/yGcF+sUXrlFVEWAFr7YA4WY7hV0oH3wCtvF7n0pY4fQGmUa6oxqs1z90h
ImN+areg2IC2chOMhie9Jp2ep5e/eYDEjbK95xHyMJU/UyKFYLaauTvwJ/MaD8do
1QDRE25xJWOtomRjtRW5+sa5B5EWEmcl/7Vm5TrwXLNFJYDO7ShM9EMTItCNT0Mw
A0U7XQ7jC6H3IWPFpioVTAZyT4L9aRYZi68ralcoVrRbKHIfmh3OF5owmWvAmxd9
ncWP7d5c/PgYUukwFXUIlrwBoOBJ5RFhjn0fxxZwYodF2ukhMYr/YZ2aOZBaaMgf
oJiFg1tc3zFmTYExzyZ7aobMVWlYKSL6KfDo0E6OX0VHXmbAWuYTieM0oldE3WAT
I23toxLhNYpeyg2ExYwqjw==
`protect END_PROTECTED
