`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7wQVqsUREQaZjpMLX43e0YHSfIbhHQo7BeZlu3+DjdCGD415BwQXan+ggSQrbNQi
PZzGCMW/veYjRWbS7Xjmj+kBxBavJyHHyM5kpAs3SO6bJVpQVmtjF79J/F0QG8An
VlkV7E78FdOjTI3kZq5mmqSwy4Suskqao/nvXprmsjmipxb5PMXEIk8cBqj+is1C
LOSe6TN2GXLhcL8a+9j9ZjeRyI5du0u9PXp8jEw2FDM8LSDzRhKDbh+BD/5kLx/5
ihTsFX+85Mv9qL4zM9ZwLjVqLyz7MXLyng3DoRR27w4=
`protect END_PROTECTED
