`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sx2x4vYM86IZqpr/GpKWcZgPMmTEiBRtxotUlQL5OtdeejNAfsuXhuH0d0RjRlxF
4sf1d2sXnhnrGlcUnvnb+lD6qYJ+I+I8za4iBFhSdG/9Q/b8v/smkN4aUjZwtgiC
ryqlNyn8bLZ4voY8ZeCFHhtzXeNTIQzKZRIrTq7hczVfZLCeNnWm6c6NHkiOuHCo
eCs8Ewm5/47jgGDSv3UF7PTXW7k2jARB/yyd9xZKzbFGKrv/Pe/kdSStQEfKCRoH
K98bFFLU3KdPajlZf3NeaH6+yajo7CCOg0kcUK/g7xtTEGSXHiveC1viWEGNd+E+
w5hhPiX5l4Q41gNVm9xoMQ==
`protect END_PROTECTED
