`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O6FOTC5ENM8wo1eKQGfn6gPt8yW033U5seUA4+RTWBsf8xdLgrzPJr0Vw0GkmdnF
0D9t4eKk9jSjj4ty1CNINjsUBHnPmWbZ2KkDhyddBguRgvwztjOGaRj1R3mpHPI8
xiuvgxE52oYlbzQPzRiktTTKjj4uUV1+GjLf2XQd08ywFUmMSF1aFuQI8Wmr3Yki
lEBDcAOM6bViddUvudX9Ob1KAKIFX2NE8haeBU7IBrulj3wjPBoWj4/oMkEDkiLX
x+nDAp75+Z4W7b7gfmo9mhcm2prS9qCCyrisEO9jIQk4PxLEWEx9GrZyqeV8YTks
5qqhOXsS80+FgnY+7LOCTSCTCUr+z4DV+V+FrKJHpmP25oS+OCHHKGZg3oMyjNdg
3S8fD+fJDsipy+Df2k+qRAHdG+Z4cZthhqm073tYOlU=
`protect END_PROTECTED
