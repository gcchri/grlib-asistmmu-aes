`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kxyfEmX8yebMeQui+WTNDYYUv7F3DeplRHecyqya61M1oExRivaTmM9MByDlqqRs
n+HmG2WEi0WayiP4wkVuIdVwjJMC7OH58GBBBT9YZFb9syaakbpWKTGmQPZq8DC7
bZAUOyelKkcNE44OO9i1HQS7dRXdZMwk9Hkfg1Wqg3LUMYnoK2+t1IR6UCXlMWWh
OLz7s76U5jEDPxXigLu8Cb/YxFVWbaCGzDesTku9g2j5tvW+89GD8XJNfUYCzCxf
0re32nbEMWV4UeUGRHVpK9dXUvgiw/edUvuGy1ALWkP7rhm1x2DYho1jibbq3I/8
9U0d9ZAbATGOPl57u+Z7Bw==
`protect END_PROTECTED
