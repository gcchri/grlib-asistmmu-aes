`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1M+HJg99z8aEyl5iXxn+4HQQJd+d+nkRaAToeG728micpvDnSLDgI/3xDh6svtf1
BAOeXDXkQxN325GTrF3YgZz3x0ah0KkIYsv2gM3+PiDYm/NFGbn0coLL2VF30p/z
RioZbBAodIjoKsdH6Is8GmhcTyeoa77y02X5LoPpC/fDO03I7TIo7Kv/IuKZRhw/
L7slpj3LSOPXA5dSZNsyAq7Il6/Jv5vADa3IfGfiyhKzQtj0zM07sf6OKJzq9HWG
E7elYyM3HkYxW5nR4z0LN5neCf7R1IvvzbMT30awvx56hfx6Ci4rKEpFBbda6weW
Fh/MwYLXA0hr0dBNroWfxB9wUvYb5MSBhtrDosVABLCJ0GFT5ZBHrDbqkMtNzfp9
2lCePlEcLEHjpPI8A8X21/fuHPEDBN9dnqnHAfiRlspLYBvtfnIjqOV9qorlCV+C
YRJ41iYGksqhe6F5OxYtw04rIzeEwK7ZrNM0sqJ6R5XYSLPz/v2j1npEhhm9WK/5
sfIaiUNIIH1j3ILla2Th9C6w6QbTjafCL5ZxMYm29HyZZ2Z/aJkSusGxZdRtiKOi
w7zlIAR7gUJS1JpHf0sBpNiHEs+IeI56ga2J/hnTmoMo2/34U4u4ITxAuBPVaKbF
RTG5dvRlOoctqvFrH07lAhVEY8GMzkEXT2vkVCFiPQOdxV3abqH6q/vB2CgWh4Fp
0LAb1PTfovNH+RcVnL20q80Hl31tVVaTyKlKKAkYK+Wul3k3qoxJ+8ynqIP4DxGY
/hndeqFCF4/eLAteJFuiGxC7vAeakL/IAgetgrN13HPrNaB1AIJvAYbm4D3Gd6tl
peYZ7vpQoSM1TvOvUSRwEVTmsKpVkI0k/hmfxUjAVEo=
`protect END_PROTECTED
