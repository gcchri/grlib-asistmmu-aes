`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WtOHe/msue9/y2HjbdZKcZSBqRcnI3ctzFajceoBUEPilZdQ/PyrGCgcuI1/49AU
9EW729Up4qWdJr7FzpqBhW1edabKUogv2diC133UD9QvMDLmgTJkY1O4QFYrWhhe
z09GSD5bgRA5C2OYjeqTSyBBPgRvr8cFXYCMnxez7atMQE689GxITmOf1o+dodmn
Q5giAR0istxPxaE7X7fAZ7SOEBCYGoNaC2RZ/LZgoeTkYI0PU+ld8KKKYdBIJzKu
Gob97AjZMTs2T/r3Ihth8muOz6SKiku5iMw/i+jpk15P3pQvMaZEi1vCZrTYoXMu
hp6Q3R3bKC63UZ1kNgTuzA==
`protect END_PROTECTED
