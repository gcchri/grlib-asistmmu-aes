`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TutIwzkbUGNsMWoCtr/eNrnsF42xxbN4/ysBDqOyu4SJcWSSmXUEDk2INWdZQRBx
lKq/y4hacno3w6mOJ4kb7s9XwQeaYloxxVSbWEXAhnSklmIkaVLQGVboMOhuEv6R
vop1wjZYayoHrfKHOkY5ydmNxXgvUaZVa3GJ/ap4RfFn/cJAPlLm46aq2zGQm8Fs
Gr4YGORgO+qv4/lz/YuiYSv+FDIcZJqJdN+KuXDfQ11j1ejks/byJ1Sh4DguHLod
1vec0YywYxIWR/Pmil7v+aN18Qxcitd/pp92yHKgJrwecWG14LpDNE0gGx2GLymF
FU5yhvisqjVBC5Ltzz8RmH+8vhHom8TTT62802KRxFK0j1nTqIj2I1xPqBkFr9WW
jNrV+sDcW2a/7KZgtqLT7gokZdXepPbIBWg1i/s5uFRFHx2xxH9eSfEmctIstouV
FL/BcSayevaZiSJbDJdhQ/TB9eW11EumF3ZTOadY417iTXhzqscPAErA92zoY4ZK
NjIn+w7Fd42necOiYIqzJCfqCvAbAb6y9DiFGyfnpzm0NC+krrYfZ3NZa9dB/xYi
jcw3UCY0k2yFWQoJgTW4giHaQnqGAaDi7NV3PNdjMzGUn+5RKMcRKoZD2SHPNTJP
euIQCu/I1WqL60V7RC8PbdRTfCkyJXbz47qUNLhh6XatrqAFg0MwPjRAj9Lwkr/p
PSzpHjCPgN/zu86+sZUbA6obSqIjsPDjSMM8CssGHKcMzrM6DWE9yrEe4iYpcsUL
wE4scNmgomlogZSV1NahfyRxHom8IhRKaNDm1Y9F3/gSdscaDL5Qjj7t8LahgFVu
MHOvmoHaY8m9h89HVYWbKAARqIAO6Qn0rSHjypHPuiyF+XlqeXyS/0jy4FdoU8az
bYH9x3d7bcpf5S3r/UNI9IWRW36G5YGYXW2wxwOnn20o/uOTwWqzKr9icwakfvFP
tP61eaA5IZDIIY3kjYONsad5us4yrKyNaJm+gzu0v4bc3U2UN8afRlxEDYQRk1Uh
ZFTblCaQenOhFeUFBgnfYH33AvnOBWJMj+d7QTIwGI7WOtmyYcNZ+2T9LAqJDze3
sm5SRmxjBcemJ/E/f9bEEQ==
`protect END_PROTECTED
