`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CkhfsuBzkhUVYjpPfU+lrNz9JfbbGOZaBwBNdnkEcuGgYPZX+dLtTxmhgyWOqQgU
dRiK5NkgW7GLYLVlnZnHkir2QzFwIGHhRCZ5OwxgkcifKuY+L+u7PvN5RZix850n
XewqnKI9UnwGt3ccJTOQLRTbwhpnT4wwIhejcdKcSAKXe3j+On2+GwFZKthd5BLP
VfG256FaA/OmT4KqE6VGuIo3i2O+4IHKhejRZjuxdLdifwfpNPYPc1jalcybrAE3
rbLLLfXvs8HT18ilCJq428tZUItfjTyBo5ryPfvlbgoyS0ySRILba0gqWD6Z4CPf
U9VkCsfdquwShUAREigN/B7qPOeSI0infLZ0NChcTTVmswxid+V56r3INLkORiZi
2M9AvqR8JJ0AYEEQxUYkx0lr9KTfiGxHCXHfeA702ez5O2k951ab5XQw2OXrJdlJ
EcmdrWFzbjqellPjZQIa7ot9BDpjCg5F3W3Y/E9z6NETZ/ZXxkifwnfqxlMt1cGJ
cX5ueazGm0Q06fM40e165x14sw3Sm5qK7YHh3Wtkse/g24NJvhZo/JtwPWQB/zUZ
iV+YGL0+ZYzOduTs4lCgTDb6AS+xEEZt18F9czkai+EW6xv0gHsEaRCAsDb06KM+
NjRtJ7N3Kb4gPd8vYOjV+MqjqOp98MFJET3nCf6EWgtCSRuLNdyi+qIwaljDZbTM
/dUdTFMP9TT9EOlsrHPmiXT0tp9M5wFLrqt6VQKniyaFlY3rq0V4Uet9lv06mEF7
R0RTlLk9974SUtV+N0sreE2Wf0xQyuUYSh6/q7fb+M9VWvXIz18a5XM30GXsTUDk
kziuMAPCwNkxYRhtZEJ6/WC1h26i/4JX7W7SnBu7qy7to/+GYt/Ev978jy8svueU
U2NRQ2t44JLJC6419QfSg3yZRK9sfUKIXva0KR5LCM7f/2Oz7WaWMBT2jkDDsZkc
vmpktyPqRtj8MsfxvyP/nXXQ6LYjWwkh/h8ZHy8ELzYRxMNXRLMEhoqT8/XEjoQA
VoEtQFgP0c9BAOdOr+M4d/Qf1s2q7cr+L72Vt8TnNyu758F4o2WmBZugIORnQiSv
axKIRBNYr022vX5mRLD1nX49sJYxYTQYKChZXUgN0qCupF7KhJblW4khl0T8o6Pc
1MLAbd7rSBfKNjNdpkgiiQP6vTph/5S3PrY3ob2kgzZN52lh2YHGAgcuPULNAkVu
RgP7cRGUSOWtdxOxy9xOQQK0y3OKIyM02Eldhbh1V7fkV9mUrnj+d81MtTOmkFk5
94icf71LDsSHwNWB0e9qqZkp2DVaFQWKqyv9R3MzDl85/wT3ko1CoBR8GzVYm8bL
ay8bf+TxZAsAw7oOyE24MQBLDin/3XYkJ+JLmdTjcRFHl8B0JK4gsh8DPsDo+7QU
EqP6q4rzIKx4EbiMEm4qA3ehYFR77wPAsdFGagon/CL9CBbskdBJsJqM+2NsykJ1
dA8a9+T/xSm5KNw0gYFk2g4cGyeFAEgzTF++DhpPtT0uR1R+mViHMbAh2HnWxle0
Cqd4l5He2RzDAvkkO5kOqOOqNfguV2KzHijRZRIBcUBYpoAt5ZwCRQAq99Z1Gm9R
rEPH3vUtPupEtJm/H8/cpt4sSkw3zb4LryW6uh2/8qI4j7snd33Rz7xos7N1hkZU
M4CSwf/RF9puvkyj5VnEgwxou0RDFov4H/3MpLUv79eaPzn2gt8Hj87R0EDFPp3B
yy2hU618yFZUyxk7m37jklaN3Wiibt9RWqKmc9Keag+05ZPqJfVLpo1Hcu6WHlfj
J0amCqbUXAW17gZMFRjv5smSqdbVXD1XVMSKtZwDccWdm6EJxQFagHEjwfpRDssS
rgACVa0X4d+zUZlvfv3BXW3nmxhYF24aZ++fDzrQwS3b0HWA2+TXAzpDJQA2yroC
MWntbJDcwsq1NWqvLpZGfdBL7l8uXw5xAKj9qGmWEgMnPwevCRF90Hbk7OXPVcMX
fVXaTzYzC1yHG/GD6xEu2wpdDh1YYcDkskyrjOllEnYKsIYBg8U3hVWsgGpxpNGN
Wl5Xp8b4v/t5KxYjdUDlhbKgXFz/+kYe2MW7OolQs7fGuyP78AhlOCFFmK/w2bgt
pFfr7MOfUoGum6NtVAbLZulcDtqLb4ZOo0IELp3sMEnLL6oIe4KIzF7qOSbBpKe1
5rUpHr8TVQsMh92Dnz38caU3iIA0BvJuQHyQNup4RgInMcaz8ZpzbFFt8zZsJ9C9
H0FfZnL1pw37v81sj4/IerqUWoArExp80XdZ+RY3QzxI8zS/GryoPiBm1Tph6Kdu
NP9r9tjQ5TLcuCMX0JFI9vJL/f7DJYyNM7+87WEH2n+mbyNbsZ9z+bV9M0TTfLPi
rohT7mxdUTSoitTPtM7H5rFqTM9Q1s7/SFlk4xFsN0n2u10iqBJhgGsqTdJM5DzL
OIpgxzn3H/weLshiTMqE7S7ewF1hNkkdDO4F78TQQecNKgDP+Z6Lbp8yFYoLDd67
dB4rA6S+Q37RyXsgXIg8J0LdpazuxsYwO6yoBrZFKS0ufRhfp9Sf3cmhZDWOZpUr
sccy55/hdToF0L03ATgGsKE1/hNrun1k4p35U9DsFL8iAjBkGmKKBFW9W6Mk6X4W
5fgq4rArcKOIeoljw3ba+qNi79bVTBOqDRy4agbthZ99C/A4cpsn1H+QxOCNAav4
jdUj2NtOyNDZL8gI1/VFTAvabnG86KEjBGDVSk4LucKJLoQmBzbdeAFR44QUEy1q
gOuPSJfjslI3YPDo2UvcaPxBjHYgIHRgpJS+LbXPkz/YqaybMBACkRNaq5dHvbIO
`protect END_PROTECTED
