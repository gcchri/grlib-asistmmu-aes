`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ZyGrMEjlUFj4Dmz4SbZwYWsWaYIpBeFhna/0FtvQYwSO7lh6/g321DP68npD4B6
s81mQ/55fYwjjYEePt++jweLJYNQB/5vLDoKCwHP3g+qLnrN7C50egTSjCk4rBml
KOsgoCywUQvMP+b+l2kmS0Psfs3++v6H2+D9ATeTkPDCAyympMZ7+yPOmkVG591/
lGYmZmzi+T/68VrKZlRqgQSqGi9K4fbs6Oc+4CWll6IahSnoyuE2a0bew9qAfDhN
09tPcrEJ5odZ+ibHEEZcp9r+ZufXDIIAPcji3ZXySTWep6dtuUAkhEDfU24BW2WQ
CxrFZny7nRXFkktZp0WccCk1kataiDcAsbIXtRIjcqYTVgpJ+9etOwOvV7AvVUYs
a1TQ6pRhsgNd5qNV2h7ZlQ==
`protect END_PROTECTED
