`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m+fyw6pYRon9HRPBC7aqBi+NZamZpBU2aNzMHkxUnqEyQcvNlqMf/C92U739oZkZ
MvFlMkKpc4W3nC613RNLLCHNyAPjMyA6XFGIccZS+5Zfi+w/lw5f8bIUWCIzXpXj
YtDUwi7imV7dtULRO+TYagKJSHyubhblrYLEj8slKf03nTpIMx3fdVIaU9bF5vqH
6T4TD0ebiOUInsFA4C3NFXzvIYbsWCmAevCppLn/9on9LmAzJhIDsDPyYHrYc+o4
5l34YiNs+iw3qxrJIm0A95Bfmu70OyQBB36s4Bb0QOhg6sdERw8wuQNn14AgSiTb
ZEd8lwWvqB2xcVcVfX8KGS8zVTNYfby9KhwjEbKWFb8EqB9v9dLm8Uj49rwFmxFy
JhGblDZ6ZrSOiqcmf46HDRaPID3k3E6F/PyoPYJTQSw=
`protect END_PROTECTED
