`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1fHRFUbcEDaA/+NZSEpeN/0d14y19dDAKJ4zrn573KroDfypBsWCBoDH1lh7BLB+
bU6S8OKcAXd7HPITQ8njf9bjz7ICbRQZVnM6PGHOYiMTzV8bqnREPNSBVCYEiLUF
9vPQQnkLlxX4YX3ZgAsovylGTWUS2bIYVxeEYcigAhCJI2Z5d48asiHKvpAngVs8
OuVbVyi5frxVwBvDjzfRCyTdVei2LhjyvWx6DY+PEgdyJu6gc6EdkpRVmJy6e7UD
xkpoK86ghxhYGM1czmZ2LlfzuQCiTs7b5oZStpPjc/bgvGkYaJHLPubbl2/k5Z2n
AZjxTNCcCwijwpdkjqKN6XXRd33ObIa39AIIMGJhHjvQ/fhS9NYtIRjtUEPHVd8T
IGvQvMrLfCuMRQl1exz31LY6lsY5dXZWkajfQsWN3cg1VH3Aea1o/XP/NUWSqWkU
JPCdXHGJgryWDHcqlThGVhGIoO90wA6QWcx3sMcaDkAjhvHVt6my2AfXqfera2+u
WDjPPOJZ9awKz4b8GUpUZI1FOT6lUDg5DzgYkIRpe1rxyL/bk5VTLtGdu3i8kpUP
7KzgS4b2IfrRkmZAScqnODjbpmTZHVo0mBmmg05sGHOKK9+dSwWYXgXdIGudm+tx
BLg8OzRhBjdCjAaNj93vPsTA+dzA455o53ec+us5hjAYKhaxf9B02HIcWPlTiWWP
sRZOoONR0+yU+8Jq0VUKjw==
`protect END_PROTECTED
