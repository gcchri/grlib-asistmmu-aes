`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WRLe8sHq7NtXivT0g3ODdvAvscBSInTG4kmmO3GgkgBzQdSXgpJONKJU2KNh6RU8
+rFuE7eSYDfeS0M4OYWab2gn2GViVfZVvB5WCmiSnq2fJKz49RlNwJEwoNDcvrLf
s0HMVI9wzAG2g/254rmR5Hnc/wGNxt4Hlei/Z77/HP2kxg/hxYZqlpsiWwNHWXN4
xLsJuoHmpKkW73fq0mbGFnHu0YkoPa2/SNI4HdgBoxtRkik7VT5oTWf6JCHhrLh5
k+vfZCk6UU00II9KXGMBIhcGEM0MJgHAPAmkyKMY0eN7p8hrr1FGtU77I/AKYNaC
JhMIvWzvcoHm07zLPmk4JxTJ/VhBf0mLj4esh+zwWcvOI9ifXwRrAFZzevXelt/l
IVO2P6TiUml7uUDNT0TqzRrGAkd+mbbSjDqOUQ9R9ij3ymZAq9vsWNJCwLO9C+C6
`protect END_PROTECTED
