`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FvZMT0JOrreFPgFdszceUzAzyG1QyCS3KzEi11V48lKz7IwuinLAIgK/vsjzPm/9
SdS/yr0T4v32tIosHJWuaunLxiZwKB0sV8y/5n4QP7Hl2KKKQ8E7nRErArvB8oLd
r+5PWe/EcNfIxlcCPDU5Y/Ia5PRLZNDoLxUwIrm1oZwk66aBcfEQK+RAZzU6atB9
RMpapTaHH6z5YhYdkxobyY3z5VGyIr2voj5psi9pBoGM5ikWPHXVF6d5rsMu0WNh
p3QiaPpDtWyhcEfvRHa2AZzYsNONBrKv+BlMx6C/Bmo04EGWLO4y7xSbJUQBRTHv
kvjqYHhZqxG8L3qNCpbbhVBK017AJgwYOJyVuC/js9xdBsmiy+PslYtX+/mIKfbd
utZIP1Djh7QJeFWHMkPSvg==
`protect END_PROTECTED
