`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
luQ5LW+QHc6ZKyXWxQm2CirC9T95D/hHJZypznVRdCEa950VwfRjt9OjLRmuY7B/
7DPqtoYOdYZ7vyx6h6oRIuAolZ3ZMCa6BPg2GytkXjPqGjxSoVpREkA0/GUSfrjD
8cr1aglZw0bvBBBHej71JopWUqLKR3RQ4jFydeeBjVHGXZsuSG/fDn9hujBpfVUe
m0km0M/Hv/SOokzJBP+3s1hA+XloTUjMPhT3fAlEDkv8e4w3MrMWKfydoW3W0Inu
7DvsF09YafVtnTexCMPncNP2mTUojAPRrxnqSg4BvuLAD+ikuXawPr0RDhfp9MMJ
veyPdm75zsYj25Hnz8Lfzg7OIP8QzHjN/4bVqGZTSrfce8R9MEZ1c+LegHlSM4B0
vSSLGiQ7gTkMLu6eYlDcLF/LSexz2Lc9NKuEqr8NNmemcVRAMfH0ph0Bvjxj8zJv
W/nypqv6YtKYE0a+AetNu5o6xRT5rCVUDaKcZYPIM6hpwYx5pguSCouC8KV3Cu39
Y4Gz0RiYxXiwg3ozovTLPkSoKKS9XCvTXzG2HTc0ovqB1JG7nl5Qkv0+8LBY7KN/
GazDw4iGw+uyg50laTWkH9BJYPnAe25sUS/wZvCCNTofEFqUXfo+ZaGNt4+Cl/Nv
7NqPrq2r9G/tWJfz7aHRvp6n0DmmRCRZOpMzdiVmhiOlSUjF+Z7/8Yb26mVAO46S
OOcYSaylGi0DOwHISMkaKjA5D2zCJZYw/UNcNUGe+2SAJd8KMBK6hVQO5sYOqPMU
s7c65OZ8DQ/UxzovjT7xtoqfjQvcXnw+O5uUwSYDcW8lV8s9tmi+CHlKkU2TKG8T
gCKwP4ZC5rc+YijVDUnu6lAnToNe8zrQnIEohprXAlDM4AClomfHd6UzrIOvq6RX
1ppYDLoxr7oWF6Nz4eLimQ==
`protect END_PROTECTED
