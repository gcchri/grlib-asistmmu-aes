`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NjtRmlpKiHTSp1CfGPgrAmhnoWwDXGn4vLodytkBsn+irVOw4UVPZ6tiXRsB78S1
a44ZdRTVi6ee5RrWzAz2wAbxCdQK5YnhHn2C2ITGqikj2i2NmzQ8TwMWvHx/Qn/F
aH0fwJHOGTcVQiAUAF89ScJKEanZpxoCmMvLHxVUjtY9/unyPW3qsRMMJJsVWofW
nJlHCapWBCk8qIWkGffqBcfD7ttFmjjNYxfw43Rk6RMxFnG4vwvi6pyrFmNu16xN
I9N/Vy4CzZzl/+fQbAZnL7/zL/MzRPzRJia6+DMS65tGyp41fwT1Mng2n4BvuxS+
hFU0g3NzjIjOCHWCNbUYacLO9MWB1n6qD52v+KCIhC7UwyGWEuqYVXHH3u0iuC2Y
SYx+jgmmq6SK8ZyRGk6Os2cfSc/gyUw/QEmJMayB93iuWJaeABkwMgoN31unF7e0
BwjYj9QSiiOLyzj6BXFBcvK4ofrDuBCXbNZ+G9ARC0P+ZcbLaj4MHBC46eYDy11C
vwTgH12Wwki0G3X8jqp7yNoMCP05cmMqZrzF6bMbRQcmOObwr3r46ILvomJK8o3E
U/gWwmOeaFDzc/09cCGv23rpFuxT0OiboSEz0TcUMkg/T+GuO6l97ja7kFlcuqK4
qOQxHUKOgL//yV++tNKz+g==
`protect END_PROTECTED
