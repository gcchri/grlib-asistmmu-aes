`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+5OVCGfu3bj+WozPzTtQC6CVrOm2Vfo3TqCFshGRyUhZXyZ1MKddjwhKF6BLNuzy
awx6UjrCVyDPYKFzB62FOm80i08GZd9xR78zlEZhQwnzs9LKnH41HiaVvxlhxT3i
Aa1BjBWtGbyXJlDN7WAlUACijBeLuWCMBjv8geBUOcts40+8d09Y/rlbiOhAa80k
qgJbpepHOYarIBsftYlR41KCKeJYlomhhtOmptdJHHcV5bGf3/1SipTBWfyyQN2G
o/WKGrbWHqa/KM4QPfpIMGV5S0ykwR9W/oKMib2lsJNHG+t3RLSeKBaKIe6P/3uP
1POHYKu1bBAKTXsVtzuODacwA/5xe7ZGXuNGPQ7TGbUNS8ZBuhJ4ePlHrfglahCS
r7v4xrJBRaP29Z9k+CeUX6wb5nqja/WWPtY+izAyW4rvQUrguPtkSYUOHh3MA95x
5jdlNOUte/qZnv5jfV/i93XmBWVPHhUgLGFW/x79TNxp36Kn0vz8AROLE6Hbhmgl
`protect END_PROTECTED
