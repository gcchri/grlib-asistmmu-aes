`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v6TdYDXXa3JAO+BKUU3XBhTgtdoI6nXR6q/VfOankaFOLHLUEQNAWT8Gfi8Q89ao
kWjLsQ22UGhro7HAHfjEeVm71DktPEi2EQirtDgRQmORQA2l2cMondRMgyRTr+2f
QdO4gNW0A/Olf3mzqGcE4UvhD5dtLsRBJoFdWzuMJI7KDA4IcpTA443FxCG93Cd9
5nKWr793pYogkEHQjj6tOtI7/C3plUvR0WrT0SUcXZJhc5urAbj2Ty/nGbT9eGVW
Y2aEEJNo8VTIpNAYEC4h1JLtQDypPFunq/He4SRfMWcmbb8LkjeftqiBLSjUyEud
zEJkX0YSyWVZ3d+7UTjv+MlUEoaTVANNITC2zcY4slhdOdCmd3aFNPORhlniMdcL
3KphxILTyCS4oiyQPO3btHcOq5XthLLY7jAxvPwxEu2kJzheeP6qdazBpx/Jtr/7
PiVRldiD9lKapgK1QQP7wT0Qcvh2o3JwsAtRFhXUNXVnMmqscsAysQ6tdEJzHkJI
gdRFmesEeh4So539rnPAPuSi57WaAqIbC5Ykpo8QYNA=
`protect END_PROTECTED
