`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YXKo4KSM9DEOA39AgVdYC3rATrBNuTbXFE423LlJqpCJRZG3UH268XmklPLpoD63
ZxTTpntYJIQX59aeLCbtX291tsNoQiIXmYpJJRkyTQL7b98LjTmeWYCcTVwqWoz7
xBYoCg7V3wvJuIl/lZJ0mQF5u2e2nR/jsBUv8uOqnumJBvJT/dPGI7E662rpjbyb
1l4k/KDBZ3Z7JHt7yU3evFZolVONQBGBKmPQDBYJ/+9TDMmZRyktc91YMICemD0E
yIViMUvbQSng3j1IEgKCS8X5Wd8+ev+zJC9rP6pohy0lCuPiyfg0RZtlyUms7ri+
xoWhV7B0MB5ZvO1r/TYMYmldtFLhGj8c/0c4f7DFZjLf7D2GGOc7lDvBg9zBtRVu
y8+kDN12kcjrUTGFTzKyEDv/kuXsAx+90+R8C99/vDIh2zX8zNz9KrtogcOki3I3
IY9E1y9Cy3JcAEotQ88icNqYtx/Ug16IvJcDPF6vrvs=
`protect END_PROTECTED
