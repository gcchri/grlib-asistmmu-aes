`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4V5+y/aDq4cb0vW1RsxVvYJGMA/5aDZmgd/qW+9/J+gDd2g2UhErejY0Eak7bpjy
/BrpgWQD3dggQspt4uwu+la167bwUxsDy2jWbUd3NgD7TiR/Uwn12bFrIRZPlI0p
hxbgmrZ8FFJlwH7u7F4VcSkubhxqsThJqnPgCaBn+chXNe2Px0PABkZI+T3g2yne
Je9QqozHoUbsXVfHRnkJ9zyer1c0vUU6et62ZmjJuiETsZkqmSa7rl+69EpDpGGi
PFDrpmGKXNHtHVW64Y2d2jhpXAFJgt32oI9oX0xNXADXebCu3qeTP5YIRYLWv6Eg
o/NJBA7z4sS6P/lgIAOHv3PqmcXAIdDak9vbG6qDW643Yt/tIbcdnENDXbW7JYvG
D4MzHUILJskNvk0RdmA+kIxaCg81n3ag5najjwEZn8jfWjcWH18HUhkQzRqK10vk
uXyP/2+dmj5H+5tuPWNlsk6J4TcrvBmHUpSYIAVnhyZy2En/zYq3h5ivq/cjWnS3
8PI+XbLfN8Wma0QeZ54lFyINVXpezkLvLl0KniWzcNBIniDqvLeDeyQnMDWu3Hm6
UegsD+ldbnu3q5Cp7bpmS7dD8wd0dAqSaqfnQUzwx9sSLbmTtvnhsPJCG7IMEfJP
JTtCiue+IepAsg7sqH1KSTsFCT59Cvhyv3MktRj5sNGVhbqGgc69qi/O7EB/4HYb
zTGRdal0rqwjxPa7LMrjLFbiu40RgAELewdQDoIWVdY=
`protect END_PROTECTED
