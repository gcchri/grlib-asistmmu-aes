`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xpjozi2yblX9juSo+htdLVgSAW39sQMq3E+61cohWVKqJpsPx4bdqQaBhADD1xKb
EO87FRzkIebt6ENxn/7nBXHOAQTfSiHs2u3E12t6thiIRt4fyDMGTHGzX11w5sy2
Fl/dSuqPNRlRrxw9U5RHkAhudgWWvXMtMwrbJgkjXhadEotwiiiytVJI1ZjR/Cuf
CUwOVh2dX1yud5lRdsQNamGpvLvaElvj9zcD1q6M1aZOfsFRPIohNmB6dHuS32sp
GCo8cW6FEi75q6LrQUxLFG5KI2gnbma9U/bFc612IlEOCH/OhnB9GxCB8lSBNNSI
Y84OIYpyj34isRWtBMpH6qicrL3DbvpHE9Kqje8JjCUrojDmzkV+OT8GkfJvu5Ua
vGmQqrGurSOCflre2YMOIPKG1SZWDbGtIipcnxjmCPAmywqk8E4ydXXNGSgzdI1n
fBh3d6jf1ml/b+g+HrunByulxI2F0CgNJTfv0KPUWSppEGZLOHGa3Yflv+rzlotP
KifHvGcfzFRZ/p9ZcHe6yp+hlm99H8Ahx3uSAkwgNQY=
`protect END_PROTECTED
