`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xg/6oA5yknuf4conHMyOx/74I1OwUvtEG5Jq/013KAazup0tZCg+okpsQUXVfpjR
QL4CLuMAQhVER1Q6viX1zxA+XSf7tP4Y11KBEo0hC6WlKUoHKgJHnEWny2Q0YxC3
DVXMY4lcCbgLeFxF+g5WJu/01ElEwJIPnulJ0WD0hv3/qjSP2Pp/lSGI0PhIZzHU
6k6irxlSQAakZp/lmd0j6XYB1DGnkRWo68fvenDJkByXuN952J+yfaLvhvytw6ZE
kvSd0dMxp2bHIg/Tz+ldi/mymJ0mJvKTNbQnDf1AWLAZ64KXYRNTo8xTHOXxuTu+
5Bjsy5EZWnmxNn8IxnjaPqg5Z2XAkrsZJ4IqRttO/gKH+hr1BhntIYbJMxiBGVsa
NzieRajt6/sIqR1P8y/DU0w+ZwJPrh1NL0MCcsbce0AP5TFyPycocZiIJnkqsWE8
XpNNtOkdoJQvkrhBPYf+Mq7M1jNRMaYviE8sjtyb3jxhwFraBrOZGHJH1duXwh/0
IyHRK2jxpdhSQ/4dOtfTdluNLUT+n1jOvIy9lDz+0SQTvVYKsR5qJZJKhpKzZa+Q
ORcjGtgYNnmz7S3OxEM2SlWyMRpGCQKFXIvz2Y/YobZK3dVeQX4HXHc5/zp879To
VL7WIvUmIeIH9kf84B23iVbQlbCYLjHpm0Xnz7H3/dmuHjE3ZdgnHalRs4OZNuKc
Z1UTJB7OIObDdWgoOEfMR6ecsdc9nXKyR2ta6qVDRUquv+pFiVRWhvDG/+79U10m
Io3BpaENwz0WeOEuNA/4HA==
`protect END_PROTECTED
