`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+eHtE14Yyh5kOlPd3rPQG5cTuupJy+Z9Mx++2C2alA8aIDjQR3/Wfqx2p+09vHnP
OKOrDIV/JhhHMy+roJ+/HPBzQ5o19QS3XJdA87KWV+HDn3iwKM8t5Tzf/FNnqPFO
FxkN7+tS73sU/J68dYezzKeF2dj9EfNra5dIabW1menFDfYu6jdEu36JcWDMJaZ5
HH6guONo6tbQC/3yfIUnarcrf3aT5rtsr1RhP8dyvjZVwoJfsXqi6MqcswDJTSbK
Cb7QSZEeeTx72zjP5yzA2chPUuY5TKx0ztdBrDuwOAoS0t/AVwJqFHwTioDVjjTr
0G+itQo9jnaSwbW7wkdDi68kSxA2U+G5u5C+ntbvep0=
`protect END_PROTECTED
