`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HtBpoNALQGqL1rA0ZEOBx1w/eWJvLVbvMuVMVZxfbxRVBZhCsQcD3pFJdONQKuz+
4cTAxn60cg84KHuNsma1lVH2sFy+/+GvpntbwbCkOIDcz6Jk2NHkG+zTAmKyWK3X
KX9iP8r96Q764JQbygE0GdMkJnhbBQxpJ9UGbO8KS/HiHt2YUmJ00F9dVBEBwlCi
UPhVrTtfmPNF/85EUygeRPOBTLdBpKHg6xtut+uV1S03Vqjpchg22JOHEVuhuwzl
cIXJNFgve9qPagiB/UXlLO1xVLKh+WC+oxLvhsF45U8o1ENuAPfDTKGVLsfQKrHZ
jyQX4z7e/MLlcaFaNkTueHrfRDyFZsLcqh+TQsGAq5TqYjhbo1fm689g3uqBsZTF
Md05OKUD365ymOE3EW4J8xncBAV4F0r6UdWP44+SbQE/U8c4eGbCJfcWtz4YOKER
AlMaLUwqKfkgzFT3M2x5sNWVS0ItT2yUybJC1V2+k1zrgsd0yVUP9p4wKCzlAR6e
gqwz9ev9jQI+9E/LPfRx4Ua2J8A4D0F7nY0SqblQ52pPFF/G2Ncs2gERvRFOE+fi
l9sr+tKMp553iXM/3dQvFrJK0LonCKrp799vt4w7LR/dZgPCe/8bYdF76xaflk5a
iTAOWxgChNgQ2vyFq5lx6VfFlMV3FB4EB2BTlDmVFmz7e3oOZ5vzOP2VqIbrvp0O
59j7wSyvNEnXYgPbNxBVeoyNj6tMJKU9NQas95ciOgEf1vcbje02Tb92n3Bq8tyn
gMwlnPVFoYsW4A2dDz2zNQ==
`protect END_PROTECTED
