`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pb5U4RQhXe1N+/IIciMHAPrKZ9ytqVV4SQ9l+d0GRMMprmjr0aiH5+Z89I7/e2r3
n5Fd6gLfQWEazrJuOzdHVPf+xKX7obWnDTZ1vHM3r/YEq3Aj8RRJe6tTbI4ZL+7e
YnHxD74B6ONM6leW/lZuYhgeH8fa7haoYY78hkYfWF1rnhgIbFqdgfV1sByJyNk+
3sX+BmqnFs9Y0602Ewth9HV3iXli/fSLlhY7vES8VEATY8DAkLrWvSThtIQO+ibH
20XUkUS0eEo4nXHqeGzVj7KSdyn8RD5QmNs79Pm0OZfcyvIg7IchpLFIgXyN27LB
JULOQP9yxjCDEbDPHnl6bTCzZz1BPX/gcckppIy+ZoMjIiol0JHRQhzjKDMsDePu
GlCEgHEVfteCfbj2lxlJLYwEp/4ryOS6jXjdUbpYJyDtaCvT77HqC4yXa3jinid3
tG2G3J1JiA8UnkaE6w4lLa0hKXq+GCKkueJDChLYY11Y98QXs8bqOTSTgJ6LrPSz
LyElDA75AMIMwyp49b9op6hTNvA3JaEETGjhoZnC8rwOpaaaEFVc5sgdJAK6S37v
9vptCQsiTrAPzH1swlQSoawNGZQPZ8NsLn8YflVIsLk=
`protect END_PROTECTED
