`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wF55TjqkZJjX4C2Vkvc6r877pcfgS9qTcrEY2eMWPplYxNd0cutgGo3zycTBi5lN
+3Z16aSeoIYmPhMlxxNZzyHN+zZb5HhIjFP90ZLJULgqlTLniSVHmdif5v5+gDWv
6WOxHZKxFvV16Zaj88cGIzr4lB7J5vGdnNcN6TJS440XDCXe94XA9kMSLSIe1ueQ
YETGoaeInfDh/UGNKMOhbcdDRtrXWfXrdyiIGe4w4kIjEyqRl5h0mZeru2tJQ7L8
oW5BjEdU+x1neGftvGOFA9IEIzmkuNiPmcQH39U4GRO/pJH0MNDon661s1d61Bg/
OpDw47Tr78zkDxZqvQdwnRg1LipQv1BFl5/wzCBtk9N/jwvjkVJswP6XgmJAia8c
VSe5QX9GyE6HhnXNG/BZnCsuBPYPY6Jx5Sj1weuh0NVEo/HQO3Pa94j1CXE0+dJZ
R2340oLN4WYRF2o1LzX27N2CkOQy64HLddWxxGA0T3qipHMWVgXMu4Jd/YAra+SS
DwwHwpuAsJZ/kXsAkjWinZCrsoFCyj1vLSjmxeDN7zikRxaSOaqXH4QWkQQfoikH
j4nDizNAV8x4rVCXH/Aoe5FYx7JSg93tP3nwpw+6K2fgM1jN9bkPeTVM9zggQrjy
ygwnfwYFeMk4H0PzHcHunDAI/r8WnXTy7N0UomvWXTDSe1OFu0kXTiN5EZ08CLxo
xofl6VCaxmextB43mCARuPvmDV1EB1eT+BEDa23npRFrypumbj6YL6fFnO5onK0E
3kKKZaGZuS5zCo481MTQwMQqLiUxlIakfULiaULqlr6SHDA1ZRqjaoMmSa+SF4s7
BU/ep5vLowsDyJw7HrtDYYZ6jIixm+p8NDhrd5fcgYe3PHqmxuuWwMJ8NKaivKEw
qQao5Hvq6NHQVeqEY7NfZw==
`protect END_PROTECTED
