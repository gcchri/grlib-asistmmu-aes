`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aHGKJCCMmJvBW0f2ft8FQzPx7S1gmSTMAGjbdhR1dvdeOdMgV13Ul3PSEchJNkgu
rH5zUTuT6+P9cVok4ue4Z/WppqKtA57OOVoncwkh0hWCqTER1gE7TLzS5Ae0JzML
QjzbnTGbxJ2fDboQh4DrPWGAdAOAV7Ya2pDqO3LmlDNmU8KvqqKT8aIa5YWyFBcz
5UM1eIOEiCjjfQJgzUrNFjaCVF2Eg698FNtnhcnlDNqOzOrYrpZU5+0MfFUHvhlx
xAq8RWVQTgpjWMyrGWuQh1okCPOuvZP0WKHmuO5TVtmUpYivAxXUXPGwQDR/wcsx
GXCkj7QmuFcavvAJL3LfOK3nmYsXN0f3rKG8B1XD6YvgxsofI6LUPnsROkNQO3jQ
mvywcUVqoSQV1C0Fqgb2/gaHKBh9Qw/2CtmNkjtJKqUoIJHDtBxgjLyuEdqYYW0L
LNSMrPkzfTppv+98FMAa3CbVot1X6rgxtS78VYL1bEmzpUWL18IJP8ZqsFFFPIjv
TWstuu4WJZPSNlDwzYPKdrbqMpSZFkfyvpjm/JP19KXSDRWXgE4Hy9L5zBAlhSBF
tA/b7/yGaYPbOzeP1mBJtE2jHXjHlsbJz8Y06/bzf1JBOTXnOqnPexeNiSEu/cOT
dEEn/4MXpiw33r2+fxjBnipo1xlzeCJCTSzTEAHaMV5p7opsEUtKVVdCHkIY1LRc
mj6o+J1c4vuyMA9IsBh+c0T6dO07gp7cxyJHpT3uQNwZYo5ixSiueWgok9rUuXvw
4SNQUW7GR0YW6ai2+WVY8Qz3YHXXQwAGFOkPqdxUJgT/UpZJ1Ns/i2JSGpaxYEuz
Q9/IeIKPleBf3+vejqUXu8W568vRT72qAPvEADa+aHU=
`protect END_PROTECTED
