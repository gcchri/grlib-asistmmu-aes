`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L0Woc4LIe/6GHnKvjlg9vhcc8Dr52J4W0AGruOq9rMoxfhzhmUAEfV/+/3ub6yVl
C28ikI2K7skms3BlHp8ayrvqoGKF5QhM93qlrRD8Ta/EUsyXicRPrBpdYjjK6+Bn
u4CJnYYbTc20uLOTGSImkdImIAvZVQFViiCI1vvno3Q08UgFkGEdAQKCrpbWYJem
pmEMo4a0ND5K9j7oCEhDT1QchbVjdag089C2ysqSUJf3CLWLh/lplZiIQHk+3SXQ
zbNERItHK2weMu7LS7S0u/9VNV2RkpbhOyHEPazt9QSOQVW6UCUIH6eJJ54bpfja
5ClIIwI1uKA2s2pZnc6tqBiqpoW22bG/Iq4ZVwMRl9gAUEc/FDCt2ivsaNos6XGp
i5TXggfkJwoU1S4rvOYHdA==
`protect END_PROTECTED
