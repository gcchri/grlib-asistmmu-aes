`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KMJE3pW63F7rYxXviX2OrUBMfvtcVJUXx8bCwpSB92X4sSNlwgHVQIlUwJOkl54L
NvwltfIoIMrGwl1TFQuq5qvTbi1RGCYyqnwgO/5KlF+VYkKfDdY9xqd34S/AK/jx
WJ50XBmYn5ZG4/EBbBd6I44kdu08Ysf5foLn9HB44nXdSLeUk8aQaiZHdWPWVZVM
7jGZYxok8mom11Evj/9EN6MB9HyYsodBGxQEBVJ0ziTu//K8TTlZm93ORszPNY3E
+nKkVPfhDfkcn/tJfAv9RDzKGWLoq4r/WqKwZKX18xetAv6H93PhXqlCVCmKyCol
sDBsM6pPfQWySlrR10hVbuzaZYylmFr8Tw40qExmohQEK6wseI1jIid15PiZvh24
R7koO9yUbRH6Lvsrmqu2zLi4FAmFTTX2tgYat6u+pOL/D3J5fnqaLPJv1sAyACf/
xsCmNc7/XJqd5nwzsbrfLm/ijktZiW5JlT2P37pAzBWLPk0XS5RmtAKvMWVDQYDG
wjr3UMtELUKFbF8uHa1NUe0ksimH43booWbD5EEY7ABdYCUv/gEdcnJx3p5twSnp
eHCrwojbEZ4XVUnTgtOkYa9O23H85t66nvi5XXCxv7TZ1Cnf3Lfbu6el/izDbs2m
`protect END_PROTECTED
