`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tt01/KFE9l1WSLME9XRd0QeyOEJSO+0Y5oqpQ8vez/SjbsYTXn2ae2owPF/NX0Zj
W52tRtysACD98XUO0jHlg75mNGnEW1y7iZeNfU1fc+uMKZ8NxfLqz/rWD9yjALiZ
N28v4UaePHp/VuyKpbBlWmKGP0mWBFhobS76emNSxsgQwpWGNZ1Yte++JQiycj6E
fKZUnriOM4ToUhfs5aVWrw4RT75rbTcMm5s1MhRnC51ISjqg+AjtkzS05wpDcI7+
HXWEdeICLJPuM7t4GaBCAL5hOlpcop7TrBi3Kax44Kx+6waDe9hCAOsUnoTWiK6b
JXJKE6AHIhn02Kge4c6qMQcvENSTLQ+INHF1VOgd9g2FPw7c3Ua9aNzoHyTp/OZ2
m4cg3ZRmtbRS52wfcc1GPPbMtmrXcaSnzlouhcUmd5S2CcEQdBwqaBa5w44ITO5I
lKY+xuqlOjF72GvtlYf++lwKfrplYCgDDuTMkQIEEp8pbblQoSS+Kr1hRjziqS96
zPNoD7nopWmiCtZfovJTDpZyrZrvCPL1l8FtQsfA34Ts2Cq7spC6aQVfOsNfLkyM
hdoj4JmevgwdsOmFyKpyp33D30spb+fHoSLR/vdWMgDFoOA6Zk3k+AzYHKEPa5iZ
wTbH+1ZYoPL5zjwDlq4XqIhDcQYcvXQ4muDahrImADiRfL5xIzSlpzVoJjRxheqG
xzH4t/k4Onps+lQl4DSEAw==
`protect END_PROTECTED
