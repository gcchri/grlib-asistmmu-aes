`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0brQEHy0SZnspHGuKRL56v5hnaU3b5PIKEESvHY2I98cZbSwc9yssEzk+BSoEbi5
Zom+RE2WMREj7dm8XreBpBNen99NZ7DmMwE4lQoR36GYDAI9sJmJTaCTKhlT1kym
nBUpBUdT60JB7n8lfDtS33CE9aUqWlZPmoSKToEKN88GXAegZAZnGYWh1X8qTkof
OgEw4osUyHGuC8XbKYmrwXMJHtzRmrdAHA/D7fCpUnrQwNn+rKSOgR2S3fPjbWZd
SXi9e5VE4nkdG3gz3lPjPEUcVg8P/kIfeRalt6lS++bbhYF2tveC9PyPAezZ7vCx
tjwAapS2t+FRDLRgKPXBBYtTBYFpyJ4IGrNGqiwJ8QaQxlueJtnkSVb5aqEfxGQi
Vc3EHpjECXYYxqMu4egP0Qmt94q05PQmeNvKAaM4AzM=
`protect END_PROTECTED
