`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GB4LQErUlKTg3ABKc1GvN5qaDP7GoVD1rICpwmJ1sqaqVoxpTG6MguAFu7v21Z5b
Zmt3rubAQLZrxEjSINpOQLeChTni4WamsWlzIR2tvVrSswvkZTYMqVu/Q/o7uxtL
BycIVyE0oxIzNm2nONgFtgxthoOUGCtAqMt7Gx9XPRhcafBPNLFEubwgs7coRkEp
FK/6lxTHE48YnGoIEwPGcHuUK43MLus6/ARFn+Mii+Yr2Ki3byVSTi6UP3rty/s0
QHfyIgF7uA/l8GKPUjtL10/ImG4cFYolSI3jbfu7kBn0jAQh1R4y4+nDlZDgqxTp
gJJzY/1a+OULkx8CUE/MGYHs5WqtpS9DpnvBba1qipk/Yhm4D40Pxj4/+Cn1r3LU
HHSBRtKoC903y/OLCUlEggh5n/4WjqjxExp/onmTZXCmAdVYj35RlTKnOpLU4UHI
1utGSULSmlcJ7Op3loV1jeJQD9tJG4hrGBFBXtBHSc7qTAAxcKaH9rCgawk8nv2E
VwJ4fszK+n5WnA2jiK8pu0cj59TC1zEikpmmna8KYhZq7u2JrGMIknBY1wZtbe5i
rRiu6KW0WpPM9tfNziSnm3kVmjYKlUtwFgAXg8oIAU+XVqyoHletucnPskNNdTg5
I7ry7sIOcIwkH78JGgyzWu1PP0mmcCxPbcXwSOw8k3efjqZMsQKE4DNDcXBmOeyH
4+81o5wCdzmZRlis+DESamKNrOYBDiktVFVx2rmR/I3UfoLU4hGBxKTUhlchgJPN
278xjkRgUYADpnbrmJXIDhLp+6kVhH+6DeH+KwjauFZ8ymG7yF6QtKBI4nCqj5ul
6JEwY/51yfqNfjEWDmQ1qdA4A1lOjppqwor3T16crGS76T8g+Gp0xYiejUXlnj+m
HNz+9pYkBCi0yRQUr6uMjPNfqBZviqWjHmK4Jqk1CPsIq7XDSUHDkkAU9Gisf7sO
fXklYLFOi2qEBbuCWvs0e1c71rE5uFwvETljS4XLLaH9fCUJueNRIuf8UXJ9YQch
ulfyojylFihM2DcI32U392aQph1vd2qTP+lcMX9QGV8cFmm95Z3W3PKa6Lmvt+sZ
RYkHe9Vhj5FWFrIkkZU+Krs2zurpgiOozD3Ge011oGlmBP/gCJYVHDW96NhL0gFW
MLjxC47pdAIqU9UkiH+/MRN0Un5+cM8jQKiH6h8FWs7myrAB+ADddaUK6bpiJxY4
FPzydCGfrl29LQA+ksNI95qF3GzS7fC70EX1TLxmDVw=
`protect END_PROTECTED
