`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SaBp0mbVfN8c8jYcA9lthNoYJZhXsob3bgGNoJElQwM5q03UCmKxu/yxxY4bZjhl
IkSBXKX27PnHS54gPkJ+elz1a0xvkZn/SUh3niOk8E+1uc+DnsQNmqABQhJaeI61
0QHPEphpv4GTg0A/+gT1aHYhlhgR9xA0DMcGveGKHCtEkMVHiXCTrlypJahsRNIl
ycIOCtXofI6rghFLCD1ABH2MRTYMlLLYTmSEjyrHSgqdoyKUiQ9MBWNjfN5hor3n
92k+3GfRUrkwLzc81fh+7GTDwgNdgLCNj6h2+G/MCD09ESqcb14oB8rwpNX3T69r
SsOETOAFHqZ1Zw79Z3I84A==
`protect END_PROTECTED
