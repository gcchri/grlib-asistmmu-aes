`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4rz3aZRQOM51SYHwSdcfgLrAU4Xr7gZWVFfXdRs6qoneuTeQ8e42P+RitwIfM+lC
u1ZavzaT/puyCzrKMcnZvz8dXq70XremQ+euPVM2DWFMHrqp6hTxbRkBibR6cMrd
8E1nxpCLp2Cozdebl3LOTD0Raf/MbpXGoSvK0ZtDkYLxitziVcml+5PvbMnduRh1
cJfEJkniwZT9HdOZGYwUpC3/1aqM1m4RHOwZGogY2bXAyMQbjMu6U/oE9owxBOBx
/cp6iCsBKqjWWrPHA2roYVGe1whJ6jTPDrIQd8HnMTU=
`protect END_PROTECTED
