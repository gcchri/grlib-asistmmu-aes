`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
geKFnRqL8/louaiiV+Brvv/W4SXZ8nbcKg4bAY6TD1GbeD6cnDJbtvqUjyKmSMu3
uDOLXxK5A5S0J4mmb/T0EHin/l3P9KwxO7wvaa/RKG2zr+zAaRze8hpgapclkWDf
lQC6M/vsOBwHvpc5Cn4cLkk5z5iiYqwZgykGU7zk/jR63otyS33iGJHM2BQsJlt3
zSZ1YeIsUslwZ+wdeRz9ajwVtKFr6Gkj0o0hUFdsqYr3MQAQoceaGLJ40OCuECz5
E5bLiGQQIOZ3lUznkqVuwvoLU2PCyB39cj0i8arOjnfF+mF/khcyawEh+Bufdcwe
UxibzS6S22rgu/2PgtGHUZcRrP1SrencrAxahvt/J2xbTVxjxc6VsD9fyXLVRkBf
`protect END_PROTECTED
