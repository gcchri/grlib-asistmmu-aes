`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H8qFghbOAoQ5r7leLdOrBV/xA/4c6nsvENqBnVU8oPvO9A85rzOxBjgYkNDRt+1B
QfbEYbWEnnT5QKlyvYOYF5hHSPoK+4CIMkUdruAjEIMl0raPBVRL//Ok9J/LUEAs
p3U3lw1JayYfEYQO7G3mlMnClgI1mJA6GlpfEKgx84Do1tll5MbWegf0BRs2u0Hs
Q+Op9KyM+XAd7soZ9Op8gTseVQ/qgcYSlPWPRaa3s5FUJj8fwCPIKzPJmN4ktyV6
`protect END_PROTECTED
