`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P9B20E9N0L+6g3czD/VhUOpDF61X+tZ9pzub1q9j0qH2FzUsJVEXsyfpdmvYyGO7
l5jYHrnIkLp1bIwIGDC9suRDf65gcCapjj1kHJvbgdx7fSQR7eyluolzjN1MGWOx
317nQjkx+5ifrhJ7cyja2ImPSvIaQll+2yZlsG1ujqawebkjBhBAuu0NQG0J3tgn
lHcTSn2b4JClac1rzJrxZA3K9tMqFcUnlofmrMRUovcJtfNgqDISQxk9fYWIdrKn
dtO0lM7hDMbGKD2gVljz16Rn6GKBUIDjTozdwSmaf/YsHaIJakeIxMVPbaKZg/Nw
r/pvqyabkxRdVt9s+c0bLy3+n8k2hWNG3g9HQOkyTedw0ksW0nrRS2Wh8Jv1oSsF
`protect END_PROTECTED
