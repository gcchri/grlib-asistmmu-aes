`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9F7BVQzvlDvr8NTqDJ0jyOxyr6EYM/iJCBhuJbeZGeQALa540mcpBLKDKAf6KlOP
FsQEfycFEJbdzV6P9m2TSicK2mt1HS2UaZ2jR2BQvKSb2+su3/5mqV6Cst3wscLx
Rpq3RLxiHAC/oqhl2a4yMJL3cMvjLzPvosihsrW2mGDLoFdu2j5vbcn3hf2kBAY0
kqieQ5Ai47neokf+zruZ8zSKcOU0Ni8GVjKNZxivsfb8uaqvwCrEO9+Y+fI3/Iap
DuFR7qcZF7E9xoN+9QSZ2o8zhgjmJsGmH0b0erytb8dy5PGFF+Mx7QiAcBx+bYBe
sOQk7Z6kx1OdlWUrKchcY9h1QAZ8w3YBU+A57xoYXy4u11oLZ9fmONb50hgEHh76
upc550IsPdVBcJ4N0BCfkHzT5ToLvNYRkGg4dPkVdLGLZYwyK2+fPIfUN7hpajiY
SIaC/PXdKNvqAvWooNsKjs0+sMRcttQPcJGMD7wK02x53YYeLmjjfA+NvmRj+aUu
qjihqZJNXlnRdjPTkwxvqZ9ltRko1Nczn9wGSuO/6Q3c+I+9N3F8zzJWiy8LyS5U
wurd7suNr00XvaA55K5k8V7lc8szgrqCp1tvzUoU6Pvl2hKrK/wcUym3cT6Ee3HS
Ona0kwdrFP9bpVrNCT5zt0rWx+ZaYd3P4HHf5YnWrsYUeOwsOQ4HccZ/Figjt7Hu
06GQOcthHDKL2srwZaWAzfBwCt6xEuuqJeQAdiJ7ZwAkpoj50B3wXaoDxYMeF3DF
nbMGrcqUqa8M1/oCUIipcCOLBlhuyM9oTp0Qx6EJ9/6YSlP/WfJ8S+TXE4Y1sqba
vzYPoq0evPI9Cc2nerODHIWnIoEnjd7xb0wQRAnRma00vgAcdqC8pRXAMHywnjMf
MaUXXiHD3iIDRt6TkzmGPwSsTxRj0or4Kgi9QSLUdRi8Ze93ofKJUOVtcJ6Bqbbo
L8hP6Nyg9lim8jgtzv0plobjqLk9v/iMW/lvEYVL2U75vczyKassg9BRDbbvJDwu
2euImAz0xkpvF+RmDXIF81IkjpXhyM6veD9isMgBiggLSCfllph1gc8QqI3OeFFx
JNPVYaetIJSE7ICHCV4JrHruYmxlw1iXIBAcYeb4NT+9dkaYYDU53vS+FAdCx3BQ
m/Q+RC441GzFFQwPdRtgfCCdS8sA+Kv5YcKSBLreHR4g/Tvc46WC4DNfNMcmbGU4
`protect END_PROTECTED
