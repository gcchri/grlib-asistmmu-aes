`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TjoL7qZWirKE7K3/Sc4TE/hP02kgtoYMV2TuJcj94Z9JKjvm8EYVwZHNfwt2UoWH
Syalx6PVcCuheHNQuaB7kFwFmBhcjnQCDX4K53pg3Ie+XDjfuHZp1Nfm2+TkzamS
LjNRVprFOWFUrX9xp9nFKqdSgmT7aKhki9YBXzge9Nahj37hDOji+xfeZGCWM/9g
NybOejFKURduyymAwWFc+EtWWBSHXlKPB4NAh4KfHAZm+O/sJNrlf9QWKrN/bJW2
3jW0z1+l8ejhKlyPM8MuDmClDrH0+mJaNG6mr+nsTkoXnFTaxHcW1hj+dLe46spa
a+0N35W1ADmnDsbcJWmyOLOPjLHUhW824WhM7U5pcjl00DnaCGAhUbwRhJvoH+d1
vHe7F8h+M3qrUlb5b/xUAVI4b284aznnUMaawcBbKWyQMqoDY3lm+Xkk79B/P2+1
KnfqKxTDT1YbnLAX/exd3Q==
`protect END_PROTECTED
