`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QWj5zdjyUt7m3Jq50A3U89YZ5u46DXgDWf2/OVa5AbY09Fvtho9XXWd9itSLp48T
MMqMxaiOrDc+BJbQ2iUilQs4gAudllOxv4kLRNtwqVa8uhvOHcyLEszcDXBsPxFH
sLBZC2HBkkOtp5CrgQfjl7Abzl06UCOeSg7zRZ7xgPAIw9gQfIHBkapFbmUNT9tO
WYgLse4Co+UOOLcDrHGTH+23mdNmshJterzIVaBim3adviKSlumDmKkUJ/kFXRmB
L4JcEq3DR/J5rOCDJ+zN/sDAAM3SURGnN7Y7oPEjREeNp2Vp4F+wX2tP68knw+pl
do75mDlMdUXwpbNsAIVJNKQ6pA57gCdpwxbrMuEP/St6nLc5LNrueRnm+QgaRp5b
DKVcX51PihCCMl1Yujla9g==
`protect END_PROTECTED
