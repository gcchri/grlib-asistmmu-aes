`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PI8wBA4kdVX6JnRipS8yfUA2qmfzfuLwy5/uPmTSOOUKXSd0xN8weOsNP/QcK8gB
FZ8tF9UoqhMgY15Lg7q5X/SlE+c+PL/JK6SkmyzkjfNQnasV6Kpq8PCupOOsCilQ
WhBD+bGF+7BmVS8OJDtU3Y2tMWL/O1SloHEM5Q2/s6wAKfU7/JfIC3IyMS++3WBz
YodzXmiMS2Nctbpd5J8jlgoUZiltWcQdr3yHG4FIiEPtKaSbHIQchXeCKDawEr6f
DSRdOLsOfXBqugPNjkTKMaj1Ba5mmAw+jrXOlCv7z19VW+epIVRtG2agveOSahR4
ZWqokXBCVSyJAu9rFGaMvcWUiCdqPCC+mYrSthxAMK462oDYXJta2NrSWg7bNgu6
V1IohvD4yWYxRvPnM1lo10W0ISEmAG2AwbzJeB1DELIu8ENkV7wAye4p0+pzFzE3
0ul5IWCm/C3tyCxx9YRwZSZaXmplrFG5OFd/zk7mFrNbyDkl8W2SdmwXjcP2cElR
Id4r5ZmMUO/mdbCdsaaTFGHotk1KKdPozkiuMv3tv1yvk3rCaKWBdmzj0F0W7LPt
2HLQQhiRrXmMkYuTNCxNb7+cq1rzTd4vqaj1aoirLk4t+tkDfVnyb2nkTyAS+xC/
9kmjoYAcM6SnVn4gHvXFooCN2Kh8WtYrWo1oCp3IoGbsiBOFC3RNoENa7RdslWku
WAaJXBKA2U+GdRJr4QVW85AuQAN1lxmE4f0cVWSl0lkZ/FBytqEfEGwzWzkykX8v
MadVY7V053uKqoEr2TdYHuToGFlUMUwgEr6vB7ABWAhSVvJCse3n/+mO2xz//CXP
MlDfRKgetyZs407c50xEFxDwW31b91v5+BRQiGQrHrlxjHv8PRtICiO8HMYTgV6j
t6Gp6roFXyKyYn5jh7XBrt96cY+1TDcgtEPtVPXHlqNk/pXsbnBB1y5UnBf1DKJi
hRLsRf2K5IAB2QG271rm7NetrtHmxwPSHmHlRTbiHBKHbMAJgk0fx0DgUiBQ5MXG
doDzSIJNZZDE3D0TeR4/+KwKP/cfw/Vc24rlrJwbhDzd0D0n9dwCCGzqxnyoyt7z
b5SfFascnUBt2Bg6TOBzBwFyCXrUu3wTUl8c5lWuCd7QEAAuZ8Uud51IIrTgtGwk
trKSl3kKCHDd391FINoUaw==
`protect END_PROTECTED
