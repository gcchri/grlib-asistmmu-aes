`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8IHz7eo+mjEP4kGmsqptlCGrFvlrqsSahjW1HkwVDLI3+SuIs3RcqOhUWbqb1GwS
/vsxn30zUfxDyZqLzAfoN16mXI+jvopLt30FvNJ54JjDXxTPeWWhx0vSxzf1aBmM
/LnKSY4eKFw9EM5ePjfyFXtCcHjIDgIlfTLBZ1HtlzCuB2SlGoSGmF6vzkVX9PNf
Z1XuZk5qCSKei3Vd7SvBlPHU0vdY1PfYMDkDrUsxjlXwxzcAyCKCU2yroMT3whG2
Y5dJDEKsMpoJIgbVeHAwVhl2mQcvh7PV2p82ZL5T+WsekX9JkAJ5pddYuqo1NB6l
dIoMREoQbC+H4aNbhAjdijqgMFFOCqLpUPbIGf+jRpDalWZxnTx822xLEkjrNwcM
P0tobzl8hjS4V0aHJLokfNb4JX3tUsTryo4gOecFHetvO2ZGFJwyT8kVtVa8/Te3
k+ronKv5R8QQhpo1tJGg2+zEXIqkiZwjYq0+bOvIL/siQHb3OUil2mZnJxQ7+zb7
nhyJ1Eug6YNewJta5ISDFGvAH/OlOucyzXP7k/HzUavRoNglT4T0lZbwNn2NlcNR
QXYhw9pgW5O9fH+XU+QDyvOdypqSQ+dF17bNwmlaCFggxBwumbcvFNL3U1xMYg7K
OljJPcfH5AN9UNpsmjk3hmVQgyeI3b3FsLui+jpPk8dMEfsIw51J5xif3exk6a4r
GEVXlS2XD/cxfJ5KEZKqXy7IkcooQOd6SC5AVhCP8iy1Mh/2kZZm60rdBeVcZrIa
plz6v1w1YdN7N0JtlhX6eg==
`protect END_PROTECTED
