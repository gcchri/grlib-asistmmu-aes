`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cli33jeZFp+SETv59ljeQIr6UlVoOf39WDY9Z6VC81/yN3flW08e5J5r+4RSDGw9
jDNR/52C667lH/+sJsr8+Qv35+Q/FXmWbAdjLCn0/yAy+l9tbwyUFbEbXa9zbH+x
YBtOl9lZj5iol+xNfHyy6x5rDiN1I39cKGhTwYgN1+sgQQ1eGS20x/Vlajah8Gus
2/BxSZ3AguqP+cWF/TvOe2CuV3Kh/eq19VR03fgFyJQkGdrEqEERto/lpH/g47JV
bxShIu9215IgOxlHJ0P0xJylWNa0gJwUEzW/b9qF8VX3LWyTsKDrVoXJ5L7K3kX7
mB2DyzaknF7FGlKRv8gGFnIFwFKQDap27b46HNd8ij9EYSW0M7imTtCwIbifuBFS
ftoNmsnyoy7h/b4ufZrUtB8BG1IFx4dmnece6K/7UeuI1AlyMWLKE2EmY1fRt4KK
3BxDj8cL+y/OCXdsqDyxlByCb4O6GJC4NdajGlWStW7JW8EYUXdIDu8eDgRx3TXe
8pE8G+lSn9s6ojPzNLd0tYMWVJl82UQf1pf+Qziml/MrAfWwvU6B9Q8OkJ1JB+W/
8wJLshUMfhHVzqCzSiyZjqvCgINME7qA5eTTTkENH8N7w9KuJAMuinOd4271XuKg
jm4lCXI8JBi5C0bhl4qAYw6iKlhKW0P3BUA2FQX88QTSg86rXX5tOhcdQ125uaXN
GOmZLaXCJIebafHobKtegpsTXk6gRqyP9Nn1k6ITwmTpjCxa6UKJI5vNNPouht0n
qjLAp2T3avGmYue4eJZ2fkhw+1oN62FCpAefQFFqtY8mSD75rgDxPo306ECP4WCU
f7y0MfQ1xr3ld1NDq1dFhrmqOdhCE5ezGGquGA20wiKZoksJdx1YzCT5altwdtWA
az77D96IbCH276A3BaNc50up5ESOSzhOyfrT1iZw8uNEJKyESy1+B1LMb+R6lqN5
eHOWCpMyKdwKhL6q3kRt/Vx4SYDBT9XK2GEozW699AhKZeycqEx2AdZeWli6d6bi
VWAo9qWgmOtx/UxW6SCoMYPJwql1T9xC5J+9+5vdcZJ4ffrXuokw4KSTzY9Kyczy
ne29zQ8vW5lW7zAZSNerEkogCgcm4smulHuND/lXeo5YALlOJMCtcZ26E7C1fiCk
YL6I221w9SoOCym/hf9beqMckHUXCX8A/FarHGOgmDNq8raPRH3+HZQ+9ySyS96q
v659wFli9PV/C3bLIBpA5zKcwZcCV6CWYPFY/cLKVXGtJ6z7qnvAuRjvpRmCWnTs
Q2LwfgoD8QW+1OXR3C6B0PNXd5tpH3AYaiIDbcEUq7zNUIjrDP37TOBIW4qo1RyK
Px8OPn1FT5aAYmAQAf8weknt2MT6+a6KI6f/Nuoz+nmnXXxGtuodfkHk8LQuGdHV
oie0ML2AMiVP+Z8KviWiYAu9yWOoWGKbziYYkEW7dznUbBHYfFRG/1WO96adXu8x
w04XAVDIQKix/q+F/azHb6TGLGntKRzQO1WB+Rnm2kQ7xXWm5q3qd97+iMbKb+Q7
x6Q9LGbxetunPZHqLFP7STGHzGn2nlPSQghwtzPbf2e5wmFNnMeo43GmCNrCWS0R
rKkhADSUQhLKLcdHmnKkwwaq3xcQcDrjdtx2U2btGnNLv8tVVA8Jjna3wmUHYJFc
BS68G/RqnyU3muqVhK7khA==
`protect END_PROTECTED
