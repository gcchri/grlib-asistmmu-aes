`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cVmM0himCct3YJcKo50yo+GMCmQwPbpUy0Oi9bwn8QJww68Msv4IFkgPo308ZmAT
EG2Rrzci6R95GXM0xRaz8wWH9Up+TQwbM7o2s6/DecIL++RHV5uylLedRCTXkQPD
wyk48ea+zqNvd4ioQW612jNN3Agow65hTumPzqGnLTE0C9lbUicQqmt48uansvRF
XO2Pk3QwaeVuFQzDSry0YGq6EiosVn7rlvDpAbL1TYC3lXpcKwrd9YnCvcONV19V
LHO534RLZyw8pVB4wyNi8vPKpEXPP0NSB3GNXSuGEM2/CojLwDevnIgCV9zpZE6t
TtTTNtX/q/PmmYEOpT4+4laWxyCy9ar+1hWa03oFule7NvsTPWG+hZOwH6j7R9/g
g/rtoZeNcL3EpRDQD1thQNnppWwxKTiuBYSX81rS9iwdtZECylnbtyLvoky52v5p
rNzuvdEtSLSQM8LBZnnMsyI0jtthONoaf8bMlJgykNbVDdv4/EnCmyUceeIiHSxl
I/ONKQool22dAj8jgQ1bxvVAFItNPXZmcxfXVDyiNKVVmEYdJEOg+GjWt5HDO4nQ
moCl3P9pXJnBMzMBX64FjeMtEQwHfIfOJRb8bwB9TQGhE0ptn+ttnb19kdDVXYUH
zAFHWKWjFteInvxssMtiuwrzVS5E75Qi/wdtidClec3o+d53asKbQ4bgCgbM6HRR
Xtfgds2qpVU42B7h0rl79lRa5OyxAkiLmw7L/+wAYL0=
`protect END_PROTECTED
