`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mNXRXjahwFjYVr693mjrb8mZPCseRkBn1Yp4yNr+z75m0CoAS1PQRCMMK/f/76HX
mbcs/s4UUD+CifJvLNXg5bLUUeNy3KJE+0Gnics2zewFKway6bLbh7n8YK+m8ekN
y/EluKh9jNSd7gWsTQBfcFElLaGRbEkPfqajR51a2WCtFd8AjOB4mjeeYVA8DNB8
c4rK7WZggiQQcyXoaiMx4a1/TvDu5tzsm+Bmkri8JqwuVceD6DU+RHRvd6sELUN7
aywQ6U4115DSna4GuodMx84D4NKCQPvYdr/7Vo9DqMBba3e99/pjG3EbPXucefoO
qq8chwSdbctLsDAJ5ookHb2Hxz8tuYsQn7zmnRk5dVI=
`protect END_PROTECTED
