`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ntjGVtY1cq3kQo2cziXyGblhhUvlBIsd2iip50hY3UELI5OJIBcbMsajUeA1fblV
jKmVTSHw3ouVndUplSWXEVlVO7uN12gixqj953hKo76PorsCSmzB8NnlJUBDlz7g
FICe+8/xYAoSG16wyZThCYMXfcBf40smLKaO10QqkyGmUHxNeUs72dsaU2jSbo3P
2en4rnBr+L8J9LdK3cg1RscgFClirb3fAPyiWEBQ+U3a3CrlxEorkN3y+P2vkU2r
FRXYVDst3v+niczdvHZiL1D/bJ1LWMnEacYLIJlotlvDgAWqNL9Ixc85+9pQ8bA/
TpZQ57ivCOtAiTcQf7s+6ok8/ww5QKXmsJ4/keLIB20WDCClV09X5eo8agmxhOEC
Sfl5Fc427xlZnxWdN/fQ9vCi8ZorFf/C6uqOw3FI3nqg6jbM84jyvaxtaWzE3Y7/
rUiHtwPM+VncWDAzFUDZh1taiZsmCN8zXhdl996EsrY4A7bZZIu6ojAqFnHoF8JB
XcUUrB+HweNG1w3DrvcRyUHdPBzwYFZwCLwgkntzKaFH88lUBswAD8dlQ8Aqdmb1
gQiMJ34cgXbJZDTJAD3C/VQsn42pnlP1AAfojZ0shHLsjkz5Gdz7NRi3wbVPPZLP
nw269/D6J9wAlaCwP/bsovreHNjNdTVmBJO84zZSGW8pRSuFa7Xdl2hEzOJF83zP
PplNzTOU1R2wVRcVRnRUnXPLpIzPDjmt69Zg5DEV87TGg7jFEDXAALS0+1GYa5X5
LeVP5tyRYwn/DXJIEmtXIqFbs0TKWAP5QlWjBDVra7XNwlsnYJtvNQ6uhIhX7qHY
pFUcKtnETG8RYjeNaGC3O6lYpmlHEv1vEbLdat8ph68=
`protect END_PROTECTED
