`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/eRNMgjrHttlhbUbil37REihOwm55INPV6fF+WyV/Fid4bho0LIWvwMwS+6pFa2a
jJsW1VqxII7I2PjGWnqb4kxy4AuCVLsXIQc6arLddfIRrHofYj6wn5bf1fLKutkX
l4ve4xslWld5HbBwupgDwR5qu3pyxYFQ2QP2pU4ZfAXwhL/4O6Fp3QvrTU7BiFKu
uYMa3XqqD+exc7iEReiA0f/RuflYtUNkSmXMMfcT/Zjffl/Om5dlHdTGJhR/uoQn
hZyhAcbQ0UyZSA7dZU1pJcBgkKqp8cApZH+n7sJ4MB+DdRkUv9WUBSVzI5fHPajc
GA9udISPTpwoLqE22hQXmYBy6xz4AZmgdYMOdr/1Jpp3fMePOz6VnPhSSQojgtjg
/ODmESdaIrfmeMcmyYcGDf+9MWqLld84tExfqrtngOvYUa7wBAtGRFDu5L9ciF9R
`protect END_PROTECTED
