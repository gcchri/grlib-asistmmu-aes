`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4bgw20kN3BtrBR5htjnoC9HW3sxnzeAOkeScJRRe9T7e+WIp3Rymh/6AWbCWA7FY
qEmDiDu3Brh+JITcmG86w23GAgShHmewuzcPXujJtoZ0h6t8Dz5W4DIt9akzqyra
4wR4KcFvt5gmG+FhETZbqsB34MJt0CsmuzrrnGVXpnNnjHdivFe/WzqaicbAyTBS
+JehoOMNjncAyk9q3uF5utFdR8V6hIh5SdNasINP1rqfSI3xdor504x4Mq9Ht9XE
LY1lIpDLR/K+OpF3N1Lx0lEBx9HWU7J8aCQ9JTtLyDW9rL+4XsYOBwvFF76qB4Qa
hohkbsor00/PmzdJiwUjJ5llfMcZGglI2oAWYCz2j5TSMkDQtxqFld8A7lOC1El5
58sfs26aL9wrkJhzx3kMI5VgLZUXwZOr1wm2wFQXLMM=
`protect END_PROTECTED
