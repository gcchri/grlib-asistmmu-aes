`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PtbWEPFjMNl70CMu734R3/QJBNaGzFU4pIstxVPZT7EG7PNLcjrsHvHHxmFDQt8b
Ln22gCYVRZ6ZmrBKDFjkB4cFuQCen42tzkqIP1GY8yTHftEiORO69lb+hisgIlI3
StdxgPCn8i8BOSbXR6cv3kQEELVZLobkvSaJu55oRZcXUquyPPyrdkTLQsU8B0KU
WJqdv4COjClD/eqFwt6ypZifPrL7LVSR4PzILFg3tJMFNYogxv+AQ56nCqKAkVMv
S3D691yqllkfbg8mr/y+K1MnBMur63mLToA+KDp6ijM3fAEmgbIzNNAEIwlcvBMz
Od8LXZZZcE9OYDUWZDVjiH8KDlRXlaCY5Itbg5EzGrF86x6h/qPhDajPaPce3Bfb
6Bt548jy/LdUcQ8N17zNWT57DXX7f/7/Z2r0/27elCTXNrqfyfc3A/d7abFBrmby
lEy8b6Et5T2+h/NKQ5iX1g==
`protect END_PROTECTED
