`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MIOMnd0LWNJGX73O1fqCqGUweHYZibYJ7+5lpMo7mMhr+PlPfDoDxXQoALoZp9e0
nigYXfo10AgtwS4g9dq5KYAu6afsvd6GFjVS7JvDRCrY3V+vSc1n7XpmIpZpQp6v
6dKNcWaobxMUl+W6RD4dADwzoD6pldZT+PECwEs4HoqYcc/Xy/NHxIW1RfFgIYhI
ZBw9ypp2Bi0PIF0sck7SpBNo8Pd0W9GqAPBIjowE20kZR8TNFKv3gb5cnIInzs62
UlauosgaaIUXqG/YYwjzD+wdpRlN2K26OS8D9xsl80nH7Ekb8moyIqNyemyOD74u
HqBWeVksILxPzjC6qXwO4NhApi6KZlSE+ZI/hm8QoRuwI2OVy6ZvmpYIif5Pcgi1
aGHM5nMMbIkmDMjcV00NtN0h6E18/XE5fvuej1kFFm5irLn18oREOQlad3rTHcG7
9WCHlW+rV6ePks+95+Ry2EG/RA2I2OYMbGYcSJAJShK6ADTOBj+wdP2L9VigV3Y5
JvQPJoj04uWLZvrou7jod57QGzQBXuUoYeY1c7Gwdfkkz3aUEZ70Suqvj8RNm2xf
OhnRm/Ju08J5gOnmTpCIRzFL69qpLwKo7dWIWhHpIEPI7E668TACGbgg/v7+mOgH
b34ZmU+BQZifP8rX9Xy6L+RF6CFCnRA07CSktG5eZUU5+tQGaX2SPEoYQ55CpX5f
Yd4mwhW4XEaUXh9sCbzW2VykGxiZ4m2zO6amxQQOnsZRNetqfU2g6FMSQTGV1uHI
NgQIeo86BVAZ9m/39MUUvBM7iM3bRCEayzIZQQbyroCClSfm7yMDrx7kui19s9jP
7fT9ttzh8KHEmjrEzvWyNifU7yIT9ZkfFzuqKq+b6Y81zMHs0phIU2gtjE3b8ZQ8
HajO63tis2QUaDPqu6Z8+u9JN59QW59Edv1qwGZzaxhcmAUWYbaDsgl4CeL7jNj8
NLNL8il2UuQgUqvmurSrZxq5xF7n2ThgRrwjzwjsddGgz9cy1sNxGh0KQcXJzAMt
0uYaB41ndU2GfoBgT1iRrlGc7h/gVoVsHD5fCuE/2ntUzPppXbV+mJehcWJrR4zD
GDuwty9DvEVnd8Ql1yEPmFTVDLouMKs6hAPcPUuwdEl4/8J5kB3gXESKDfRLGO4K
NBqzZSjpvuQJ7ohnMUwhy3ZyYPj2b5o2Pv3Iwk2dYgyS3T7BzZ7dj70PdUA6UmWG
JM+C9K53ytLbCYkYk0hnF7sr6WaQ2cPL0ChMejZ7gnAZQBU+e0TOHzgV0WkqLsT/
dCS0j00XTl8pQdowEyprHmVzEWEeeDTsxx2DggippigoNNmgBuTwquu4H4Hd4jC+
xrN2373U4ahBLiDkNlEP5V5jW2JnUWMY6NZQPTeIAT12aIdf03VrXHYDom0bOp4H
mVj83etU5X69Yhufq9ewB/LyhCJaL3FPrgn4eB5pzrCw2ykVt/XKAJTfjCK8+Dsj
BzEI8aNQ6DpUaXr8rdrpGENkAtTi5pKJg4rvLQkNP6c6ofGUpB24xq/ZvgFeyDD8
YZsKF3QFieSKVxLn+ECMseXTya+1p6v+ivesLcud/SeE0S+TCHZFLgq8+cFZ74al
kGjDpAwif5edqXVb64iPKqALt2z4FvXvxXDLmFQdEFfrTPI/by1fZhp7UhQPnfRd
yLpFOiK7WvjPzl//hns+ioxHN/hWWU6nyMiXibxjelzM4SMDwi3J9VFnz39oHjCk
5i0xap0+3m1sbGyN5jtzvyNhXsLDTr7aZmsT+bzDCweiuXyu/OzlhlftucoRr030
r0lNU9o1+elYlghD70KhwKcxDwGJH/RIlW7DFxh0d173qftW3lwzpniV3Ul5iZes
Su5/aoAWloyhwu9FMr+QWJqY46xTeBtoGk49KhcIUXHo+9tNjaVZ91ror+qEV07i
w21wZnTUakKzRtg0c5Wg+0QI69ly5kbKPXhfaCRCe90p8iqcG1UItbPPNbulKTK5
nFC5u779dzBuCAoyKhX4Xgqxs/+cHHNV+GvWTEc8a60J+KhNkFT/LWOgc17DrmsU
t3JvuguIARFXO/6VXaqyLrsXwBDJxEElXYcu4YX1W9j4OVAa95w/BLXT+ZG8UigE
nVUKgRGlHQtGCTMAYrz6M+Bpnlo1Zaj1WGfd+j9w5A3+u4Tx6lDexlsCE+Ru2Vxv
KleEXB2Ost65ygxRkJRvxkwpxMIQf/OWB0bIcQS8hSSXKIeMoyy/jIot++cIGxFe
3ry/oLvuv1SPb+ZCwE59IyTPzE+WRN2aDHjvZ3k2482GWLkXJVESf27N8JQiy/5v
4gTWM0qygrJrzOnnkXunhpaR9vxKaacsQj78s94LTg+Ry6QYyHq6r46b0l11Y9D3
0Ihd1+bbdC4K0GlDGmBqhL6OScCwzexLLRAp5x01ZJrKOPOR0Rayo+gs/IHu/G1A
VvFonvBNdyi/pBUKWqnwxXhwGyNCXlv+QsyClTixSRE+Fqse4ro1k0keDL8WzlGA
G1iaJ98X1kYmxrr35YwhgvFfTnbBh3I4rq5t6gZ5mMW/pL27ltnd3GBCp0UrnGXs
g9w9Mcq2jxVLKlR7LrKOOTgGduLN3jUxBnay9gmWX5DCUCfP6MjxMSdKR0Lz33k6
Kf0Jeu8YZH9ix+26qr/yUia2856cg0q6JaiqhycHe2EDZ5f3c9z/vvpCGJH/o0Ck
44If7ZnDOwvZA6TTq0STv4lW/Cddf6Dx/AES5M6XFEyFNXvhVZGqn5po5a5Uoy2s
H6pSj9CtdyTTAMAaamfCzISEhEHzSkpEqA6KnVjKewcFdrm6m+agNtd2wlW+8GUV
137yXe4XHOHt7NDYqbGJqo8sSiidQ8ur4WrPCTxZDAvz3fsVIa6idfv8zULeR6wx
HG+KDmpx/XpniQIwQTU3MdDrkl5rWaTPRyOSfHHheX6LB0+D+W/k/d0iP+QlXxNm
MnkhBFRaNFbyvuaBBI9Fou0Zi9aoP142ICEFABwy31953403oGCuB8nROgSLS1L/
eGSwIFPec9kXogcQIumg2Z6VCI4yImnizmunyhAhUB0418uDRDCYeVrs8WAlSl/S
ebaQFt9LpDghIOh3+7o3x5O66WPFEz62WB7Bz/dZ3AJtrTBZ12JQoNIHNH2xTIhD
/ywepRoNlBIt/R55e2WtMLsBhRLmSKHeRyTrjIKMZVkiAH4vSya4osj4W0yP+NRW
QumBcYUfe0822BLsWyk156uZRITun2trniUnSKC622OM1dIo3PyaICrPX2K1eqUh
g8qSSXjt9g9PENzGk6c36ZOAvMy0nGn42d+dtOZto3KXfym2acIIFH4OIXE5LIhb
reYarnpsJrHNgmBBdAYLbylz71dhy47w61FvWu/9QvrbkVEdNDt1vux1tHLI3jXp
ip04QHwW8dickTnCZx2MbpuvHQ05zp0fkV9VglPB4GH1ZuH71VAZpEiX82GsDZUB
DxL/baOJ1+cNV8H7OboJOgoTZ7n8o4nGq9+Opj9fTZiPjnYu1N4VzxgUmmmHLlEq
zGAA5osAJb+cQvqbt622gBz3S2V90/H5eEMJ3QCaNvhaFFr4yas+Gs7CDcqNLsCc
tw4Mj1tZP1QRwRTy/7XW71lkStzn83apB8Jpswn8I7bODqkA6foCLmgxCK96Zt+f
hyzAHWYUldpkcww7lK73zQk9oQhKpefZPtGS9Uy66cNAL8KuYL8cj0wPCz2Ac+hi
qlkgkyenYgoEU2IKwDRcHM0odFX1YrKNG8ykKGDlU3Idk3W22Yy0TQKpcKgZFoNT
tFq8vkcdUxpcPPZq+dbAJ80rLGh8v9QP4Dvi4maQ/jppS7sMt38EaMSFDDi+SQTp
3w0020Yyo14ccHYlXikqxjYoUU5gedZ5LjaPOge0SLq1nK9DXSCe8iDly/QEKYwl
gUIkoVz+GUbGilTQfbCSQx3fNcMF5+Chzf0tCHppZGzreG8HAM5O7+5HHdnxiK1F
Y79BgZGCeve7R9yE3mabJOi7+MBFYotcf976tSkG6wScfbYUfvFl/DzPqg5ffdFS
t6pxQ1FqHoD50mSDsbYcyEjzqnXpP33awPceVuXsG/0d1DRy04TxsU5h0xpDDmkT
Z5HkWgZ2mj1Bz42PHXmHh/CqZuXqYvDA9yMRoZ/YOFJpR/MwIahtEQuK+B2vD7p3
FfMThSVLvTre3enXbwfiBEQzSmNdOgJZDbwscG1sZESzQyjLPBFLlEtBLEgSH62V
+MISWaPEhWo8BiKk4o6K0tJGD6isMiI52lNq6o8ywXplauDIaPQFh+CBiAxuNafd
+XYz69w5juK6yBMATgklAYZigs7yRGd/eRFTE3HgVF3XDz/8+GIr0rUdPRvTRGsE
iaTOmwjwgfiPrOfLJRChQUPmL/SE3aMfQctrzmeCG+KLnVlCnKf1yPD7EpEae3jG
c/jt1Jr1TD8nP8LP4Fsy0aqCgNe1mkunwhMpThFRTmuTrYZMpStbcOnnSjMKH7ZR
sCmEIsKpY6vHJO4eTOYZJWdIJSIA9kX3UUklhTExEhZ8L9+0x8SJviUKPrpDGnT2
muJjlDGYXJRJ1Gp6hU+4QdmgNTklCbBVN69wsG5FFk614L0usJglqC4Mz97WYffc
dffNcIssG5rD1185DTlssx964M62uJpGjoj4UeVraMYdlSy81G39Xg7Uodvkbvsz
s+wZdMje2seh5vm85GEvXtCR6IKhXZoaCVpl0WO17W9ToRbLX3wyOvWPqUBOJIKG
oPiWnnGDJPog+apeHJlkNWtDXSDZuxfMsMOa/2FWC9TbTL7bwAmm9a2MAVXij9Op
ygDf3+MjlWBzl/mnzmiMFFfqjkUj/B2EG+17SkeYPIRh2+8toHjJmPYQLmaBYCAr
Lr0e8UKG2HfW/YTUN0/tHUPb7RI8zynSJkvUcfbFNvZn74v9f71jxUo5lEIAx1Gi
fpsqchOX/pMczXIYnQtX7SjBylKFnXm0vkczFxfjx/jJliqQxMhtdn9g0Oy0ytDR
kr2uR6RDaPmQA/VBIefh7Do6TvCMgJlu8tikLySw2BCE/ey3QYE/tL41Q2HAKagS
B8yQYKgM8IuAj9ECp2pNRyfH1h3u40GH8NXh7lNXFdaHP92jOGMeYfengGLPkCAR
l3Qd3h/zoQDt2Fec+XbfWfUICIjenId5P3ddOnwLa6I9hTkPkj5892GVL1o8Nmop
HB32giOr7uppmmZEwa42vx17PRwc2AIhNzJUG+TiJGGoHHNQEKmnSQzgppaJfwCy
M96BkePOQGn1d6cedpipKY2+oiTU+aTSYAQljWUOERgQ+ZVEjLlBMtpxJUr/D9AG
z2DVx166u+VLmN+Hl8c3VYN7GsbXLUQZxebBsyPMIdYKtU3CppgdMeg+mL+XDrQ3
rmwNB9u1AvMyR8gYaiQbisCcjroXVEMPNSx+xTNjZbMPtyobUe4fdQNSMHy9dBfu
K1RAtYgyxB3p/ie8Es0CtNxKCYXVpjqIKOsxyAARUIz19smjQ7GMK+Y5BC/9GNTT
B7dMrHBbjLQJfDY1FN1rMKlDudm4nmXLKN1PUe7WN3Q17NS1kNjH/8fbIDELa5S4
U1yrgT+Cv2qTQX/DlgrWBnurMNCnQ7FCrUANXZXEmieJrZL3PkhNScD0v+FLzKEb
pjdtskAkyd4KoHLEVpTH707BEElLFWRn91CF/Cii6i/UigTca44JHn8Vc9uI8bCU
nWs3yPh8dGo9fA49alQ0Zq/1eBFNpfQO2JoyWrYqbRq3coLPpa4Jty616I+UqLhu
liynxmXkpVER3T3GKi1i4Na8UM9YOZwhvoZNWQ3A4vTUGmuG+j9F/hxA5x65pj4q
g7bw0Ce88fiR/V7G8KXYrJJ7Rec6ZQ/vO74enf/qL3AUDmwud6FTkQe0NHpRf70i
Q5X5ytzfuto9bFnEBuUwNlJYp6REJSl3jaidbDofki2lwclbeIZCwjDf/eYZ8Imm
UbD9S9359k9km8LKYOeHyxSw0IWuBnkRHc/2069pUnFWrn2KAs/KnolDx1iS0Pxb
ubVvBprLHwQNHV1meki/akI4Z1wJgW/v1n74afEArP3SxmKkBjMhXjdBg7LRMv/c
TQdwe1oYX1xGqgAhc1oaUbSgdku0Y43nqrRvzQPcSglprKaNXmpkaa5nBXR48bos
PdvLF6O+M05a607M/WvoV8PfDPz+iqduyg9RrjGYyYlE6xXnzHQWMooKJ/DFrPuY
AXxT02NWFrHqSNYmDYZC6DdgOqgpDZN9pa5VVBH7+7wP6DtBJAJFTLJMvFRip09n
XtjcV9x6rtWDaFZ0yCbIrbiAezW1e2yMOZzgZgCtoh+5wI/GLWT7hLaWOOvRVMmr
JzYanKQQBMMQY4/0xjUscK9gTnxji3REQrx2T42p26ftRMkV7xzkP0JY+ywSbqSt
WgFSNQSnLYMDvkfvZGpueb5Iru6IvZmSNT1J85GIKop+7OJyfRgokUxRs5HBgOZP
NNaUqLkHN3UAKh3/e5388LCTraryIswQQlfJ/WXQrn1YF+Ek1KMyyWSJwqRSZwQ5
XB6nIQEwAUSK1BsEGroEXzhDvImHrAYn5PlaDO8Fh9l1HMUHJXL/boYihlVGJM1G
3vt/BQB6c4smANV0pdgsDe9kv8ffbL/1ZQ98QmAcwqPqETv8ZCGqv4CQGp3/Cpw/
lCEv5Tx6SIOTFaDE11HI4ydCv9Jz8GLjB1/mX3VroxcKjUAMb5BhBtseLaznxnTw
50ICl5LUOPlTUjEGhN63stBJxHAI7RMNUyKl638/86SfYk+EVcMPXBbxw7cPl3O2
52JTDYzCfp5OQ+a69/CxXyOzrpsePWBGPND3OC7+h1Mi3nF+FmSVg5MXYLf4G4OO
ar0Apnz8oclLO9oHx9tNjSZC3DZuJ8qQp5Md86iiAS+yqbsqZofBm+uYaWvps3HP
acSVsC5eOrmUPLWKPgBPQu5WnMVH3hr4vzgfmcVUvRnCKYTgsI/PKm3suClp8aQZ
65Ov/+AuF2RyqK9HWR7wwZlG7e0yAghppwEqr1Cm5WRK6AVP+PWn3xaTqV9PS04j
KopvBBZ6ZNNYC7vBuKMwkFCxU/v6/YpLuDjvoz0qURvLJOcaXD6bbJWRegnrceRT
v1vwbyY/po+NMSKVxR9iiNNUL/HXlmhLJ8GFvFQ1uKoYsgcepBRFb9YfrYrj5IqD
eLYDyh/3dZPVkEfgWyb+vm/x9WBiM8vEPFLmrNFRp8Sfm1X//E3a8gekOvX08LKr
G7zSnrGWalUIjMgquwCpqus7zV7DoMtUpkVUCzlfD0NFmhEVAP+MV6x0USEOeuIr
LSUVjD1eVZ4pOp3WAmh1h2CHXZ3lr3t9sruG4WunrmZL98ebDze5iUSYfWBeEo9H
8L/NTumow04/Pwfcq2BQwv3K4ufqp5xLw428m1f0IBbjOYU8niurjXx+T3LmuFkf
RGoJWBN3MQmIHOrdpx+OvuknhSFMyztFJMuGqKDlCAT1nKtn456EOfgN4dqf9MbK
nU/4H7IWQNKIo7iIKBoHCTmYzk9qpYdmja8cm/Wv6qbCZTos/d2K0CVpy4gjjAKm
QCjCPD38LpK3x2BY3rHFepbkJNdvVdlPLNN2qwWFwNynkEAVvQGucTDoE5aN7fwZ
7vG04YlecBEgESQo+ptuYYw18FPXP10Y2XtJJ6t1DSCYMVZ1eKwTeUpenJ4E22TZ
rxUE32U8qmtN55eeEBkHsVDiEATMd9J8b+w2Vd5ESgCgbxzAmBzFDddbQ9Vy+klX
TYyqtnNrTbwXvhQAoM7gbXgr0fxOpOoJOhMWl192r/9puyrNeWt7wT0kiyf7xVsD
J+kpq/3+cAsJhnFXDEIbLwY8VpgIJSxw3jgEfiW/w4YUgroiPaTYTJ0CK3UMeWh4
bRrnczSgh8Um13PvKTuMaW471hRS/JgEIioMSX3gefqaSbJPwDevmd3GWeeidn0b
U0EiIIP8euq7f/Kx0QZPRyyXIjz52joHRVdQ7H3k9GfwxQVxcaIyNbcPXbB092mb
evsPFmjD72tR+HicPJwWyC6BMPeCStQQBNPHPZw7OABHtdTdWS6tC5LzY9lCzYuu
+K9IapvpFNlhBOMk2t8qNgk+YT8FLsKDAna8q8HUdOcA4xEgBDbmiDD/vTZenVoA
qy2iN5azi/PF9A4SSzIRceIPLXhiPMdLhZ+YQ9SGiivmZy024uRYwLRfTMJuXq4H
heU72UjMXuQwp3Jye/DGjJRB/O3G6EOdRl8Tg3UKu4AnwjjJRcWdYzJdigDtFo3v
SHx9n7Htiu/A/LxItTQaZQJJnD1SWXMfWDmmLdVoGDFxPWxbTMD3/Rllj43YNb3J
c21FDdv5eS1zyOlI3l55+j1ZyXCn7VxGkpTmZJV+7imKU61RGjJAQjtOlP75mR+G
dFIRADSNo1dLO6c0B8B1jnU+19hJ5WVHFw1xC7N4WaVgNuCc5iTLvFEmyy9cP1fZ
Zz6iFk5cPvpZdKY4/FHRb9DrXyfrDPT7Kd2OtFpNFPwBf7gOy8Tzp/5U+SjAx/r3
jyOxfrh/WLjelGfdfkrM+rHvIkOBMtVzU1KbauoURt/JVN3fegS4lT5sAAIoAWTE
Ak3KUk7ReOkV/zwr4lXqafGWHlFvXnMtFNkjbH2jEKdhwZRbNEVms5PS/Bxsec0b
whSKeEy6cHqD8Nr2G6Brh/NuLxlvwkMTrb7nDa6dgVoOHQuVD+X1mImfGU8+YR5R
kxMDVBoS4/aHrRdaDED2Lf6oFynYcLCO6RBwpCpVDVVGq4MQuZ+6XgSo498KL+7m
0cCHHIM+t2nRmDJi8SoSoX3VGkXm50+lmALzFRnEv14W1d01wMbVjVTITnKJN4Zf
8p5byXCsNkFJTWA0K9PyTLaqcyDaLJ0IU2/FOn0+35mw/WFPBuqPbDFYp0mr7Abt
ZaaNuMpmgCUkBOAOaT/tm33/9e8JXgYW2Cxx9ahZHtNlcVFtDa7PgpCe8QdeWeXC
iblHry0O0dGm9JoAESfPUh0P+PiFcVCsuTh2xr2m4PnjKghejhB5E1w0ga2SEb5f
ROwhoC0uVkNFWHtstVaAvTOzPgSTPsnTCJ2Pxr+rqphglpGz8+4dbcclb47Hjn7+
J99YdFlEdHZTRWMRoLmK/cUcD5cQ+1kzETEvYgrxkWhTbBqKBHMeHDLLXh5A2ruH
lebmBwU74A79/jTBEgGNJUkrO8mpOTq65dDldnqRbhSARf7k37UGOaG7c3wG8XR/
OjfgqBdbaG+NURJD0RGlfkUOHhUbdG56nJNAY6FnYzG7s7Yp89+LddgGsqiOfZ/h
d4CsrKVnccowCPY90I8Yxv7SGht4AHnNnDBuXEYBbG1m5noeBmiLZPvs8cXSOabv
LMgYzT2aN443RRVvSzj3dWTXEJFQ2ScNF8FI+Q0t4htmO1YUIFbsbfDqV0uk7cNf
D9JJkNenW/d4VBmTnNAdeyfE5ZwS9HSwcQW7emD1oVNDKyKLQGTQlvtFsuA2OeBe
ikn0+jw31EaQv0cjnMVZcFQXK/b9BHwmhTecnLxeeyTq1nSVG52tk+T2dzqB+Mu4
N/OcSK5JTFlCHlNEpgi/Mwk9p4c4TB5/snDgcFuQyXtPL7FOYit59cDlGmHYypNS
sQ6NzmR8r2d6kiopKRv6SgDeJqqVueBIrFUEbxcRJ0HqmA3dJotPuOJsI2VlSEKC
uRtd8ZOOVZvEkHTyzUFtkw8PMp3r4+3tfLDVjCoDurJHA+TbRF1xCtO/HRqcLz94
bGKQfjJcNxXDELvPc2DzrTmwmRcOMzgWTBp9nlEsr072XBwGxCbZswtaff1gNFru
FTf0jLytHcxyxUsCjUrhZhCDBItpbocBgDu7e1wTjOCot5xR4HVfZFnPzCNDqy2R
C0D2Nlh9ChdTRSY2uZKVy5rdXsE8AHqSyP975njz5IA6ZAXyP9KYixo1XsQbJKZY
oR5h6vvvpWf2tMwy1VD7802a45RRX6buzaHziGyYmu9lL5hpFSJI+gJDKYWi8+Ow
sPl8VbRKTWn/hV3mYUGrNitUxf9woK7BaPh2dNOs9gUKS2DS0WxnsHX49/WF/mPd
KkjHfUZAHfKOl2Z7yJpcgFt24uIgLvL8cu5YufEJaySCVNOZMyR+o2Mi6A/Z0mHx
OxEhqP/dQPWMxyYLwYl2KHYli1uAkA44d6DujuDoKa1Akgl5XHgZEV0Hb8GrYpMD
0q6Fc3k05WDWtR02yq9mWyYxswwiDLriCDERH5aimPLFMqvgAyG8kt6HJLvk4Hos
y6cQO9d6MCBzaGYqKfP4uFdEKXE2Jrg4TvniP5TwwpLSCe3Zm0wRDpSkL7CMfvAM
3PRg7IFbbxE8XWpH2O8Dc8SyZJ9r7gCMZ89PXwf3ViUe6IuWeMOmCXh98SYj+CtX
OM/5LK4t81qvxje0cD3D1bzJTVQP5QT5fam+D4bmcvuCC9/d9pxOWhIPOiKFwLnv
mxxCveFfATSfTZVypcyMC1WPtOIq7eoqjQpEdU/HWr93hEAzKAwj3IDjssp7785V
JcaO6ikhp0rs4IuWqlC6ETwH6PD2i3m7CyLFax+T0AX+mHCRSyrgOShIeEhyKRyy
5PiwgDS7OoyecSrjNogscFRujhvE0dhtyMyIt+jh29CN5tC2Zk2NnmDRKBJKIhqt
q9AII5pVe6leoIoaQruGnb6fwZqzbUXBeyJ9sVD+Dea+0XGXAGIgI8MysKACf53X
hd3yOBNcatHowHkTW5Cl5IrXdQXDX1iyWdEUmJUPQoI3XatFZ/I0T9/WBXyghd6r
5yqfkv0NGOMs4REy4jPQMIEQGjOzYNhJSKjvEy6xmSugpAFNTcm3JfaxkV1zH2TO
+zMJ8Xr37TLtFJz+5cCeENk9wXEVxFSAC0s2JaKIcKcB11RoxAn+wDvFMgmDiZ+O
qSUjLbDloKmF1GBKeDYJVlmt7+0w8E8nVi3/v/bbeeiu9Es1afbWIyHYsfFA2MIm
zWQsH8yCANaX361OTZgirgxuPc2uwl3Q/7kvAyQzRokcaRqw+1MFHWbDr9MUfZsq
V/fO3zs8XGUo1WNzSEgdkKtgh93e1qLApfw2FbYcn+5G++ZFWv46yde9mOUuAY0g
mV9Fjj7f+NG5zaxGEK7tsrBU1cfkZQAIoahr62D6LZVXANbbAAeS34V1WEFue4S/
LdpqSexsYK1B2gk5zMs/o7KTo7Sw1KjH3b0VFfIzTaonBqUEoAxqz4ZtSEGKz/nH
RgftRyh8zOkViSaEO9+w4V0Wo469+t9TAP2f+Zz3B/TBzCYEW573H3bTnjWvK8N2
lHrf10oJgJ08YI0VcPeINpX37zDQJPAqC7dWfMazUs4+fXudRdqV8q7vT1W+MyD+
d7rLLWPbpyE5vVaqhd3HaVTRSM/1us19t/rmroLipN0Pht+6HvH7dMZnbEC99gHi
4Ilt59JKdeUHkfM8N+WbyQres2ByXR1aatGa9fbXP17Tt6U6eolTHUnRp5FH6WgE
NOoPFEysJr71oxljcx6Z8p8kMBnydeudi0NgWVKcuqAJ4nB8ktTq6TWHakqz22h9
9xnfMh++aVsvBNi6f+nwsclfakQZ2J8QRn8xudA4LkTv2M5bbjCtfk8RF5g0iVHs
VYbCYj0n+RX+nfiLG88NXieKLXz8pcDZr07luubpL7elMqJ3xcpLtFx+IfX9oOjL
BU0H8+5RjpPpUcSNZVWm9FGzxV6lGwWuCRUSWHie1CI7YJSym3P9Daftk9aW4D+v
t2wXW6oqD/9IstouBL2/fCLUIdooZyiTtumW9Zoo22F5MQ8OgX54zkKiZ4fB7z3r
sat8S2nsbR1RstTyfFryA6iaDzbyoAmxYSui/nN1cdu6K39tnIgL1GZC2sRWIJ7y
hBXnBUEtDYxm1StnOJfqN0IIwT3quOD4V+MXbfmV8Drnh9CpUtU+BfnxMiIDN1Gh
2cF4UShAzqXijjPthKyxTMWRgURoLXgEwzGX03rpKZinVdG73Buxg+i90cWpSSUE
e1BI60AT+NxWzQnUttmSHWN/ARr287AbOuuc9SVmRJ0N+17e10Jcs/ojDXQf1Ij6
BNDsB5zptltKtim/PTE9yQAnvW/eLH4bfzTsNweUyQR8Gliu0MQzKwXUILjAPBaE
xtHFi0igYdiA8X4qFLQ8CSH82QQHxc6iik7Pc9TJOSjBccW88ExD90CAgzmjfeWr
6R25pp9TqSr1oyvNZqJ7MknKtK2xz66fETLpo+f46/7cx9YTOHM1eZj2m2j2pNYT
d+1fFtf4js433zZQMRbHf+oE+upS7y7yZVgAFFwQ93KBNHOLySrUHPEqXBSQiBRN
Xf7TE7CfZiUL6Dw+vtXPUcM/w5X/rDnUneATyVQ3zOOqQT3tAYe/g7f1T/gblFNg
sNEn2x+xyT4mtWaxYryJ0o9B7937gMb34H/xlKHS21zolQ3Y44xXtkW5qqh5QV1a
dS/rQMxAiYW4iX4cv7NAvq/AYX7lwnjaPRMj404lYORU3gY1Dvlxy6Obrxe88JZn
3sp3W9mbB3wuFUJmZnbarOGFXcGg+NO9Wxxr8+mwEcmtuk03GIlyk3+/9baI0ojN
XGIHFRn55Futvy9phewc0DVUyJtTQq8KZJGygn691FQbIVmlD+wMw6/NuTnMl//B
4KvX71xKw2g+cKZVooVNBHsZlSE+2j7SU+rgGEhm7ArrxpEsYF3Z4rBRqRR1k8tf
OAyIU3O7KO6FnJ6BHjvGk+Odox6/3k6tj6iXIxpN3OI2adcwBnHmhvHIJHEMRJ3C
meWCtn/Qp7z70lV+WuA438cx6Gef9Iaw5pa9Q5T/mQNprq3cRup8i1r2LJ7IfAQ1
NvuUMPtjJHCEPZpkOonOuPckKn33m1iLqbbQNxyuPxtEUPlIsEQLo2Or3xqBXNAP
mH7X3XYZivpIycYjbLdyvL383VP3Dqk9GnOLRXe237+XS1l7dosPRjcmf/iedM2Y
JN3dIjaGRz6Of2mIoGPXS0o6Aibt0sbwwJ/4cxoENnWCaGDFxwcJR9WocgY/r+vS
cUgxRdOwsX1WqxLZEbZBXQDs5W5Yr7mPBenWmzkDbJq8l49kKmK83Vyk2Lr9ND8N
iqYsZnKRbVW5fR5yUaWjSpdJzpWfr1WA9wC+yvEBejt0fA0rNEBYkdQDDRx026zh
p/D8u4SQP6p3Qvub9PDt+1PwR/LLDJQftoGWnvIysNnA1mrPxpfID4PQKL70HF8m
OaPcyoMhrkcPHfqGQJyAZar9PtVyzGGk38DVYCAGDvrtTrtIx0/rxIVXcg9ng4hp
AHFXHsU1W5hlQT25RBRK+uon6Eg69QAhpmGLyP3uxaNkZfpgS8OXbozg73IWOmj9
H8FhyZVGdxGEXWEH1brlZU+0aKKLi1tvTNTJMs4NHMRRVUM//KztblpeG4WdCxKQ
LGLhRNb+XuY9KOSxDbRg2tz2ZapiNMMe3U1tsj9Ly5D/FBY6NWO4Pd8OzSrulkS6
wPCpyWQnJZ/V7FZbZhG3S6na1U9a3eKNs+zrl4QevTmbKHe0xQt0uuMxyj8iYyE3
UmFJ+bmuozUqijYlaotPFSGGwMO/rxjTtDbxr9a2udGDaumqCbclfqKVQxBINZXu
XWy/q045eOVJyrRcCWJFcW0Ku1262UmTwy10rNaA3Zs6A9k0VXGZ0E8uEuMwumYo
wGlfeRguyfDfq0DIU76ZyKSvovnXaMSRE1Hpue/AU/VtlngeGHis5HqO4HBW6o7V
Ji9HeGqRvpFoh5WDkodhSykX/L5OMBf+vHKUh9rHxAeGwrnUpGfDjZSDZl9KsoFk
LyAL+jpibaPZUFoZCcAa4DgnPRNv0sNqmEx0NjZZ6YnkC6qAI9+gGflanVW6ycQZ
iBr//qzbsjyNHXbfyRsgaMMr1vCDea4oryvfSHGr+rVnQ66g3s91DoryGZPvc8cI
l1bKDKhp1g4L2Vmk5GgIJUPYZvSUmysYNcgMehpAiq3rrRqSBcOF/6fsnAlkLZHf
s8ws8LiMzRHC7utWcWHFlZOWxRUEuxHoB2hcKSSsTF+z8O+4rGrROTtPV1lGKFaN
zBNaxDrx9GpsTtcEorDEahwr+091JFgMb1rBfUrdWNu0jOgKjCPnxkU2SIAGWRO6
P6PvZZ395e9CwRvPGRJsUoa1ZSJaIfFNWjZ0QrhSgEXQxfiHUv4pWc2aOsyQdy/K
c6gkO0swkotcS45loxytwQ6UXVHxHKxFl0xPGn9gabpDRcq0CHYMj/dI1U5id9Gm
nmZDgnxGsR65lj7S7SYuV2m37wMGEH0ZZYDOTtzNbDkvRlQmdDUodDsE+pyTHC0P
IN0pLbBuv4CrvYquBD8pCvPa33rgpdrop2eljh2ORrCN6zlj5nFpU4LwC69OQ0bz
E9R3qiKiCnVxUURRJL+WFea9IlKEAqcQCrGIpWIycUYftL2bo1WhipQNOZjdry8h
Z1GhSyLixJs0BBMe+cQWqyRn15mcSdBBu8WagtKdpfZKap5R5nSpC/3qbS3vREgm
Po+pPvJ1DzuxNihPov0XNlL+WjlxYrQ9PTuhU9EcPfNGNc1Kzi8fYmv/GfelaclR
ybESr/8qh1lN5ORh34xD1rYCH9KrW5i8wy63LYtvyo4E7X4luEtCTYxt+emUVYgE
dCSqtEWDTdQe4fw/D5JoEmpcL92oIi/aXaD0sfi2wk4g+nYdm2gMaPRUU91Jb2lX
1/zfC8SiPKzz0e48wcnUbsWRFpZd+2jPTvnvnI0tFHszl0+q3W8eQ89ZrNYEK8x5
xnHi623Y+8YAojttkY8V/0Sw9G/5kxZl2zAfC7FhDX4AlZcil0jSjc76j9X/wuw/
hJLG1OyQ5YQPbGwKX3yJVEjrhoQlmCxSgX+ggJaR2VTSyKUy5yLQw8TwVaAIo/hr
vJrKAI8BllBt5Qln7lQqOeSF0jkrgSeh3oWEPBkh79f+eTUkeQTF0hLO7qzCjDlG
KdDEvU8oQSCsGXMfu1QeM4T3YXFj9aFFn2JOzeLWK9vAGCNXOqH9lIhAppX83OMP
vMVeOz0qZvINjFrWfR/gLhsUvh4E/M7v2b+ZPs/SnuicHtbe/rr8xMK/rMzUU2Ai
W/j2htEk1g3ios7DRkIx9vtfVWpJ5IHgp3lwvWBe78msYDTJ2CD0vjS8SYauIkY8
HfaIUstWmMFR0TDyp4+Sn/jaaKyceeVp5JzQlbiodivtWzz8oIRckYuzF0OezOEN
gdz1hYwJ7apU+CcZmsm3q5QaTvRVZEawByUJim2ASPhk4xD50SPm924BW6EJ+YZA
aH5PNNpwXE0vOAXaqnXrBMg95lCiJWaBTy6QZmZyqslAOvMgUKBf4U+COKIqqaDs
lJekRPL7P+JPPGli0oThvNZyLrxuWweqawaakYm3cB+a98EBZ9B/MmXTBqgt5L7C
OOLpKp8lQtp1T7JYHMAtbP5NRyxaCPcn2UrSArxui6YXMWitIhlmBhWffdhVWTig
TRl9lxyroEQbZ+yT3XPkc7l0gV5kvQCrOhD2fmzEnvt0+zE1TyGWJjvvu52T6guD
yoclL9R9P/TmVlihvLAGyo6aIfb1o5kK2VV3rgMLXN+BLg6tsWKjVYXeC93jGp1+
G+O1WGv1E93M1ip3GYmBHPJgYsiPHG1+6A4IXoAe2rx3tXkhwRaCB7FOwO2lacZt
JPu/lQuV5UHqluN1b13B8IceHTDnm03F3BqOPQ1gGfxrXM+pr0ytwAsyDQ4RdW/l
VEiiOgcJHrzqkUHLi0Jd3A30J1eAB3VGT8VhLyLSPaFUZj4tZYa2iQb3KyZkzYu7
9VSqdY4oHykNtx0h1QHfbd+KD8yWxgudJwOq79phLYpsGMsR9KLxXMqO8k0qI/Ef
iVM5Qnunk7npOl2ekObXpRPXcOkwm/6OwP8T64XFwA54NYP6+tcH0drP98iFs+Qx
54koKx1yvDf4HalqL8VjLRDrcZSACVp+FIcHzTQJOQdbYo3GZnPd4UQOkbElrTtH
h23aYLNE8jr814ljhWpN9nc5gr9/zRQ79fNUW8ekZoe35zaVcU9FNGKvtr2uyNER
s6u/dr3PvEts3c+G4/OV3d30GrE4nh1lsO3d80xKgoBCWykhGoxCUIXosPXVeIIH
m5ZttzXd00pAGJthbQ5WbqxjSJCIEAm5XtrI074qaP9/f8TyUWCT3M6LEcE5j3nY
lLSdyKrNFBbzIGE5YzijVP2LprUK9LU1U1XnTu471VUaO+EYIUCs/ot8yIwlq8Br
DdbDtmRbpnD6YpEGmvTOQrwBfL0xqmHI5XG4rrclC9wzHM7QhS3PlDP6GhQZzrfl
CK73wN/Uu+PBW5t+JGn0XYWgQOofrxPOTZKa4buEsN9ajdPvdEifNO/LFfZlcfG1
Ff2y4qWlGXZnN/I6BDcu2y9WEZqlMUtEumIp6VbYL7mN21QysZYq6jAMpXmMcGvu
q4ohm8Q1ct0YTBRKIfcUfclJb7TJM2szmnrOV7JDuVhBdLSz3YEOTF8gUOJAZybg
ZUvjyBknT4xRrdtRW/dI2j+PF4Naq9kpWqPVn2ate7P7ntvHnkYT3JqgwUHRJFYD
/+3R3QFJq+/ZrG+sZmvu4DpTHtzRYRQp502Dv6hOw0lxYHULxUmwUtUcDVaXljIt
KOHGKjLlsDk+o18MwvAFwEEpotEUkvyoByAtwIXB2KiEdMfuvXnM6jgmRtk0bypD
bRr2tg/BRm+DfnktF5oC7YtT/ck2C/Ltn3KJg/oXn+4JXebwEkv/bXLr0DEnbPdu
+N03vweLMUdob1tvr7pEbywn/xmZJyjaD0EbxphsYK2RrhiwFF5B0Ymj53jeZqIA
3e+hkk9UMYiun9tX7w5rOFFrZ0IONrmGaW6BKzTVlTpk9W0427oNNw6rQrYT+hlg
9DSjxn/foF9G6jP68PjMrbAqKMLJRz6zLD+kW88kBRsqKkC5fFywIjr0AsQrUkjQ
E2toBVADvr9CdhPTno/02SHle6tEB0GhiVVAu5IlkliEdbGj+qiUjXRBTmfhPKJe
ySIJ6kiJDD3yTeUrUSQB3XOSGNlwgFUUHhClwzM8klliERzLrMIAzDKC+FJXMwJ0
+4uiOvOFnMZ5Q3xNJg2jCM3ETF4HgvXKp3h/auZ6qDaWIsizDGpMrKAr0gr6FWRa
1p/PR/+/uN12t/ZILT6bcFSM4EOCixWyMAv/HREZf5YsHo68rNpW0+Y+a+VrI8bR
q2jV4q5m2KVsrw0hA9PY1rcwEVEr0N5RM2CuhbZqAWVKbankZhQJlwVraKvr5Qwk
uG+6t7pdpK7/GPf1agGUPF9jIe5r2DaDpYxJzqKlSgMyH8KuEnNHu/G61MxSKob/
FBHtt72Tbta7xxQ+wEW5rxWwyl5An25yprUg+t81Nx8/Gd6Qh8kkYsg/MJ/ya2ne
EpPpXG0EayvFYpqlD8XyP7u7n9pH5a6kFq6TRUdFaALZxI1ByQBOwW5FR7uLR/Yk
OaZe9yFAZjWq3p9cNgqVBjz/D2HoAun2QY19IXDvCiZUYWP7WaZRMgBkqmGfR9q1
O2cuYpq4sS7Y5wwVXAMLe7NDlHw1tPY62qiVKV5/sZQrpMvbD8Dcnh1+KvwDmfTj
vFkERZqCFTcjIQnCdc0MkM9iCQdIhLDjngU2CzitYWcn02c1c6NY7ChZd4YfmAGa
XsJHRSkOetCyxDX0GBjGqp1Ne8fqGrYw/MAZGF/7401/4oV73s8lJuay+xP9rhij
0AzqJHcT9dpjQfQXtV8QirapaDJxKDamuCWCzBDKpZNplZp6eXqfXFEb4MfREHFn
b57UEb5ImkyYOMa9mjqOiCwa3Mw9OvUFpHA9UgjLGQPA1hJIePKww+nwW5E7z3O0
0NhIUm4qil3elg6qjtYM8mnxoxKgKyIpSWVtX6SCcCDyP8CJFq5zjYC9sqe3JFcI
cl3O6vlweWcPt1uP3N07ndEhz9Y4SX2w5hkdadkagsMNxVQIJoH3AoAyBNW8Zkwa
ZSjRDy3AWrsdjRNPK5w9ZbgBxNHp9NVatmPAWWrCGmvmndTueOAeqXWtajrOIWsz
FuoqGIh7VbdZ5iJbhs2i4qIWxks9ebWsVc/lRI7cZjxCjFahyZnXNHpY2V3/ymRM
W8Brsh7uWR1wH8fU5ZKMSkFJKbSJjYiObTEedQAu1Ha2mEo+SsEnGt0rgvabeBaj
LTm4GcCMRK/8SdZj4Eg2hur8NN4PhLkv6qu7DEudkL8p/8YnangeOeHyI9vtesvp
cSzCsVQfWsaZZtoMaTkySc460DIsxFgwYkz9jAv4emQyjgYFW1zAdjGJmNr7eAtA
Doi3ygjvjkVk4yDFXJZXIoQSmHwkiCIyExqQ2Jf3Rxh6iKGDx//Am9xSn8S2B7qP
jlU5VybzvANtiSbsSOGOQ5eyFWeoK3lrzA1/VL8J9Xxe8nQ8flb2KJ+T3y91II37
yxO6Dr53x6PlSlT5fX8dbDrvOznXUJG/+C10v0c9YCMLWNG84TX1VutvDvm3Efw6
KaOZKHrsXlC3Ty3dIXP7t6aGbYNb866mapQElsPvv+81h3rXHrD1PxwtZAPf5pGX
0u8F7FxDCQ5t8cbuv+n3eOmB1GMQPDqHfwqFXD+zjuzr5DHR7SaVzCN9Vmw+L2e/
g/FE5yB8W/BzXnEQKPwe2k/eJRUL59fsgnWuV1SrWkxsiip5jiipN4soGC+OPu9z
nQjSSogHLWDvuXJcT5vrmwqtoZ6HXuWnXGdbGUcwgpWTF9v0HEhnDN26lV5K3njS
6n8uZEg2H1F3b/FxEYfQ9SmDV/hvYcJSfEz+s/4fid4YzTyHBsWszhduN4Ftdw8y
QdRq3lP/8vHOCuYg/cRv+M5oson8IShpXmiUzjfcUsdoC97HxY6Zbiuni2wRz8P+
PrFyd/1/TPAiy0WQHGFh61cPAipFnq2LOrIOr/zRLQK9tQzmicbxnTKe+N0OuA3+
im7aZHBk+aQuUJPnU43hdJxqfihR/Rl0wyvfATF7xs2MFPv6juGIxsYvFc7W+k0K
Ec0RPnaKrliv7nYmrOfhB3PnkL8Am1gG2sVK//x69Oz/Tl/UiHxJeVk5j89JvCFY
paeR8T/sojeV1h5GSM4quy0Vg2SXxS+de6grXCeHIKkllqYAlU6sJLvbhd8N5lk2
A5tdT9XYwYGF/MiKArvwZE3NVhaPgSWXMacJL7qsL2U3YPkry/lhrWGPOYEkmeKC
41cJ9M3G9TXcXhZhJrMGkmQePZPFVJQfnZLSxdo5MsM+0BTzRxrucouf8OJo0jRq
7kvXw/vAZqc94e4v69/ygJY35Q3K7/nDshH7G4Zc0iHS1mV7RXhIzeUZTzPBePIw
NHPhbvnsk4rQ5TbQfmYzO73leXrAaC0HzB8jcS0akTqMvNI0BF4NjvsIFi7wjowj
f7i+hnmr48PUuH/s1g/iIIM0oWDJ3TLIRrjRPA/T/V/OSM4qIUhNGepAA3F67ort
zD9QW7YB4PPOsyBvmIWEVkY167nHfky7nppMKwv9kWo1zMYOk6/HbYs1qPgGZdFE
WVFZ1ETgXqiKWSf133zAenwHV4LgVRcmNF2GdLQkQP/Qp10vz27o7/AMwAQ0mMkO
4x/csFd9ZN9YRkCTM+VxYWJtLmeDmWTl05EFyVAL918yiSTPIDJNn1905Z/tnvvi
DFUuc+73ajFxE7z+IoYuBCoezWUsnndaaKRvnnOQgLUVOQF4s4YjdbG8y7CC+GkU
zVUNMDzbCL7jmv5QDUqNp/bp/DipMfvvtc2wPm3++pILH5FBS1UdbhjUNilVvAfj
KJlIyzXcEGPIOUBN1qxeS7zKiEBs15aXox+QKxoWeWEq1VbAcs4Jb+MiQsoTCw0k
qlco3qZZ3jHP+SQrVl84aqCylxMLlDatphbB3Qwn/pVfCQDEUUSt5XlucGA4oe9A
AKqkjLdM8tNk3cssIYV4Zf0sfW5d+CATYKdnAI8fOHesIWfGZGFU2jOQvyUmb8dW
As+Px0doKi+JcW0gLTjNq9j1DRv3jAkfsZbQieV7gwmeahbnobYctdMhE2GiHJre
9EW6g4k7cb1S02y/z6c3hWUfupafGiFbTXx87BCUQkXV8sWobaKE+CMxCJCgOWuZ
Rq3pNwdSVwbc5hJlVxdcB7ye9Ya4uFWekktGCXJgur/sj5OJlTPfUrIdqPLC3cJv
q+Dem/Irsoe7mT+r3rvXk5sp4hvsXDkj2Rpq2mRHyc8vobD4V42apCDRQzUDi96n
AAJefO9wZZjkvEoEk5zYihHrW8DLFHeaR6FM4HqRzCRAbi1wdgj0AsRHMN63geB0
DAgLSgd/aIgTQq3nCuyhLlFD5FyP4oUrHBG6yKoZKQJUKY0U2B08A3T6dHwIVIJa
eXrUS9UxId2+8xNk7cjym3kBWbYDUWjKV9mVSz/JjbWXnKM1JH3Xsxxqfa4CDNPs
hIVvFwdSn4ZCGl5VkPgOfaP52WfToU5ySItXPZaND8f7SZn7/tU+N/oZHwtPynIX
4l7t9YqEXSLKSdy6goT+pDGHGjRq2aBk7ICFfU+ILJa23eeY7JlRDEUcHTfK1rHC
aEe/vQhGjgEmdPEsUQK20df2s3d9ookAubohbq/uU5KF0ba0d+By+C7IDECIMVgA
7RN+oeh9pYWacjHZhxPw1gg8rqtAqo8MBF7ITZOZ0PtcNXh3/QRHj6LY2HKu1RuN
cJglxzT8i6KMflRM0xn/LYp9WE/REObWhWumS3TfXc9bxMwrVdUJvKNbhCb3FgOs
gn4Va71edxMJcnI+6VCS6Xwq8AN5JpFEobazpHm1sSDS7Gvw/5Jgr/zg/5Mm96MM
NIs7GDAgVVjRjdvYg2ejqgBQUsahWkQecpxiMAQHNIQ/1inLG3si9QfQaQ28RMnR
H/mvhD6wY10dcOu6I3uEO8ufV4qNvUtIikuaLJXndtI8xPbpqUSChO9oayXqH1rL
YJU+W4310Skpml5Yu/P3wUkMLeQkdU7uMFH3lDBmoljIPBFbM9uFhYeWScfKmAhh
cm7pLOV95XSW5LywJl36JLOkV6Sh5nqdKq15koze3IvNgx0sEMPOQMhYy3C0sjmR
OTAKITj4m7nCFfJ4TVhKqqke/NzEQ1p1sLSjdFsYOPUJzaJt+BJuIaUgiFA4KYOd
+p7Fp586kwaQCgcKpWpOC9nBTc3yZYLF9Za70gSx+SNIoWUNjuvx5Ir0t0MQPni1
Gx2L4y0fM2TJx3fFP2S35Abj+mZOe0sq1bn0+etcgKhzi3pRH3E1s1h8zyNg2N/l
yDFbueIq+hdtvbLBfr/jYp3S4v3Op+NpctHZMalwsOgULTuE6HIoLJxXQ4lrLGe6
ckEiPxxIsHUPjBTKsJfHGxhBBv6l/+yNE7+/EgdN3LzTAi026CStnCT86uQiAXN5
KclGdcyK9GUVX71FTA3/JgqQ5JmHt8q0E5VvFwdUq2bi9siHl3O28Xne6LpF36qO
9qNxTGXXpVqV+u126S8Pn79tZIbT7/lX1T6EslQ5Pq/ykLjSuIhtGfZGVxxBPgtV
x4KN74lqBaz0VsOb2x2iwTuaYGdzY+w4vfvMcKVq2ncRu4droNJWz9dAQ7/CHa44
XwDXwYNWpekFrcaKUN5gMBZTHpqmISpEbe2xJJXL5EUWQ+z0LNn7Ao8pe/VETizO
F6fPB4DG2nXhFd4Tjq/WNsKJa1STos6a2C5rvnBhZ4sSuseoAOONnLCmj/MDLWJx
Vps0TtB6P5/4dmTiHTq615iPcDEGI7rgzngUiOc3e7HKAqmQGm6SOehCrXR/lY0z
ur1G3Cm3RN5wSG2KcouxOiYT2eyqPfKtPzkCDSzVtWBE1B2DP8l8Ca031S7FUUKy
RCruaj7/3XHBY+92qGWCQSSEWVfpApwctATvfIoO1YVOPlIWNTKXlZvCx9Vbn12v
osWo++HY1jNFYbMvj4qu/HM33jJzCUssBJKq7ijscPHRhZqOhGNDIV+ga/X5Eam6
jhhJz95AN54P9PDut9BRvOa1+aP1kPW4CmTf4xqXtdDYRNNTaGxm+HtQtapKgTys
bOaTIDCM9dGKQxGgxmIMjEe4DHYcAL2hBy7Mg+mQ10lB2JC4jtPROmPq4luyFR2b
TtIBy13LXB53ZoZIQL4yArikn9+ANAohPkYxmGMO6tZSGESSm6b6DqUjcyndtIak
/o7hScOjWLVy2wPOz2AHpWaZCRuRUKHdNbrIdgU0tn6AGiPKkwwT1q2eDXa0Gm+l
RZFsBuS4ekz7RO2Gq2oDuFVit0TuB9uVPAxsOMEhZ91T93ZiusMwcYtCuXz7xsog
7Hodx1qiya/0KRLZtx51QaFXV9n+WU3pZ5zwTKgCyNQ/Q5zNDaI6QIB7tevu4dFz
EXezaWjIG2xva/rhUKNT+63rXBoUOOSzmtlBrWlTor7TSrwvjEDg9UgYmohMvrff
hxOWpReDC3GgwQYa1HhQMld2pbUFFKsMH1nYc6FC+hZas7DTDJyavI7c87Z3Zi0s
o015WxrhS1+ZC8CR7lng8IP+MtPahfDEy80jOA15aCXdNC3TmMbr9jeOTQjIhcIk
uEVLb0cbcLfo+4MBYMKWdnF5wD3dq8pXAMiVZpzXIrlG+WoTEL+xVv4TaoWx52p8
8PxCy1CRq840aWQjC7UJScDrlksqT2vPphEk8qPoerrb1taFAqLxbkl3uUuxTPE7
kMVgVFcNxBOOB0g34ITug93sKnQqmCm+GHcWD//p4kIS8eXBPqjT9TDaZkIkWwdf
CkZIWZ+nC7NCfurr/ys904OB1Yv95gy4PsHVF5wKZEWFrjd+bKi2lbCKJyso/6RX
+cIgHpfDsYcX2j7mfcE0UHFAokr5CPhKdsENbnHZXORaNbxLTfmV2ajcL8GL35GT
Y/lVStxFFcNssvVvhf92vPrtROVSkxxzU25etAjEgMawMrgQbbqF4Y/m2LV215+4
xZALWNXjYYNYSEisUA/nD5JMOUBfDD8JrAsDZuEvT07fBARHYzQAnRzwdJeNJD4c
7YL4HP8DLkNd/5qumbmXEZNy8tE3i0hYZPBNtSlLF4JlWHyd5lF2gXKytQm1k/sq
ZyYLKMdV4CFFfCJ6MYwdv8obSq+G3S9DnSspcleZOztlo+DKv5S17BGRWzSat8v6
7FVh2ouUAsPN+TagW1Lmpjew64a7g9OvN22Vs2QMzGrqci8I2p4iTbXfQFYnTUdw
RhitSCihqmRJcpy2nVUUv0aj3gaytIoalmPBAXQ81bKAUyAV5INwqxNbX5E30PH9
0wg4oOGtBzO5Qrsld4wlVymVK8Y1HDnoAJGqrm3SBRc9yyr943RE7Jo+ycMLENef
X6cavTkVck9VxYgiF6G+AUobROqiCPqkxSdbFBnvOjZlwMsFuuAVyT1VjxNCxJ9q
VAnHzGcT5db85Ri/bPe0ASu6v3MkbJL/i734vzA34SSffOE0y6NhOh32jJVThtiP
+gnDIF1WS7nbSfHkCT2bpOxQ1KU8yURQh4B1RoSBhlHYvLScNlfqxNPuauUn1p15
7nn/KFMhok7PTXhwxIF4/uUqFQ6ePKlnma3wxPmpwWSSyfmPpqYbFK8DJAzipAWA
nnIdhXk3LwhAfcg+mJKXnzyMsgHzOrwklp7TrVS8L1DxnKQeD0O/9hQc8tE/G2+z
J+imT9H/IZwW16yg3kI8zqohDiOiT9uAXOFLiUF7c5Tp0eRn02uHATEhmDyyf2OX
m0+1dLTb5TF+o7fRsDPVAVKgWUMH2sCYUkWaPDw33T7gjgxTv8hGLbBy+BwQm6qH
dKTT1oIwpv9f/5sRTD8F9+6wu2RS4CsotZOVdh8+whzA7499oTpnVCovqGdhLRPb
uQgirPtZ3hz1QrYPV4FhdmdovUN+pNWU/qf+JiLlj5yKMqIQ4dzfJUcc7Xg8l5dl
yt0bamcOq4mm8zkgZ6xsmX4DudNUwFL62MKqFUivI9eAkWeHnxFCcjf1aMslk/cc
7UdoTk6FqbBonSzTRjjs83uhOwj1KxFCGp3tPBfqf8n+ZRxo4a4WwiuHlihGmrHt
hh22RhcTYYH4rrXI2qKkR0Soj+fT8IQorUdI733LQa92CJaYpo9J7MlDotKdwsMc
F0ZhCrB3feCuzT9g/oF9TusA0n6PAQIE8tMBM1jS+WmE1qZVNZTWLe/uM48/yJvL
zUsTAqw4JO9BZfdn8Op6eT8jOxj8F7yQ3XzwsbAPNYSohFOKTwcbKcnrLMppUKRY
ScdEHD2jvwmjlCLO1DnlhJVr5YnWkWSXiwrXNYJVNYvrdTZgnQ1jJBiCLKr2OWRK
uTaec9TSVUXlAAyDKwvEBFcu//Ejk1egmEhAhIH4mbX/f130C92jrt+wtsm6QJ8r
f8aZIJuqZzVZAZME1OkQ/qyW3+iR39RlWsDwBk6+vQVbcH7kJG0+UNKvoGHeLMzy
PYd87fR5NLG921a1UTsgW7bV342oIrojUlWMGrxL0rmF7OWTZdRgGlL6Qw179wX7
weWSRalQYITE20MjpuOaYtLYJmFVEsPHPSmcuz9WQDUXQLQ4w1tkaTBr6lc8G6vh
HWkN18Mu94TQ8E4brr13sxUHlCJTKy22Ugezu4K/GHuNq1qSYeycGtqqO6vIQ53j
NcI+Ba7Fv+63lkvdd2zoUKOOZmwXeXXme6/wYq7chM7XuEXBWuJ9z8GfvziGjjzS
lnSd9AqAo7iYFn8rU2Gt9ZbkDISluPSAwVP95eYAbNnXPFLn+HHDPidbZuDV7dXe
BmaSmLlRF1GXd7hcgBFTgSVgVZgLw5NYkSL3ceefEHRGPYf7H0EYoDlbtZsBvYyZ
DM966eYL5cBQYNvBeUZ2X+f3sQ2/2NN8i3cOlZXpnyv4v6F2dmgcIQjBh0yPa6UB
GX/p5qtDivU8QkV/R/9XVq+R08IYEOTOFyJ1qDQtpxbcPT9TR4wvAtnMpLChK6hE
QSwgn66mbgPYRQKDrTts1gc5YsyERNjz1ko9lJ8PKk66W4K0HW9OVDNaxJsiLkmE
fimS4NH5+dBLqWRqzI7v3pTOI9LhcDBK8oGLNTR2KXqMu2wsVvm1k4jnBrxHuovi
kuwS0bBbUEF60jpglX3MJ3wNnzIkmzhBMOB+4aoFuB3DUTgN/0c0kePiaJBgl6qF
qGhV/8hQ9onHmni058aOlmRKFW31lF/rBDiVufNr3rJlb+LN8vfaEIpphjIbUpjK
Qs1fXNOGRTWRD1TBIzeB9rHOazmffvEFxlN3k+5n6BEVcnpz3/5heqWb6ILrtNSn
y/Ic2YAPeS+Wm5ByqppAfshb16PZ9MqYkV1PyxqDauRZphFd8Ndd5vzBu2iFt/t3
ROOpsRx/QRp1/muBwneh+EQRKGnmux/a/9G4XVRrF0ou8wwZcMRGi8TJEXXUVqzA
UPt7AXpJOzpCl74/tbmfl+KcUyRMdEls+nVqB3Pa9pIY1o/azLKIiAcRV4NldAOL
TRfGM0zd4j84n7ib0zeqt4AHRzFbtShjALYrINGd7fKwWVMitF80o+k2B6az0oia
yli/aI4reXOZ3DOrwfNe70Sk+VQH+1jGLw45SJvQjrDkFSDoTdazruPu+oe+tnQZ
2vHa20a2Pqr8aO0vBYcg4Cz6NQA/ZPpIoWwdwkmVJpkjOWMtDf0ul1UxHsKu8S8o
K5Tk9gzDIKh7jgz8t9EjGG9kXqBSTtqDHLAlPLRT8eL4+CZFG3uAL2KbRqpUpfHk
Q8iu5iLRjM+Ej0b/DxRXMEynBN9NYhCJ8lQgVv2DaYke/zP/VK2ZvsOnNjHLfMXl
q6GwrTCutZAhmyiZy2w7Jjb3zpWG7ycFeQKEgbwuK1I5fbBKnI5wQT1JOtIdB3Ac
MmCPwxCpIuHHB4GbzbcGpoiVxD59CI0uE0D4zVhgnOKHqg0KzSg0LSsMKEJOf7do
jaQ8sO5hyy6JHIXGj2aFi0GBEP25kouwFdvQbg1AbB5XAAHpSiYkaNqMjaQvCNxp
B8Xg579Dsq0gRFupAGnJx/uYZ5CwOyvZQBUsIF5z50H6i3YSGiAfNx2hDNKHtU7r
0mz/xNS4cHzc193ilqvUyQKaX2xWywtpfuAzLqYaQ0XUFZ51KlHGTTCkCHzDDv4W
Qoll72JXpn8m0X7SWFRhA6Lgx5s7P3Nwl5B0OtD6qiux3CFdPdjuwSDS9wQxDYKp
UIJt0i2Bp0iUnvw3sLOROGJ8f0s/7OyCY27+OBjvqU1Y9wdjIyq50+kl86aKg62R
yT6WBiM578ixcu+n2VFaYEuoC502hRIJJFcClvgX6f74tUkDT5FeVxrIMeh4cdPK
tBAWcVDW6lVZ6pxnQKcttzo4edT20/uz2dHptuTZB1ZaOv/qxy2dUso23qocDQtP
TVAGT3rfWDeEgNRYmM+OL1cofUiSkkyp+k1bmPbiFvAMLJ9ZqdWlaR/ZVFWTGOEa
jffFep0aZXxqTkDOyiJKzVbWaIT4ZjCIs9e4xMjfDkVoSQDsdy9FTdLYdgqqiiVd
2oROWGu1SScOxHTXvPfwbn/gXHRmcaPfyxv9+ccZWgW5dB8Z1gZLUJPactgIIZie
3jc76Er02R+WMwRWbzOrPwe5qJzXGbQZuHnRvixQdiUcBGJEdpVQW3BHgZrMba1b
/PUUR/2SmdLxlk7Xv4M/qhDVMesm+ID9YFAOwvw2ws+/8sTKO02MurDSN63IEFvD
8+651lq0cWl67uxfl3zgghnUmT0YLObr4o3IV7+7565erodKHA+3w4Yd6plF7/DP
QuQO/izGe+nIf6vxoUrjCpsTRIq2c/gCpULF0bd7DCiPsp61TqTF2l9oQLACACXC
kN3cxnLP4Ks4T6xVeFgZUOZXOBZxBlR0L1UQ6sciz0AOqhf2qnVn+T0FOu/IGFUI
o8A//hSl1KMkaktYry33uETKLuBvB3Yl0rnW9WBpEvd2b7DAxEC2fPGGI4T1ErsZ
yA+cu+fGVkwUJ+5jwJQy9JfAdx7w5ft8ItELpU6iFsXOQDqRYMnPf/jrMknXGhRD
PukmUgvPOuqhh8xl7fMy3feLdF/jxb9BeRYhJRDMgl0NQyfQxWclYKUl3NOCgM3P
cCMpR9Kx18k9/rjUnirrb1YEPYmQFIyS9Hih9xV/2Gf3j0oHTuLTIKZEsB+Bg+Ap
yoJfrNsFdDQXhB5mNPMkY/gTRR3tjU9Eiadnvnp7ip+U+AxCkD+2NiMvnN4V61/G
uAp29IPxTDxkIy+1IO09WrXTJ4Rh4YK4XPE4cSECbnqeWw8yHwKWUfBGMeh4QDfM
3JyfRaOuhgjqYdtM6yhZEsXgGgnwmg8xLYXvKwh52Vf32o5Q7PJjdO86ADo6DDUs
15j9jtaM6/0hMuU6EQZRlNpU/irZrNRH+KM5TcmVMo+zb619gE3pBWYooLvCn6tI
FVFImAqNsaYtyVbfQ45lW309WaxA7ZhmkfUzfGhwC0ozsgURQAkG4jmZZ0Kj9ObR
znz46imGBUCgm1TJWWnZea22UiQT2sSY6sIzBFUFsvAcus2BaZIByO3qSUB6c6E6
mrHgHDkbf7IUoVO7k4e7xdMlfelQjtX28D7q8ApcB5wVYN4DnvQ7YJrU0NsOGI2e
Emy+KS7p6kPYnPo7yxArj8kMY0lTUOn0j7xgJRV71//x90f4CcHLEn0jBiwuwSKY
MdwQ9PUMFIwDTRsERzlfRRUpD4+kjdIsejlN8RTiiA53dslMBDMCbxobUuvVjMsc
NWXHIoPqgr20DmhFnaqq8/RvXQf50NGBmOCvdHr8aBuxGcZHEgzmn4EfWKLbsSOa
8IvsB3zO2Y5uWBDpYyBZlZz+xh0yn1Ci5WPHzWP1ngfSXIzkdgpRH2P9MvGnjIBS
r8pV3KZKnuZR9aeit+lqQ/NleEtAOhasfRzchnzCNn1cjxIomQvIu5bJ1ybMHtTV
bB8BRWYcTrijfw67+6aoPdZK7Y1wb31qEq9sHifrYIccagm7uPyRy7awcGhehNg9
UKaw9h0MV6ViLCrkRFYJdQFbkzhGUGisfWGl38/XYK6m/2oE4ZSyWnpFXs6kRGId
UFIrerPR7X5oEFYl1v5Qa4ND3nZCzQ97UyK6sCQJiT3xQuQIsNlHbcNkooo0ncP1
uqQk6RLEWQFHhJ89R26mQtccD2Wgo2/RLlco9xp1NhOvxsTRUq5L+5nhQV07EK8F
aKP7fZizCRYlY707El746t8CoWAPHrFcajRscwlq2/ad9ORpSPKbYXLhOymKcoaf
0gUw0I/Fo5hOt3n4gdi8dhhzJukgexbS5nI3wpyCKyMhZbq97FFrlf5t3RrgAT2W
O/qnrrnfsS4/aEm1Yv5yEGXv6FvDRamUglvWQIiJcc4nDSYzkfMVbN5wIdlHXtr1
9mjsWU6TZITkyG4rWh8s92Zd/2YY/ZV8Um2eZU6H3/e7yOyA5TkTXQ8H17sIaYtH
gMrlQLZbuRu7NgEXsHKgIF5UHGGWsZW/ByzpqyUs/eY+90JnMi1Cli4Z49zeKjsI
AoHAe+Gz1zvGUimxzrRRijvlRvZKu5qDz6Ow7eHxGuIhUOvCk/28FUoKFDeD5FZ5
Y1K5a76DDK37qOGd2SOeWlOaBNvRXdhgH2XFBd3dN2ktxJb74kWPvajlZ9GBpQx1
Uk9CbA8pbflXHxArKmBdBuJuNw+dRSSlVvJvPzLcimlkoCoGVEMbTL3Q9bsB9KDD
Ce/YMWx4SVQxzTKWh/Xr3DNOtRRAV7AEIgafwZ+HG17k5/FUQaxax9Njb+jKE00W
yt6HKZ5puTnutx45n7e0pNUMnXvbIctC9uvG92fdQYJTik3VoMnNMNqseA2jJC5w
eGX1SiT1hzrrmeJKxtM5afkAiQrOicxNm4ZYcEazbiOLkrJ3hqTlC08LsnF+g/l4
f6W2Fvq/yIhAoi6rr0ayvjngInKxNrSybXCMten7dGk+MQDvQV/iALgEaWHvUQxX
VZsfjhRhkpr4LvPhDVRl8GTyeFtYS83tOKWs/e/cCid2Ah66p5aq+cebb/q/mcOE
YYJG2AhsRCtc5XT2LxIEYI3Zh0o2R2inksLFiehm3EohTuwZiwi6JEOvEoa50l/i
5cqJFciXkEwtYrpZGHQQKEkd27Op/sbzxmtN1KyYmnDl91qWY6KJQ51eC6+assJX
fDgqwE8fimW+cu1QPUOTRNV+sGreUENZB0KlRJUstR+4pIZlam5856N65OGuBrOw
F3BKZYAKlmNKiQStPKH680ra9UQz/pXuto+Po8pkUdfhjT/HI1OXZVNMqF84TcWz
4Kx3bzk5aeKIi+eBpxkrAwGxd2YFiXEgEYX+zKCVkonGaPJJ+ZaNVQXwXnsHR+tE
mHJgmhlTsAxwmD4Tzon54EFCDGfhP6OTKnU4mSeX+ZBy8hbAJ32HYICaJaRNAdqB
Y8/NeysZ2i1WexTR4H2F2EWSgmY0Y5HO49K6AGgQbJ5REJZH+4LyHcTXG4iAS0nC
pllBkzLMAZz9CG5Nkx499aJpQbNza7/qsy8S+wi81f1D78FeeJXjgwk9M4qGmjpS
0A92+xuG7MNLi2D5nB9uZwpmCX5LwQD7NTCRV5FnHTKEHdpvCrqUTCD+AhYIxerc
P4aDqxnwwgAj3Bn6B78b0onfeOhz82hagvHRBVfJch5n9q8bBAil8v2OjzDlkax6
0Hdu8w8eA67Rh/R25lcNKa9NzxZGCvrZFhyScI9MSWVxIlDirmABsYprYwKQiGg2
wHDL51eVHWJA6CV3Z3jKs56sHOrp4wae2KiNwZxOXmW0bZkb8AFnexJdb2e/Dz3X
TLtOwGTkkVutHbQKkja7w7LPIxplP5ocYWsDRi5eYthyW8D5DzRjuDg/JO8VDkZw
rHexhxKehs4omYUaHC9ss9KAZpfA21PTViqA6vgoX1i3Tje/3vIdyv59R3e8XoNO
iV37M/ibDLXa2b3LJyDSn9W9nxRk+H5PQwcoFWNr7K8Ysy4UrgEXbRoPHh6csEMM
hnXZumxeSMsIm55kokTRXCN7ouveJbLaipPt3AUWMogxoEZTC+zsx3pNFG613sys
mbmtmDptkRto5McSD0TB3qbq9jIbil4CrJF9orPNEhah7ZvDQ4ZTQ/hoITYkZ+kZ
5EB0U9fBNslkgHqCCJDgCwc/wayLZ+QoTQIf5W0uedBd/D6c0blri5KdWWqCBEKA
hzqg+0t7tTpqCuW/egjrtpPq/5iTNfP1a713O3/P/jj3ASZbZQO2tpYMdVPfssK9
wcaNQ2IG8IeObxv7pBpivXqPYYtqM20CQwDqVCGJE0BcnE8wFEN220qfYP+qwxkJ
YTcqtIpQfk4JiTUMcptd2ycFT2Y3FndHdiPfl9yv+ht/L6860ZfKtR8bC2Xk1b4y
o67AT5BTvKmvtc4EvxF9N4WiESNzIm25q1QEIvDXkUONYDJcAaJ/LQiYIrWzywul
vJLTWT03NGjjbw0FrQo/moUCIYujkvf1jKDUF3drXLASOZMLlPNYEiwT/QNo8Y5a
0pz1OeZuYhNKefgljgFT5kPEKNdo48rgzHtPOdf0/I4Yo4yAjV1GVA+3P+DB3/MW
Gf/Yx7JqqXQXsCfpn/P7xAa3RxzAuTx+C0bRek2kN3LdiY4FMDmgzdXKRK2Ems9Y
xETSfQDInsLH4fSe2vVx/ZoFos1Lf3UOvm2uMdZwm8wgu4vb+TcjsfK9vwIv6rpj
i/r8pb6YwKqcNl7x4PVKvvxthwALhGm8O9gX1cn6uTSVQMaTLuPk0uFMwtdXB0V0
ox65cIz6JMyVON2H37p4q+d/ssjLsfjXhihBIdKz/D/Klq3aDJH3yO83tC4gDsxv
n43nrMuR1pP9xE4b4AQawkgKEmn0JbE33HnkXkpsDVPAdh1iIYNJyYoH+9fR//Xc
xMVTWxSyTGxTpaQhcd5vX58/jTW9LeE/3vvToCg04NhDQD8p7vpcG7yAL7emjEec
eBR5Zfg5L6pKz4Y5e6Ec4iZWuAgBX0aNri1VimXFow0KUnrwfWbl/Z2iT0TEWeN5
SB+3IFlpl5lGGFmK9ow7rkXwDIYFosp9A7D73/KzzqLr31SqlfhZEnNPqPzUnYH1
Z+emqQf3EkZDelwjJBFLLXqSpisXVkQgD6HwHsYA/NueozXMnSzaS0kthT6EdE39
JMLBBmakmnxUnXrJ7HLh1ex/c1SQZCfx2Q+xZvOdJY9+/ieSCHUFTRohfBG56toK
O0Tgy4SY8bV4A4SdIb8yv92R1Gz6oGIgi7B07aFeH9BIv/zqytdPGn2sBZchXmy8
p4rbLEbqlELusfEOrrwKpfe48p5LY1Yd2UqYO3JMVggaBkmBBRCHjBsFBTt1vm+C
opsWqF9RRHX+ZwLpeEIF6LQ0RBApYaNh9Ee5e9bocPU/7NtLwNczu8APKL+YQvhY
kY4wlFgdSJlSAH+dkIXM5Th4SKAtBYRDwIpTEpdnB6J18Mdk/z6U5KBKFqg2+s34
HnLliyBSEiUHteEiLh49Sajm3/wldAcgBuRo9qzEGOyITwN/b17OkDwmIlHfVPFF
MPlVRSfMCIDQ62XD6g0k41VFXdCCYHoBZll5NWWswgt0XorndzcjOMwXcbMflfDx
tQ26dUy7///I5Rk/vx1EDfchQJfv092aYOR1GxBKIyrT6j5gWEcvIyfISxD6rWmj
4Bdtae+tC1mYKKhFh/oLO/LQaOSqMTpivVkCUeiphKNbneKQ2/bISma2OLS3bM3b
Sv4wr7tpWAiFK5Sp6OqHKAUbzoDCAyoODKAWtqVLnU6nvtkRjYnchm5oRvbq1O6V
+wjvf5/OSFAugjwi6pssnMggYiWn7BU3kVCuP0ppZl5P7xk+qcJ5zU/bthA43F4q
WponyM/0bNaqJPpse+KeelyCmDKWDKIoigaeQJ4W3LhaSEMuAMjOF9taVqhzpHB/
CbJLhjQKN6WiEuOfemj3wFDcGsj3GWvfKh6sppxS1G4z+keEFAsbgtvZHThTIQlY
aEHO8yrCcYf1Mzh2Tkq/IvJMw1WQHUy8EpWKAmpICIJs3ymEnpBHal7pwA/1fwjC
1gH9fhgU2baW1wL1Ysfe1xUvXpfZqyAZGq9c5lxkF9JP/UQuQ5pXr6ePHvMbqYTH
xJBoj4qoHvpnX71l/P5dsmjI6dkitjTg4nzJBYdX8nvMJFGhJa2OOLY4FdwA6zNG
Alvmb8WpRy4D27M3druC0AI78ZOkm6lFQpt8cT+UgFWgFo+FQ6PzTamA3b+9D8gJ
uarAFLnv9BDoOyXDldhO1x8DdX4iAxj3RnJRwOjWsitEHTZnCnw+z1PfMzKFjar1
ru+kGmCqQlCNScsNfikOkor/9YhH8gq8gIX0uYJIom2DBW6EIxKp5r3BQaHPAXDB
xfxRDtFvtbP6uiZQ8cMNXO5Su7MD/Ds8BTYe/ZnK0CG2katXf3ZlCjG6YHICgPze
W2ojU9bc4jfyK9FR7UKKcCmpfuzKJarS9rdKkUsfT0Yf03/q9nYLLdqFM4Qtpxe3
/Hr5g1zZT2AzzmOe/btI+rGkbqpVXroNfoPa3ajACEQT17BvEtyqync3MjVz7ZDN
UvYoHP3tZtqyGxPKWHrBmQQG6Nkz0z9VgR6hW1a68iIHeL8qdsMe1ljIUtACl3Rp
2uJtBxizEpO+X+DuJhQMRTwVHur8PAqRIHe3b89jMQIO/I53OZeHbSqyAnOD9wjf
dC+pfyfzKvVZq3yXC/5qmj3yhX7t3RFVlDcL2cdV7/nqsA00Xcl1f4432BUvgN/O
c29JZxCWrp86r/xlXsAT8z2KMN+TW6eJG0I8ish2g/p4DD78bO5zVt3eEnYfHF7A
tKfKuv7v8/fo/Wdbt50GaMhP1CmBwj1NwNE76Ga7xy2/BWhTj97Pd9D+DENlovvX
HyLr6lDtiQ2Yg9JGTEZMgWQEis+Ho11uwF6F7UBuT33jBNis9NeWz34GgZyKUrP6
uumLKs/g/8KTHJHLuswhIdGIjaS8/G+/MDwOVlN4YL7iHoG8XR//As5Y43a+ARBA
VGhqcXn0z4vkj5N6V2d+z4taWQU634oTWzRPJ/tYe0J50DWgVbOx1RBr41w7+5VP
bSvHuEmcjPj893qD8ElZfLmXEgW4/sTmnjQfAeaDz2gxFUTO8+NvlNiayE5+UGt7
KeNFAjeevql+RBoCZU3n/ISWdpei0pE2HGpuC/lUsmFSFvRhsHoLzTBpuJBWn7Td
E4rz52X2MR2zKid+6cjxCIZENOegwgMjEYD7+Udj6vzRke6S/vbPuYXyPMLIPxkz
F1fQKLKy+Lan6nTnCay9xrCXAHmmZbJfHyCgMnIQiGQka1Idx1iTMNsq2NFq2sJ5
Qr8vP76xEyE1kwHu5lrJSyjk09OfDVIEePLvbjOs5wY/HN8ISnZVHiX4W1I21SlS
G288qni3UGjRkZByjRCSiyHJGThzjSzlfMWXIRuFPUg1S7eVwrn5yLwu8fosl1Jt
j/gmkvmK+XCVnhEraPHQQ46qxtb7PiRLa8yp+Rj3HhuknD/nE3KwUdOzsVNi3wJA
Akq4omh83gLezirZotLxYl6gnEtsL3cEGbC6/X57d6vaOftoZgSUrmMc51cK3/TT
CQl6bpW3ZBI2bOTM3gejVgx5stz2CRPQJaIk1c3s0dNhIIhjbuXbS8EG2+UNVl2P
2wA4LzlKL7ml/ZPMkxWBnrWNa2qS2y8ddVB80XcZ3fyfOQwM4u9DBQXVea5xN7Vj
v12MuHF25CIT+c6pEK6bCBPYqgantYFsD8UWseCj6mar+AQk1kHLGfQzodERFJUh
bKYFt34vkSHhutsWDbnitK8p8nK0X8+5xGFEcouz6Df9DD/ScA2DJU54Hcc3Nj2w
Hjuzqs2Trh9HOYxkRURxfjPVDH3hz7WobqLS+R0aVdl9rzuVvwOnK0+/CaUKAIqU
uVqWScZrd16bhd4Y9KqDs1xWlML8uaff99LvxlVyhNDEYxIXieqXjEnX5wKUeQIp
HieQbSQST4cwt68LVwoMrVKSxcYpKzZNfuU3UmFri7CRfrqnk5f5fVSYgoMHbdMr
9UjM2DxaQaOw7ggm885tcNSdRrL1xSUi7gHJIZjeuHAcNgEhCvvL90MRgPj5igZl
ZTLPNTPKtBG385pmolQ2ADC8ZzlHr7ycn2aE/UtIS3lBy6bO31n3l0SoPQ9yHqXi
iG0WtUt4/A1HuKUVGsD0Q9GnoT9LRmTwmFYYtKalsRfVEC6DqlwaAkW+JaXkH+2n
Y3vqxAyafPzGMryuhFGUhW24gW+MKTs+P0mTPhIPoSevZ6r2fDOKWCXftcaZ84oR
bjjlTbkt9tK5giy2DIpQkCrn0aiBlONb9+ok3OpvwiJIIy+AsJXkGCPR49DLtTjc
Emrt8iPXGMRB5NewL5BxXto1+9kRGgkqXPIkoBImtlWucCqo8vLsssIxfrcqPo4+
D2yrp7uKQtkHGONJ3XLy5AB8QFpqQH20m+BC1GsADMpbfW2/t1ohSdl+QKRlVgY1
Mg1yo7o0+M95KDqXLm9ckbs/LnQj4G4t9FYhx+ObV2xemZMS6lY04IsULqEtZ5R0
zcmFma7kBZQDpopPU5u6cnh/PNEK4ZXPQR01DbOV1YaAC9YthH58lqsGwOWiYLMI
rlf2gLwkoiuh5K4klZfIGhnKRmAU9ix3efDdFOslsI950PGo0MA/NZ+CsKEKxmDo
6J6+xzQXq4ovf0qSf7gCZngCkiOSHWm5SiO/u3ls2gBmNKwXV8tnqy7+YHgQe9ee
1n5XWGPM8F2LFvRqB4vg0DJCfR98ZZp6YqmzANYpJJM5htgCv0kCGqou63BQlh2C
bdygVF1yvQesCqALEc9Yh8ow4Vrw/dZ9brfRDp4ceNYRwn+l4u1l6RABlS5DAE1v
AB0vm48OURy+4RNF0gOdZY1cQsCUFI+N+BHX6iDvmEbsVj5Lgci+vkYGB3amVhSp
CJy4IqbiIo49IV0IfNA3GnzUjQdnGsL3uvPHm0KRHiG2I1yDSWNT/gVMwK0rZeD9
RnWLYWaKBo5I4ZSYQCwPSnrSOMm2uj7mKyxwjO/Hs1NY2/UrHojWcOwVTBkwgOHj
3xtd+P3rC2r5mAEhWQMBNpVnvqzWOVAK3ymcjl03CQx+K+j0aels1ncWhcwhBngU
yyvtmPx2cYSxUTihpE8E1kNRcZWadPpQPEsP/lm1P+FBrB3POljQTKB4mwhFi/bL
pDzRvGgdWLghxjzM8znNJcYa/+DFlUvWsQ26I1ehKhcviVAdL0cz/K0S64xWw3ki
3NSTaTsSttE1W/a6w4KKXMT/1wMlHwN3/w+BVT5DS9SaPwCQDIQGs88ifY7eynah
ltnfz77O3eWuMTSm4Nr4BSmbYeFEQtiPelLzQl/is8J9E9JZM7O62rBMrH6MQ+NF
j2t+zZJO3GwfMXu/k+i2Y2AafD2g1y3wyD22zlAuDQHRmK1w7IuAs7U3IOCa8JBi
bIWNgJQHpTEWMTOrMBRdBjET7wD93cTc34IN2ird5UJJY17IAxHkwU495nxaWJDX
7H5nqaDF9sW0wwg5ZsFvOKoEGCb06qXFHlBCPh8SkRJiqT8tKnBzRjehnyyLrfrD
jN7qcOUztqXoGbtw6MyFvHNt/tlp0goFyVxZjBCFXqaRcJCEFFsH+dr9oAqMC2fx
O9qJ+5/tiU+E3cVRDHN8obN5Zjs9XUNtvv22qFEgV8sGwZbN4JaOLyYRV0CyrGE5
vPlr85eekfuynlTzfy8soRuCqkS2kWxkziUvTbyyQxHxCHVqJ6AP4tQ92xakNB0Y
smi/LuTPX8Vo0t9Di5CdFRu7tMQFiBocG8AKL7roIA2GBcHSLYmxW2zlU0VEZxPb
YHmsTS7G8FURBxvw2LHz1QAy8tWMyebtn1U9OGkRLFeGOXLE3pj6aZ6LViFFGpkm
xJBhgMmhA/F58TMsYU4VA5GcFM5dI3InIZa/+4JNyinoi/g+OA6nkmpBJiozJ5W3
198D12frY3SM6oTJYJ9Ijzslw3+6pER20FXwbpmE8nwnoFH9q1GYCXUryz6ifENo
Iuj6wTTvG+UvyhaMA4A9NARPUEKewDyuJN5Y3ATXd1MeNLfQ3EMv6XsEsQBUWUQh
aCUIBAbD/F99/297sqzrfHbdl1+YhApYcgygyEdYKSDuRrSJewIqIvshg1tw3R3S
6X8vnKjfaiWbno27OH8h8rsAqF2FEA7BATM9OIqpaU9ZKhvj2L1BURmhv+r3pl7Y
tm9snrCLFnNDZ/+k+kZK5/7MbRFArTaLEu7T9s8XHl4xQFrfUXHbzxuigRma4V/Z
krCUwkMKTbMWW2a+3fVd8H67ZjGeVzQs5tkFz8rH6t7rUe/aX+qDRrt4SZT1HBFA
GAXIMPOpSirA8DU5aovByPtGWzC+/BDkVauNm7PjHT7b2KCm+KoIy58MIrd48y4s
Gx8HHLEiHk26pCGCW7FaCmkQ71KaXik3HlHQz51Lr8ylfdK2NszraN0IAOD6CmEV
1mSJSixS3KR9wA5a4Vk/KY+i5gimlC/yOnNvh+e7er2Fr/p85SOoDHYwdNMMDV0t
wxUCnbyqquMUvYzKTrbzPqOHuhMZpazigZM0SsNr5m6SgOXNLyjAhYzA+b8Niepp
+afx+7/8cqhNlo3sb7v5YI6EleebjHas5qOIG7SzBnVh94vf86zChTENFMEo9bse
MNi/M311QqG43gI0Hx2DH7dpznCkU1KnCk8jkk0cUvYeN++mRKI5ES3SuqzpFxLn
4DlNq6voMyuKwne1UbdRn/j3q7qJWzvQKXCdf+VTd4ZzDRTEPi8j6RzYkRFUXatV
PnX0xiRJISd5gxPCYTr1DOeUUQn/KSAmA42B03PdDXqk9XBANhPXD9o1hkO2CRET
XVkXf8nVTaPxPy47FM7aJwxlwKNMe+Jszmv/zGd7bPe/9vEdwMQfb1rSow9TjVsd
2tVQzQwbkQOP5r1GRPERdJmPbmzIRyYk1iGWSVdO/ZrpqKeYq2uFE+9bWgWYgoMg
kQL8AQzj4nzPXGzEBv1r9fhGBNhdCZ4KwgpkzPV+ob9QodhxX5UG6jbohrLhe12p
uuyOvdsGgic62kBBlftodRc0W6h5cFpewbDnmjEY7Wb3kJKdAfdDzOiYls0N0Efn
U7/uow1JXnNtnbn5d0KalYkRoFYrqsNcmi6QRqEbfCK/GQsGL4pmPqDrsgnO4lDW
zP2DXUNs3UfrCgkgM76d4JAdVZXy6AHz8kkzqjeN5qzp2YFWwWTkpx0niZJYdrdr
4362dYtDP0IBR2hnXbLr7KJujHFB0EdT06KI4grSYAgDbGK7sMwyRyuDHZQT31/G
fB4N0wBzI0nD1vdXctmCeYKk5AG4cL8Fwir2cllot6fjefMS+ah0PYIWl6v/R8EE
u2yHaD4IDTl3JJ82+vbA//nGWP/FYcAAy7jt37SFKDBvUfoNtpc/ZvVzs+gcmZNi
gGHkmfvev/QtFT4CfoQPK2b+qKrT+OrX60dJXVxg3MCL5Vf9FKTc55NRMnQlUs/M
4Wuef0HyG57soabfARhsiIXb3vz0bHRpKfTnlVLavxPhGY/EAJuxSIZGoxp8ISnF
Z5ZwO7FgDwmjbm/tEir9VOk4d4KDyWBLAoyq2FSfl0aST2IeyEI5dSXrCsjMAAQO
isnJ2DeQJJZUTkHJkEzizPWmVZymOSO7AvTonz0yuHe1sj3EkVajwcPvhEi/HAPi
pdcq106qZCB9d9FzzBpdcSJH+uR1FTKfRc7vdgkwqwV0HZ8IWJsrDtOD+UEy3pdn
hfEuoPyPItRGBlev3PiXecR8y+LY33LZRk8ijbP0oMkGZq8QKeT2+/0ROFH6k5QF
BeayxtUFoipRY5fyqyVWdCTlAyE7vu/31cn1K6prbTCOkUySr3ESDRA/1vHq1DGE
1KrW8AqxpxCKrVGCr6FXWCpAp2x+uLzmiZwhqO+ZUB+7eFvPbQD/RQBSNz5tvZLM
FoLkGi8IMyaUOMk8CyrKB0f9mDl7EXQs91xFfP7d52pZKH7374NUSKpAYBbkEpiU
Sl60QKDO6Z65mt5M2EfOPFasaYw0asvsvBrhJ2pl26VxMpZaDHUtgnhVTyHKGIW3
bP9pj9U+KqlEmbThBedP9r4wCS1oKehHnV84KqUBK2oKKrodnMRFUU+/bh0PDlNp
rLAtVjktHfMspEiMPolVtlqoddieoEFwZmXGqA0wSAJ9zZmEuepgnD8oX02nPi//
J62mU2bazjXoRpiwXXk0L0pJurHIINnZvZXtnQg+bpSswoNYeEcgdhjoHCjLDw5G
VbyJ/eRJD8Rz7Q29Tl4ATfo5kNvRN8f8nKL1Ww7c3mXyAAhxxRr7nOVDFOlPSHtu
fvOg24mtPkOl1+mtrZHnNurc1STagMnIVSGHRKdxUAYoUHDtrb/ApEBYTrMTIOHN
r2hkqIvVJXZhvYVZ1q+35En4uPL8fzEIfYykG3tGtaA9fdI+6vJP2cDnY6k34of+
I8r4BYExhHmWYqFHDdpwBr+WXx30O0Jt8uX6DQ/JsVUBp+b3ugyOsYxXGQSD/Hql
/FMTL1B+f3XARh7PoCNeNdetjUchEZagEhIJTN+SGt6sRL71FCWrDw5pHeW0ANOD
lvLCgMN9ovFxqNbhM7T7KJax/vSOD3dcbPRv8zSCEbWKa0QClDb7nTWM+VYdjCer
ienOZLVE2zTctSQzOvE9TaIH9jhR6sMvnIBOQcmrdVD5mel/8c+vatGpXwgeTxKv
jSsdXZKoEo1MwzkotksEu0R/lqq3UcChb+fkEtQKHrkhy9BuuBxaXiuO9k7o9mCM
b2xK4FQlQnUFWw9UamJbaWp9HXgOMwTC9qOUEMWAd+AQ1jfWZXaDoL/BhRqlpSnW
bAeSbfOd7/aDDfJ+5jKihPReuP0BdKEAT6ts5B6j57kh0Yd7tTPl38joQJLYBRfz
89SZi/TGLOvSaWqXfaaunUmvaZaDgMC8ghpFBaBoSfNF89KrehisY9RtXSMWamnH
4qLFZIME78uNf8fgE1m2zfobf9SmWVsSNhheoHG86E3zBaXu1nyNbJHp5T2cF9aq
Qf8K95luxB54BzLPZtl69cKAmbiwh/uimmnxECZdQ4DCv6hzsWpRP0qi914+VubR
VD+N/AWbLZHsgctwMw6wt2A/PvP3NVX0pWwkAVAuQpgKY6BAZCP0SS0jtp4zCXz/
HecTOeaxEOMg1yuftLCHfZnu/bTUpBG+sxGjgL72VGgggV6EJh0KTts8p5WBCcLc
4z6kwBbj/JXfbWOxao+oolDbaYSmMR8QRyoUvbhet3YXN03tIjzJd13uzOEhY0uV
lEcAq8NQy20Zg6hp36V/P8xyPch4gVWH+AwPEj1jlww2B5b81TFEs+TcJcInVTXH
sFEon/Y9FzaT45XIbjzELCIRtTzrvOgGF2QxGvhuQckdRg9atYYomjb3sgIXMgtv
sKQhrt+AWxDFSGaOR/r5n3HUqw+wXLxt2/L/n1pPY+RQ48poIiXVqTVAN7kGx09y
8dixJDiCx6iDx60jK3M6I/kjMOzyaVKTV5rYPHlIs1FRtlhd5QaqSm3HOaats6BA
D38xUSwHYm+rXPeDghSV02qRkoEnOvJgC+Y2dYDXe4iGlTFv0rJSUh2eNieLUmLT
VHDRJPuqWXy9k0QfPZOKG7JLiYybUFNZOz33/lUL//QTOUufjuODF7+IcB72NCyL
I6nS1quHQppxeT7zqpeUwOzS6fTGZm84nIga45KssjlofeNG0XcfHLAG1T9p2H77
4iOZwGmFkWzJpdKLM5ib2061n4Mk2aGEmeG/wspneASUVbxS5BO4+2M1KSZjnnwy
22KemA5KflVDL7bH7FaEk8CpxV62ceymMPuuDGzejA7mqTWXHIjN3RkfX4wL4Z4L
r/3j67HvuTaNgUt/66Z0n1gPW56GDmAqCeQJG2875l26Kbqll4X9gBnLFWxPCZY0
n4wE29S62fDlrNyrT76hjt9lPTzSeNJ8WwaMagfD+wjUms/ncCU4mS53nqciQnfO
TVmB1QdNrG6VmLOdZdFT6AnJ8iIWIL29ve+BvdNDrU+9womBFIBBsQMyEPQObZvD
qotzARddHrXetPHu6YWQ0lqEkWbFnluqoOR/vgZhW924xFSo/ZVTZgVZPCC1R+Z5
ESWC7m+4lo9oanM+P/kdyR+mUlM2cK21Is9G2TWs/d0TNTFTdandoRGnBO9cgTqU
3YihlRyE3hYj2Ju6S+oXZQvs2GOHqM/N1sSkAw1O7bC7dcQzA6BsM5pShLq6auZJ
PuSQz1/8IqQzFXiPt+MeY5LozvioYS+Jh00rXKy7/3NezgyjrZ60TbETxwc6h9kz
WNNDHeYScK+vuw0AsyXVHZOwfq6a6zrf1Ys3StdL+zoAroYCoVE8u318UKdJA1UE
Djg+a+zf3cSDgqOvpCHdch72zu0neor10QvnmFgCQbaqJLwTpSx4PZFaP3NKA/us
6XtoYBqBBTQHkV7V9NPaoJz7kV4YD7B/o4HwrKJtyNEHEFG99TrbLvooNTks8LTw
CdruuE44UqhLWED3CUK7MrQtReD29a4M0ATBT2neA95MrTPfIvs7090JfNsC0yIZ
227+ZL+OPBzhJJVMJM2H3ml+t/PfOFlUNImBPLlGlK8Rg468JhoWXsOTaWr/B+u8
4BDOjXbg/0TCbwwoCTSr3QKXSoekfqVBl7ABdrRMSBXeS9GojkxnEDSbbKby3ige
ejZHFb4uns+X26HnSuI9J2d97IHvmIIHcBtc3RVNPdIT31bjxJ+HSVt+c1OR3N87
nWBIIP4C4ZGpyHcsSP39XIHXR9cdBhrxQiqczNR4MtXKptQEuSSuw2nUQFKqziO0
xyBOdX4r9uN2OZ77ifpwqz6SfUIlGkH8Y+LZhJ57HTAioTxcE+Yc2AQuCFAWRw2c
xk+XZYYM9n+QIZIHh3iuSX7jWqUrEUK3EUevWgyrr0nQlG2nbDKzyGozovzac3i4
PkrlEUvOHusFNj5YDcw+N9Qz/AOIdK+PqP44ie867sFNt19eAJX0JIYbz5g0fHVi
J2ThYv/3YGigEso8gbRPWVx8pzXMYTZgHa/Kd7MVnBpgsZnf4BR06lUZelKI9qxl
EY94v6mdB7oXmRbfULzNOuGWs5zbo55nGqLgOi4AGS3JzNe2qD1kWw7E4ccRn6uv
DEXa15VDS+ZMzJolxNAp311XXaQwSQNJuGYWIEwDFIQP8nTFsqkMh9IlscXuTyFm
7z7vcSa4ivoDJuy8NBkckrj5NrsBHS7OoFQ0yBQ2bSDkPOjTiyq1ViMVppajwaE0
SNsya2zCcL218hSqP4RZTwiC+yplttEgMFTt2m/8rlx4xuaQWKHydGZm+wjyAqFQ
fyO5PJ7bi68XnFqhDzZGsPpLy7ai6/yTCNBGFVoImRHe5z7N3zKlJH2zJp2ntnBt
W2zoaXhjElGZKTCCd9Cl/HJmocl0Vq3y8Uo9lQVkxEKHxPsdoub4PUJpbv/JOJbK
xs3stMflglh7xsE2CqJ70aKUsPRChf8wKkyOca+xDN7a7UAvA2Tc1p3eJRyXP6QS
yb1OU3EZyk/X8L7dnaU/u5Ox5zHGbxMg0b3wcb5Yc/xBlyZZMYrZCFm0tk+kcPNa
7G1RsJHmjuzzzQ47qPUP9GMNlDMAl/c+nfzvogKcjzHykyHw40gEr6kI/bczYs/d
xIGRSpbuRfuvwMEsc841oRIWC8XnjypEI7CGB8M/2PtAq5DsIZ4RbyUx69Q1rrPt
p1nIhCcP0rAqd5A4nqFL2JSflUSu4fVvVk0NKU9RUu1Fjyxq/n3b46cFgrmo+ty2
xPgJuqks/5iHOdcGQXbvZcyB+5NTdwbQ+cbuF8DnwsDpiby26Ondl55vNuq15Bg2
Y4idBWCYa4IapE7nL7HYAlsubw4bS+t9Z6W3OalWs7vEsN3zSb/DPVWI89c6R/ov
Uxzxs/pQ8P0QbyKxAkZH5aT5HVLpZVe8s7ON8gPcAn3ZEuE10QNQ7qlAiXe2yGEF
HK8azdQS4j3BJDiAyE/0cvJeMKE1mVBqD17SVZDfNX1nyXbgU+HNYoesd5XW4MCm
+IEEbQVAuLX2aNkVgwLOMOBtab1Yk5q0QroQYKhgero4xOsls7do27CijrHj5MH8
RK5BWj6uEbr/DkieWbFPSF+7ZiLKfWEJIE7A1FObX3ff15E3PBttkaYdPGigtJJW
s8KI8SCxMNhckv98otS+1dB+Bho5qPPF4BiGA4Y1gIFaRT2xp8cfRbocFY9ZpS+d
hrvvPVHkqzeTVO8MT+3TV1EPSo87ydX6GXDbX2XSTmWWRL96eEdD3nPSScAia0Ps
rFBAaCdS4R9409DbjNBUQ+z6ukJE+jdAOCCfNdtQm3WMz3koNuedk0A2FFoOEAKA
gQKZNqqYUd9g2ZOecUUS7F0MZgTftWzyCX/NVCoUHxhR/Xl7wbwbzEizySApAqNM
d5jP3vs4f8JreHZNA3IaiJbVQtMrOW8nvBauwsyslrm5WjgRLGrRuvnYQkwulPXR
6fWyUtgITbIs0E5PoyhRlJ74bLz5/s0Wir9X/kriq/UM2MYjbB+eNsHQZ8I9aKdr
e38FQWyaHauby2gAV5d5LLSY4J67kSBJdCCCwswUKIkZo1GSD70/AUlAKLSCqhrO
yvw0tFVmqORA/QWZ7UEBQa1DeT66df2R/3y4Ko1yfaDXyXQuKojB7i+YqKJCxW8D
Awe+ZVsef3BqtckJJUKvFMmHWxkNGeT5jnqWGljXau9Rd4USrgS7j6chdT96IbSz
qAprUW0SNAvIvQO4YAc9kYOSDeTaeASXdiS/TVfor2xGiEdp+z5rn9cSgD76x+Fp
kPo8xryeVPcKigK5GJq1n7nol1X204Lg8yZdVUdJyo9SiCjwY2M13v9ZcESI3qX+
gYw5XQoEXBXD+YFA2mci7jtL1GuE95ykt1SIs2jQapJZWOAOiYHT/uy5SxKaMKYY
PqeQ1+UMkZqCWMth33CqYhvXykXh9HWb0t4R2Ni2SGGt0hGrgKOkL8s46ZsXKHjP
/e0A+mfTTNML73k4sOJWxkJqd1CARJoPMe2VtADKiXIQX5kFNa6VMi2J955FMvWN
OhtFFhUJEk5doiHaf2T6sV6+pxfamlmwYDDzXEHWwuJU1Dm+tpWcuh5zQlNqcF8b
oU8til8+bPdip5bnbm1EyJ0HlzyM/JSGZ3tLId+Zg0lbmSurKlqStbCtHR+B/nRa
L9qYE6L2J5ByELOlNaEtOFCl8jnj1kgnbmR+3GFOiF08ugPeY63g4x9cqmsais7X
gfPCbjWTemnd0qEeAXyRTrQ3pBcPef7qtwOmGvBpvkkZ3Nos8sPp+7jRo/nz/lXs
KJYITVXwTvWkgjyPJCmlVrj8/a2KDhjnTK1LnT9jTSLwOkdqrY604nolAsn9cKXA
wRB8pBMaABHrAskoDIjPt2CxGTMYTsvsaJCm8E9ggmyzCYy79q59Fs9lgwjBRElf
EHWCu801vhaSOPimp/o6fOXX+zTXAvvmkjbyxqJLoe0+SiE8ZLZ5ihwRyvjVH8hG
lnb6IjhAZp7F9TOIifGetb9R1l69+EgwjP7oJWEY8Br3VlAW1IVy4W4NkzM+U28E
telMGgSFvLdqq4lVLYNiRGI2P2W75sQg0uGfdK5CR2h4m5j76NAuiwXhQpEfy/xG
hafFVVJQr7G7vhErpFpJ9IEnDhC+vmVkKX+YYDd7vwmsTWU+iIJGPS9gNdqbl6OI
fYdXTuUoBltc31JsMUpVpjXD7pKsMcdFaTK1yGbcCYmvz9N0o4o7ToNf5oS2dIqD
8Q+km+NWXXb/xxVFbn8cS5eHYpMyrYV6onhD6MtH/CJ+39flRMfld0+Zgm028P3X
Egm5gZ27O3ZM0Pn/j4niJX0IIk1wdxIO1d1RuJrb0sBzbj9Hh4z58C0v1BZnB9v7
IdSnbiDoKfM2uPeZhPxc0XxIO9QOP5R2wPVC6HuPVBll+UsKkyBqLZ/GiEH+u5Tc
2LLOOx1LA3I5fxnhQAwBAZbCFkdmwpxQgLb4iFU880V+R7kToF+i6CZKTk+W2r9U
uuNa07Vaa4pJNLZMMKsAMaTLA/4guiB0+ZSHWr8zeyibSvRfjx0l2axLYtp/BP5e
ozEuvdogKhrcUEDyw9jQ26nECWJnfRm7RMeh+v6QjncRKjIGMofuzYv90vBiKiyI
3xHMvjr+4vCbHHHeuJVsaY7JWfzw9oXVrl4VIAm26M/BKQpG/bQuFxkRjXMuzBIc
7xX3P7Cf7ec7E/3VF9CGpYgNkGa8z5hU4wbZVGCuXDK7LxTcmST2MFvUZq6SKhav
GbqG376CVLMvNMLRxvTc1etkUSfrTbVo4PLMXxnvfuozk8mAbgVEw++5n5lzwi3f
RDdjN4YSeCl+dNNUV+HlVdHQckQ9ZyI5f/AqmfGrbedRQmQgX5x36iqugIFQZSzu
Y4ZJ9WxMFJWnYAk++p3Vn0N0m50A6p+DAhcLMxPmdz38My4kYC/hUaiLwqV+BrhE
8y/nh2KepyMAy28fsK/bo3Ued0rUp/Cz4c8Fe+sPP+4MmtJWZXk8gcRUAgkO6AIt
J/TEzA0nFcQee+0soHIR3nFjyz7X6TtoYEdW2gEbAR1MuOKoFeNi06KFN2uOAvXs
mov00TNZa2D8VDSCXreBMDR4FlNXijoGy0e6p57lDcOkGxeGZvPvsLIrznir/D8w
5NmgDWFqUFrvNIG9s7Uv0VbC5hPH5CxY+m9otup3VRu1R7fKYzVwF2bnzZo/nNxD
Vo0JrINVtTq9BfUGKhOorNNLO7TcMpKb1tjh51uP5E0obwJfyzsRB+x3/4UHmrAu
v5NlNba/X52W0qJP9XSqdhDu2+dnSgCX9kDoaEIMXzIGSsHTxnqLURnEfmBP8mq+
OhEWTeAUxigpNhQTlHofkZlSJRSqBSvxzsY3AyWs2CFmexy9KW5tCzjCrtNOmZFT
b3LqARyWP6NLt3K8i1201a7K4o41QOkC3mEfIDEom4b0Ead/LPLMoBKnNzwzg1h9
5MAqSIoZWCzSxjL/lYBrZzuDq+MHbV0hOkwfyjBy28OzFcPO4TApgdGaTS9WadQ2
a6o1xnokZPlPn1r6UxSXOtBVzG5XImYm8CTAYzK1PwNbXaJVhTv3efv3eW0PuJHF
SbHrWCnogAwoys4h5/SB5KnrUDKFa/MoUUf272/Inggi4kNeLlhof2edUHk1Mvv4
XJNBv5ifvtlRz8PaMYpsdw1hoHAWbMDSC5mGc2CeMllqpJPdvUwR5YanIP0lYVmV
rcIfMFPQNbHlyDW6tO1GBqypoj/j5Vv9JTjlOrPFzWah9kTo4AWJR118oDgYZFor
1a5j13pk6Mgm7/hXZV9S7dyXDrrGOvOtwccW4tFZ7p14iLDUh+iTjEv6UOj82lHc
ddsuaEIKh1oBLnvKVOVkBjuzXKU4zS6bfp1RENfsE/x7VSIFiW63Lc9iG7ijXlzm
yYGG2Q/hqBK9yMNeHFOawuD/TGXMSEqZwQmaI5FXrWQb8X42AUoJ9QtYf7H8UebL
NnmtrvcLfIt+FEsC6rX8t+ANrxBncTbv7RZfKLvbQ5sIQaHCTCN93xnrStjavZWX
zf8u9rBsu3+kf1iA5TUvyiLUuwhaZNVoUQ9X+xkiiI1uiMHae4AANu/M83zbxsqb
62l+beRduaziIakAHu+Ooz7t53cHhVTKpRaVCf1NG15ORHH/jRVvTsZdzQxfxwoj
WnyKe3HL9zsUKsTr2ODhgdc7J3sXPk22XvhNWJiTYWo05U4wsL53jgJfWmHdEpoS
oAp+gCHYuuwX7+/zawN2rKKSBL7iDXNMAFhlOFya6e6FnU3uuQcOmFfD0uf/iBkP
x+xlp+sNtUKLegv78cLYXi/Ve1G6UgY23jiSBCsY+9vr3svseqlSUPQ42bugX1FC
WKebjFaR8e/62YLDFG6tbQ4MxN0UbaHwycfxb8RnlarymKX6xLNbGE5FUXuCpXUT
XdCcpe/3vsFiwBn1aK8I6vuGVC84w6+tmJt8GS3qooGJL6QqMRKJlhve7imAdvCj
QUyS2238P6qxLaKGzPPBuIiHaIaLq0LJwzsLdgUIcw+j/d20NHgiD/i1ld9Xpdk7
GCu5kFrzPtRDhJ/xdwsuwm6Tb8Ju3ijxUx0l7hmjIdi1j8VAB/TeuMIGPqytDLVh
ubGOWy5nm6eocdh2jO5D2WyG17jywrGqotlmrSh68/qqT9MPVDNDAZtJYErUd/be
+dqWcsuAMLx7W6oMeIF0V4C3wTLsgf92e6duEKTQDgq0jBqAnRZIyF+qcKhLjwCD
9WsCNaT8vjWHBucwb1RTXKP3vRYFckiAK0VhPoRgTARg2+d0phVzEx44FUx5avkP
xxSuBezljuOEuFstoEvCimIWTwU7oJeIMlFhFIYiLRjbnG+DT45K2bfoX61Pblob
d3hLV8tP/cDdWdLD4W6HgWWgHL4Dky8nZopwNcPTIYDLJKZCt/Ftgcarg7ZqlAQX
9u7OZTGnZU3nyuRXtlVZmbzpRnXfNUMTFVi4zG5guyNyDsEzbbJnEMPpKT9/8rwd
S9MU6WHR+bjvEOm8k0wzb00PsZgzsVEvwjXWZOZkuB5F2I9ya+htJPSDYRA18Af6
MO9Qqd2wN0wnt+q2YMXuqGpDm9mMHiGNi1ZbPKTMC7BLPLTzM0SwEVSZexdQPFJK
ZNUuPaU+qVz9SGMaFiUCsFLL54SugKZgqXavxmQ7+0kYsPtCwo8G12VTzcfZ0+J8
7TX8KayKDQE7Zos1+E1V/BjdZG7zhg7EgOWOeOBMBRrXdvBDFpqhLZ8aS2Ig02tH
RdlcTfAv6eNOVLk5ZK0v7VwHHjDSC4wOed+at3qbY12Spg9B0+cgZhHqtKJFnD0l
DhgqoDmoFRn8CrouOn9PswPDsfrW6Y8PenjCt/jJ9Ee6cA/Ci8x9xjPmZ9FojWOO
3INNsP48o70BMQbFWx5MOKozASo1IVz2eSrNDikCuTYUUVJqBjGxTRe+9PeSpk+u
EpbPrHyPCUjD0eweN2FiCen1ZLCt7phT31S8tv5bJdx0hFTqE2W1WGl98nE3/56j
ShXyxcqp2slH0TUJVTVGngFDRcR/GPvQvf4wK9qEVfGwTc0B+7h4fxVnpoBedDRO
z5Y3UUojSnRJfZXXPK2qAuv+iwLnA+f3PNExjub++PybBKmH8xmOauDeYEONm9zi
YAJraGK02tSwUk5fyFKRoHFisNKcNVmgyb13nM9A314Acc9zp1P4PAKY0hMM8g5b
utlqjL626JFVIq36tf8cP//gR7tPem+BkGc6NSdGkg4jPjkaHayuW8BIDvpUkI9t
k2EshjrB5ry2jk+V8b/gOJ0ZGSQ8NG1tTPsoKkQi0VUIGPmuxhEwF4Qjs792N/7g
FWeVLca6QeNmOCkZRgMGMsnlYRSeGZEvwstlZdytf53PLbtbiASB/ugoy0tFwjju
9rtWc602BnYjR61+AMFyhVL1AdnCNJ7dVvm1nXA8Eqh3T8OtObZmLSD1Rr7+zsUL
+RUoMtRPcHLg21fbfbQN2YUZpNgmnufzcBjBLXbmDl3KXZSvxtsRsDmhLuGkwd6O
MRsiEXrQJvjaLEjTI5vSgE5wc2NapyilJNlybfHoB33X9EaYskv7K/xE+H4vlzSp
Ewt6rzXkuXrGQnN4YXL6KF/6Jtbu3Mk/1x+8JeV8Bu1vlpZrp15OxgWeNOcYU1PA
xVQ4u5NOZzjMfJlFsHsEUxfMJX7N6942H+b3siQVXSJYpXXX6k6Vky7B41lKfYuu
K3otnZNSnoKPrL7iTkiSr6XKLJJ+jdxR+TB6N+oZFvo8Ict93FIKcn+pZe04TL67
7+7M8j26BeS3KHRLRFKnc8XTX4Bqyvz1GxeerKaoKg8EHLftl5oaGmA+dGTK19Xk
+72NjukSW6A7HymGwxv+xXqh0cOUr2rop6IqXIjKds85+DLshzsxSllDzC6fzSVt
swnnDQEeNWKxJqcjr9AXtZ43KA8wOQJMHy8zAiVLrpdMzjsGEoJkT/Fynxoo9qYN
sHEHLJYsunFzBWrdIMvUcwmkN4mrWIev/TDH+8vITHzoGazWYYK87Xq8mAkDDoBR
8sgNXca3cE6/B+Im/YQU2NaQ5BzvGLKwrN0R+8eIz+r/pW3aASgG8+J1neYNIGZn
t/TY2eNz3KNwhoq/9VQhanxuB7df5qCmjaa+T9bgu6q4N19piYMpIa/fnuKzmvNA
gtPfU0TVmf1UPaR1AOrOADUWnkCJZL7qtUxgngVYgKgMtPfpMqntXHdVlFfEVEPU
B4DKz8SE6eLHPizP1JMmlWcsurewDwUtKDY72nW+Th4bE6CpCL65ef76ZIolgWyO
CJcK+W9NHXUhXLjeJ2jwrs+FzvMzXBpJB/5BvyLKaz88mN7kXrUJqHrnbCs/RnY5
7IIM2SitBlI2/3EE9mDvvBcd2fCEno2GdXs7/mOCkrfx36IvqY9/UzU5hYA05WAL
nbz4JyATkd5g3oG+l2njF1VIJTchWvhPZh2PIXgL5MT5ENQzYIQIgDwZFqGnFkQu
O4fqXLfQGQxo4CdtPHEecI/rUAKvKtDMK/l1guz/e9xx4JO9B8mK3WKvxTJsFlUI
MHCiyJbCyazZtKFKr48ThVgOVX1t5etrGN1vuKEgI5yhmg38NAVW5bpnNqh2qHdz
eUBHB42MuujlcLJFafzSS2TVPOY/CfsmKjYfMJG8HfUfTP7tzXh2f4RmN9ykx13F
I5BTwxyJOO6IuSnWFpnhuJlAtsPMMAfD2OXulr5G3q/ZWUK2YZ+7rrne6a7z1mkp
zpOk6uMDNspaSAWxTq+YPylbzX6/kAzwiUQ+ut1JxZZCDF681r+YMNRWQ66cWey4
rxLH5Id/aX+IoUL5vQMB/u8VjUyj/+sY61MWbK39Z+kNDcZ8sfB6zr9MEDqCgyIw
SJ3POSqiG7Vr2rN6dlqeDE3xuYkJlbCUnJRiB/IahEZFgi6BqpCMaWnWZbH0BBvG
enkjbaZYBP7my2K996bIfbV7mzoEXt9zGHBx6MzCs/FPvB1mkAUC5x3b5ms6cJ5+
cYEl8gv6kig2a3gPkDEWycgqDKdl6sm0r23R/aey99TOj/6rmVMonpk8Qsqr6Ik9
CWTP0TMaF5dOz0h2NY18Sx/glHD/mMTDpD5z0Sx7GM0Tb2IN1/YJ0VJJUiJN2OoD
heKcmTM2AQzfPXFZGSrSiuuB4qz+tMuOo+fr+DjDyd0FQs7MZmKrPIMp7fFG1xGr
xIMfaG0bxm3orK1aaNLqs8J6L7Ehu7aGjmPghscw3Ae8pbWGnMbQDVFCwcFkrF7J
KMIyA2kaUfWO1c2jhX0v2ThNPc2PR8EM5Fo8i/3yg5Lk2rj5iZ9ACb6Vi0JMCeEr
fyE5umPkdn4MRQowmCjyGFEIZPNg2ZO2zZtWSFCwJ8egUq4Ge52rYqjvdEeBKois
tIUcQxtAF0IvMTYeO/AU/+OOM7Ed5Rs9O5yFfzI73HoZDsnOpxUZnEOaYKSxkNjM
8gL7K1MGizTiwrxY7jD71aVbU8lQ4I2GS3zClJXYGHaKuvzoqQv3/D6fSy6BhehQ
7Dp829j6P4q9la0M/yFhGwTbaE5hkUB6akAuYzNmffz6un4OIHBhLuKqraUeehpW
iHX03UNa0CuJVQy1ozVf54CMzyjyLuC04OIAIMcgmf+k+l8aTrFyi5psCI9lkT6q
d+jCB5z+GLLP71lkSXRCfAceFE+ENllUS+IHbQggoslj1Q8KerNf1rXUmNeUT5Wi
fih2tyM+8FkS3lLxjGnoMEt93S0du7pDDznxqeHiRXF1eeNP9OCrkeADqtNcWKPQ
WMYgV2ro5WxhQ8yMc67eZNeEYJJjS2mpI81Xl1RORQveWVwA/A8zPrVzFRc46+1s
RsAuw6f3zun42Vt0W6+u+MM+1IyoXVPlZziuMicEIzpmg0nqAIeSLOzSiPhrMasf
l9XW4IDoiKt8zQaZNU0gwgKc0nH04R8MfbyaprVhxfXJpPfGgCCo9N+87Mm9sIz/
Bt4q94C4vuan9NZSsihNcp+59zytbuOvXHpOlxtGgLM1+I9mNg1cLWpYIF9x2Wqg
s+L3LORsp+LxEgSi8vNs3BuxnmHG83BZf44k+Q9YOKT+TyLISZN+bsVISQkS/J/Y
FgXyAHKRqlKHSgiABeHLMT0O8JCCuBNyH27gZr62zLGGSjhre2efc6Wtqd+V4aBE
yLZ9uTE6jPwAcpLzYPYqt0ROMHbveA33AXB+K9Luc5HSO/X/9/QBUYrbrIIP6Dlq
2qG0nVAObylyEJXKRvscR4Pl2NsC68hMUrsGW7EUHSp8zzHBMNjUdoe6dZvbldG4
KF1oi+EaysaQLNClxFmOled4byZU6Um0LLp/rjeZFXHYlyBLwQK5a7V+3iE3smV6
UoW2TmLm0kxZHCBkQTwtb/lo2qknjObAwYqU9kD9nJmLEQsefNh/vayZa2lyNgbl
qeNIwRRvVdjFsbFAJa65eMCwObX0fuC5RtKWY7Fb7JixKuf63j89MOpENEXTz77U
XIATPKBeXaHU7fjFTV6raASBo1HTzECutz7twJpXatmP3FbdM/mwIaQW8y0WURW+
NmrUOIpYQrLOL0mYcayBVM1MeFi+dhmEO3Cdi5hihDGNEwmxCeUqRvEe2LVlAtFI
GKoUXulvnQzqaCFAyLA+LVvn+FAEUHyiZp9GW8GIqsrrpI6xBirFOM0YY16/6zJi
mRLNXSBHAn10R0/0L5u4u4D1fBRdHJjfBDjV6TPXLsfIQd7s6g6nRNXV6sMIRwXw
ub1NcTCx5gcNhzWoOyCUxzvirP+ZkiOjypVyThg5OqvbFm38HB/Nc/J/W4m/07nQ
zaV69MdWnt8JkLk46HBvTQSaXqknoni05I6E/7Yb4G187XuZTvn3As71zUGiH6mY
/eMPNJXVsvFKdSJNWH1r/ntiapdJ6JD3L1gKzmCUxhwU9Q+hp+pO8xjoZcEj6lbN
iSwWQP3O5sWhD2Ax9Hvow3kznrw3oicgkmTWPQFuwUvdz6GA7Unahv8m2TER/Zjn
HYr1tyTLIspZZ/2RBqPUqTmF0WnZa0rvRfvaeIh9Xe5uvmvMRuTU53BmEHQvAxex
v9woYWk4EevrcjuaBGuMmlFg4lxuhawddmgU9WByJ80wf4eYMQGAI1p0P9lLvkCa
00c2nM1aneTqzxg8ZSJQ6KA3F+/uFgACW5L71qW00UgNybF91Y4e/bgjZ+KNBtWh
Q19GntudSV5v66PTJkYx6cWz2I2utCFAra3rrq+AxHADxsqay5r6CuJYuKvEGqMG
cGsdimoNcNWAFHBz88asVtJ8AEIAcY8dV2+v3RN+ZiFEHi8g8QR60vqdEQEG6iiP
kgJMzzAucu4NOaFlIa5KKfmsVfjuyrnacQvImNq+W0lxBcOEtNTc6w70EYb1piBw
adku1Jgg6JZhubdT6GQN1buJZg11/yFJcN0PkzyhyBsrdRp+jZ7NgUD8/wLTCR36
LTORXrFByhisoYALU21N23bHR6UkV+BJyIkTc8w87DEYMrqfZBpmOnN/O63wFv4G
tkPMGliWx6D0hIDFmgGeyxopPm9yqPB8BWB1WsUPvx1Vm3uO/WmbuC4iVepUKWfO
YILl5nbrepJrVS9qOHNE9VegyzdTJQ4rQG27nzylx2bO85hlA4Ffjw9P4P+7zYjx
/KrSs/EHfOdEtGxDHPJQp25rdlLV0NSWR0NoEIyq1yL2iP85e8Fhtaf1Aax17odm
nbBZFrjQfH4GC9jduJynp3XfH+k0aLBtsBNb5M+RhrD1hFB42BIo7qRfA4tMBNqa
wlRO7q6s+TpvCqsS6LseUne74WXdii5nQHI+VR+HGmN31czNGtHu8rrGR1PyVBXQ
VVdWYVbLUYUq3ExsnsSJGt0V3XY0vfTMSM20LboURMVsBUl5wpYPL/pAUqpMJO0Z
Q1aPv/2Xq96yeiWvGxobA0ryDVsEAGba0XoRd8o3iZp+bVyXezacv52Cpdj5UPdG
BeGOsW5RbMHCVMu7JYMPsNidqlZoe7gPmB1a0oxF2cLTh7Jo6MOybL2SwYUd8Goo
YSIJX/RwQ0RN2cUzkdBct8QI8TSi/35+HwZpO6WQIpMVfRokrB3djcf8kEGXyz0C
ZrY7mStyPh358MzlECilFPTYhEyKErX+bF/eTc5felRKwEd+fndDHDx75gH4iyKS
4tTu6Ni40tXKICPJ2J79/zyLBVWvazSWbKUy82SS//IWPQ+XPvwzdFJV2cdamSA3
EwA2xomkoRyXgP/XwxaI8gjtLfY4mPtSs+R9cjxXTVIgcd9nKOjV57sEQdcFZlHg
`protect END_PROTECTED
