`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iRZG6zwJYGwh5uZTMcvgsSPVKCYSL5LM950mrKhU+lpFYX7g45s0sip4T1CqOYj4
Gl35Y6ACEpRdZA/8/XKUmweqYWf43v25I8Pna+wyg2j8BMaN6aYBjG9pRq54Y6qq
8dXyG4XmKOlDituCQaODMl6BfTIWjbqY0x0rAYGvZ4wGp2TWPmUpn6Y3HdloCJkv
46ddToDoFgTvAjDnHxNpSeMdCStruPsiz8fX9455RjGuRU+nbMadXTMDQKFFgfox
8LVf2depOc5glxpPCRQuP42tMrQV2JlUMZdtFxQotyPvhNrHwYU2EBLp5qDWejTt
apFu9LYFStkGkFG8KrqgmsCj26ef2fbNUDfYx+p6PnmebeBfgltQ0KDEWVqmN1h0
JJ2YxJtJd+z047mjYgF+sOnazGZ6+BtIUYML+ugNh68BEgno6rDcbHQA2Qrm/Syk
EtzLnE26iHy8AyyADI1jgLeTHZ8XpXtkrJMgJwwgKf8=
`protect END_PROTECTED
