`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Za2KBaRJAUBbnukHYaXb3ddaiV6qU1bDsU6iFwd9pg95QpC4xi4172wpVJ35S8kY
UAjRiVzSRYsqRVj3yvHqmlTDL6mPsl/pSzZPss8LbmTZhEqJndSjYKnHbzT1t8v6
ZOaJk2L9msh9V5uLYiY9+FbcgpfnztejNkddoWz71x075JUR/7eY+LLiuOcFh4Hh
DK2ThI9xWiJASvLxT0rWDrtpzv4Oe1PRfShc7EAVWzRWpZZT3+yn772jvqEAshwz
KWTYT/fZ5vjuun7AZNJhZuuBeFpft5qzuRGWcP/cLz7gcOo394+YiUSY4tslI5uo
LM5XE8bYXs7aYlItcVDkXQ==
`protect END_PROTECTED
