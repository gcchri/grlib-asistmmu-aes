`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u8NStMx1qLcCpFynhVNj4TKqIhYjuNI7hui+dW6RFSnTn24u7MtxHK0ikD9fjlJ6
HNhk1lU7Nqg+t0tcXWLFDY6e1OXLbcFzGvp5Jn38XTwm0XmIaN4949/UrCIXiO6J
w5b3qZ2nLTTaiM7bnlto7XgfxmKo+iFmpzfUfQsoXWog62t3tCVjnU+klIRqwcSt
+S4K1C7LgBVNufWjvFL6AqlkOoCxoCrPss9/z3q7NObCVhcy/SvXnGvkxdyYwPlO
pgzdYGafQGKHwW4GXz4oR6FhbczIhg1NIpzVpb0Ilan1+ZL2MLe8YRAEdtowagW5
jg8pH3NfI9nWYHSMr8aO4HKEEJoZZiQrKs3I35mqPT2UQx8ImMo9dy0JBsB0KF5t
pvu8rKuc4mUczNSv9kw8hcsfpfGflztJ+pLHRwayrsRuVM5pBbhCqq18JuN3yacT
2SpWbI0gwiI16PjMPySlt3qN6SQFc12PeLF+ntPOa+vZTLyUZlYvad4eexrPLKm6
5f4w+axF2U0K40PYTPqaYg1h9+47IiGdQLaKb7WW3HtbjywcLU7+5pbLa1sUnxqC
oPZ67u15CaoLSSury/2Ci7+27+wqkprhy7Rorm9QMrfFY0y6Hu71aEUvuzpcX6bj
oTnAJZ0hVmLp/AqkmV47O7Zbnh5RXfZxK9XPcr72AyFTSBf05obbCY+IUKLpcSMe
sYkh+B4/hIq1/eJPcH4rN7wZq27+ap9c9mdX5OPBEWvijPJy5jBE06zjckdiSk06
VDhUsK0S/emKuMK3matDgQ==
`protect END_PROTECTED
