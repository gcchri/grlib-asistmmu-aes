`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wZwMxV19QLrh5+Y08OKQ1/rilaBEjItO7IeYd6qTprrEcJ/ARjEDVRp7/EzMxWm/
V0MBZv5k8U9lxgRMdzDAO7ahUfQMFmWTdByREtwxW1cCLPgSU97I3qO3XVMuHBWV
elanRhP4LBPUa652RCXRC1gusPqiSN/5+CvoFKLoHVc0g2Cm3G++80JOWYTyHd+8
E2bi3AZs6gJqIRCoDsjtplMAHi3bmFq/B0UDllPD9bSDQLBHaZ1lK+gYQg7IRVYU
jwHIDjyWKWnUmHFo7zyDD2F8WXyrMVjle3naKENo2XDDXwWSgbYK839IBs7qq97Z
vvH6WK5EabmsEZqGr0L9V4z8D/7TlDgIeZ3Xcm8XC+8XtgbUJ+iLBoI7MID2P0x+
OnQ20ZIAzemfSRAOEIGoIAAoTxpbbI1HKLCGmTkNyhQAjKZrHW+1ec/lXhcBYir4
w2PMJi7yq1C/4qh+PRGghi6btCLkD9VoGQEtSl5a8GgngmsI1sMCEt52KjSvsrrN
p2Iykjs5cYW80OEpQbEb6BZ9kpFOnXL6dLNKXf4dKYO8TbV+R349X2ZVBQPUhvED
o9B2vG1RmX6lRdQOQKD7Yn5jiki7IleR3dhzk0zt6XB6TqHtmXYCBk3um+uYjIno
8efRlhsyQ8RSIyAVvhGYH7JeQ1bXSV2QTKgvBAPBsXqBBXqRAjNwk6m8zMEYI50i
yOSN53TWhnbuVrWGPMmAjYwznzkf8zVZ6ycMO1hkVnKyAS6NpeOicZnXw+3T7urB
puagK7zIbvjcs3uNBkhH/9Zp4V2rotL8J2cIv7yYjheCb2H6PleSlGR/QNQDUjW8
ICFykDR9HCL2cb+yPiOYmx88iiVM+vceFD0QPmWlgO7VkYagqNqdqWyyceWRUk9t
f6HBs04VkjqA/0GvsNppJWZXVKg5xj/T+agCb/eCzZ99tayYEjuFgZ52Ex2vBPAe
Gbv8yK8vlh52HGuOPdxXc3m/Ue5x+50gDmbIG7BNZ2Pn0VkmLkkn2PXjCmctMKcN
A2Y4h8XJnwEfm2cxkoXBqVrjJ/hpibYvo5EgpWh/nPWo6hleS6f6uZiXtv1pGzO1
OAbuN4KTP3tr3OJipksfV9yIdtJal42VXGIp+PBcQ9o0B9juueXrnQbp8GCV61hH
YMU6c2AvRjviqPeRRy5yFBtVXIykcxiGeQjYh1A4AWnkQRoXkECwU6lC0zAGsdE9
FCvxYoeTkEUh5oRb5BXFeuua6u5Vz/jE/XeHTRINpNwNewkhVhLJUBSeCWd/YkJS
ghQZRl3Cl/QDRwWeTixnS0bMf+W4C243Uv9C1/HeuVWfWXhbq/AHh594IMuzlrJ8
TSVxDd5YfJv6cJM+cDS28OVwqzJJ5+GmWPjbYZZ8ZnRS4upzNbvUe+9xN/gA9gTt
8xUD9p9nkElzThhuZNx702qZ3NvcjEwIiKEoxZEax17sX9PWU5T2Jx5jF6M/NRkn
m6vBId4OPzIy7WvJU43bcnJPjzkq0ZUOKeOQaY0TKeizUaPap5Elzb470JG347rs
yqLTVXUqthNjeEQr6lP1m2U/5vQwLJCSNTRYMqc0+8KXskhfnNYaT4I7shY2aD59
cfEvfe5h7XCP5a4c2hF2L6QR7w+orhz/jhzBYSR/N0rohSVlZ9H/g+RcjXNAnmFT
dea+plECTkXLfsM1kdnmwvtHwVvZnq8bEQohBol+zpBYh0aO0DxvvVcxdB2TSncZ
dO7DBIIQPa75TD9hJuhbK99b/jauOdzmonMB7akvQ5I+qeg+L60odGL6r89wZBq5
Tjo0Hr9NwNfgMqkwhhuswun8YEqqiqDYKSoAaz0s8m+IekgelUfOJUI1a8WecmS8
VbmUQyGhMXT4MX7OB9mGQuBfIXjTw24WXWIpQOAQqPmpeYDO2GxRQAV3wLONrcqc
ywZ8Hdi07Ktv1nv3oF7j8TMLUoUjqwAxfaWk8pOa4gtgGpQQPd2TB6JnZUu/16Xx
EjRRW86ROGAX/Q3L6eiWARzo9XrBrBUUy0qn0Z3Y3+MBUWjpWQEbQ6iuZVJ34knV
HKHuRW4dR209B/oHYCaDQeogxg3UALAkRipuer5IT4ixj4suIU42wyUM3PljjtMA
92T+Ak1Kcd4E2R/I1LQ3ZwuPbVi93kEOhTm4vdapPQX0JAsaV09VbRPyy/1QbDuK
jWjGpboQGxHE+1gbFOo7fgb+DEO5VbAmvFOMlBSPqAwdJiQ3CqqSEZfFlWXsGKgL
svsgfMNQFdkEJplkXdpc789cQhpgfJqH0AZSr450fxP1sZuPsKDgXtKcngIpe52K
11WN6k5ftgr9pEJmGlOdDfa0G+Qrmxhzr1X/zTrghEjXdDsWUtCyUqowcR1eAEK0
eTBLEhgKz2FCWhel2RXX6bLR7Zwz8vqVQ4DLZDg2hdPKCv9SN8OTHrXzipNKiWUt
MR+Gs/1GcbdTPNWHbGnaO9WQVqZYfOgEyFI42vc6sRhKM4quNNCW1JtUXpAMkjUZ
vEXDPyx57jdldBR2IFu7ok3rkvhthPJJuPNgrkQicqJRrRQBNRN829uMDyd9o1BN
LXu0VcfRM9jBF9wcMXJXtkqRPd8Y67hCGBEsWCjKhPMjbE4FEW3NjHhRlmA75TDu
gT4vlnEA7hbmiT2jB2IqiJq/J0MFBfSCzjAx5JU3IvFjOgOcrfAyDEM9qUNGuR5j
1xtltmnhNiRTeh+dgVSmlP6vn3hoD6HeBVOteRC7SGXIY9pYjmDyM5ZhGxuAZLup
ge2vvE9uPSM3radShCIAwJNhtSTL2z7/l/DoPKrcc9jjLc5XfVTmkcSpUYNVes2Z
EQAplMAHHns9HOLhMer83dxZu+DcSOrgLV5PZJyJAvFrdf1HT+NLHIYgNYFmLkve
/zgraVWBCHthKq17HGGLnhSrqGcEmzQlYAA3Qmc2g40HoOPQRbLeHoX6saRRJDsS
sOrIfdzyqEUeBETQJzmLMguvUDkgCdulazY1A/fKUjdLRwy5lNsINZLmUZAAlNOR
/+QsyuYkMQ5yvgiZEn4Vyv6mLN5DVRDkhLK8vD9xy3Nl630c3Swn5qPlouX7D2YL
j01VlD/I2GDvKL+xfESo/4g/srUFnKhs+2GrTV2UQtNDwFdP3kzdEUXkY0FgV4SM
UVjTxPB0bQ5CGbHVoiMrrr5QthrCZZuxLxXs7x92Hdx7Wbp6BW5CQ3/pq14/G07u
0kwBbffewo0d/fWFPv4aErjQiLpOZTBmYhKMabnqy7enSkmNiKx2EPFVr2wEooJS
xJCz98drz9Zv8v57MCZwT6N/AoM7kkJ7GplCkcOJFU8vVYHoIaSKMgeWEmcWg2PH
fhrThD2Snn3iLfB+NXFocrw+eKe1PIW24ZsWk362TM3ciwg7hSbgeQ8x3Qhlgcq0
N7xjxw0slPo6sUdbGAtJIzb9Qllvp36CciiL+K4fqLIDhkTEhJPM/KYaq/pF5/Zn
rS3kEo12EJDgrrRuQ/17spyUp08I6rVCJSzB4p3HLX2Y93ZMwUT1A1gMgxOv1Osg
1hGIAXbZyp//ogytmvrDzT6AzPrGgHd5LuieoUQMmrEEeIeY9RorfvqAd4bUo+sA
yr8SS67r2+pZcG/0qcghZXfAn4pUvmOrAe0bty4njKCviRlPhHIYRfGspr+K7tIJ
g7GkIqk0/30tBibHEFNPQXRVz0R8emXuDGpY7yRZEYQ57Z8CgSI8g7+cxq2C8YE2
OcAn06CeW/dpmzPclrKdst0BM2YskzewG7AFRB/CFg0s2k9fpW4bgALcbogEQNp6
aW56gXo8NCzSQg+QtVYoCtD/cNzFh01nEpeIUwU24j1SCAKo901uM6awqf50iOXw
TWhiZg9PsGCuMFfXSCjClXF096NgSpUm25LR20KSzMw4lgIWRgszjKRIVYkR5XLN
J1DiRjx7Ius3uVZHhPDOJzN1Bb61D8Ow1f+BdMyo0xWXtmajRBMlMHqrh96B1Jtn
4bbSJ1zzgOBwovtQCJP2BG6vZjBhKH3fLgTdPPx+C0zsbJ+yjrWy+zGijvus1AEc
RxgkcZaOnVjmPVPeDGLKVgyaeHg0N1/CnLtY/k4SsMkKKaspekpiOEAlOQ3FrzRA
ok0S1VVOlnzutCGWEYYCBm4GGhuBbsjX8o6BAD+NP4PikmH4D34whW1dcG/eu3Wb
p6w6fM6CC95fzhgz/3WQQHtkwRHZpQetLtttrbv9NbGcRWcwyRxTHE83XtIwcM3t
W2Ffer/ReiMkl3xNXMgd7pFlLoce/+1eIhvROQt8/bzSfNOm7LWNEQx9HbqsGvpX
KakB2ZOhe5qP7coDXkUm5FdasTtws/CaTIVU07ktqfYdPLIByOuOpu7hmHjb9Lfj
th1yL8OG1iYEerZst6seff1VdAWm7iYZgCc+IewdJ0dn7bVQ6unPFFPvpZXqazeb
OhVuuUU3U9+qc4vlnpgDmOyzxrRI4r3/ucEgBsjB59O6iE6jKlXWsP5nT20yGRUw
D5si69X3SXSUzg7iNy2GJ9OidiT1b/gOcTGxmgp6WBxSNhrdckfAMvQCbTuBGAfK
psdjNGXvrDiirPIX0vYS8zXpwC8ZtYddnhFkPZQcf0oLn3yU7IIgki6+/w8364po
7+76MzQUkYKetekU3iQ6/5P2pqmOjX3Z1dq2FmDeGZQf4O0IWVTRIuWJM2ueNsYy
tl8Q+iPOg+8l222mImogha7S8NNOgziB+74lg9weQp8YAKAoO3xQuPKW8pm1X6TY
rGbrUvO825B89dr6ilOit9mZ1YnjWHUIwjcF/30kbSnGI3ByVcg6JKFt+ahELT6+
KMnDvmx25kYTkkNgyvYx96Z0z9soJcbFy+TVe5q7SAOmEE8ZQEEyN18XCoi5AHWx
0lXr/1NbTyT4HtaAvIPYCgm8jeoJROm8tp4nwgJoEH1FTd7qwWPWfaMHRuHyjO6F
EaTWMR27GqCF98vHR2HS3kJOU3WY5byqjKQPQD5sp4/QvjlFdkUAQCVpyQ0pWVjD
QaIjxs6HlwUno6xJcezG7efjsHrz3daR6HTcjHHAS5ZkNaHlveSe3cSQO08R++rn
t8Jbhp31QDuODTbaxBfCRmQlG7jHcz4PphbCa1BuXgUWZkyWl4UYu1FEf0NjklsN
N9hR4JfZuwfgnG4sh+8hL0v9w90+Fhgp63Vz2azoOQerYa5nf3R9rjDVOYKXNH33
SZwprfI3hxCES6DA1FXbk4TZ+9US4Rw3kOEGBwZXSYsjHSDyfkmFzg7qbHdrkh3z
Yd+Wyhw3XrXdpO7lAw2rUpPapmm9Z6zM/KyzsY83Al4KTVZfd5k1VWdb9se+1A4b
ZNA6UZUoMWW/OhkOeQUMpvCowuZkNJFq4jrE4lxJMNRaBlAxMxxsIFfIE6F3A+2D
WvqHgQf765ze6E1L37mmanyo9LdqUT1d+6qpRqR6MZGaJT5dHoDTvg1P1fqktu0o
ykpBKyWRSeWY/zTgvrbsI4j2e39bub/oJvTNE56J/fvs5nT9hTtzP1n140wB0aEF
td8CjOlEcgzOGc35gN//Fc0zKYZ7EO8mGTyYDzfz/GK0RHhGia3o1u/ImK+3sJKX
6QwQE1GnsVUm7f0q8TgEh2IqrUH8l+12YTJR/NZY88glcuXybMvMXU+StzJVyXWo
tX1oqzupqhztq/4yUkXv60WTTSg3zz1jnWofGzL6gFBMoJm+mfGnhKpbw0AkP2Ew
PWPeVd74iLz/Vhu2y/jK/wxe6/3RGl2fDL8686i+fFGBSTYL392G7g+eLmrNeX24
qDptYcXVIugAHHugUZb8CHIJdK4XWqFxPLgAf6DlJH2ZcXyYKxs3xKh1qcTgAJH+
z5gALt2ATv3AlbrI5hXr+XCjcvKNguYNuCiiEQZJd5cfd8zGMtNFYTGF/As6OdlQ
twR+7rD/MIrwulucYerp0RwZ+oqRuro8teAQNb+/9w9pAleLtJPcZr9Opcmys/qz
u9O/6qDI+kneeUN59z0r+WBZJneaMTyi40EwtXL2Gh0lKlzD2fTbh99TNKP79wU1
x3W5KmNXlM+/DBhq0MWdxWqRLSGffY1iUmHabnrXoV9uu61us4ylywW6kJIVe5Fy
QAcbJ75F4ewWTyj45XKNPw8Df6IrlCwchI4YCUFxompKv/UFPKisNuAdwOzV3j54
/HVu5XTv3N0tlLJZPtu653OrxkMTyBFNPKNYSckQETvGV6QsILHbL+R27+f3YMmh
8PecuvyzjCm7XxuQyMAp6kEB8pOOLrREBnCgChC9gaB04wkL6sCOgcpfW/sFAw25
GGsTXJjLTh+wLrazTCjwh2rLXuAQuZJJyEFR1eRmkI4px/DQ8Agefi+obMjg0MyR
xV7dQKrazzj0wyFbXc1wdd+cZXwiQLYBaNv42bHqD6XjzPTOXz5FyTsJRqFNK1n+
halnGyjNB7sblEuxmh1EDWcKkuB8ySpjH3Id85HJOHDlj4tD8ZtXFEEPd7+JnVt/
GbYutNSP/0/ZWIgYG4tQE6pvXKn9x3WRFEDrUP1hs1EHyOiHeYpwj4F3CJM8wH8x
wu0+JKR56Wljf8EITfF4ZKDyLUm2xB6cbfzrjPZlg4Gm9R8lRigrp40SZzkVkNOB
BKRAqd0LlDGmaPTR64t4Iqukjwy6dCGpWMDeJpozoYElCTg9PIuKqEY9hIPtGxG0
txdEPvAQWzuX2FzxlAiH861b76Onfxfxyw+CjRbjjbOxTC+MPm9mFHcqeJiP11dT
TDmL9WbIQ/3Ak7sD4LyJbIhgWwoz+pUXzhCUqlUnbgpujqQyW1j8PvpjwCm8FW/4
zlfifs/vkZiV+px5boVGu1/nLVTops/RG8ClUbRQiNY6n3BKtris/7phaORlqdok
W4ity73GWlYC0sKlRLB/VHGaCF8/jiAVa092d8giDMksqkmPPPQZgebVcmmMM82U
SX32wL9uxjrOA8gaNP/QgeGIP3AK7xHKoq8JqY0E8ue+SXNP4l2qIksjPCHGA4dk
WX8eYeJuQEkfCZlXqVPcc29fLUWP5Z4NIADltFrE0v01v0larIOqS1mCjvjZ/NjQ
+UlV80m/jFLqhFUmMYVdm5hPbaaYv/S/s1NAFdAb4S3ZE+27XYhU623luRyrG4cr
1LSPa3M8EEkHoWLeyXUz1PAMVN2MmzpdQfCmKp14VZugBjvM6bpn+awuzAozos/t
ZlV0DKeiGAP28UpDM0BOQ0ezYjP5gbelFkAJ6TKRcyCBiVDG6t/CBHZg7fzJ+v6I
j586g1jGwz20aPaAmKcH2CbLCy+z87OEMmlXfqpwxbjhEgDCGN0KgB99DC1sAYMP
h9uBmZt56NtD4sBNc6ik8Fawr44n1VbHuz+9oJVODyvcB4sQV/M40dlqW6pPqhPH
H5u3sA/sUbjerWwMiTBoHOMqYFX8wgd1gryHOP3vhcuh4HENl8PydwzMyVpTidaw
nTb6HjIF0VXS9lH/aMW80VgfmoRmYvFyBcHPSMCHZo3+jM+3qgebDHBOe0J/+MqJ
bGJNZSnvLtbScWZfnhDDymr5d79UiUbx6ZDrKtNSRrysc5Wrgg4G5UsM8C5wdiBh
uzvZRb/nOT0kY05OV1e3bZMw2Dkqv73CqHzePIpQ6XG7Jy+96QFClRsNQFEHsw2e
mPJK4TLwCdXlEeZifbDDmN7vs50jvGDzQ3lhYHOq4JIA622oasG3cpa1eJHJJQ3H
48l2KQMhSsIIsbDq+DkyQ3V9ScNWc4sOoBKk9lXlbwr84lXHYiSKW0g23PfyTdDP
wfCEf7ISCDeN71sRnsGvIcaG7RmnqGEMWqBksJ+YwvFF2TfWki6I7Ug4tsEUGUt8
9KsttUAFo5w0kYZH99P23A533LBLZsFXyq7gUzpWdvTS37WchbJzmSOtTSuXwuJc
VhROyPHcvhrrBfxqfW32M+K099ffXSiGgEYmhlVNhbIEEmxbF4L5JQYyUj3HIP2w
0x4gR1y8+SfucuYTR2Y5MfJ0bI7ME2NbMOysnk74R1gQ0q9Ghpl++lGdHnvtgIXd
tsMrlTFie5RMqcA38I8kk3v07t567j5dBQWkHnfddHPfZ2+TtUNUTyJijfjLkf8X
+uElfwKPcnqX8ppcyjng1fJOkkI2s25i8GFGY79O488JGXIjivY/xlo9J7CdsUCC
NHBe6KsKzwR6SQl+t82DM+Dr2JsCeIpGxsiuFm27GBIsVDzv+3TbMiIUZp7L9nNH
0RgGwPJ47+DWloca5hRHUva7hKNVWzkNbf+ajwGGrdFfN+WdAk7G/ILKWpJYAvQT
qC3VCjGS0nTvsbp3NKxOV6qhRsnYk/MIRmtEkOAPoI6cXWNBih4p24+dON/YNf8S
eZ0jkYOnviUQKDXHL03p1ew98IG/wk+yTe+vxaS+q5WDyC2b0HvRwqxTtc/8EsWB
WtYOEoG/Fd+oEQ3aD7+Vn//Gjj69SzKtIRkV4dRnXOOIOh+XmYsoNm+DHbsA9wQ+
dEz8gNxVE1RIP/+ro651s/PhnLkN34EgBp68KsTldofhwT5cNXz9y55L6DRp1O6i
+JHb7GSBw/bhTy/oISGlaAd9en+Fhgd1udGoliqfakRJlFMp3AV/1nvXDcq5EnvH
+KjZJ/7KEuZ99/ZVbPZhwyFuSRWF03d+jYjwrbvNJ8TN/ESpzyYYX4EiFyEv1QqT
zyRQQw4UlC8wgrtOIJs37JxzWlhobOWUME/rYEUSd28yHSfTOiZ/IgH76Vdai/1R
vGnQ23pREyhzoH8lgFsJo85/A4xHz909T/saRrmOrnn2Rt8pXZYbGzqr5dhy3xV0
GU5f+64hIYNVO5GPM1OqyBDidN5HRpyIMPVUsacw7IKdcKsTODqfatAh59yeQJNd
hDO6Pv3ifLsZFNs4M8UwMAXSMwwjEOuTOhKJqfCtHm2Gur8hCr4TmK8LQTuMoB6y
8ViG1qJb3riuckkXDPU+zKAjVuej3WYfM3y+Al9JEidx/O3K0uki+rE1xw8Bp4TB
47l3mECsTs1FqpQWiSuphyuOnqI0swLJ21rEkgjPi3ip8seXHb67offYiWAbrQss
s5O4jf85lRxzcKDy9f4VEZwA9dWG51x4kTBSdtwdE/gYhRjGdlW6S9ThGuxKJ8lM
rBlxElAYDGPG4uRDRgFIs2XSqKy2u0uZiJTjpNeEox47XwYV0xVyBnJEuc2kn5PE
nULcTHkGRGi+lakp/gjvdEWIEagFOO8/AoRXTzcPwqYdKODSWcp5ySAe4Bt8BbMU
p0ynxrW2ruaZ6TC33uGTWT/VGRVX05tBKbpJoRBCezENEOYUYeKiKUkTuVD2of9C
C9tOf6Er/TXYAuHPnXfCziwtmlPYoHQ/327RMilTB6FV84e+LPfRAZYwITTnwjyo
YGcDIzoKw0ucu9z5pUaYwK/uMSBDNmw2vxL25U44FTdoDVYcgySsj8JhlCGi9V71
ANO3KZqUd5LskbHRWxgPYIXpRy/lB8hqG82oIc74YORQ0ONhUsuP33CDpE9zIH4c
ZVb0ylPrKJ1MXOUchlfLKcuRAGHGokw/CTNnwxkbQQXqoYt4AxTflW5SgCtX52Vs
MHxF5XaYkLIpftOdIfGCSgXtzNvcA7AF+FkW6vZ5xbAogU+BUZhT276GmEyTOteX
bpqT/QpstQnW7nCDG8UwJ0PS3ESpPySE53E1EYt6zf7+s7CJQySfDgwmLOfdxOeH
Dprxa6sq/D7X68AfwddA0NhGD7VlYGRY3eeWWaNMTxji0CJD7/cr25LJZ7tG7/gw
sNqc0R2y/TAP0ea4COQz6Nm7hFkPoHHujg/dzMMzscZCthEnOw0dcsDPwsfogaFY
tp9o4Xl2LTznl+k8sGXeZLGLS4oOY5bNgfrzBMAdI2oeJo7o5QCIeqGABTcBn8R0
vZfjGI9WPXJfzGq1oxOyJLugGAYfxaI3GvFQ8TE+HJTPDVUXWRLmP/RS6gb20gdm
CZyMX0CeljnCFsvGSh6D/GR1cRq25e8SzIns+twzRrYmpFZXIcRriFINzxvxhKhB
FoO1Z/DZ1BRp8eeH/tCa1A==
`protect END_PROTECTED
