`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZFDZ5QH3FdhRmF9hNZCn/vALJR9pGF940neXbrOdiV3u0SDtb5uSiLNI2WVR7T5P
7BQPI2koSAbvxJBcVA/u30w7+vo8FKIOG1GzsRyMNEem2Q1erhT7Jf8uN1E9CGxP
RSZ4YDa4uTQYO5OisaQ1B/Yw/3oCL6d0lrBu9HmVpcUwRZjBHUhNRUwde2ZYo/xj
SsXZ1eGbrGLG44jr9LSMzS3bHTt6DwuWarLeU0hTGB/9MpmhHoGXaZtHDO4pCLBJ
Sgy2Vcw4ho9iOU4V9j8m4XflDBW2pwH0VFnjeO+hHXMeKOUoxhsxgQ7QP7nGLpH0
fuxmXCax7J++U/2Pje4qfjCE4OhUtakChON4ClGsaTW1YSR2KdZcXW8ro54pN02k
89PpDg8ntG4twUb1Li8plgEUeTpEjaiVnMPGd7PL0K2yO1y8aSHJrkzo6mRE7F1Y
7LWz7BeKLZfBSyYHzGa8oEdpfXwh3iX/ZDf+XW+QTzuqsk2pDGsuNvb1dvCuIZ0G
2rSAIqHuLUlK3+Gte6QHaXpzMfxpWhzWZhIVVfitHbXVr7yjbR/JLfhlNoDXSVOm
vboybhHDM+k3R9iYG2IkBOuU1ri0Y9KsZ5rzcG2ZwTvTv/hQhoSKO4g3fDYkLDQV
fgslhr1pRzxneyp6GbwZe4hqgOO/NwVvcacLr0CrWnRMYuWSZ5zRbQPry2rpZqhI
d5aspRCfmBvH6DdTRzc816UWrqOTOJAbVLgmBHqRpImi/0m07O31f9Bp9toxa+KX
gUT9MeGja0TynRM2/nuY/djlvN8Fvl+GNZNwyR9Wy/ho8dFCnLSA5ac82AhrxG0N
7cCVnUGEq6Bqe11f/WNyp2iisfCOGNvsf1RIyYqR66mqXenSQTEZCRnRl6OYDb/z
GlM4TV3GjZuTgnIZYz23093FYd4ihd8/EwscQPJUXjagaabqcvFtnjM8fIUSb7vL
6S2YUh2+KORgVIUZ+3r8gKV+IXlRGZ+CzzavpEUHJKUR87JTdk/aIG4hOkq/MYXH
5skLEwyOb9hBvs9m1mWvleMmMBp6Z5fVJ4kR4uf+6hCtw7Kepv+vhaEou1rR9JSK
2PpV1RXTG3E6zVMtsPRFx2YY8bjeHfgpxxN9L8hpWWuAXHzM15k5z3H/ucfVhjmo
PHfhj5MKliR73bDzuMj/XZWk1tIx47OUJB5gRfDJCodb/e+8dr2Rk9q/NhEvnPqT
4RfIevVZ7nN/Wfid0MMTs1w3LAj+LyS7VSMuRdHX+8XqdmVM0hS99BrxzGbNQ2bv
Zl+hZxbIfJqYCRXXbC6Jyr/qHoW8YI2G/wfE0SiqWoGDyUb0VeQCYYcuJRlPtls3
7Y9YNknv6oJIKqi3KzK7coFaSRZFubFr/3PzvNDlLlAbZ9CRd5u2RudGuaoXKyx0
/6Ksi9jLKxjyvUtjP7ooJoVw3NEP5BO/A6t1KEeXI9RD9XyxeGuOOwt4i7ip3EiV
cvLr78nCjjXftAACZxIdQPrCAeWEVPs+wyyTnV4pt8HXfrxjwv1FT07nxb7gdmZR
vNejJoIaICiR0l3rUOo92GAQQxekwYZdGdsJRMybP1t/rLcrAjwHBE2WtlJMJsrC
h9NuOo3EHgPY8aNbPY5saY1n2qJMKY+5FccPMohhQAjnI/vkG2bkohbQTyzVJZiW
TKmZe+kMIhIlWcASJQvWJ/JGytntrjZG9JNUu0+eO93FJkbQjVA/6WI6zK4phls7
sdeenWoBnL56v3EEhWjZF26lt6RLMtHvCqUbpDocbaU8/2R1Jz96btuBvtHlOck9
tEcenjgm7r05220EOrrM5FZaUQQXRXI9B58u5CyQvn/6lTdetuOeiIYUA3Wg/Ua1
ykhTE1neAHCpaH9bJsNemVpDuNUBlq7KVKagNc2ZRUx4+xvn+R+sp98vO5cSZYkJ
VXhcNX5faYr3fzXdE9oix+M3bIncZsMtdX4mMcF88NqLo/hdhVRP7wFwUtE3KdVv
F8Kr2/dDTh2ICSJM45PmIQd6NVhAIeX9ugMSje6/wezsfouuvjuczdW542dAgoeY
TMPXyGMydSaXz05aYqQQyL4KucDWR4bOvH3LLskhVG4tgT/DYfXGmfCCI1yDWGDb
dfCVYmtx3iEE9eAP7YVlr5dd7er6sp+5i3BRnvBPqZH0qmjbmAvfJlq3KQ/nq2Mc
gbHvHI4jlIRaijYBziA5lpb+c+xfOpzDoKi5C4WU633lQMGkLlPnXUQmKyvsDHIi
cGc0ukmSRa2tos3YYQRPVQ6Nk7kgdRzCufcIwEHp4Y/7Ka08SXOwdIsv0YTpndsc
XPlJZqz4+nUFnwZoQ3VoTFYC6jgovMUEruiIMujN/uDPw9hpW0c1M0M+yih/exQT
CJZofFLDbcHuRvTAPGV9uwLG7OEdto17dmMxn665NBMDLBWW8w/EL793PG0bxisc
YeIFnZUYJBOqALrfaedVfw==
`protect END_PROTECTED
