`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PXSPSk4q1RcHodTJqXYvaei1ZYxqb67ozcq83FTRVBlI5pXvSPCjl4URE9GK1L/S
dQyu4TUPzPtAOdK97P5JnWmeUwp197m9Ubup1tBLHnf6XX8pZTAafv0JwkYrQ/Lv
ib7JLhQwdu8ZcaucPJs9/2CwM2OhQBZ9iTwjwcI44lIBtEPgaELqazPO5kAFcBvg
NAytrz2sT1BZh8MSqaXNGYYc5VAutOVyc/yWfOwT3nmxiX3vs+U61c2WE08SWCZV
myMF38vP9w0adY4h34lLIYBs2fS2zhS7p6i5LV4tmBpPxBUgazy/+84bRD2WRzoo
8/fUuJiJ0Mp9qHXIcbgcZVARUpkJJPT/uXG93sO8aW0Ux1Ol7ld7ELYQ8YXJAXvs
c+UnrfQg39WG3PtbKGqh8WPlUS70c1cArfxnmOGSRbfZlM3lCijLOAeuO5Q0qTTi
Q83oBLlZve5RM0Ilt0JxMIGGB09Y1xbDeifGTKufMwoQBt37PE9EqfPtnMC1g807
sMyyn5c/sFXzNGbS3ZdSu3w4KhC3tfo1kxpiE5UjCJKWXz3Z9qguvoTrVeYA95li
kgrFykwz0vt24KeNaPOZ4yt8c7baGsxK3z4qgxUFW8bBe6aBh+CVWxzznyj/6zAm
V2klfWM48W1ySPjR2u7rvDFyd4IWqymrp0rMiRFhxIvVD1UH4lgDizTD64sjU8Bi
D7RYXz2yI97FUrI/scWw7MpRzwk6u9yCi1mLCNt5vs5I1my4yLn7S2s6DIwWnjCG
LgosL+NDSTIkWo5qr4nS7dNN+l7CY+BRz1blX6vi/L6/owNzcRjFKip3/T6R+tKh
jytr3z+OOduqlSlrwfi7ves8mxnRL/I64gfDOqH3FFJQfe6s4HTXizI3HGa4TRkF
8/Kv9qPQcoswIUR9R88pQp0OlYKbJn5UlQuvIFsBJxEugFxAsD9YdKQr3oxxtTsw
8jlMlFdyuSDUsU+iVvn+tjKjKi88h6v7yYhvNytw4G1qZs+3T8knHGYKZCafZ1Y+
aVxLs0VvoF+uAGO06122xPMBkNhKLFPcYWsdNZBMJYFIwSjra2ZkX2qOLyOJancQ
CAYH5HBOHJNO//ABsMNLNwTlDFK+ObqRBOaAnJC7Bav8dEgxaGAk3+Y+TvFKNYYE
x6ulBTqZ5pXzSPhgWWgsOSDDKTdLcDLC1IdEMa2kT5OBfHHQcFNPZwmvwwQNwYIV
K5gzn6O1CzaCLmOebl0Q3HERcZ5BA0ci2p5U83dEEAP9Dv8Y0MLMljsE9MSnPhs4
ThO8bSKgX2lXIS15D3uSdCTgvra3LQPDk0ZZMkMDGwLF+2PIKREC9xsCY/7QPK7R
92mR/q6sfYvuaPRvF9w8dYNGMFbYblMyrQZrLJ8Xo5E54tqrxq2/MKfOZd19r5w0
WNb40gNjMqtiTUC1/0sDrBItvrmNOe+Ah3ZKCvsG06DpRqnbf3zrLqsiVlaSDXa0
MJF1UuFsPpd81/ZRCsVDan0iBK25SXIJaMTrC8/HGmafht0VAudebcyYcNsEBcCy
t15AJwUuuHnEuxy0F0WLz/IqR1jihHdjhIyGfz+rzGElGBhteVutWYDuicELl4N7
o5GBcUdBDbySPHMq7P5IP4eeAxCO9qjTf1IqBEwla4LJX/aLeU8+jtMwKg5qfQ7/
PUjBhiGWhoGDqKDVY/5j2yBcE8xCQfg9kjtg/1fKKyUiHTxjCgRDkN/VCTd4uKVs
`protect END_PROTECTED
