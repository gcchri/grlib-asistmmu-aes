`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0yrAtqvfwgDGIh4Po7s1UXcjuW7HoyBWqcn7z4FP+LMaHNuyVFMDw7IOjykLyKNQ
+SVqhoOQoLgXmTlIHd0QePJ4zl/GJIDfWhUZVwWUMmEuw+8pb3/PQ7u2RJw6rGk7
u6Y1hx/IZNomYT3EhFduRw2zW55G17KzJfiZWR2tEsBwxyk3Y8ITeOvjKtJhDHUU
S+rRrxajYDpjXg5k2RSkV0d18RzvLpnibIWxgFCZYzO9KMzjZGhPcaC90Sk1SAkP
SGrmR+c2EmJNyR8ul2OX+ZnURPCgFURLmWbUMbWp6J0S1DDatu2naDOW1i4/l5EM
MeZdYRpDHeYeMFHeu9bOP0hUxjVV7R5fErBUXk0PdkwuNwoG5P7jQYpcG8BSGoOq
rUTD4K9QaBM73jc/Hvfl2WVMTAtd/EAcKB7ErPauDd5IRfqgieObby5ExOMhE885
DlGGb1I3YS+p+hsVcyvUmzt+0ph9UDeogTG7UoYADackjNaNXLxx3SmuJTJpOiXE
vHbeekrtrMcwSYGMJhAAA8xoh5r/7OnV7wWDYSwu87bRfeQzHiNyjAtDPsLCuKLg
neMxU0pyes9ANdi07tURvxxxGPs0PU3xVMs36BHW4TGdxtN3WcX2KBNeZn13gJs7
UTV//EBMorPNWh/QNshzynhiMUsdinj6SlJAJ3v4QssKHiM5RSjfw84kmlPkeF0r
3Kemwe2UbHBA6EhWzLPNOL/Bc/MwKS3RGAtXY+6NrhsmJqm8wWWpn88jztkSUTdU
1DjSI+Oec41u8O8x24WPZgYAQBdYuyIBj5rf/UCfh38EHAmc6d5owSkOna6vY54A
opi5ydRzr8BWi6U0WDlIZzrrDmjoxGcl38xuhi/I9Q6VHpna8y43TADq8/rf1KAc
ZzfxboRwuZ5xM/it0OUHH95yk55/vub7u98MSzElJblHxtcjDm58Zh5oPUp7fDT+
`protect END_PROTECTED
