`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4eywOkIpiRn5x5u/lxBv2NWINsPf6jDiNib2QbTC6PcBgPCHetS8/Zc9zpetaOeT
Kf2FxwLt2anKJdnGqAZ+e23W1MVVr4Az2QUikYjtnaf3lbLoojgAOkObns7hjUmp
Jhy2rcZCQrHL7bqs4aym4FxjKt99L9F1yPeYh0EDWiXN5Ra77tSn0ZXjLThxvaw/
Ejz8yL30l17S/Te704ajwQr48UtB5l+x9WWMcwmVRYIm8OJMTv22gSQ1p0xc3TXW
XWXQA5ropvCUn0h9e+xWs9x+bRBl8eWaO/vpdYrwkekvlAMetb6lWqDyZGOgMn6L
QRRTlkhJWRBdTWTVw9hBaiKYTWpIqAXtNbsqrXu983j6cSFJZr4XqIU/o/7nGbr4
DSelTyeJJ+rZDMPWyYRLWHy+I+mkqx5XoQW2CpoUNseEaCI3BwM129xmbhjx4S2O
U1XP4LEx5KocOph5pF8H8LGWtyoqiLNzak/gjRYLJeoQ+mgOcmxf4shECPnCqwgj
`protect END_PROTECTED
