`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dh/ExAJjp1jHnBhkEjo0NsoDrKxdvcRw8RcNfyeKnysjdnNgLqMxvAu0jUShqYNr
nHmtu9ksTprIXtVibkQkowfCSy5mcoZKP0z3UfhbNmXigl8IodjCCAZInlF+qydf
7PueJ9vzTjLTCbKKM610trCs6FGmoUe+SXxGc/kKNLr7wfxwtzljpHFSUPPYN5LA
Yx8PGIoHvqqRwZczQEK3fDLYdujG3p99q9Klb4jPNK590e/xJZHPMV/9yDo322fI
9SHsogqodLpQL0O1ZgAfxXW6+hYxS6QikYBc5sIsKu0GfWgrPqOXJmrMED9f1s8g
5ncu5GUwqefBKaVAPEdkWKSusIwEDKsjzDJR7Hmfx2RjyTEY0JIiFqSkmAerujLn
qtQwv1y44PQdmafA0tZst031DzZRBZal4jy3Qhws76xzZ8TL2hY2YANZZ+aZQRqW
`protect END_PROTECTED
