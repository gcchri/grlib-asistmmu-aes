`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cUEiJN0bIZwy45Q5QLMhmbAymlQnNOUUVgij1UvxNQwbbh1d6R8658fd94xgXmj+
znwveTsLtpSULGGKbD12m8PWcbmt40vWAYQjIbub5pXRexc1GALZPsCdQaBR8HkN
3GUH8yGfTdw9+pTNRbN9N2quojCu/FqFQOJ8G38xsMYJriFFGdjkqC+EakH7D41d
QuNNLy4k2TJH50W9eaL1vNQwjUQnafIKLP4mrMlb9TiyMd/qAqpmOem7so6SM+Tn
et3CLahY+3KvoUcm3AifZE1H3VKg3YzXWU+OR3yyvWKe1Kot6J84288ntfKsamBf
/q/3FmH3IhKmlSA+kOXb34/l/z8+3YFKlRGP2aRbqep0TwHPYvTvlc7KBjZ3akI2
ZSSNPs/WBGSRuvq/vJR991nLz6Fd2vJBZmxiKKsOebU=
`protect END_PROTECTED
