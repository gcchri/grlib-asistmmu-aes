`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SnTr73Sb8dhSsVJfquJMuMEVpkDOsgD+Lg/BcRBWsmZ9mOUwL91jFfiIhotxNBlB
272zUYMpNcfwwv90Cf/bq89wGP/LbOEo32700r3hZwPuJURTXZvzW8zWeaOIdU8m
3vZ+7BY70X5tlchgovnmNonycG05JWamMT8esIxbsjhApf9W9k7xMYTbHXjSlTrz
CdJQ9US9UXLb43dnROUWXR0OeSPRv+6rUJQUflSEoLsTMwDr2kGVV3CyFjGz0jhs
yT0P7UKyTLiC4etcIZxng43gqbWc70wHbnvaaegD+e0=
`protect END_PROTECTED
