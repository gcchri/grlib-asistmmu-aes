`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x+CjvKf5gOovAc3i7G6wN87ZItdLKfNTDTV47XH7zHZ7aQEiVXvuYdig+id2S73P
kO6QAH4FezQeIIuIbhJVpZfngeNzt9Z0nSNwY9A0kdmn/SWDBsDb07tWSrbCbhib
QuCBQhNiC6OyJzJ4Qu4ZR6aJvjt6FPUUNf7+IDyE4gXrIlD+e7WDq3iWxl1I+ear
pUEyXsKukorPQXtRe52IfXrmdlM9Y4V6qQO7lDbXkxqR3XcYTvCh+QKx7VnFdTVb
FaX8QhAb3RHHCOTi59qhFqCybeVj/BavBvbO1aqSNkjLeyy3LMExuwWOWSyu90L4
Om6jA//oD+hUPH+/Z+CL32hR/BnnnAa06VA82ej7Cu+gKwbo5j+eOQVJfkMHan1z
LmT0tyoXRn0sTwIu29WWQwBUam7Y607m/1IsdWQV/M7cQYAZJb6gupZUbN1yrjGC
CQTWbUOz3eEf0VJhPMkF1ixjPLlDCmRmYnRCeDhCh4jnDc0aUMHZ3I/zcfGcJwgs
W8NnpRens2eimglmb218EdPuKRqGPITdu+N0F7q9IOFqxKisMQiQ/spKfdRLpDgK
Z/1vY7juzlo4sa3jXzSRA5waeLiYry9/AvR/1xTXZq0=
`protect END_PROTECTED
