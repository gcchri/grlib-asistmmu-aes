`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BUTR5diCr9r7rqTImcMvy+t2VbEiy2dMlr3sMBIHwr2sM/CJklP9/c6UJ/exI9WM
qqvHNbbjqfvu3jeby1S5/tsusdg5RD7bvNz8rHUx5ROMhRSq3ZS3ghyiykEaXNF/
IADK8JB8xBOr+YW3uqGyjwfJ3ktor8LAwoRVw6xhdxZv43l6v+CSfipzVNX0lsSA
29Glse0zwtWQtECqyY9vEdfYXLLjsfuvR87ZG1ULcEut7lHORvW9tByAGVlPFS+U
7mQHVvMcerlqhkq4NxfJ03NhjTHb+Q87apsDlGv89zwL2JnHe2VAH5/M6vXgoJh6
eP+k4aR+GLG80F/f3IxwR1Ta+KcRheCNUTh9Jvlp786tvoTIvsrMeV6rY5SQg09c
yV/9kxDIq9osCkijCvz+vC0QoW/ovWwlZ6aKXr+TbZrr3IyU1caebYtELUZFeipP
j1qNK3Nqac054xK7Gu5mbcFz1Pmd1zSdt9GoC0mH5aFAApnz6/K0mMdhFjJ8fu8M
U5scu9xhB7Pe73zupve9rpCdtOvfr+c9u5q76wWgXyRxJ6ApHm/eBTFxZ/JCRA7o
y32+7z50aTRyRxoIei9msYj9zUqMiweKHHx7owGmNpVVaou+ym9xjcI5cnWhDjL5
RfTOX48YcJu8ATKEC2g5SrhW4tezbGSvCrG6dLPJ3YE=
`protect END_PROTECTED
