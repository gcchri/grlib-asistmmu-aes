`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qOjH5PUH2Jr9rhqAfvv85tq2MsHXikdO6xpvZrTgYK0sO+UKo6D5CcmEhBV52DZT
TcCTUkyBFkSE6LHfvGQOO2HOwH7nB9Ybeudx2sC3PTMC94+uog+e4/J+y88V60NI
H99yNCpdFRKS0CL40i3QguIbTqSp8CLRbFVWx1MLf66xxS9R5mZGIsMMFl8Vg5mF
nkEfZxkPKcOhSqI9iEAOtfGwYJrzPV0ViXZ3WDi2soHZE1Gfk9kVo3XU7aJtRpwI
DC8D4a3AHh0blyLq79ELT5rhnK9/3RTRtV9JkYOA73e5Ep9mwTh7itMvF2lLrEMD
UqUcBKF1wfF1IHjQpNrq0w==
`protect END_PROTECTED
