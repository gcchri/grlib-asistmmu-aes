`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
taqkLr7NSoMmWzXIBZ0Qg7anlYOmXxF6iZEwD/NYp6fB2KKz55redTaXrKcz/yFv
3bIp40lyA2Y/9xZaUGZMzVZ8kXe0yTGGob4yODy6hubPnMfbxUT1xBAuo1InI+tc
zyi4BZVbS4bH+qg3uY8K8XF3g4vYu1GY9whQHPqKQm1vWepGUCFNmU5pfalhG64/
f1orNJ61D/sNSz4tlUukxrF2dib+SCcAW6dJu/dkj9iol+3bnBzKkvhw2NmqaMfu
+OYtxxU5mKfOsq+gcoRmPle2w9ld8m1wsJKmmcrhozjVuRQpFpn3eFGJViz/UdWP
lHhYePrqUY3osb1tlT8HZtu5V0age95B8ownuIU65utaByIUm5tnZxjCWPVc9BQE
c4QxfbZwP19HoBOXh0gX/NBwGXMqRKDiu/ZS9YcKMtD04lmKBagl3BGVztBM+zyr
OlkIOf36ByhJH7WssQKDSYIGaFvVPlbdQBytB/CD8iK8uZNfzHCfeNWogfSHlETZ
MUi5V77Fubk7QB783XEggg==
`protect END_PROTECTED
