`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R6UVul1lNBxgVJ8STJ4z2PrONhCrVffRf9gZ0LlLST4PY/AlC9RXE12xIKoyvk1y
QTNVW7sV5fdJl9uAB2DxGy/y1lBLIlapf9lIVsrAJHtkh5nrk6PofECRDLjIFIBh
hm4Rzn1fgGtN6H036S131LoAMDfBeNHwboW4EfXPjJs4kv/YLdY32hHk/RPD8URL
KYx9b7qMtiSIdFNN4fiXTVNya96qsHgpCjVIxTuy32xTstpkPi0plNGbht+I4BXg
HV5zKSmbiG4FWo/8YJRNo/3ay0CcuZtJ9KD7l8WhUf4SBjd1Rfi+uiyxYonA+n8v
0cUno+IELt2L4qsPmYO20xYMAS9MJzkBSOo+okwckBoHTSTf+KxWjkfcCq8pKc3J
0HNPltaNRXLVR3EIAszq9auPQ4FfcNOKUckftQPPkV2cEbXg2ktnqcCf7OYdhiQP
5HE4FBbKGpNwxagQM60gIDdmPklvO3eS0A7KjImM/LlSC9RerAGp8kKHoYozLm8w
ARZ4j9ZiGPrYxMt1dzvmg1FnWBVYi/YmuLUWfZ5B2TwIouUoRH1QM8eFc/jfC7O6
ZLjq5jCyX9KVFR0U8Py4fk5qKDRnxvmFswNdSjfFxyBLG93rKnhLrgyd934sHGqV
JmIxqAI1r8cxWHGykx6owg==
`protect END_PROTECTED
