`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QJ3hv4R2YaweiE2/BLuzW+Vbj90XlnW+9rNhJiBPT90CJPc1Tyik4d1DiO+SlLzg
dv+tYpB60qUHqa0nHwjF4wWwdBuQdJeW7kzgcE+su5wHALRyG0c9YWn9H0Z5GzYb
ufdBPWsvlYCZ/Bk8dlmay9VCE17bFL+7wVrRF3HqRAscfDlHAI0CNxduxTeWheyn
pB9O55815dB2W9YVzTy2GApVrpQdhBRGjOfHHYHlVRLZVZr+jlJrEwRiE4XIVLA6
6d21CeIvatjKOK9zg6QQziHP6o6kys/wptE5/wklgyht/Rvwj4lHP0t+Uhn9yClf
j3DLLkCJNUudPK0jb7t0bMJEu4ZXn6hvOjHKdav71++xQuYKNOExR3dMGutKfx3L
CVvFHMhH+kW8Ahi+Hk4f5YmXuQ8qj7QPFx+OlWpZ6IEo/Ss+DN+fZXjFXMxCXfFm
kSm8Dl1K3xWX1k1XrSJEj5A3FlGtvzi55FNRJ3d9m9EDwWaZbpxS1x+41w8ems5d
tjQFw+mvrdDU7UVOGUBykFaSd5ltoZUmDKKm1TNXnufNZniLTsdyeEYIyUmyTR5T
3B6ghwj2/U1erOUBhA0c6BuO5OORn71GMm6yANT9xI2u1g6sU2TwsBOlnzMdsGbd
54saF4oCBQfovjfUitjdJbBGO4YgAlvjQKgtYLdyxqvbjFIpCdfCYOg0UJBKWTKU
jA6WjSOyHDeUy68vw4xQTg==
`protect END_PROTECTED
