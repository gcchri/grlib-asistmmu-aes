`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
So2gRI6Q7vwkJvZgQhsDzAXY6Xwca3d7xfbSwTh5tBNZJCKZUPA1EYrCZNyGtVnC
MQ2k0jB2fUMLkp9V/lo/7qU7U4k+ZUhrO+Oua7EWIko8zOc1wUOSA2+m7J4lRrmQ
E6FCTjFiLqomSsN54LSydGp7qQdjAqbAQjnauqSkg2kD8hRINzEgKyP9TMN/QPU6
UUEkXxTi7t86+YVljEbPd94abcqszlyv+mIHuR0Lge5jM4MRbH6WHw14r1U6BOoL
dPayi09AY0l7miEj1hWWRA==
`protect END_PROTECTED
