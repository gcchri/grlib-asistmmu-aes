`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kfAzM/mWrMNZpKLbSps7TYE9KNeRAQXUOZytGXAh3xrKz24BmFX2vIckySy/+kJz
HOePlvyaNAcL4ND44VFh3D36LEeqSjrCoNQVslPZf0qxgOaYgJZ0SxhdjS6s5nka
LWKuAq9J2GePa/qQqWRq81OrTz2Q2HBsEIFowSlY/z3GSp7KxI5tyViyi4owVKs+
d3kSY7NkMuw3rEYtntfFu3YxJn7fJXEpDh/aRHl4GGrE7HNUTK39VgcqRKQMAupi
zqXqHZIQWgQ9k9J52EPIFrhsNfE0LzFWvae+KmPLm0SR1FBVtCIE9RV5U0LFQmcl
au7QaVFNbLqGgqBYicqoJVutxNByUPf+W9P3KCQdHyMHMSzGtvoPvloG+phbxqiM
HUMnD6GgRRz1yw5UUTQyNw==
`protect END_PROTECTED
