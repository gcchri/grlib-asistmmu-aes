`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GAzTG7p7XdMprFRR1R3/eyO3s+otT5DTeOiTA9DHpN4mk6cUNYA50b9XZsEIp/RK
gCVAPru/ZCIwa+l8pZ2qrk+A7kb36vlkZGXGUsM8HAeHkPzTFBDLeFtKXSy5kwuV
lIkGYguPzaetg3TKNRII4fGn5uXob9Bivb3jdtrwsJqJxdDaLq5J1KtHbvz2tK6H
rId1TWPOlSNG78DVd/f0zKESfzQ050i9VseVgjTKo7f8Z6VsnI/TZ3BoeQENvAaR
cY1h63438cQO+xQAdUHN/HptvoyZS6Mf6oSz5+TbHEriyRs+rPLEcelyI3uVqpvB
vcKGcGgLo/+yDFCTGUavadpjgc3q3M6LgExz5Wr6iY9W7ohrJA5L0xEdICRHzj/s
ht6Q7kdnqSl3onKUWwDxGBj7BDlIACe9qY5yIBOhtis+XcWuEgR5r5GGexEriePc
LyVf5FkW9NeStLegmp63v6RQGHwjlP97lF6gv2wQbPbKxTcPI/ZsgUXDXNVDhG22
pF5nmr+vMYbp9vfM2ZiQrD0Po5NImPOc8KmbT2PSE0xrUogWqFjjSC8idDP5arwc
9CZL32Us6OMpD+35RS3REEZFLail64xmYRTgU4cHSBEf8PdJzqqBI6FkobW7HzA+
98BwIzo7JB2ko3U2yf2WIaOsrT94ltqTnUJN1HImtPGL1W7act6HfpIB7Js5pLrX
xQCx663l7sS+S02qYFTkYHkVWU39c6XOBoZ7Jv2ESJevbXpCzNgC3aUIp5jZAhjZ
D32uGwp2JiGYb8Kbn/ThQhRNcR1hDjo5ycoB1QTs09ZlV3FFmAQZedrKAK6Kb3ol
O9+PywrPujFfr9ehe/E7PEb1rekVIuglDMZkhgN3bW7B7S+BxfZkEkoqwuBfRg9T
+U15y9CKHtjK5/SAugwbNbkqsGy6vYvyEFQj7dmuNSQ=
`protect END_PROTECTED
