`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p3KuppuPCrVpJMWCX2dZX2oyJLlvYT8UER2bxBDoGeStJUdeYBRCXlhUnSLNKg71
uj2/oxeIniTvSkz0oNIZIc67h8W7Pcd9y0nakwuJXkzZ7o93JPr8xaJjezJ0/+YE
GOFeJmZepqGYKGR/k9YhDNSYC4i+9PJtY0bquXJDsL5ph2IOJG3RQsp4jz0hp6rZ
WQoywCLsOUGaYvHc6dnGLMjPSFCpR4O6UxcZUD/kHdMfgwxOfaSUVHA0v+UnplPH
tlGkYv7Q946k5bvZVDqSabCx/sjabKLgKUmawdgXJb8RNUUT8/Wb7DEu5JWU1COD
eoyrCQe70oJwMR1fH+8Fs9UM86JkVvpaC9vhGckCHQnqHTzdLueWJKT7L9m687G8
kb57eoTugZ2hsdyYeVJOZq86DZXGG+5bcQD9FjKU5ljl5/dLzRGwTOjiFlPHUoCO
vDMUlkgApxzZ6MNETyDp2KNhYRr6UYCLS/Tb0fzyUKwx7dbEnreEVARSnJqQoRH/
fyOfWtSH9JQgTKCriymo8YXnJvXl1CcDGkBR7AwELNPLUaEeVQao/3LTYhgTodR4
Nie5wXzo8oGsPGhzGYCRjhT/EOBVPX6FrlLDZMM2mmU=
`protect END_PROTECTED
