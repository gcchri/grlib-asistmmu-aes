`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qFrCvW9Cnr+lA2Y7xGDc7Trs5IPkzX1NJWNbrbNna/r589AR9wlRHcoEigtrGddd
NpkvITI/YNyNgmu56/DY357PFpOvvNRUf3mv/B3e9oWkCfkxz6bvkqSZEhzlU4CV
NkXarxj5DICtnJBDsZVxIdwWT1/1uGQ3VgNkTUvszyPljbk41E408Rz9IjD1hMM5
/M8w4qVVD3hPy9yXCjLTJTehVnkde1+aFE9M52BxdmFouo4X1qtTsu9NiL7ay+me
nUiwj/a6dr12yKSshHrk5vuuIpNuWQ4X6PO5yrQPQs7tL9UrWD9wPeL3wLu8Vj5d
ji25tz0mWrElb81MGbwa1w==
`protect END_PROTECTED
