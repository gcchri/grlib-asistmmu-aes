`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9YLHh/3fttUJnFOQ7Gvvyg8jkcq3SntjpMeKx0+4li6BSHLr2W+otyqpLKbQSfuo
XXfd9PUOFX2kggHoLETjnboTNzat1KRWTIRYIqEE2Qod0mZu57J+C6ur/LRqUYAy
JZaTN62uoSrvbyNz3ocC9+D4pAL4vOrdnELi9F0gn75UTs4ltdjya8xT9HeRQl/9
ULcdB0tdCP/EdtojZZKxl34qadOYpz9wieJTSpJkUXQ1LPFsLsDDwIXYr/KUv6Zo
/vbPa4vWeirsTCxVEDix91eg4SvZ4+Q69QSjj84t3VcPI1SExnS4PjhL5C5lJHak
X5h1ZHzZMngRUEJyyTabebhsvf/MBl9AL6LGaBr/WQwHpiAa0B2QoLT6TTQYuKBD
hIwhEAtaAo+eTNJJqsm7D8rDVQLGhONsrR2/tZ7E0A+8ZNlaHMfhC6ESngSsv8M+
zpn96kpyAQjgshdFsgzYWFDyLLeL0gcdtZJkYZ3AVJY=
`protect END_PROTECTED
