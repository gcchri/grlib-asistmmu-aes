`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1mQQOin4gAg0t/aOliu/eQ4Mn/pVsJ+jrwTeoYPrD1VrmbTYzCl/u8s6zpC107H9
i9IXAjowILwfRHhexyw3+hBaEzeGDflzlSQpC6oSzxhoc1ioEjkkRnofff5shwJo
f5Ij8aqYZ2SJSjwLoJ/qhT+R1holc8uV1OioYK2e79gkNC2HA8kTIAIAn/kejbBY
EXr5Qk8uEvYMJkPUl6g/0Q==
`protect END_PROTECTED
