`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5gNwabnRd5aicXUxee6F18M+d7StMOZDTkJzoauKjCfz3NVFk95QlrZEJ3v87Be0
4OMj42PIQKHoMRz3ynVb0Df37cfOW1ZSprq3qXcrdTB6tt3avc4S8QBSWY1IMV+t
jxCBmKRABeRlXQqnn6rJ1q2Aq9zyrvvHNORaIA5WiHg+RifMimBnxQYSAcH5Urka
+ZSTnEBV7tV8YBxlzCAaXpyYFPqci7UWBflLd4OdZ3x184etlg4xbaOXpbTv5Zho
HL0QcFAdLtkmI0QfX4+ckjnmAuHYF7plLtbqZ781FDfjQ/nwHOx2PN3KY4hr+pMe
aVHbg2tJXaC2xGf/qqfBri0ja4QdNWNORHJT3uJ7NpwKhUn0vtIQDWsUe8j4SIUF
cUJ9Zll5mUCwQEuVCKjHho+lJOQLHz+49if8GMpH5D26WnVcC6Io1092e/XRxyNb
+AHLEVtSM1kPDdyQMbElSdToN6yBLuthDJpGGgafBHOkjbPbNtB6v5190S4x/7XP
CTygBPkriqvvQPkm0uqQurabNH/w49mang4dqXW1V6TfCny3AJZEeI4+f9d8ZRNx
RqRflHclSu4uNy/NtjdE1fNsay2F4pNkU91Q+vMtApoo2sXsQBp7q8167J7OsHNu
46SOzPTWQTinOe4Kfpl3xdPYLN5OGp7uKhOyI58u4F/Dm3QmcLEJQWn456WecV5M
QWqidP5VhGSFoiE54Da8M8lCjuXkdhD+1KcWa9ZgR1pSQsNOSobaza+iajIcB+IK
Rb3jiKH6x6pF2piI79UQwTc7hYiYUF+Cy1/5n+Gb0fuNawqD0BCKHFYZ41CTECif
1aKYAVsVdRTirA1HXdP/hekOCoRUmDCyh8Zydk+E5JIBMa/UbAmvA09PSGPjhaCC
jaIJMdigZ+k/fOaHCKcm6Uzq7ubETg58BigK2SL0XRDbEkvIwPewOPBKmVkpriVL
kL8iZSYXg6n9+2lWczBQ1uvvLWi7H0V/P9C8wLgPz4ZvMbE2qBxOn52mZd6xQRqp
mPdNuq2oghtwvjwwchRj/D5X/NnC/oA5d1fS1yCVr79TBko5ZrAI9qht5VjVzTk2
TGqY3yR9HpySgPocYNuEZvvlR4G4fzcBN+0CNQRuhPAXp3YH4GA+qsxiLWejGFmg
u9Ffr9tBv8vj1Ay2ylC9wdb+Dyozxy4AgqhSsWYbZa9grLbsljyIFdACgrwNgoxI
xlXrlsJElzjg66nocBb0JyJfXSoqXE6mSVZFD2SpxF5rRkAoHtbcRoGPSwwjqnHD
dSTZO2vi8e8eT6A3JEoKXmKq2ypI8RmKOkcJAvZHeLmeM6E97U9lVBUx/Sdi7eul
P6uPA7aGt9wvd8LEz3uvo+a9AdftY8XGtFqqcfibwDk9V1bQL82bzwSjPidbO79h
vHFBTLhqU64IDpNeGw+/n7TRJ+ZPAEz8DaaBjbXQf2aCohPzq6cg8645xUHbj7+5
iJMEZza5jzc50LNpCIxVB/jP0/sycAy/aZ58GcaE4+1PEFTHxN8w344hwJlMIZuf
HsICrFJx7pbOoHkS3NzVnU0JshfScAYZ+lRR6QUfVV2xr2XQOWvSDD/dcv8OrZmr
6IBZQD2sYPcju+9ntQwRfrW0YeXf9DnFw/CZpXyDc1zaqNxTrGa8ls60RowBDmxZ
tylRolwSx22ymGxZNTSH6eKvgnNG55gAs4ZLQTUJwsGlLB0TtjAguqf/8qiINRpy
QgWSAsP2kEYGvN8MxAK2Wny3T35CJC70LSuP49ktrlu7w7lmp71epkcSySgoQNUZ
LjdU1dpnM8LCvAhe/JHLC0mQnc9Uj38Y7v9Q/BaXCNIJKujKBkymUoaGz5LhD/p5
ZGYCfF5ZnjrEht7q9ZsFUCbsV84rnSjy7GDKaGTMnexZUU/meUOmEDdLgJJv9dbr
X+U2vyFG9J7qikfhB/Twli/VHrYu7IeRo/n7eVpbeFu/8ZgBSYuUwCoBdrNpypRp
qobVBgqk8+Gdpi5fZ5YpN/XpKc0C/47NgeMxWtzJSj0Akkf5pdSH8dpqKDqrWYoW
MlDsXxA28z0QH1jZCEbnq0QxGKR3Uaab5JudmlaQTEK8fsTsaElfze0DMZ8sN4fD
8u+wMhTrZIYbam5HCIZBCEyHv6TtENYr91caR6NycwnzN95kGZCTPfXzPx0q4LVp
pRoS00GO2OzytDgHwxXkFyQgtJgSFJAGRAgI7WRkFsXLxqa+Fa4bbdAZBsKUqOOw
gjY9SBaaziP9FhudGHHHsjKNoid/XAEesRP88eT/M3s9kk6xteWN2khEskg09A7x
Px0j0Kj+1Ze4PLQI9SgZYtsJG9qE/Rq0BspDGVcbJcwtgzO0Zhdr9xojscpbnPdE
fuiMDZKLVa0cUDPp7kFe32koawmVZ3HQnG27nfZsT3ya4WN6XJwmlR9EAAG8aCHO
hS6hwprc45NNPI5vzbwZEaQS81ChytxH7G4SPtdZIE+ZkZ9+NVBGIaX/AB0mmOsv
xG3mzLR+043aVxK5LAnjXz+XZHsD/Hd4Rkmb8ppQfzmpAV0eu8R9xYQ57dQfUJaK
TDYmN3wbEQLXHcYqKLjSuYlPyXzWE2vHlb7wN0cOEwow/qgm+px1IwEgenjsPg2j
YgSB+J+KxxflSdmJQMw/diNGmvuK28flv5C+yxohYImzJFI68D7MDktoeRY7WsIS
bO+Bwl2HxyaIsVX08krCqMR9nUrKm2GgRkmHgiLvJ5CBkI59WW2eZTKlR6h5ojb7
Dqr302nm+8xWdiMV77Ivcg8xafCLvAN5Avqtp1+3V3o0wIzaBdSm3kFNE349c2ii
neCF92HIX8rOnxNBrHtNApIQmOSQx1P9x3tnjgLxLeGTl2pgtBoZyXZaOAk6gWsL
90aGmmdbrxdCcNCijyxQCAbipBBpl/fnwRZpW4qmWvYBkEfX5ckpHu/wPuQzPqjS
0jDmjBryo9BmI81mrSmPIqZ/AembWgwiFdQe6aUdr9DcEhIvYSGQerFfZfCXBLU9
Icqmu/5DTvK91FZvUQvODPOL11DmRpi95zpUAsopMoScYLGEeE7pPxxrB6vXOltn
d26aHzI03zSimoXPeHRCchfUtca+f4UONAH5iVzgbgJMcIQSJo/R2dcMnQcWltob
Dc8d8/3lDIi6QYRcCGbyYzOKm1RCyCvAH7pIcSYvOqAzKwbeKDchYPDB+q71Ivad
0sNNzHb6Bx82goKeR7tF3+NoMJLgUQVmd1OoaHL1cwCQpdMW3OTOQMgL0dHVWGtk
YR9WYS52H8+nwD7YA//Ehy4rIl1D4uRJv1jG/fjXqqYuwCrrm/m4pvdS83TArIaB
0yGrc+BLPBFU7yqHZ5P8J/bYiqHojOx4i+PZ8bdSp2QlFIRiILPb66ThE9TRTK4Y
tnj+6WLoZ4OFDo/WEi1corqiJhErtAnRy2uzOQkNo8x7A5WgkzHGD8u7R9B6aeKr
+ck5cZr8v7DVVE7Dcl5zrw1Pjxtda+IcBKoBJ/SWtjhRPCnzF7aqeZvR5+avRyEd
3vTV0hHEfZslNSDsW+Q8+/A9bf/sqMp7HGoKqyTTU2KFEg5lDzdw22Z7qjrG1AT6
aBrLc0kje6ZYS01ovxj7a29usHQzkGqPROGa1LESv5ZrSplvkPAWS1cBvyrKdZzz
SBB6Vxiji3uUGFc3bzkfkaw8igpmrK73muENTFJeQw9EGbueleiSyT/Ef98gyHFF
s7G82ItGHj7V30HAQWOXkiE6Q3WZZewy2BjsnFy3EjwwrpnlPFW14TQU1KMJHirz
gp5PQgYey1QF5gqUitVVbkBqZu1nrkvHWiCiymHky6MRH4znJFDLlnzV2BGLEQHy
FdeqgN40toOZTTmqUnirsFVEYdDLaOtdFERP9Ueo6R1SihYloWTQlmyTD9KxBJjz
sqdQvajAKc+hizMXF5pMC0Y4VHnIXRszhcWXGYOttP/DcqC7q5ptKnekCzw6zUQS
CBgeHiF9QrFJGODsJjgvq3NEccwd8fvyjk+X/yl+zwHDHAZYHkf2e1Knu9TlisFQ
1tUs571IiXJV7AnTGCq/UNVx820dHF8+Tn1zlyhf6EJ1sb+/G/I7IqbteKP1JRw4
MjhmPHfB0Pnyl23GdQ+gOCQvVU9/4wtGHnHpPun4HHgN+T4ji0jKEgFdE3dvGLEl
qrinx9fecNkmFTmHQK2hqhkJGUDEPrcb9MyFlCqbOrh5Y2SzDSXRmYWIZS6BUye7
VZRUMX7YloVrkm15ZewPtzzeSygjNRT3CQVxfJLylbvikL2pE/pzDTNh/HgHsA1Y
WJHAkHthKVg8aNQNv+PbinPlpe61OjkxzbgmfKNk0MFOO0M2FSKSLjZlAY4GUOxI
5lLv2+NZSAWJ3PDc7qN6Zf+EgVmpXjQZExd3hlJSnigVaRLAbA/27CIB8qE5aCTU
vixf3ZLSjnJZgS6ByLbF203J4Ld0Wb5/ehTE3pVTP09ytELaMXxRSRB8snkoTypJ
LJ1BFKpkQ2kW7qs0cvLhv6ez/eifhd8zWBSjBaRROQ/rE5TIWn4iPn4KpWMckGgw
4Q55l5cSgQi68jD5jRNTnITPrnbQwT8mILHsRhDDj4p6vQyWeytbUxUTTSdhd2Xs
8e9JH4bFQpTbRPbMtngzm3fD9jUFFHDMkZIiR/pZPfV8gUZXTP8AlHQoGNhmwqMv
UrLvHNFSpJL8P+Ha/cqeZinW+ezjDfZ5xt7EC0y5vMPGDOopEH9CDtiUvaiFqxT/
jiFMNh/vFQMnJiMquKvmbS/o4U35oVefsd3+WKRtF8QsVeHgPB/wobeKFJ78AOFZ
5kgEXdDxPfoNfNEbYIUXMwy+2Sykxn/yVMdyCSAkoeaviBsLy/Ds8mKda5Cb32D9
4ZDzHBjhzl4RSNXSXguN5hDVKS4IlIHFqsLcB5rSIV3qFrxBidRd8n3dQde0OsQ/
0VlDWxLW1KGBdhUCv4alkZ1RN6Hevm8rVhrmy0G7lOFSBv8j/Z5Y/GpA+65jPkzd
fyTwvBqCuhPPoNGeUZwxwD2EsBgUkmmTZUDoODzJPoHwBE6SUJvjT6ftwn70IFes
DysaRzhAR/f4BGL85ejJVNA35bhgq46q9sfJZ95yqyQIyzp2r9E3Kh67LO6tM8XI
vLsyWdXWx6lqwiRMUcss1N2H090/VMCGnkWwjJ8HCKuoFVK1ZqIsOJecHWCxsLdg
xqyfCDHPLdMU0ZJuwDz0aYk4xu6lifKJFPzBwY9GMhjom75vbD+zEJugsaoQzeAV
vyT0CND1r3Trcg3XBVjCN99vtAtclSkMY70G3LGSBluQn3JhL+fyE3bTA7CQovaI
I/uK5XjOL1OB5quoArN8/kyQWZUrdgOF3vGR7K2n0RoKOKETabicjA5etHSvvnUK
0yZOdeZJQvqpnt4xT2gqnd7Ls4zjkZ0sLZh0B1GYBUVKTLzzVpwFvbZ5LF67pV0N
hbZQy8ojU4/2HgdQrhb+d4JoXZODPg/1KRIHeye8IrzDR5v7B0RJ+7tiImB8JDkt
dUJukZstTWOITJH8bd+MpnxbRfhun+kb/y7o4bcQobtMYxgOBhMSjs2bVW/5T4qn
UJjGFV1CiEQlm5KsuBD/wOsaikpe/OaWEtQ7j7vcz+HvsRrS2YdEMD/q7aeg2ofR
YQik7LrsGuCk6svbTQtyVKBYKksBR1Rlc2kJnJSKeaNLOmcjPog65SX1ZUirU1Am
O0jAN+emBDiN5oNS5fhWcy76QIIIje1FUenIaSg0pKu5Wls+tS8L2+ibl6+3FZpD
PtshLAWZlmrD7vtbbWPYHWjCjtcpGwYBUID2ZpGT7FCRutThJLU7dROWuebLCWew
fUgQDNeiELKCtFdNQbJ3F4lPvWO2RWfSroek/DzF1xrDZggMw44GmM4l2Va5681p
1l7UAgFvRSfeVs8i/pKpmz/WcDkZoNGkbd2WE2nBYXfconanCVhAQftOyTlyxFl8
s61FbCOQMFlDf2S2DahglYJk8gv4VdzK3RI90oG3fX/YppfDRmLBF9n/PQoqVDIh
Iy/3D1V0zRZPN0xGWTnI0vC8We+6VBlOdipX/oPzthjZ3QMMTttVf8mvASwFWP+/
J7qt4daNxAWme30w3B5DIgs+BYNRPItp2aMGWUB8kfLZGM25V7vCstmk2UdBxu6X
Bdkf2qx9vlPxhDTqNoxBoqeQ1Nry9tzjPezmUe0kcMm7V7bzV5+ct+SNKWBV9hdR
eLISrDC9cL8XuAOWeRTcDrdVOSgXWL4xh6IuLG65RoDciJt/7oVS+jYx0Jz5tU8Y
hdp3h8WXBQakyXJWov/qM+iDu/UNlkG+XRUO9CZGBOhHMTng/LqpW5PqyUuvqAMc
Bjg1TnkJQG7ewokWTFrIbI0FoYwDSqQ41BrdtvqwDZ7vmFUAdLSkoR67HEe8E027
89yQz2wU2X00FwOXrgLOSDm8PB3JDfbCr7o/EFeUly38wKcDfMx4uB2f7u22fMVG
IRo0FfkL1xFmGQPZgkpuAsJLpKOwunvPZWe5IWPxdmTJoef/7H9ZKSGhbnZUt6UI
DL4meEeEot50+K2VzxD2vHORIHcUTKA5eGjgNtR9zC8STqwtVuLUG1tRpkFGEddG
Jcb8gDq5lcd8v391nvZ1jho5bNn0QuOXLU1FmG6jMq4eKnAnvqhha6ahgKyyAYEY
CBN7FD+KP0BaM3+OhmDL+Zjy8DCJphdRs4l6vhdLL1ei1NftGf7DxbPtG6gzCQXy
EnMEgXZ21UQl4hDY6hpZdAxEB3Bl0Us/6DIXDBe6EIZDZh+37K/KEEMplHir04qL
mWP6Cptw03Xv82FuIU8iheqFeTspPPUIKLMQANXYYji/xIQ9t9a9S4nsBtPbM/az
ULrGW5bUVTomMcPM/Uwy7iS8ta7xyV7HzYRYuo0Oq/s1y6MYm7/O/nbpwYNnc577
lzWNHslrv4RFd8FHLJI0/lAt3+8Lz6dyK54GePhxuGZZJoCzX5V3XB1Y6DzfNvGE
C3kZBlLoZzgTDBpsUw3Y51ahawXEFq6cYHuq3kJsX/a5rqYIpodtdEWM8RJUCFp1
QeiIZZ6rAeH6gcxS+EXlv6swNe7OM04aVb+VjXTzMcl0v/wal2noMqZfiGFH+y7g
WqFvpXw+S9vGndDD64Xu2XjxM61GwWBZA0EkdspacWW+2HIspEgjhjlfiA/W1FcS
/t70KOupIvRBvtG7dh+8bGQ/pnBQ6vOiuM8QFEOOQjpL3WZATHfPO/vijJO/12Ud
w/bXuqV6LWKe6h2/vPuGXe5NgENQseLSoXxn9x7f37hyGJ1M/THRxfS2fasNNQdX
30/IOzGWmh4M1Ik4DZV0Lxep6hL7Mtx98GV0GY9/WRduZEapp4yujeD7Z4KJjvL5
tVTrUOaHm21ki1QFAClwwmEL7Us+wz8rbZrq9tGVm+k/2PS0Wl5rLtYd5OlxeeGh
aWV+WrcIPG/QYb8KB+CNgDS1c1CHiRJlG3VRSvNGX1FzyX9t25OTZhPFUSlW8PbL
dSuPX15OJFXiiiKyQIYjhP0+Lhn85VmFK0TjYByZuPqgUBW4sz0k2j8KdK2pqADE
RszP0Y6gj90vLfEcwbE4ecroMooOhJkTEQGtl7Z2OE+gWG+Xv19W3tV8HCD7Kr2U
bgdcJAg8nJFv306ASlov7uB+XNp9tZJKFHStDLoL6i4AwYo8aBgE3URdxKWVY7ds
s5m0U2KBpoEb2zTrPimnfavOfxSzfm2eHKQrYZ47uoGEOtn4hfGwio4DlTsG0KVK
rH6Gh6TikzO3fUlUdocmDmI/SL/cgY/rxvRpLMxmBHDFI98ofBolKnc199azFpeq
NC+QdQ0HA2HLx04BwhpbJ5sEsNEwsayKr3jKqd9ue1NB5nZDa4y98MUqKqRwG0x5
hAT7gLp3Q31PAUBC2SpvEjOSolbU6bfwoy6m6fqdtMKlsOr+Z19npkvm8x248NZT
rlktVPzuSBbttQ2HTmfEdQhwB9ux85ps19A1cRamev9b8W8kP0OMdgU7di/awBYw
zGTRmgTSMTb/EbsW2jEtdk2V/LewKr0lQiVH50X9NVU4QiDkPUzY3QycxGpO61dv
0Cn4SCgjtHQFJ89a9tQQ++9uqTaMkUEHxxZPG7G3uxui0H4n5/sTR8xhvm4RSGMD
k+mbZ3JUkMAz/M/R0fq+IF2Hyhw4DiIcY5p1Zg94oTWutPok+UJZPXQ0jN1B0DcY
ht3KtIpsAOdmmFJGS/pV5QAoNBLXaR64v+nZbLO/qBg5loyf3JkzvDvPRQTvjjxH
k84rdDdAKW9Rblg4fdybTMYSPbQVdbMEMDbbVREy1XSab9v0rGZ2FGqzm2Kku57F
iW3zj9oyWSooK9A6aCEoDkx1z8sTsArfjdFxc/h9At4B83kN4W1EzAh2KKDHcgXM
3u/Izibdqgc0m89na1BdMnH7Gh2X4Oo3dX79pX8GyEI29+XJcj+BTERAW1xFin10
wOLGJhcMmkcCqTdQISpIMiaN8CwrJpNc7IKJT6EeNxk0QSYITCY5XjxmevF40W2i
qggR+JwxWz5LgMyzctvL0k07XNoJEFAAS3H/NPenHcVaZOf2gnD/hEXul83T2wD+
5+SNlciPJC5jqWimbps32xheFWCdDH0UxrEo7mN4LQ/eHRqmhy5sNQgbQFmB2vMh
XRyVhXXCjXNbrMtkIl93V94tbm1rWcpKTlSTB8GhsZVA+m7m0Slcy1IW5qq9gUba
GIpqz6OErUv9zrQ9VUwOna/MQ9tRv7+KNWn53Km5ZxA0Wd9gdAIFqfZi/mHpKc38
cgcYfObXQYpBpBx3S4fJod2bFqANJv8DMVyJj5i9wi8ZRzPqxzuwjEXo/t+nm6NL
HbCFKg9M4NC4GCPVpdPM9Yj2YHNKFGy3riIQsxuxAj2F5+cMw0PbPIQsbtyjHSaA
vHtzZxPJ1LpM/e9opOCN7Rj5cSArCNWcjxFuwc6VCTv4W06hnxBC7085e3ns9oAu
b9HH/FwOV2+JKtjSkU5vBEeRk8N/YQsY9tYqE8uYCtc2YGQdNaXkMWijKV2Nj6iL
xUzwYOrlyHFzJwwqFVFl1kXQZwa+3UD7Mzdxp7HqLJKWuK+rs10Hfz1FXRwcuJXv
Zyyx7YVgpLUThLsBvIbZ+ckjjAKccPBrFrbdP2pHrZxns2twOhMSZPN7dpQr/hWE
Vkpn820MJUDZj0FX5eIkPeHy6u1EO6EuiFkHoHJOEW/Dm9ICFtyC49jZ7Z1wT3uT
IHGsDm6SwaX0+wpLDTYxFYbER8WfNzxpb9icZzpcO9NgamE/IdQUvXo+vAAHQtIm
6FalK4iBK9iGFW1/1w+FNuUMDDbVyukLfpxZDaDn3BBHhShNFOGBw+pRmJOAqhAR
Dtdctraolmq3yXS0v8dCTcXFc9E/Ga8y7JFBBcRWtjsHQfMUDVDE9jq3zxeSBE0m
CIzavErvVxsHykaMmem+nsa0ZpjTLgExYDlFeG/xKb0OicVHKNSlRI7I1VV39z+C
iVpGUYNzdYcn/arLe7H3uSzpEXjQYaCOajZ5owXE7YcBMe6vwOjePzkmCOGoooat
coCX/POKkUtGyy2pv7WQgMqx3V1x97J8GLKINUhbIUZ/FqjDkCM06wzMpXvo9NHc
mcnKpI6CgSzz3RUujNDPR7ikcRdF/2LnrcqO9H1W+ANkmIrc/Ou69oCEBCW/Hod1
Qdz6NhjYSTnkx+YzfIYkz7GqUP10OHlvUo9sQHLHqXfWBkdIS4wRa1nCr/Z58WnO
g774Ib6OCpYEM3MRAeIOGdBiI8oQmdhFTzL/LM4OwPHyYFfmwvYWIBq7Cb8faP8W
CTjU2wceUfo4pbXbjNJalALrkTJvKU04zmC0TggbH/CwIILamdi+gco1zvykGCZ2
Z4JJtmvHf17wfnJfNCWjY+xg9O0k2k4ZKa62bBl1ix8VgBz9INQX9E5EqHt/hVby
wMXMFHdz4F7mXSzQMKtukHrU3V3ghDGkBc2EeqRUdepr1nf2Hln5x0QIdu9xfPsC
H92mdPTXpi9OIYr0BQ80CRMPy7BxtmqdpZer1dS/KCPMHaInhr5RPj297X9/hxT3
ENoOWEArAPI1WULGqoQer0lZvc75UmeCGlESLR/iUEJfunm6+DwOtBBngIzOV00e
Z7nFjzAeRNzLC58ng0ag+5rB1g2OcfxELfgVPZr0huNRWxHAwOoRrcsrf9m32tm9
Yjs2glsy93+q3H+dOvYjok82ClIoAjEcFbu1ArFZVeZwhWfs/pxpI2/vMIjht8PH
Y6fS6MY1+KYHcEwFw9YaHmCFA7n3nWAM9DaiBnPugh2YndyC+pOMHvVGndw40q5/
zXNmUbaMUWFeDmVAQA59bLmo+TIAscnbPH0uZh3DN0hWaHVHDNVZhLJzDo7bfIpT
ZAkWW0YJtm974oxigQG6w+qteO5rBGW3qOsXjOWagU8A9JtJuuSltyoHOyWScWhO
/j25Re2ctEeeJRnYnczAs2c11A1eMMD6O6UHFd/cAGgXlBLh/+BJZcJP8DUXcoKi
sQMd05gcaxVg+uB8AHGMeyIou1v3nHdenmEN+8YYj+jJ6sYJ+gKdL479xLASqijk
4DIZbtYSK4DdfUwLm+1RoGInb9Z+Wt7ZXQNem3Z3FxZqDB534g7D4dE+kXFAKG+3
vzGuVbTpFT7eF5QedWEZbQz6PoXDWplzqhOo4Fbd9TJ3PoW+KwB8FDgLQW+X/wWi
9t+VxVK68Vz1FXbhKsMTsneXg34nc2+IRbAH5VS5ZpMuvFpU/DOD6MCkdVOOZly1
wYnaS2D9080sT00FN5Wq71I8yRLoCvYb53IjslQpbuifBABrJYKrsdMT/xLloR53
pjaCMtHGdIs5l+CwY7rVgape+7NgyKIxXGsLTwkNMT/9gqBdbjuRVvo5DwotowYf
sI7Hj6GOlMZnyZRX8XsUqI3xOqnIwIk3Hq0g2tzgsAAayUgU031yDEADU1iEhOZg
tarun+W8+xnCxrk4Ehdf0LLjNMN6hSn3IQuxFXtFSDrkX5Akm4GUdP0o7K53yYvH
xaArMcSnelzLqv1o1+lzEtpFJGpa/gZmtYqTlflDN+Vz98VwUXa5ztvI3VQyWQ+8
L4TqrPlnf8li2O4AeYQB//U1D1zJZftXGVmZi+9s0rZyS/7zJ9sVBH4TJweoaSPK
vZrJBlBbe5slQOhIO/njNaMIdDKLV063Ao9VvYbjjLImlm3UJ+tBaKpBMBAHOUnU
3qeVvAkf+BUhIGLqzA9ZWwjRO0SuC5YVDjOa7paG6SPVxbs4v0BsrXTYKPZ0lhvz
OXFwyQIN9SOYqVjUFiIvdLk4q7KD7YVMNR2JvNQ3VLuCAjLNzAiCxMGwXywSpD18
qLddlOLFI23BnCe2z4PpidkmvhDhIrwOIKU6wQ5cxJN0r5WyHnnH0zhpYVaGH45r
I3NVhP24YqVl5zaeR/X5N5wYjl6N951uprHiBVht/nVxnnGxImz+1BGz/rvf/H/N
jza6FD6UNpqGfCtWHZxK//4XcBJDb1zmpwp9W7vEUyBfTruKlj0Hwz3Oh5+zZ4Sl
2gXQScjtwZ7PgNmv3POcHA4IZ2JsKQ6DHCRAKjObc1GfOCxlt+g5wijNmXNKYPaC
a/+apUzAaOs8/I5fBtf181nHP3Mhhw6gxRZ1lVEhzPjKw/OK0JMwrIhNVxuFhWLV
x6PJreAbujPpnFyKVjenbpld9DwkNnZQnPyo4vLKBiw9kA0PLnRsHNjbHQk0cDOn
5SjlRsTWECjF/QTxoWc8N81lNZiVOwlGf7N8CEhgv+1tDRssklZfnx7QMsQKGGg5
h1aVv27cEpc+VrzA1AxfTJEQKFvF8zL2C/NjjDshdVrLEL4HBCzDc3e4LkoxCnlI
GeqnhQsbTRQfw4Xq1vWtI48vtQqAVnJxwtBzmJg4n9NP7DrD5AuhXxff/KeD0uDd
9vJIWNEsI2IGWdo5+sMK8+t62xAOTrSK/p4Pel2qW8eVm3z4THIUL34y+inCZVLn
RjM0ZmYereIL4dvvlcM0EsfmpE6IniSKHeOQIG4ZSz4N80RUMngiOrBK9WjbWpX2
8AbD5k4TrWrdBwSZu9DhYX2qD9uDBsqmdrk6kAgMMhk9STwXddYFuMjIkr18Auf3
f3wPWMdDagZN4MzZ4eVux/MhDAnUV0mQdDHINXRmyWwbVz6/XvHDR9lFWDQ+oUjM
ErqDdpqUSEpPnjPuHzZNluZc6Ylqdy0CINGlMpF0Caou/W4o8Fw7t7iqNBPZxuci
uSkSlaCGIJC/vby8B2W9Yv7qHL43ho0NEOsnFI3+JzCfPt4WSfsIeNJnPgatSXo1
EIMi4dF2CNWomrxm0W4V5Bdd5W53WRW68ts3S94y9pRm8laHbtjAjz+9gN7xgLxg
xMVVWEhX/3URfKf7kh6vpUWJsaZz+MUQVCnxuExam0YS97bF1sDEXr3mOiVaaBMU
93cjrJtlwXsGcLPgpRgEFZdyqTK2Z1h0P7Hog2fd9Wh2ygrpeyABedLVM7fYofuB
B+WPTuBkgfV9PpqTlfKdduLdW5YLRfsXMg42CtXzaoFr9gKdNZ6Dg2JkFKNcRWii
FE6GDDqZEi73k+J3Hzk9JL2a/KsZrWobD6RLDr4WR3C62oBO1IETao/QUCMEEVic
geujBgVg4DRKsyRLiAjm+cgoQuSIZorjj8XWONKyd5mbBjyOJTe2JXjAtV8dC0WD
0sebRJR+D4cnx/6nq5fvf7uGPvi2FCaOAHZM0a5dcETjuH3lzF+VSkpNdaSJobHx
FFKx3wmK9FmJ4Gc0PM1X3Ry50KvmjDj3t9g1xbWrL1zRRoynR6IZw/15iHObdFgG
/Pz1QegzEHOA3eSXmGDKYm0OVFXIo7xJ4f4T8/uvvlcWyTem6KYuwyX8PLNbULt7
gBKUHRxAWz/H4eZ450ZtZtkZ5gsWU2JgjZ1KRg9gP0LBWxb5Qb/b+p+OrRHO+K61
uKGNPNWe9HlRKavJlBuULPgnp8LvOxSoTAcyfe4rcqgOMAYKW062LHZlADVDvRE9
BgjW7n3l5/0e6s5Tw1CC8BdOy5DhpC54EeeLtAVjtL2FyfHScqwOEA/qEzCefuvF
PBAYmnSToAVVMmzi15CBhRNfbSCXUCkVQt5+4+Of3O9ft5qmS4JT1lTlS/BXKJ9H
4tGKSfQ4anm6tgpso3sKCouETyH8BpKNwff862OHeEkLCnzRbPTRWTs1odcSw/PN
o0dKuvNjf6MhEweyH5lzotLyIustfhfl2xsLPynQWunTm0eFcsJubBHglprLGRGI
5a5XEKISlCnrZewZHFpqQdpvBevPhWztmr5p1/iuztRHBFzJd/BlcU11LTOT5F2O
P4R3/O4AxSmcj0fGV8gp+MQ91KztADVHKaxOBZ3YZfNIS8VIVf7R5rXElKoszNTw
KF7TVd2UsJv7e/tKtgh8GNVCrbvx1UPIvhkzGijFnLBMH1FW9TAEo6Cjo5pIvEoX
FhhSELCKROLmYHnkd5DLSBCfa0xeiV+rH2BleK13aETK1lSfRHie63OI5qgs4SYV
hRGBA8zHNCpnflnLPpMoR1Mv/HZp8thPIHgUF0lRh874clIHYKuu7dpjWtTl5SK1
PHM2fVJhMhzJaU1OI+atlpC7c8NUvdDfnXVnp+py8i7HBNI0/COXNrrcY6BULud8
FUqYGLxp9PBHKQ8WJTm90to6cpQq+Ve10JDf7fOl4ynj6HcATakeHmVuCG09KA7o
ZqsZKWlUz99KHRd8kmO0zv7Lh7xDId+LW+1TMoZFgOlYA68McKsJ/N8foipJMsOI
nXphhmhnBvH1wEiffKS2C6FcdvnbPUB7oS5/yTgMJwLCoqP01B51oUn0GxC6diPd
7wmf6gLWIMFGIG6TAnmmyEPRGI5eP088TDhwIOY6Xkyw2HRSs9SuvqOX4b2qr5JT
BaaSlgvN/pv5owTvOxwaPwTBNa2vV+BRl7DtOwSh2k9FnbXkYIuGZK9fcGNNPGgK
oryMQM39/BGr8qdOmwEmOrWEvyHLRoE6lW+mdojZJa1PPd7NI+07cK1aAARBpJpL
foDqCOF6JGxpxtaEjb5XMskFw7rDRBkZkRyaPPDuuvhwRFq/nsY1IdeM5wyUf4vi
i5uKNULSj4L+5Sp/guftmL+CgK5TG2YemdwMZ7aGpxSaTx0GZuic5R890MYtQrF1
VXhqpN5WIPIHh4OrYOF8+ZilVD6DVqQ7zCBJpMrNGHpH+aHJaI4Mx+OaN5tVh+Xn
pfdmn3hgT4/bj+wmxcwqzUyul9j1XdVL5/64RZbYQzNJfTzBRm2mErR1uTnusmov
h9ourCyjAva2AEwuMWSj8W/vKgwEV/Xk+ly6Z//e8P+bT2lPxcPS9IDZVpP5AOPV
NcSYJEqeOeRx/WJ/5nEfH+j1MWZqAccsBXFhvrJ1nfDG5ziC9E0IhXcX+LQstvEH
TC+v3v6N62WLCrEZhPGfKef1HYUaN6fneN8opr8LcVr8ZKB0hDEaAyYZ7LJrEDAe
llwVSkAmPuexKOWVOsF/+Ms3eXuRloqAL2JWQLai2v8AdyJw0jGL2pdHZZXQNAx4
szdz+a2FgWjqBGi4ihYEUMM7BVN/orcjmJ3rTdoYo4+LZVdfr4AiHUEwVi3eAte4
Jddd6XqRDflSQIpLd3+iUZC5XQUWSgqHR7YxfAKQw5ufR/1JN+pu3eH5ae+9YZKn
Xkw2OxWyGPCufJfOW0A8yujZDfWMyV55Z6H6GS8Er/1QGzQxeoUJj/isHLaLoVUQ
UJzFWGMWF31N/b+KPVy8iATw6ohvDMvJqpr7w/VdHTgH9vJ5esURqD84C48Mf62p
V29GR2DMW5dRRiB+2hieee+82mjesS5h8f1rDLQJV4GfR6QCQRYCH8fDpHzJ5m0P
vokMprq9iIyT7glw8a8jPUqc2ldpLYBGiBeK0kaMvK8LVVtpLPeJmk5pv2q9x0GV
PaZET6qkizZ8/YK744kAdnsI71jySMok4VgUI1kWAYBXjo5pEjchMtWrX2uHSDnH
7x3Fxdm0qvthnkawyjvaJlisYW6Z0rnbDyc3H8wKiduJ5Noc7j8Bp2/3h4oxV+r+
Ve08PfclHdepVsr2Jwf2NWyWJsOiT3mfq1Ygk6zhpsOLXalkEyYrWSiEfU1Bmsjj
tNZUPqOr2xCBtIIq7ixrGkb+lJFL0S0VVYLylaHbrdc8NoExQ3+MUakGXLYql0ZW
l06Bzjp9l+KekcYWE9oXrg81iva0NsAghkRwpW6SlruqE1Qdg09uHPad66akZ3P3
izVUA+tLhicZgZGa1lWbS0xT558Y23uaHtChSi9M8C79fMxaP6Navoy02YEVPRrI
3m61G5rZJVNkC1Det/2za34A04+O9SIJfLvKksfMQLDyafeX7laYOx/7LaLJ6XM0
tEpc4NbVwJ8fec039dlNgO6QDNAQtBt9ahEOWc6eIzT2MRz51jIlRVfPRCF1hLpl
Jrj8AsDpRdZCt8+HGKatUDaR1hlo8LIBobUhkrMxcVKCJ8n3j75nCR5irUh3q5ZU
ozuiXEgaCfZDaR0aH2ysWDbmU2yuUNSar80+7PKPHbM92KlJ8DdqRovStIA82RbQ
Kom2nHQzzgon/cnKpB2d3uSTtQzcQDhN+7YmS5HalEwZY/RkglVmDzgGZ7vMoobj
octFB9pCyJpMdSf+wZ++CrTCm6kUq0QqijbnQ1jIHa4vVnC5B+/zWXWbX3SuXboh
6RiQU4QB+BGhOAFv8VX4f5yVTK3UQVwai01XosELtmawuFU5j6yFfsgmeycdfDB7
20cOH6n5kQtKVAHvV1yAPqYyHrXaH31zK5bFLR9ifFpR9cZDuKRif/5JlQo1XEua
aq0MZIrPzyuFar+cPSfNCjEffsvp8w+JqSWwfMAIwGbOwkbJOiUZHpG/qCE2LJ+b
nNxYaYLsCT9ZoPUk+D59IsL+zrAJEwxI3/Jod0DGbNBXaHRFE4PylwqR055EiuJK
T629nkNiFjOJEkgXKsDjxB5oBqVPIBOS/9RMwgtBdC7oBEVMdFMiKKDn/gotCiHZ
vAw24U84PSiH/bl1vRhlaZmmT/L9ddB3j7fR4sbaTGSCKXrnT//ETGePn88f4xP6
hCGCqFkTSuKa9NjOmu/bbKjp4OUTijRq4JuOXjll96e7BoEbuYJI0E+O9VQEYiiV
bbvOyB+HKGV762hD5C5o4av5lulXnQRXyz1pKl9S/JYGa0yVQnTI9kPB5AVgmcbD
r1svH7XYGhnsgef+1rggi1yrVM3w/6yeaqZf4PH0CiIr+ebKLqwuGCri4n87Z43A
6PNdnFOHxjEkQcpj2aV4kOEktuywuCbpoXMlzyxJXPXEBGTsyRZNS2J+g55VnLQ6
ZDE6qjlXPJ9/z2z5sgeby2jmz7sfKv6G8jB80GOYsYqHeDXOZYwic2cgHxZ3lVCA
gmQiisktG06zED/O9Srn7MSTdqx6LFsIyY2CSC6VXvlMwZYbpbmxOSS7fYD7/+Jk
FP+mV4B1FQo44kKs7bIxbiTq80XbHqz2WLZFxNcpOd85D/xe0BPVmLM60GhJJ0AH
6Nl+EPlWZuNVm+QaJR0bjU8R+kolbRTwSJeBazSLAkpihhN9EqCJLlEIldsGVw2F
lQtn1+9AyA/pTZxGeN1m77CDSYAFZ4y4XYfg3rAhpvjsvoMfqqVpEmaBMRqbvb9z
5E4ZgSZdEBnyvw8LK/oOEFKCD/BpbWAOcHG2LoX7tHaMb2obaw+GIHffOcrH1jUp
PXrFMOHJpy2xbbPIxFrDNHHowQIXuTD5tdjNZwzUHeMlEV285RUuLS2azjMONcPS
KtM5z2anz6QlhNPLwjfoV9xije4jFTLHUePlDIYOjaqFxO6oozKR1loDO0R3mqac
QJWtDzhpHCP0WrEAqqBWhMyQulUnZSIgPz02m2D0BW4qDbPDhcPft7DqToA+dlzq
SJ11dnYNXIrPFmzTH3tBnDALrwN/7LZmC/MHQLZuL2fAer+JTxm6LP9pNG7qe2gG
yseJD/zvadAEuvGcD5+lG9IupnCZ/wen6kgcaJhYDLGTyf+AgJFEaZHu1AGW3AGT
Fts2Q+kzPllNXk7sFX9EhK+WrusySs/GuzLqXU7ZbZxsNdcj0Ub5Jk9I5AONVp57
LsncFlnBum5ylqMbhTZHpwwX/xHxsF8qliFaiWU5MbYzvJeXz4zDm32P4DbPRYLa
p/ytOyTcj4MXs8EsLG2bUzp0le9m2BmyrdLRJ5Aspi2kHfexkLsdOS4NhDFt1fvZ
0dE5G9E85GA59uV2X0s12tCCCpsMI5rveg+XCxxTWKt8uRgx6zbJvZlyptIRrjsN
9chKPmvK/+d+svZ+KcouPVA9W9HOWYTEM7Q7+jf7CBNLjyYjwt558kJKAr40YxHz
lsMjo1sKlX8IHA79vgBgfKKz2LPHJC0uky/3JJc75HQGWAlPd8SnTuhh8g7zChjm
+7ChtwXm1p1WlIhvWyKhhF6tisu7qLAyvMZtTe9bRCVaQTAIGuEAo3m+JErM9/Dz
6YELfGS80cMv58WHLpf/3v+iPwnWYZUEY6kgenNw8fRbGFgbb2VHNYBIRe1Vh6EB
bxqA3AHLKXdNzwll1BaD0NIz2FTneNYZ9jZ0G8xOy8jw7ufAIi5QoBW2OLYXFhEw
a4OTrlb4SN1cqXSGfq3p8JAR0C4HmwYwCPw+NpB1QhGF1swVwld75zb2kZnY1VtC
7ctxUhstMwAEowdMsIgUCF6ShATkyEQvNKhmW2CveB9xHTAGOy5eIPUkuKTdme56
sbIavwYVWvuyio6tHBcbfn6NTffmfTRGMkz6wVhu7lBcHD06YPMHNPFIZu2sr19v
F0tK9hpf1E9oDCmBVR/7KwrwK7Sm7ckbE5pWDDR/qZ/nAkfEq+tk5ylwI6C59esR
1Dclh/niiSSPyln83EOoFM7QWshLS8sE1shyG1gK9mfi0KZ+kOmRlML/9GCwv2zw
XsUk6/upTkZwJF1UV3kZe5XrRWvkJoDMlCmXsW/cgZdzsxZF4KKaFKwQbbaH4i10
J8u+hdS5sW/2obmJptECT6BpHf1OY42vfY1afrudYbkdzGr6yUC1Xn5/94mD8MHf
lSjtlwU6VjI1ttk3wONrOlM8UBIPJv/GrX/kNX/gS0qgxPTf692/q4hGyWpXTiqH
lVA+w1Xtc9IbYwVcCqzQVxH+hssgA4v0whHGc9YbIC7QeV7sAaOSwTocd2K5bv/C
R9n+risjNbuMqKjMCaISJtHPlVVzLaNDBgShWAP7Ab9V31PUyv/kx1EVGplWucaV
LPvu4yThybARWYtLfOnLiP+vzhaWlBejC1J/wyXLZmnq0yv+eUvUObnR+T7g4nra
ZvVrsYOnEwIh5eiltwQsPYUoVO0kb8FtFyltgq0TKY0O86WuRIzU8++DkIdeKS++
jERlyI6wFGkgu81j7WzktfHjvGE+oyZaQeV1Ry0F2HHydbCdwtQOv+5UjdM+Ltu+
DxzDJDkuA8/dt91JOoprVCLapewc4y1VrffM9dtaRJsQAGIbP6cvQm8pu5ZsD54k
I02NhRJSgKjF1UuFfPK8JYvx+HldJ+oL8+MIgXx4fck42eAyUaSKIHSYi6MfI6xN
CWnQj3oPed2B2Xo5WryyT0MemTkVtv5VibHN0Vs22IIscj7G77BUN8w9GZwOtaLZ
6XklH7zKPM8YPzXEP0CPFojv7x3j4sVtm1ALh6Tq2yRZWHiI7UGTemRYQDXKPUR2
GumUCb0wnVeEPtpjs+SdjcwD/SqDn3vkQ5rLM1tQXU9VGMC7p9zxhdGKUrnI5p7k
NIZwTWBWQJSel5QLKxhrwA5bRyp8g+TMtJBes2DOtcEFcPPi5W5YfmCjPP2SCTdz
6EHVp3r59C7OBgIEqhtplZQKIuEKIqiOsilYc0y0V4cuysfi5vIqJP1OuKYN8Ak1
N9bQujDp6rrJINP+1C40plLQed4QQa7wWTmDwX5seKfhURNUPiZfzWatmZdEtC6S
r9kUfUa3Pvff8Cqji64FzpWdDymTOgXF4WFjCRpEcyjsQWtasKoeXZedVmD8y40W
5c0SyPwjDmdjjFrJQc2qmtaY/Ad5U6x5GKJYHxC+dz55l5weiVw88lNV+UEnDR7Q
3BAPLg8/UeeJ8CycY1TwxhModLf+UAZ8fDONDYcAGtJOQTlQeUwpBkcTN5LoheNd
fb0WjcmYpyjwyKP0ZwMxj0uESUPia6BpC97Xv63yZbEeqnmx9ps7W62g2t48MbVe
bZIRTCVF61RTmK0/ZUR4gCCwmUjZu0LtZuGxpSN7HZG0FuZwzk0ng6HU+ataPp/v
Cr12+w/eGGmsBjTBGZ3Y5o6sWxKmPDAP84VOfvmBFi0uppgYKenDbZvpBHe+kozQ
R7VwhvKg0tAFpL+wIftOKDg/kgVU2XLa151RB5d8yIpNlata5ptG6FeP2o57KUgE
yJlE5JopI2qVEQqj9M31882PwZXqjYv4qQwqvpMTbcNSfuZHmp57ZXR5dMPTsXKq
uBfjI6Xw34EBiXzmi7B2TWtxQTh/BFMyUyI+e3NU7DGf2g8lK9Jo42ZZn+WT5tD4
X2tehX+ao5oZBEo11bi7GYdeABmHjHF8CRey5RnKQt4NjOOMTCk5CpkHAq+Pb41f
IsE5+khx/BQIHTn8t3haxEtff3i8e0xAAr2njlwg/oSV1M2kIb6PsZJdGeaBMyQw
yo7JA7HbEzOZqsVUA2x/WjD8GlRClrNZL5E4fjls1VvCih2BzCdmfPDGffJd3FF/
nEAKAXlGmPhXZ9Pm6GA/poKI/4I3sYw0lcAVtnj8TWdUZSjlnN70vriqH4IY/6TJ
1WlA4ejO8A/0Fc3C9jiIOnvi37YIjVldTwDbGPYyxiOTu8n9tgOk+vd3eQ5kOG5z
8OtUhMqi69bfCFUfu8Bl5n6ocEQuIDLdNumRbKX4If9QGIgwcHWbDYMkNxKGu2qw
PJqRPt9t5muBkRWdBjNtW9BKRvKBaZAFzMIClimVh1YcIoxbFVFQFoNlbyeu+K/y
832xQhjtKrj7FqEK97p63wlidv2nF0g/kGfy7HDLLuv4phtAIm2hWBKwWjRSqRFh
Xt/aKAZk802/R3XVsfwAcs8BaeMqCswKlilkKJR9UoSz/cVzi47irSqs09rlCEVH
qBGwua6A3vupLnpG4T5/vQYArByNUmfK3q05OO49sUo/FDxyPFlL2NlZcbqMNcYL
d8oYDS+a1L+HeVa9vtD2veeUZBM2u8w7vU5hh3M9ng/K1nnu8uIH81WGgSCxiq97
P5qJom3ies6wJ+4FhfYUv6KOulW0F62jH7AsdFFxxsjGz/yKGZTNYceSLQwj97iN
TIRCNx/za9cOw6dRFSiQh3Lv5taOZM6smDKSPkgQ/mHZUatJkxP3LlIG6iC/fn83
J51hnZhxXM/OYvb78kxNRcRXBnS6/yNk6BF0wFdkFM8gnbv6UDOjZ5kaUHHBTkK/
nOGR0mGGZaWPQx/O7QR5ZMxB1TqRs1TIgb5sgmZuJ0BAxYdb3nM85uY9CxxOJgga
aHCSXPLy+HS4sswi+NxLCXQfgWUE5uwRI6V4oYbQnDOjryVT9i2DUeTa6GGYz1FI
TOOJ+Ve8avuKrKE3JvTTFD6QT3QsgSdkIIvZQ+v45ThjxCKCMzja+bqncTsL0j0E
UNcv/zlLZbcvUkSjr8O7m9BD8VPZ0aECKlEynpMArN5hZ8ZkZyuGayjH0nvn+Xc+
NmEUlYLwzt0RRjckiFDeAZhHom9KF9VxyXMBnZs9szOdfTBdoe/96XIl9B6Iv2m5
K0krEh/E5zjkeJ/6CAcxTxW5QSWrBZk09ZyPu8s4qYvCfeumsPZHz0XxFfZikyO3
zcWeDSCzWhuh6X1KsnEHTQfSdnn62fUlZjiCPbQiNrpJJSn9I7lZlRd2Kvdj+hyE
0luoJ+9NZh9inwZj4B1TcxIFD31GXchStwPFe2e9ak8Xc5YWEkdc6aHMRPmqREid
K2CxfQxNw5T3DL9iDEHvUCspW6EkHRCDuKnAsypGwx96XlpZShLo0hmn1nUlLty1
LKC49N8stBaHNpOVTs74AXA3Ed4JmfxOz65xsDRLb09EicfygCGRWV1Y0T9lDfwp
AcnRvdZrR8Dp2mQ0LYC6R1TcxKgd8PsytKgwaCjp578u9Fu1FWACVbgzA9yCuSh4
hplnh/407sjDWJYkiTrWHIm4mfPBRC8hT5ksc1kUytolo9i7ormTT8oGXRjNWvRt
W6eyDqNh4vFXnX42HPkDdqG4lgfT01ueDq6siJAmP5eVMS9eVt6olGOriZXwZNT0
VUtKQWqD4zlvPAUHlmyRb3BWH33BC+/xGLtKPeX/jU/unEK84ihsEoT+GuJ7B+vL
0zmQZH+T9EtBcNkTbZCJvIm5iDraGRUjZ5sG6XwyabHV7xBvKGqDMLW8FvxwCR6p
C/V+JqDTIccJoIFrqGgRgIsmzRy/90grPY7X1e1XRYsiMROkVYNGPNgovlB3UxsR
OtTHYG/0Zd18RI79WZB6Iu3eLsmfAGCTIFPhyKytVA1UBevS2ve3rNFAAJDj2vb+
GM0244kH1hJPXCmj2VWyyPHK0FT+dcdT/Q5WFyCAplT98KqCxkS4rIdRdSoeMJhn
yTUW2Nwz3x4b8sFo+H50OZ/BYpP0cyLGqndnlnSamLYufe4a8yw1MRhMOmiBWJ6F
mWQ5E2aWNwR7MCJorNWrABymrz6cL2Jc72HiR9Jr/ElBkWft3KWud2TQ7sGEcqMR
lj2i6t2pRmIMFQNLxjJUGIhWnlXW3u46gTrv+5FxdHY4Yb2WNT52bzG4cjHPldhU
XXatLzSuiE2GZl+TMjL9vO5paqB1QoS6v4U3VGcDLuM/V65KpmtZaH0NMDFQFG5G
btpKKkboYrKIqv3THdetsQwlx9JWc8SzjOib7wKGFo2R8WIdLY1yI0uZ5OSvcHd7
6vlSziHaVhK85aT3b3Lvpuu73qGC07/TBd5YIz+LIcqbukV7Uvx/4kdoX6jP9iib
Z0l+FS0N9/S0cO51j5vVpZZ/93y9YbOWIL6oEA4U5IbJH09WHk2gMfzROi2zs5iG
q5YzK7NaGE4UF0LVnebj5WQvO6bXIWDf5IbzZRUrSOz9YOEYjTFUT8G6BLarLRn+
x0PlqjUqwbu9VnSDgY3lQHXaBJACLbtzzjq6wrLZn51PQ7Ql5hAHv5oT69s8AMqQ
1/e9ELmw+AlVe75LS+H1+546aFgJB0d52Y3Pn6P7mloeuyfW2AGdKvuJZl/pD/N1
saLE0LcgMiM74iJnPj1KXlJ/AxDCQ/0RYklCBCzCDu+XKbxjO/cM7FJeSeGJQbqe
Vp9cGpKPfDYIhZ88gphlO47QIUF1kEwt0o0Vh+fX/6GIZiMIaaNdbrtJQClxYc6+
Ibz/OuYi4nht0P+TcJVZQlHOi2P5uje5aQaS/1zW0pEKLysdK4iBgG6OhS7oeGHB
QWPzCIJt6t/+cVn6YwJgBz2+9zfIU+9xKq8bggITpw1JZTVaKY/y/x2mBsMAupbr
CZDIGUmx7jwG/rnqlaWA4p2b9ZfEVZ4gv+PNf3+V/ETGJiteSldNmE+EocigGLK2
E3lrim+SPKi8MfNrFwTcsx54gQEjJFiY8hJbq+lEHqZhX1DbEnSyjeshOs3wuEox
URLKE8yrYSQlA2c0yDWvLP3CpW/CUk5jiy1f7s3aI9whuh1f1KXwNGKdGSvazS9W
2+94smq0nhdchxlLxa6uKpxQS+FfOrlROv2MCUVNonA34DeT76AEy+W2XeGefprB
NyRy1WDmA0vB6fKdglWW5u4gCuVk5yrHESRKprbPjovWn0dDQPyp2PjG6GDcvIxI
5jVQBapSXPgYD3sMslq5RYZk467RDM+0nVXos93dL7QoB9JP3SISon9SJfzpSwiN
u/3FaqTIbYsgaUa/kJ/kinRN77I04slMgiKA2huNrJ6FsrDjM3xGvi3bbvmOYFyO
e3xHLX7hlDChZQX58EfHY7a3NkmM7242YT2xptVAl17V5FMv3d8xCGAxrPpjJ4gk
/vsdDpwBKRIgTvC7rtLg5QfVsDoqo5ilNr/BMq1A3HpyMBEelQtfbTExOa2d4Zgn
EU1PxNywoy/S5Qfqc+VfEmmLSmfoBFn1K8jKPz5KHciaZ94rj96b1zLIn4VaYVXE
uawhAwNrLRtK1dmRwGD707508bK0ldKJVmVVuKBGPLT+l0+R4rBn8hS+dDDA0YkX
vvp0cZoKkWnQa/HEh03YYeXbfO/DmYe5+e+bXb38F695AtJ9NoxE+gs/q4NFxHTE
+KnFv0y/hE52cXF+Il75vVpnpvvFqWoRjUOHgPCaEIyKxnSCVZbDqrLx6Tah/XNi
R8X/NsqV1tRVQt3A8oaUq5yEkSRraEbpQur0FRIkzqanEUvxM1jlUPdAbQb/4E8P
0U+UsrTYb66Fk3hFHEmjxrJq01ZKzhNN+ypxwu1YXVn8OmaakDuMDC8SCRSW4rOm
YYUerHUPU+baJbEA/mYQw1MkuGh2nfGyIbruO/qcsh0ucj91/jw+4+m/Q80LhEZV
LcC1Y02NXneKPQhdJ57aDRNZvTjx9jLylUHrxhd9F6TXkZ1U3EHKMMdgldesY1eJ
rwlWTxHS/fu0OI0UMl0YT3EzwnQOtdB7HPSwPUzX09DS6HeKxa4APcH6IDyog5uV
zrWzlg3n4XkTm6DRfePwKmBC2ZbbjrzP04lIh3sfazqFPDWfg4up9Y9ls69JPiMh
kzIWvIhxc4TkQXYBnlljNMFs0wW5kLyapD6WJsURdMEKiqdxonX89r3HLARZpqK8
L5L5/8FrEhkwKo73/yhofAJ//6YcCNe8hvbeVuDT7R0GFzrd4aN3iOznoFvlmLlV
GTwnqCGqfz2Gr+8aqecB+LnYuYnrspd8t6kWKzen4nV6XnFdHvjQdRdTra1wnJHw
maav+6EaL8wFLVwRDZTkHyUksx27mNNHoQ3KKtBkLHY4GLlkRAaCeBsHHz4R2Boy
q+V+NOVVYGkP80jUePdoiITE2hnXGLczXc/a60wtOAAcOSFeiyzZbyw0Y2+7t3fI
zb5zcQOSt3jSqhA45/8ah3i9KNL1QsI+NLp8AhmNh3gqJ4vmNHuhUIIOLY/PtRv6
BXa3TYKXZHFFjh+31oc6tsSH9TRs7LvHjdf/ZzrPxW1RYmWZdVloCb8cjSQcNT1b
7u6wbtqYn83QWmox4QGxexXziMqS6d/PlWFeyl3IEpQsitCXUjMmLRDF1p5K+N/c
RzfcQpOfZZfF04m8wBLDw0+F1VmhjZGrKpjRaT6GegbNCItAwzYyCJfPBh5sL/k2
rTv6Bq4fq4Nm39OhEOTdpmXgP0ochRyG2yw+oCVtb7CTpjCSTxI7RRF648vx+mlK
iUg1la1820/T1BJgSyVSK17Eh/AwhFhsGAMeMsy68uNJYCUKAjfkZIhQO8ni/pfJ
nN4JFxyYqUcSEJBOPsh1w1v7mRKI+D0tJcKVXRja5tLlAeYi7wy6DtEzA7KLB9+w
R+YxaRR63Po6lNlR6RjP4+IPYtr8kr4sh/loH1NmZloTU1COctZcfRIt2r3k3iJr
rZ/A5+tAgxkelg9EXOA6vXle5xygOSSVPbLIS/9p0ws/C4LtrKf2FGm1dn0jFaKB
bOWkFmynyhWVdPY9Q/E+6J6spXeJq8AvdLa9vl1TJQR82zTikx6K8Ae25VxF4Syi
K97HfhF2xp5BQbi1SrWUhCYNKtGCZcwGTWOJzG2GJ6QR6eAzGjfuZqSAdgQ+dXGX
HOeh4tTiIvijUlYts5KMAtZxPTV4+RL7suTCcxptdRQX1zk0IfNrk10rRByAuq81
98bVte4p9fmnlwR1XuK8+v3ZCMTcNHzo+uQt4ztKP5ipKD0Cf0BsI9yPaBgnMNxz
uROFw3MpazrzvBzPtXPkcLyBFpT0U+lJILuge2QfiBTTpcVrUTN662kT7MLJftns
wBf693gNxloR1w6pOurtQzuBAgRfeG7Uzyonb9TWAMknTsD2EA50fSprpU/rA16h
6trOEctBMVuh+/wLK8uLBIYcYhqRt5p8gU9i+SplW4wSz9jV0sZNFlMKhZvqXSh9
zYsn+p0kayijRMefwuqTps12wp9cS4dVWy20dI5Le+wjmDIRX22V5dsw4kLouZXk
4+/ZlQfsPCrhlUc4L5EQYM2EBLksXJvdYElntJ+8xQESBCyoyVCabhSJjgWXUn6W
cLmkwFwkfvOXeNnww8fvMgttPbm0KI/ZMd0V/YQEWlrBV0pu95DtFMchUMvyfX0S
z5OszRumpDprS74QzT0TB1Q07xar0fC4+MQ+s6xepMWcJ/9TKIyEh8INh8/fwjPr
gVEdZNHB6ZZ9gaLFJUY+8voF83Gn5gQMMc12xlUhp7DaP4yCmyBXqxrClStLnlQ1
nGDgher1nMuHC3c2TzEeBD/RFG3R/aa27kjF3KhVKA/tnVvQSWL7xPYTxp7QRDoK
r7ahWJeVCpzlOoAgik6VBXOS6H9Km50VUCnwurvpKTKQ+XQuieBQsNCREkjTQ+jz
0fs8+maM8nRxHgaex51hEuf0Du+xn6d6eSca6DjiEegDBMfVsShHJ5nsd3IWFE6J
Qi4ET2mVRbB3qRRhCEnYeeBb0fmcxIzg67bYkHBQKcFcXaTFkj43kk0656RDTTyS
QMZkLozMsT3oeD4sFBYS2foiYpmEwTcy5C24USlflXMCtI9qrxC7r3xWcJF8axuY
R8eIGwoPiMee4t8BgsYcZO9Qb4LmVQHjqg6fZ9YDfqvN++P9tDrfrLYIrOkHL9eL
ZnLUjQAAu38gucvZxCKypG62KiiqHoQat1U4X7fqkTksD9p5AmVf2YDDNrSOTvpe
5+QkWgSyj6QHSfNqFtB4zts6xvvnPkLwBZOsVVaEJtngauve27P/7Mym32MccQ8C
HIOGKwG68ciRGVfCyxGjRdgC1PJvzeStDAsLULvnjHpjAV96m46kPYYUMrq1qToK
EKnlHXoSeJP99ijIR4fPYOKA4+cVC+meGzeJJrw5cE9eis9og2t1E1ioj1Lknmx6
TR+nRV6fWUDssM8XX2YdaSMkb/X9sa2o30Y+Mv9KXr0r/ygt5ASdWo4KUR3bdgWd
hokIy3Pd5r0KM6wc7+8feTpR7dTT3ATVXm7n4LByRW9MHxyip20xkbe3CQGqNOpP
hsHKjCSpqEvpuP/uGOpJANGfy3Xwbab0Tg/7BwODcdhcojO3gVaYhee+IHjLxktH
4KoGH/6cb7VFRxfkfwttbyg/r0bi0JtaVL6cnlTR32+PP9AnYsjuZwdclQgdOaqq
uMK9W/i+F7RUCtH8CVmNfyusj+dCQPBCG/pJc8AEcJZk0HCklPYImcjQPckRn0Mz
TU1cXb7+uDJUPRQooc5lDTrxa9MCU8MV5euy1O3fxinrLhIHlcQYZHZjGTaa/JQM
aLBPwgyerUmlEkJ3W19NGEt8yrUx6oKWXZbNcsk+B6BAa7yKfY7yF0ByxX7dImjz
D3fWkvhdjkSmYVwTNCAOq4s9gDvYkY5WdMkBG9mMTlVkTRbWPQTa2l3cujfvhC7I
+FB8GpPcNBPdHW+hZpz3mn8/tPRMbHxbuSMngeswdNlZcU6ZZ2cXPuw7VgoVPuZe
iibo7EjoMT+3Bd7ekn93wQ3GIDX1FBAlW1JBPUGQN2WUSH/uId+MWaR1n5ZxvqnU
d94/QKIm1UlZQgs6b50Sl9uANdHzLm0VqCofTc0fvRBo/bmZu2soQgjtbM9eqymO
Ps5XE+cNyMPjeSpevZQeNjKJQid6rMSE9p939TvA6VEMJ0YzeY2lS7na0qSMHg9E
n4kE+xdByR6N7VM3ph+eGtW94ldZvYSm3EAlEqw6HSQWjE2RrHtWBehE/EdFNx5y
Wb0oA2tqKJos68gEV1njYhGX2RL6ESzVU8JSKnc0PCzj2PjUee9R+1NU6QuxdsvI
65RSqaZc6j51Rj7+/Jbw9vYXjmgYN1l1un17g2UefMlfY8156IyPB+tZurGRoQ41
efPBOnpsXpibWM03EQIqlVlcMKx5IxfIKk+uppYVMLV4pStRIe03xIE5A4DSKYGu
mWMu/COcl5zC9fwBNwTGXdqsssU2oRJtGGJ/ZWlGtT+kIQzGMjUFPP9eFINTbFFs
xdBsQ5F79N7OQmhoBPPiGUFq9ZLi3tEcARBWQKhJoklZC/iqCpe0AbpTgqlqvZRp
TgO/nA2+2tVqy95yItmaATCifCbMDmiQTHH8Aq8hSlEx8DYSpL+zN+5cs4xQ2qve
61CfPHJ1qIEq8b/aKXpTqBZCTYneL88Cy/Lx434RCecPhbGHSWpXWbMeSUwmoPvs
pvcDzBIsHNpXj+Xy6pajKkZG9aNjSQx2zurs3Vkveo8S5bTHkP0uNXCc3sp5oBq3
GR2t0V3XYpQU8pWbEKQM767GOqxDIsdfomepTn2hz6Z8GewblvUadxmr0jo8WlZM
SYfvhTOD63YUs5AbYeOaLCUnTrrzh5wHJ1oNgbgB/y33Hs16VTEStqoDOS2XhYbz
7rd2XeZlsZr5OeJU+1i8Ae7+rXWXpZ7UX5ulcFN2S1I5GhxxZc4skw2sPtshRDpK
h+FLZDB0pmTm0cvdwLxrZKpvwmER2p+uycwHwbNrS8k2pdet2IG4nvVZOOfEd58V
zAXvzsIdNVxr+zQBguvrz38Ut/cZb3kNfa8Lhf2Ej2y4cOzIZfoLAJ80lfceMlBO
Jt1vkcmoUunoQCrMOHgm2H6ihkihYZzFSWtmNhchTOHODpohZHY1b86ntmBPTl9p
gqZ2Q4UXMk7+5RVHgRVEH/YTjdNo/DVTAHQ/hl/4VlkHTs+VRf+rfoY2JNT/uaSn
NtsgXbcmfc1dS2ICdq75Cl6+wjNE+d42+1BNk7wmtZiW0j+QRkO2rVruvj1T+BPh
G4fjVP2hW7QD5lsIfgiDIKwZ/k7KsYdTULMgx6ld6NFHOY3kzpX0K2Hz6rkbwSkU
+D33GHbvfHtZ+8hlc6NwpoWPKGwBmRuL8qKOGuqDCLWIRfBrgYvRvi1JvAYFGmBy
eE1rT6cZWS1Nh2sN3dNQucz2xDYXXhYhOa9elouHjKPn1kGmUuSqXnYDPXBnWiI/
ltcrhujl8jHBjZA4Q9QoV7LzJ29F4JYWcb9RyN826QQsZ+poJ64i4uTkLO8DGC1S
EojogJa2B8QDw88mp+etsqkwaGVUBO9UqfzQFzSLxjpole123Zo0uewngs3yuS+G
kXFtqgrLN8lkxe1VRZtiyLnPsia9VD3hozS05J+ssoy9DVZ6+kMXjA4et6GLBULu
Ox1Gti0S6y0gPoYUnq3BuhAw2oGvwRk55BDhzAo6jhRTzkEpKPfShrumB0sEUpwr
rSRBTkE19WkTiT03muXTORZ3NphCaWZ0Uo7CeDyTsN4qdCZa0omIajIgTjjU1ZXc
hl4wSUpzwGpHY8KVGtmvhnG106fTkkdUVZf/+EUyOt9vODVa+gDLEjVa7smnjlLE
m90/TfFM6UtLV0Q+KoR2nt+v2SGtwNkXD2C/t2efm3t26epJq6uV4nrmJtk4X8Kd
90kh7dp/2M7XNxn8KbpgvWyEcfCxrPAUSad9urRz6u7ktUWL/Uibw+vaPmiyQ9Mb
X3ygGA9MtbC35KSMGXpp3VN0Xk1UmhgcF1DZNzB2zoi6pDPBDPSsbZlzp8puJ+mq
yUY69nsrWfhLShoNLJFtLePLokV/yF78TVyBzQZs+ZwwUjYKn2VMAA1dkzLMNoIF
Ljos0BsRc8/Qbo9eq22sV8u03PC0JFQWbP9x8xsIim6I8i/7bCPOitdMljHQrhAS
PsQdmF46qXxss/ljdWlaaoJlroMOW0IGewuL+dUtqgTLls2D7u8vvsXZm2tppX3e
ycvS8Zj4Be9R94orImSdoRa3RPD8olHfl3x1qpW5n3lxZGkhJw7o58sUdBYDI7Dq
T4cp7W26Qf+C9zgXeH32xDlDcFGb88+MqE6hAaduQEe4k/Mq23PEUB7stlhmirMd
j1hQPHIZ84TLTjPmOOd6yGs2GgP8W5PQQNl/B5SyzESEts5yrmVmyyBBM+RVAyel
M/JDhlQ2g5OMSe6aDAhae7ruIRemPHltlpRRNyvxy0VJfgWOvUjBbXpQIqttFarj
pAzLXCAS9VXzNuAChzT0HJhmgm9mbGrZsIv1QRKpqBAZIRU0+d+BF7MUAYyjA9qt
i/h7iyQbD26YNnLDyerCoflQG0DVv/GBYPTiZOJwxhMGb+RYWkZTuG+rO90fJIr6
d08wNgW2uFzjOQwWki7JJoMKhG5FOGN+CLH8aDOY/LuU81zRZ2tfcc+vcUtLaDI7
Yn/rsVUBrojPnUL+CqY0/94mfsuD9NwuYcXb3NCjkk4VyoUHAZKzjYI6DtgdhuLR
bkO+burz5Cnz2pCDUx87fDZwIbm7EU1eR3XGjLGz1fYemr6hKDbs4Z4m2VFYcwH2
sqG7Ai5UiK/xLmnlGf2PngoQKd/VteHRlYQoe4ts0cGpAx2lfbuayVbZbP5kKLrk
XLfFuu7JJjs0MApcl0osdcCDzYlTPOMHVca66YwdtP8PoSuXno7YYF8R63gcKqGC
hKmiKRiJv76+qv4EYH2tyLyICbQFPTd1W9pRAaAXw+RBmf7Ynx5KFLEfHXyLXWPk
DbpxV9kQedw2ExC4AYQrFB5bnVbTypgtbkasaCCiuAxyjPfGEkyxTjowZP5YTXjn
kC4NF+U5JjWJyiijPNoSvvHM3W4kCRpL0QKbMQG/xfsOGm8ZHVBYlodEWXVrBw02
5Z9WtKy7tTrGWDzQg3c+FaIg//ISGtbgGRCt56/Fat0r/v4mtvtQug6Ow6LAJ4ez
L6W3KpVXRPfi8LPPsS5AARn2hzmXtgZ/MiWA7j643DE7HkCYAuLqgDXWOkadjOBY
CiNPvCX7sZFxT3xnVStda2s1cfBG+0uHijpUraatCKjES+TxSm9S5gLdxcphV7W1
UZTDKK9DKJyddMuh34f5APK3KSMoEx60whNMHPyZwG5zjzl/nnefFBs6y9soK4vc
u9MrUEUYeUuzMhDkSpxx6+kdko6DB0UoP9sb5zjkNf0u8/sIK7+Nt54lVj0NdGDU
JZRdp1I028HF8xfwBeqDgfbRUUAGVAanuf2SRh/KSrayh5uRlgPphPY03ny3ngUK
Qw8vPYB3aM6droTuxOpGi6JY9Fq8Mjv8qcHfqTz484zh9Jz3AxNjuL1/KTgNgjxZ
PiqBEi9a9Ipv+KLIlOPaiAGrH435gTA/LOS2bPV7WU4WbVgf15ywkerqzqA9wqeS
IpIzYDQPOWK//5/EFZeik41Gt+/Y+Zn6mlMDmmd/fsMAoe6ANaDKgF/vMdQkQJSE
c2I4JITUX/MJKolt4PJ5cuADcAm625caG4SAa82jVKoCAl31FyZM8eIT9LC/ZOHT
LbC3SqPakHIRsfvj52uDZCwFX9YRjBRQNk1ziISoSi697JuEqbOoHbweBS7suai3
5BpJ87w48zFCVT+rY3UhFu/iqoPGQhtxu2q0KplbDCl0z02rOEKFoMUf2dBXW25w
14WenOOSVXWvfoEPrqJnMq//P7fzEoQbebBhJWabb6AlvWu0oFKURMUvn2pltXWp
mCJQIFOoo+svpRJUFeYCuDJxaakJs7YSjdBMy1408Z0Vq/Emg8RZ2lNjWRHM4Xsj
n4jrTWWyBbb58K6YusZJxfDEt8eO3nlve/1lZ6nGnvCmnX23eduMOV3frEm42Ccc
6p6KxAlkmzcgQLwzI8gwCBJN+3MZ1CRNgnggKUTYm0FlpFOzUlJxciexENPhhE5F
awzufoXVHoigTGvL+Yz9Te0EFglOMepCXCMzbSlIxvPoIu1m1x5P9ENzoV47dlsg
QYVQZUOq0JiVJqLupTYNIphF8zNZ6PHZjs+Jhb7TGpAKC6HzRFFDPtXN72HEtocN
i8ZAWgcLJcNuHWS+wzHWbFWRojQm8PAEPAh11ahYWt21q7PbicdS0A3IIFJYBR+G
5GE4AL/oMbR+MauL67TEo161X8MTWJ6q7Y7kPbM9ugWPOz79a8YMeEVj65jImsEq
0Bhd8w9cXLzqiWgVekuuROOnExUW4uy0Du0KqyOutw5M43uAqPc40SXt3yoy7qd7
qvJiQ1uVakab8Ubb0ZCc7B3oJWaam/vEyqIioWXgn9K/lgZrvpGfQKzt2drEyzpz
jjzoOnApSBLcsJ3LUYX5v+6CZ+Gqg6CU3h/fcLrNqXNPSpiABQeKkKCIq3hT9ArJ
le1r9yFsAfiEGQxDEoY7KgfXNupde3EHWty2M6WUwuR5iDoIztWBVpMRGseLGvcF
s7jhNXnKZ1OUGr3F16GtUIZ/o8WAjxYtwl8XoA3KQFmyZvBmtHoOy6GJUI3y0Grz
LPxyO++ou/x9T+ohtcmsrJQ8TOHC+U3FE5Hcuka6p/sC8y9LvI/8A2jXqyc3CI2O
CX37e+Lok5/bMHehIiB/c9rw710Q5NevYfx+AK3zGk6BfJXoCU3CNYfUthitCVoK
5u2N2PRC3MiKGAGsFHYsnxG1r3pGmVG/k5Y14fDBac+SPA0H0+vq/liKBcytHQyo
YCtN0iPNDGUF4ep1gObWCBoiqH0vGnvUZ25D1pyKWJENLeSskvrbRYnTHex78ZON
0YFRWddf72WhvpTQVq10cA4VJy5m5kZX+kro3HWZL02aqMYPZ0pQaX6DSwnKac7u
x1jL5k9BrHBjMfIdW/mVzf84KRQmbxX7RleQerDEAUFLWh5OZuylVM0Krkm+ywp7
7SJijypTd0Nq4ZyJIoFgt0cAXB63VDmRYTI3fdMB7YQb3xYW0AnCqL3+5YA5//Zi
CA7jhIK5w6McbVBNn1KYc0SDcT9k4ZjgQ3f4bTAVZ4jUxM0HrtkauFenSMtY7LGg
Q4M9bXUijD/IZAxjFYOXINNG8WmyY8OBhYAJny1Qpimb0V0oqDdF4jsxM2L0Y+QI
St1VHuv5OlgtyOURcLbIqhrpaY3CUNbZrnMxq47zlppGoJu0OksKRh+3mllq5l2S
/jbgVVm3LnNhOnmdsTYcww3ximBeC/QhW2qRHdOi1DsWfL6NwdXwvvsJHO9Umg7C
2JsWhrEt5ZhyPYSmm2XYCy1u5aqA3ZNYly4Ba8GKK3G6xO/qJOmCFwXPXjrOInyC
B7ahCRpi6ZviBsMgR3vqmdMg7w2iWFDMEjTQsZHbfJC7Gy8JB5lmJvz75+w/wUFb
glTrs4GTdv1Z8f8WnhzSnc6sVe+IUcDQdIi9BfnUbRXVjg4Xng+qC7HqjeeAqyz3
ceSrkfCSdXrY6oDxKhGVTAqBhh7aIZzwTOeRqm0lS2RBbJc0UekNmeupuiKrSX7i
CvreUIxXlJwGdf0NzboCTG/IjzFnPoZJCjx+BnJ0j9cDlTv5N+mgzM0HUShsnbDF
kr8bWhSekocv19W1YOjJivvYSfXuqVRDrSe7CLdH+Pz5Bw00zCtBt5hhqcAWZpD3
hZBRsBh4GQreBr/RFWTMlRiknz8McdZbIyY8VOe3JHFX6KqAYsgAyw3gV0npZZPw
yZMNT+DoWkjZyJyHGBZcQcBTjBnU5M/a8ky01uHtHEUr/b+9udNP464c30IY7O6p
9jKJtutn0YG/F0UthsEc0DhfkeTAJ3b3RoJnjgXTtM8kBB0xpqK3YTJMyGQ3e04G
R/+JUJJarww8Q9N7UWYeu2zfqT4cXcQ/asiKD8DyhI1v9PQinB1dow5nRnFvGmbq
U4EXO77m+7SaFrKnf/OoVzS57+CiKKJLfU7zza7/vFZ3EifKoJch/9cEdkHIcO/X
DhExr6rNM8FLO1v+e3rdBL4LG/Wio/fzONw1WvR09bylRbI5m1OxpVn6q8j07p0u
WvB4ZtnLHz3bWqC1H/sp8pBPdeca0xtFTytc1UDB+Ayyz5MgcKXtRY5utwBz12cS
jWEML3Pzsfurc5P9IOReMMqJwFUWxNsZeFXd5B8R+6rS/DZLD1fFkYYIWfB0oSdy
Wf/U25hs8FpXNUPT/UAwYR961B+z+oMRoX3NKhvVzMotqlyxQdy7m8+Nq5BB4CvR
RsMBXR/wIV+kjs+l+/3W0w0HLex5Ns+CfKhYWU6Qm+3b88W0CUEtxziGOF95Gsjy
rMAHHHxDG9MMH1cZd3l4msmf9jieWX6AG9gyAqgW6voMBE9NrA0H/Fl6wmToTFiz
HDY8SoOaaz/TjoiwBilokds3EYNZiSICCG7nxz4lh3HXBtbJryAuE0LWvibocfSI
ObEeZ92+vCJuiOPHX4/mJsNh3C9Wq5G119RzL1+PP7I/rhlrZCCK3GJk7UNn1hOz
FytCYeTqaKKDNhaTyy7zvmAKVBg3oK4fNoa3KAa55n+rhVFHv8I5n+puAiPvlRzo
D27TlGzhKp9QS1l3SpKU1GhaA42AJi9eLuogCL18y6HBDd7Sa451fWh09s3XynoV
sy4xTm8Mbb0q3ZI4i27WB3dYFOL644YNNW5mRr0CtolSP9OdJ0u/1I4naNRxdhO5
PWy+uV/wfv4vh0S46cYq0g1wK634oCcEzCedOjFYrN1/XAr73XktPVQdUMOXeji9
+0UvczHkiLldX87ADwPB6a0LVHePb2JsW3DQyoStIgaJbgDRH3E1m9MMrDr4icJD
kHQ9TOGIMxaJxiABLtq1A2Zo1bQR/pvlP9W89vPP+FBECMgerl5yhwvnGp/CDb+h
GfW1LY2Qyh0hLSWEX+F7DiZCusyzzGS8Z7pFqtxOQ4Z6epaILCGMW/h1Zo4YRigZ
ePkcn/LVkJm/3gbAESuoEb+WRNe0nh2JINCtM5VBVIMyMzCHv6j0qKUzjdJTRTbu
vJLhYBM1P5gNmd28ICf4mcvtz7+Dl5S61Qe2ofoItF8h/MmJG6dVzq4KUf2vkLjV
kzk681FoplbdHITuDJk9sKThJSkcs0K9OF3aZMWqoKiYiwNInTo68Mm9iMxNMkXt
rqPMZHi348ZMwb5YWQQhlDHraLn04nc381De3126nb30Jfx4NSTc6QQTWTmaGHE3
+ORnA3yTcRttWH1IhVSjpt6mgF/D1Bxi+X7/8vBowSzXe3WQcWohcBNOSUiM1Qm3
izvF3pz+9WeQCrn+s8SbM3lH64q5dbwmblS6XKxOnnDHWD+NHs6/PFt8RmSEQt55
L2LL/vphJ0WnzG1zzZqxp3Ou4xdMWplcei87Zu6jUCG0hE+keGfkfDdyPq5MmFGG
Skq+c2S/9LKYC3QbcebqlWgt27l3yIMgdEBo3vJf6Szt1gViy74CxvuEfirS/tfg
4GTb5IBqxGC+X/+HxtzAHPfFT7B2lJIVRS88kBFqMWFiexskHL1/B9QYGIagXmL7
9pjbfdHJWSNqG8wIrMwO+fiAplTpv20yzAANahUFMIWb5DFCJKI8UhCak34o1M+l
7HYDn3vx/4CAotysiapTwqvKkk/+KUEp96Jjhhn6LXQcMXNb7upLvcr2ehOBjkzX
TGb4frI4AEX6Yv8g1T/twh3grVxiKbgheQwrhGvpFjdQsZdtOky92UbtglukGgPF
+v6csmnCNgj0c9lwSp0koQ5KvnkG34bCVcbqaUGkNa7ilMc+CRORKNy6WVy/Pi1U
9oVaiiOc+Qh+Ur1UxKOmw7VGhfNL/CekTELqrfW3nIqlR6zPYZHWOuGgZXfgp2b0
fg38s9veVMmOxUc+ItsFn3c9VBNZbMr/DxR2IItHpaIZoy3he4JDYUM0Jg05LTer
z3xNWmr3AUy4v3oQVhnQU35bFyPoyfcb/NXRFyCMLyS8evUcIlfxxWIh+frZdMaa
om2UOwTwxHVNJm0YVvtiRUEn7ZoLzqwdrx+9HIAj/UkRhKekED6cNquDEmj5sWbP
ZvHcUBWaS1PQ3cqtgUN8jHqffWPUYfZ5Ou/YTbn+rrxceGyB+HIErGXjt1w2RXyY
yXWLbUz2M57/324C149Vdaj25kSBivhQW2BXymUo548E8rYQYAOyPc/jU7NF1Lzs
+CmL9ibsK9qi4WmL1yiU00wUqqdTq4se4tmgK/PhVk/Isa+hqRhI12ejR0WYyeiB
7sc/TRs+EJ/6ydtWjj3HiETadh6h8FO30iO682tX2JTPzURz/ixVhqTyR3wD7bOw
c1qDxK1tTnikEskAsbX9byG0UTOicKw4mWup4yaCRDr90O7csqrmJE7rwKUly5cH
+lDUJx5vLzfdKhumItVCT1JGNQ+y8rhOr6iz5Gw7sUVfESOHtfqidamK1AsVrCSa
39WcML8bc0X2e30QcLAfh8/vn0KgX74Rp9QwDccfrkrGN0iGsNmcK12ukx0uFG8e
GJijOqg+pnpSqTVHnaPR7D9Qrc18LbtZBc92dHxz4QP9ShEwdh/z01wb0dYND9hz
C+GvQ99T8g1LEYlKlsu68cqDeio+gWQjmxO08UGKiarsM1pks9BlhGEBM59cdk/e
TiuTzNvuL8aaH9unfa9T9DUDsQ28GMSo5dvYSpkK2mm/9MQzmYkOy9m1obMBTa0q
D9+x6Mq7mu8HiuWM2bL/VP/M/9a9YuxBDxf4Fu0bq+clt1ZWx5sWwZ7H/8hb2eR/
Z2ClAZNnIujsKjxsZeU3c0MVw+vUwLZ7B+kq8JXW1DD6z8JJahuevRoDHW8H4Jlf
uzSuInoTdY8IMf0JY8yYH/rp1P6AB18bNsP/NfE9UcwT25QsTHgt4Obo2DV3f/lM
8sj7kmyjYiO0Xi2VCaV5ITjzAyYA4LKIUkubd063AACC/bYhcgH4owVlTsbln8+T
ccrrdpX85DYR+j3N4sKJVEhBtRxxSb1LxNJlwKUvkSPFQFt5EKG9xEDe/bJSUa4r
1YWmSsyA7J57aFiDj62QnEHRAo3Abe1CdXEUWwF2HbfHJXpwK8O2CigLaWtL8Fwd
g/Aa0hZhR0986dMc0XZDskTgRjTefAuepU1ddbanGerkDMM17rrFCqsQ9IM99fb2
PvhMEPbGxpAh3XbjwvZPtlrz5REFRJBKgqZ9gw19KfONm4GLBAv2JbtRPiPTRTvU
D6AVYnmK6iqLi8clPJofCYhqa6w2/afB4Fe+LgdV5iq2BPEVWohnGjDX6gWa90yV
FNd64Gk2iNNKuvY0Ojc3flP4hX2l+j32KZI8s+sv2a7H68UA9ZClhs1MRQOeeg6B
9XsLoGEd0RNafg7qYOAXSxS3FkC8dLUnIo3Ennxi/dta1j7/xA1Mat5gC2vJN0lg
678v2XuZtlMVBMMtSgl6hYEB4ABEE/8Ng3L3655dv7102UtUFK3a+s8Njis7ILzA
LldhRoQ0xiG9ImbJFNEVomv8WUKGc0yaoRnpb+XlmFKtkWG55g3Ap6iVy6f+/TYi
VwXkJ4US23HVgw3p9D859oU5SXMgtqe/3yhQFgqrgguZbVD4Gf6irmKATa9Za3DB
ZrvG7NHSJZdKlrnhLn/Gp1tAXv9jMtLfEkj56Moo8wZJL7+V5oOdDaRGcxhnV3vi
GYV+jnVWhQSZhajSK4bp5TnQ/4AhpGA7MjVI1O3TABOiM5pzUcCTpneLAwBZqY16
fX/PxbetdGP9Uqum9W4C59295zNPAEKNPpMRSs15TW5E1qKe2HYEBbK9Zjt7WHBG
3Bz33J4ki1maNv5dgWXe8CRZbXsjeDQlWY7vsJsraIXzAar/D4paHx0YTAw904tU
NLdOeDougL2YOXneup3ycEP6/YHWtUwKwymdR58oxmzbcR4T3EdLdglDhdyab0iA
AbzJgBStMoqDF7WVqjCPXi/yZFwC4g8tSJPG/zZpm1TxBy5wWdx9PW8itKUqnkEr
VKxMupwVxhMFh7CE+AwauCbnTvkOLh/t/oo5yFXMI9J9CXTNbfb+PLjwTLPEwgEv
6AzAF5cElj96uxK2BPpwsfuWb0wFJ59z1+9w1SeNrPps6lSo5GflJ1sd9evWOzw8
hNmOSc2h6srIS03pOQN2ljC31Vrooe4Qw08RhpTcHDdro1XeiPTSrKsOPcCS6aVf
K85LHLnFqfagYfz86LTrffWWp5QRk3ca/jNuKFUUwZJob2unh5o7ZVG7+S+ovjeh
4RlJ/p7moCvENtPAwf/hEgrqza6qv7tak2RJQb1ZCKFDqbAiUBc42AgXJ2jmo8J6
uz1+nFOgZFjrR2Y33KhwirzLRZaNlPRmUm/LISslHybCiMibHiP8MZUe/d4gOLfz
MgIKOuaJQP2EGOOVmkeDqT415GZnVQUus8O/HGfJZep3erqm0nHB4Kkj+zNTVqE7
Q2K+VjcmV0f8LPdLGhN+a+NESi7A0ySvtzPxKZoUGcXm+3sCz6MR/U+hueOpDQ2J
vyTPHqGM6MVZi1xH2rNoWDCgsklPXyAnUNMqF9hBE2AwNlrsGwATyXed90jbOSAT
Ak0n4Rq7t+0rl0n5WZjVdzMZ2kwk8ax9emMgdL81tcYyIUDhe9hD29np1JGf5Tqf
W9oKTv4aq11q38Vlz5aAt0LtligC3Bxyy5jyy4kFFDvntBnerUsN/76rE5ExU9zJ
HfRPf0PofieFXybfLlVasHxSNnNlQvFtlONHzd8iOrrDm6ZmbpwyhRExgunn83NO
V98micbQgZDs6qqJyWqs62UyKFUTp7txsEVr5gz4ae2BXaeSuKceAc6FUzu6PATm
Bk8O2npPqrfcyPb+2+bYdS62RuLjytm6u/a3BYfeIfnexP30KBrLFidHFCpkyR8K
Bsik0jJrDTMNu0Q45mi5MlwL4yS6awbsdzw90Phza4heuJogF2HOsZElaNi3+w/K
aw3yInEiG6glHEOu564N8j6MGC8WNChfDJlqC36IybRWoiwEOvjOQfH4QtSbPSm9
ot/nZG85sPTKsJ8tk3NMv6ixSo8eu7+6R8cXAzm0B6ESlU+zWtp4Aw474aqYsFEx
8Dn1870JJLJqjjLr4ZqSnVyLlly4qs4E1y5ArcnrlKZTUn+D5bq+23YfW8YR3Neh
m7se0SORDYK8dHyv4YnINdudH/0H9w+n4noVHQNpFl067G4LZlWFsgFnHw0JM2cC
GRxTmQnSU2IXrjgcpA3yYs9zu5IJQShysanFtEjoJnSsJ6aX1R7SbsZhV43L3jec
vtj89J4DMhoM1qFSO8wnwb/2eSn5QtkPxgibRBw+pvu9WfrzNDMHyskLCjQjwcfI
C/ryGOkrkoAABtCYhZ2ObEG3/I2UpPZNNL70s2rCw3RvX2Nt12yZzBQjKCAh+fOh
NNOkR7nMDqrh65rGrm6Vi/4ln1MbpW3gdjVVodBQMdvhbPymEyDCO8FGV2cXGnBz
ZC5EZe6FMPEQpV0hmhigqdNx9Ainxz5z2Ze3IA9Xk2uQyklNG4FvKkXf5YlonWg+
BGmrsgDzDGqlQASBEFKXc4IL5lcpVnjFmPM12svuZxLWW95ibsxZWceq0RGBF54q
wSQeXbeqmVO163P2hHKbp8SIu6bR8b8uqpviJKy6DYB7sIpyRIldHw3rUendBbBK
3MMbPAbMRBMwZ8W4v7WyhGGor0EUe6XlRxSP66Sz93M53R3/j7Tf78+QkJ3+Fsmg
PJfvxgGTMUbbVNcqggRh1HbX5jVgX5UcuRS3zgy5DUUCTfPMwo43RX1yuQJhkahb
DTF+ej6K+EHIuq+YYNEKwAQx9CgRLvFYq6zcp1ooINRmiwI01Ok4ErMvT7d2Hzhi
w0rezfizrJ+XL/EsNJ/NhQKsX6cNulh85I8tEm9fryDioJVdZ7DhScNPe1PwGkaq
S3hKO9GYm8onnbq8Ucyp+53+y7aIrRu5YtjOqjnnD8w9HXb6qbjVUkvJqY0FYYgf
tJmuQFYhCf76EmcjaZKx4T4pQ2iFx/dBsfQol/3vGJzIa+s/fNob1zqY3cAhSCJ4
jt4QczdiDXKzCiYCUz+EGWB3sSDJxwmdsEw4eBBDRLZ21AD6s306XR0Oj2gGdPcB
YqZQMQrHzhGcf5Yv1WHSRV0mnChRcs0JG7Yn+n83HFK8j+fND5BYXiY+aq02lyc2
xa7yDVEsdWsZzXxB0yQlqQ42Fl0d9NNfVjxHyr9KvfTXcdoxqROGliYBh7/Swpod
wsHL3XT/IEsvh346kmmYgiMV7ihsNGqZVXIOkN0TG1ca8uudMPN4B+iLLy2jeUyK
xcSFG6+WjlGoIxW9p4O4QV4Jhrn8y+tTSi2lq2nzZ2dSpboi4OwzHrTA57COPDqC
GF5gm5P9eU2cSw6ybXbSmxUsb0YQ9Kbgzk8XOppC6VfsAsMamjd5YL7QmE9Ktj9n
QKIWitWmGN/p3xZztiXu/QPJXEBcKP8xAqy0tGrG0gtVSMlUidTYi9erys3qIek3
iL4d7z/7YhYeUC9hTRQpk/OysSrzOqsOsZoYEcHHBcLC8cluf6BKBZQDus03/teR
JakOkaoDj8qqWSakDBQnKxmAkzivRUBVl70Ozf072/R8biqXSXGm89RTOQUf0gzB
bTBNHjpwmCmCZiB3bPIszqCPa/GvtfMgu7C9+EfwZDqMAn7lV2uEO3qEidXOpaAq
VI7fehHuUSLbPHBUMFaPZK8Ayo8HKgiNx+TQnzsUcwdHyV6rnf/e/c21khCG1Tp3
gZUkDkjDZ6h/ALEJZW1LLMHSq5oqwOiFPLSHvwJEuCopuRHqxSkWWDGYezDYYnWB
/aPPrEp3dzsp0F7jWdiKoLa3OOLnx91LUttDXchTR4ectgblUVSg9wpgr1U8Mm4z
VLX+LYpdR4ewK5t9LFhMlGihyE47pKyNNQHEe2/1KaRmOGwoudjgWr8ucaYNPqj9
8Y96aFhl3FQybFx2PW/UVsJa5FX8Yf16Hx1J8Td2FETD4+g/t4EMdrXQ4nObWl6a
PaduRG1v1MJj8l9ONSbc6zp/A2l/+exEQMyN+fB+4KO3vgj405wZuXNutL3G7mRA
rwHDxuDn5SVQwBiSKTiAZuNxMthE8F89r5NNHkuVGOH3lxthP12weRcI9t4aAd06
m6KaaAa5I7fERPWQLLN7/Nj8Wwm5kbMQZE28rw57qn6Kv4kr9ieaIMWFHtOGRQT2
RcMN1wNVWhs3mcLBDRUhc3DuQ2BNkeGg82ssVmbPOWKV7TGYX5ocy9oTcpMQ6XUM
AJb83UTTrwpzcRNKUwTTXUHjjyW1gAGXCYMFlIG6TjiyvxUH7xqlvv5BYTdNhmLY
TICWg/fuQp5jylHw9NzkDRTZkN/+gt59hLtI4XwacW0n4HdQ3vf4OAGD1t/MHd2X
fDTrBrK8DMP7Kq6pXyLSEjP+dtpk4KelJf7mi6jD06DbqSqlSDbQQChDfqUHbIHq
Q62ccXOG2lpNmXSP0QzYagSefPNeLoHcUYKUfBy4jCBJtWF8/1vX9YI52F41MYCx
kXMHBGU50Rm8tX1uBfimIR9CH0EMWGCmXgErYQrrLeOJXyqVYZixPT7Jp1/PDx5a
bfus0OoCNX0lvgR/MSyldvNhQyNMOvaVbkWAarCjLnveIGTnaNEI1isLpnV8XUB9
TmN93b2AVa/mCpBi0Kwd41EB0fd3ht8CVREt+kszbqJOHhGeJKD/73qsQsy6K3S8
qolZ+ep8jdckYyZ5SxK1Vxr6RApys+QG9dBWWAqTqJQXm6qx6w6/ZMObIijjVEv9
8xnZ6MNKtRz0jERXpmHs7/rS9RcWe+pZS9b4c3GGABpiqhbLAy9It86smWJxoEKC
z018ga5VQf5jr4erbBcG3ZhyshceF31cCL/TRdQuF+eBuaaHxBjmOofRZG0FyVij
ItwG5JrsLnqa8O3j6rKO95rfLR+NSOYeT1QbOBpVdVnElLRKrhPIpbLeVJcDoWq1
NUbGULlR6NZwj/KJwcoaTQ84hRDXgqNofv2S8em+TzD4sNRNgrM7lHTZ1U7dg/kB
gESQNev0L9OO27M/2JNMcoC5vaxM27YWhYoPfqgGoRhkVfzTwh5SpY5ndN2r1WtB
sfVX11WW9I96sXsLDwfqYnjnLLRxmPmgyLyPMX2uxEReh6Usz2I3lQJ1dgq0NmfC
RGWv0mUisChBIFlZxt0ltXMKZ47Vn9M4uKliEefCyTAJDcDkbBNxcfQfxOnRRkAi
uvG6pTg3WQKe51OEixfxbqlxRYEfTBC7jsoVUbDugMLjlgYgwzQBREHXU/tnh8YK
+Sidq5wZq/SZzNwUbFISIEsKsvg9+afpFuDjG4af37rTY9BYmq9mE1Axlz65D3QN
lkGtHUjIi4x/dMEtA60WjRiKYbP4WD8IdKviO85cSIQYYKn06/t1qzHGLwkH3niV
Rr98AQLMvjyQ/wfcp0ExmweiH6d7Yq96zudMD4u8+FFv85qahJq1wJuzDaMpqooj
H40hI48+AnFjpHtuD6Dw2QIbT0yD2NGnRxP2NqYCA0g/K90sk+nrcRKwE+y5ssWo
M585pto8TM+10AscdrggukFJvEsuZHMOTb2w9o+9gvqo14CjQ9CYIAJ6r2FzXek0
ajMfxj2JlB3ByzjJPKLr7z/N3JS628n9qAWzELnZ9WqJlHRsY2f/62vWInpyUnM/
8jZcA0+dqLFrGXcTiyKNHOTA0Tz4SfNWkFq3nCBknPeBorPW20OMdZ8dDlpdQcj5
MakVwYxK+siuR0Eb8ZzuGl2Vmg3sq88Y0dRWIzbIkpjKMhrQ3nnPdjLrtf5t6uy+
ArOgmTBWjgec4/HV4H2JDpbaSw/EdDbvnAY3ksRHRnQEBWKvzzP6hJFyzwhDrvxS
Oy3hwuBVgn2VRBYjWnmm/aBV8xB4+Z1vCZvLI+vJy7BlbbJwP8BZD+vi8eLGdIlM
ZxnURUEpDeECWHx+IkpidrWg36bsndkPzB2Ex2k81bKWDU2rvk1QFqJc2H07XniC
LoRQt7R7RtylDTan6WaHp2hE/XXqWj5aeGegxziK9tj+kKtj1asmDbMO788s3OT2
zzCvzytllO0B65aGfIQV/GOim8SvAxKvoRIPY2Jxdz54T7Hzc851ZfKnoIC3VsUQ
G4hHhvu/7TVHUFxQ5d+rNpWNj504+aKv08cRGipWaXSzxCKeDd9w+2nywU1T8r5U
vl838UR3MzDoBXwzg40GTNkzh02qU4jZLQkoUyxaIhSZyHYrsOBExVxNLD7WfHH2
Anz8BRibN2Ub9N220nvYbkGS8/ifIPstIw2WlyCpIX23YTgGm4NYWqVTFdyJrT0N
a8jdKMljVFoGKPRpUupJXg==
`protect END_PROTECTED
