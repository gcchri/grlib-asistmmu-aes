`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B7V6jkLu1mFGXrlsNk0RhzInmgCa2UaPSgV5ZEoYmrBmY/+LMplSrneuvGdY3iYz
j4vzglBERB+SBdIj/tk12sGX7hKAlbp7qTERwHWE5hXIN1Ci87TSFn00cfISkWOF
U28bOJj3XoDpX9saFKYUSdfdo1gySa7yLoJ+unxKj1tYUqHtIIl5/WCGhrCuuO2g
lUjEry/9d0EKRNTM6FbEYCA9pyjB0SMu8qmGTZMjEzsfRfdGLfScJ26JUqaSGwMk
JRfKfZWWNkN6EOaiCZ/vpO/ReY06wqJKd8R3K76e4lo+Vj6JRuuwIfGDnpkplK3I
2K0mKJhSUr85M+nA6p4B2vlf8vhvXDKCL+SxSn7zLXZwdjFfb4X0Swa1ZgQ0uYKr
h/wLAprsN7lPmlgcAUo3AQUBLKdHyD0B2/lgMqzZaio9mQoHNQPDbfeWcUy+Xlod
tywDg+2c4fCLIrbYlGgC8Xn9AJkXM3bHSecTo1iMRKFuiVAEToXjrgtv5bg9suuQ
xea/w5UhlZpWru5zg5SgxCb8jbi46VQlJTI8EfU36XdBy/ABG5OiwTAKiPcb7HwH
p2caaOsM6YZl+70Ru+7ubNtv1Tt/oQBGukcypmRaY7WOmji3qOn367mOx5SJi9Yo
v7k8x5H5BuAR3KzqNd+yjA==
`protect END_PROTECTED
