`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dZdfVClgG7rvyI33VL11OJcq6hAORMVg+HDjUQdWBa67IwyAvQstlG2OBJSLjr96
AjYBeNRZmJl/H6gTxh04iIQ8Sd7cv3+VR6DzMgiOw69JiwBgoJnDB08SOPBiTbtJ
Ny56JAgar2r+U6LSvIRBLt18e0wZufk5Kvqc1hQSsE/YGOQFppeIeyn50ma3kMPJ
rtJVKntEecK6qmnPSD2Mf2H8u77nJi7F8fa+VlxPi58xDpCjRXpyGc6dBoLNBtzn
aAHWF0WCESedX0lRaO6Ya5Me+TcVg6Zre/cAISr87zYRROep05OrH5BJaLgpIC8U
Qda49iKZ3WHE5rVLAzhaqomoJKWb3AymOzyZavHlR183/s0YTZqO/dxTZ3pvBYgD
E22wEyQ5cbWw5cQQ3S9hhXiRSBu4DQ1tYqRkMd2MWhztLRpvaHcEzyu3GZd6elEA
SAeOa+lfTY0WsBk9hzlFCEW+mYSFc5OeB8R8BONJF9oUa9ijstETgRzcCopZJRjB
Tr9eOoHeI2f8LjKGuxUyPwMHrVYDzjywZHwcPyFGePvHlSVZ0U+MQWo68ghrX/3C
yP5u3fYlLDCIdXAH/RQ9Z5SP5ZdAac33dcaYeK5isgHBNeVha1UrMAlkRdqoH9Sy
cbvBtS821lrZoAP6HRg+GK17KdQamdwfaRY38IBxN6KXC+sv33STza+msujtxbwf
kmqF69LrJWOqBJYVbqiY3z3EsbU4d32w1r7FH5yHjfftxnz5AnwR7ML41k7L5kA4
2j9jz+Pn/g3Gz3CLvfhIxugGBUzLp+jQAvCW6KuKDEDl3pGpZ89OKXiq8DKJbwxc
M/1rLQXQdYLOwT3yAoyRdEgP1++zFRcQ7XtkUSznCm9Qy9WNuJlGgI3M6a6y53vJ
k4R/Xuad5XEXKRkgqcZ+GO1a65UO9MjYJ1uIQRxUoFjMc92EiuqCuCMqjT4M2aut
7TMwwoGXQ05oOhN8SfCFT22ouA/mvHhtFJQy27oMFuRkUtdCW7KOYdQZxX3aGE9U
XUbBuUEGV1IrJtxT9ZUKP3bm/do9D3o7De0a2aEP9OUMhE1fSTyWQOE8mVARYapw
g5ItseRkOvpl8UatWsZiilvivVnj/IOcN60XgZeICoUIzF4eM8GTM8BgzO973x3O
++jD7GrzzWe6P20Zl+UJtC6GktZQZPVOwbPpyh/JuKQLF/zv/hfWTZ5APRTxSRLp
8WVqRNPjI1MANauXHBv7OwzZptVlP6oNiIDSyoXRbbQSUUTNPnl+y5RiIc1B3Y3Q
YmVyMbkzo0d7LDWL+UyQLiIXbk++DrIPM0Yr89qimROhXlTIeL58rUQskZl6q429
iMvbxaRxR1DWLmcJ0OmGLI5/ZuoxY88nZ9COBtkRepuyxUyTsqz6m0pdM1370Ddl
UwLwdgcNzYvbyEkBgdISXmRB4n4Y3f6QqBGNGgMEEsFFV2FLjclx9UMnkeW3vDb7
aStJhHbt67IK7FEslrqS/tu3vtDpK5VzLrXBHV2ca7x7uM5+ClgVSl8YnEspmb1e
D0x4Lq19P5l1rHyVz4PQ8o3tH+yIRtcLFVk4wDlfoj+1lBARhg2kKyH1mWj97dLD
b95C6wn9mNlI9/VNLUbvZClUbD/PjMF3OebcSnW0naPou1YJzlTAuJASck5b6m7n
gNXAQcCvA1gvE0cqVwmUZ0PAwCWxUTqX2UnRTgW4eGvHjxZCUOqsexPaEjSrQw0Q
KrIu2El65sRlR1IQzWJmIqQ3fORkJHBZnZUNm6chFxVTaYz+HzNrwgsBOHLB8ESn
A0ZDBfJfHapJe/RPDNy+2ANfPA1hUCrORQKX3cmYT6V1eGEP03iy4SG15WyahW6p
Krf04IXXAWjzT6GnXkqzU/yuLRmAx6nGKtMU0GcVryaeMcux2lmHMa0SIXw8tuoV
GmYRUWKknpeP1iGuEZk7YbyU5bZ+J2dx2J66tzqlsoZKertvznkDPvVZJNDjXO+V
`protect END_PROTECTED
