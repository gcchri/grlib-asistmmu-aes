`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o4vdNnRvF7ReNqanPMnD+L+e0Kb/UeOGxDTUCBiMmo8OXUOfI5l5MN6PUnDxyMQT
Ova5nNV5pTgrvOQiw3uXWjCWErKecxoZMYiEJD4Wq1/hWKLwohEI5edBJ6cOK2wG
DwsgyKaCUOslcv1uQ5pry9IF8JOyFX+dFCHJ3V4Tpo203VYjI+7aeSZXccmfjCB5
SKL0cLujexNyT4tef/gmTSa+rTsgReQJWTHxrmkCVBOe4/z1kQjZFXlSwszlOSPB
4b0WPBvJjCAJCN+dmFz6E6vFO+D/+Ayot7H2iLE78NazcvoK0iNPKkc7903NUvQu
G5QK9Q9Jg7bxWzksKPnsdSkf2uTC5nltKTP5k/UAt6HA5cvsZ38XMggzN23iHnLu
dGW1WnubXHwimf2jcFEVCmsmzLkl64RGnFwVVHiqE5t2gSP8qoI1v57yw0+qvHDK
Xv1jAlvLjNcJkNW9oDqt50x06YADbZFK8qplHY7NjhPSihuOAwp5s+pRc7W9mFcw
X6MHSWkyvT/nOQQwOtFvE+2AFUtgiKC2HiRPc467uvXu0V+s2sFJV1FnxOfQCF1p
0Xv4EThjbAwhMMp4HP/SkocIk/vfa/XKE7j5EKFEelGvdfXd6CgTvhJLPN4m9Qa1
DjsUHtPWlkNuNaKgglVpwg==
`protect END_PROTECTED
