`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HXYoY12KO1wfrxxfxGeV3Ej3iOo817RDnX+bMf9dmRybKSyNkonkaCQ+TzJVyziY
tnvk7Piy6nUSyzlfks77xnNohmQQTfSWx7TOxWuScZIJa7gQDEhjRWQVOYN1QChk
RcARTpWMOU8nNmJIyyLJY90ssRNldfC0VF2gZ9keYT3BBQft49+ZciHwJ3mdFD2t
lxBqgHw3JyIi1V0cRk6TGAjB+yRDVpJyjUWksHLaZMRmUpUfPtAyUI4qUiJstwBf
Ef0keL1PbhMnyCLeeQCruDafiPdIb7hXqpkP/tgApJOXCrmfc6V0FVpyATmk2SQE
vq3jEDy8C+iDER8TBMJHFAg4E2WuYHRgzP6BYe/obrzDXbu895EXeR2E/3wrgWaE
YXID+dqI1vZjjrQHCcoqfGPiEhkZCd62E5G/i0kA/l2ozcCSdkP5NgLqcHt8yPPp
MTs2Qwqo1pASUgShX6aagiioReGuGtRMHn83DC15RmS3fByShEvzV7l34JFKnlp2
D3kxFZ9H4RgGaOxAK6mX7dYovS3WkG5sw9Kybw8DDhV1+Qm1f9kvWWjXEGMJY9Oz
CA0+WGYWng4FYxOXrR/sEw==
`protect END_PROTECTED
