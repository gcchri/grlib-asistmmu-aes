`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9OTRK5khN1+TREUlgmmIaeclEc4eVIOLUkdij+mYNSxfRVmmqt37gVqHkezqUcuU
REintwUWkht/FzDni/RcfPItRDbKCJOyEYv8O/6sMiIidP+FrakVXWlanbzBDXo/
xXgshGjBzFzqLOEKYIX825pFQd09vToWuKxWmXYyTy1cWtIZubJqYHN6cci82Nei
76pTNtLvGtk5jWHPdebh8PsEHOPnQDHJrcHN/f/pIHWtQ5rjYkT/5GunoDcrqSeA
DNEkkMdjkkN5rnUi9BdVcxAylcRVHocA11wKQANDjRv9HICVpeRr12uIAb29wMpg
9idtnseeC8t1UAIi1mEUbGQACoestcDC2hTWYl4LKmMfFDCNrqEHnetk3FAl/uhE
ASyW/mEut50fQWz4p3vezQlb7Pl9w/uFm1rhq+AqRVMPWZXqt2MymtS0UVj881XH
2NLLPvWwx+CtwuwVVaNX+aYJLjjfp4Y+mbXo8PJr1u8oWi52/E+jRzZOdnqLV8OX
f+tz79YdsNzpAo5DuWNGN5k4fNXqZqWoUHaNbG1Z7OFcmG12U7hvPm5SKasx61pG
mURKqkJAndlr64bumUgzn5zm9qq9grMwKHzCuhzcEK0KGLd30VthkgDTycGw1uk4
PqO9NNlXQLSURk69q6jK1od1GvyC077Ifod/hdifJXCukdC7tzRR/oD+MrXB6biN
timQy9ZSHGmlDEKS+A0oCox+A4Zj5GWIOxmKk+VNjagQEfgCOCjALgGNpOk48Zvo
Uv53OBuOtzcbaP+933qWYobS8VD2PQJ+76TGkW58DRvlBUt6tNHGn6xjsDq5mnLr
VpZscyUdRJ5OQqStwmVH0vRVynCSCtx5nLx0XtNFZs8NnoDkDgZXuYRJ4jyTbngy
em81EQHsx1W6H9w6XFHPLENz7LpRrwkYu7kiHUPFmoT9oY6NBVP4IJ/MZfZh9njn
N9LL7qfsH5jGPs842A7x/d+tclIKjnPX4avgLA8FASzDwmYruOph5OKncJFU8ViI
OT9FwELCSrPjK29bH4l3XUJiNpDqaI08/m9RiNES6l5sZgg0fV+KcTKXGJQvZujM
3W+nZ35jQKTD8GbCooGO7lGqXjpbMO0rZEhT6eBcq5HSEUfEMz3Ze/uNhGp+d7/C
aZfh4oO1H623QRJl82/juNTm5YM/RkKrxIPaq3O7ouh3rbqDa62d2dZuO2pc8TGM
RmgnRS09eJS6nsrq0kwvXeY6+XMja0gGfIJdQHbOrYMQK+Vy3u3uW430uvwSn59K
1eaPDK8XDBW/yU6NfkoK0D70qGG6nWq9LZ/RV5hb2QJhrK6Fva3GuF4RhCCmn1Nq
e61nXoYpdO+Oql0Y46kanloqLRY8Op5x5HtyeHebu8wQcOzlBe+rYy5GNf0mEsBx
IvZDOooSXdmYdZ+c0BPKFaLYkbI3gil/k1meUXebxtgLQ5EEJD8pvmz09GpwXInJ
`protect END_PROTECTED
