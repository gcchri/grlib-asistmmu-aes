`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mibWGgiaP4KOzTmWdUIidSChD8yt3XtQY1SRs/BP8ML3oeTxjBJN4phj6fdExhjj
NdbzKFVlKl2BVKoUUqhGa2izQmqFVDc/I+vFuN2UjTph9HioybEUuBxVouIhJLLW
3gHpR5lL5bW9+G8LKoCg0RUb84Ieub3WuScepxx4L0PP7l074M2Rf3DaHBHGzhXO
geJM9JRI9Ffh6sIreOgKSn1TuYmFMricYlMCBmqOv3exoGgCaJmWATgxp/dUer1u
+Uim3mLrg8v4ro4RF7XPMX5q8PcuTIYlCcImEGf1SJU4NLrv8/WTDaHPDlx7lxnr
tH4qbva88sbSePHzw7o5NXxUpPxxDeZY4EQY0tkoGp6BSUOD+VN8X78vHbD1ufw2
hF5nNdRhZyNfRf6yRnDIfnzodGtcSx2IWmmJ9SADuvzmuApPcRltcGKtrOyAPLiz
R5MLeA7TqyyNXA9vwfF32Dwkqxc05Wb6tV8uTfFU2C0gwtN4WbvbcaIZGzd+I4vc
igarZsLai6SCOMbLV+sl+vynx+9w7pzge49RDCIOT6M/j0w9GjOnDx9ygkvq9oz9
aElTNrzhBJrV4AogpHcpvbNyHRFBJ/UeeIORhYePJ7kOVKYbHhcDgV9zdCKD4i4c
e26wvZAtvoFTpua1HtR72rNvP0k3zAg6LirCsivBLMLUFIm6oXjKJgc/qLYG1Bh4
h1q+SV4qbfmWU9SZfXMpkIKSJHk0LnicSTw/XP2yLvIc0HaKIrlBb1+8iK8WyBCS
etCOR6Mbr2A8GZZet0VANI0EaSSW9JlJr5emQsQ3vv86llq+NUZQsYZxP9WwcjMx
CRuHQ/3AE99+oFVzjxzbV5KET99aCLKBiea8EX3jwlK9YMmuk9SoCH7z5RxQ1kxb
p/7FHRsOcZCHxDxYJIbqPoKo4C7mlb2XbhTYfsNMnmpKzCbyhCWHPprEIeBmNOnD
wgbXCsoElkzQY105l2edm3INZQGJ+J3gmL+EisGW48r0x4Xvl0tJOu+SqkBSTmpA
rJSXxKKtigcWS4AHcV7r4F5aa1K6ucFix18XjQ/pGkRiEebgRwEfg5kXU0YdMeYv
gQCF2xJXv9pTwsDzGZ9k6Ba6nwPdOePyv/Q1ldZHV/+UtdazJdClcw2st4sSFTZ+
gIgrpTxPFz4QYzM9wS12ByVqt0ataOk/BxHsRFCS0z6m2KCf26qP4QHXzJuarw/1
aqBhUZ4zfVe6qemyXSkXbhZ3FMOVTfYaokzikisc1CN1uSE1eaI7coqu94LQVWJ1
m05MJ27scFkitnzfUgc8vLlucv3RKDQuF9AxYAMv7ITSHa3zYxEN6je4plotFpBt
wNMt1wIJYzrP/Zv4zsGGTfvunczQjf389fR8Yusr0ikNll+P4egbbsw0lO0G6R70
OxH0v8IdlRZhtgc1KOxfE7lEhC3mfKrMYtxKkS/wzl9Wpxeaj9ufPa3eQjjZaTHb
N5HHYKBHza8XJ4pRL/SeCddE/M8uPR4sp3RvxzGA9GSk5zMNWZFZ/+uyDVqXBNR1
eoFbk98Hbab7kM2cXLkGjBuoNvjKXr0W+Vl/42XFV6hwCGPCnVrbEq0qiKkqr4e4
3bvH09/lJmy/XC1BU3sC2oCelrBT3JTMUINxLGdpfiQHdaN6AasZuhTXHA9JpF++
QKrLtI5g3HF8UnY9ClZil8+tbApL+OlaiVumrVSgIP8K6SouL+YhCCG9/PNRSglo
YesFt3XIyMInq6c7XcMvSv0PWUGd0IrZi3v9ualEPef7T6iF0HW4F5pkCwURKnKy
WrLD8pG6P3rtgNt57LAUFhfBZYOivXSfVDRyIe5ly0oVuqs8SujK0bXFquXnKIMZ
KlT/kFTks10f9I+tghVxQ9/qmYV2h1NZDv+ViFsEwRwvod3tuPyjucR54OzRJ+fc
12cnD3IXVbLlefjeSZM5LVszOdZyRs7CTS1PoeCwO5rfEVo4xw9xBbj8nWbgDstM
AM+tK6FUdVPuOLvlWt5kOlWKvAlcsM/IkxPDtyQjJUxb+VFwMKb9EPcrhFRsYtgb
Exgd0PLOlZ+glRKga3aZv/JQmZLmc+H5uupzvLc6aPWNMksfPM5pEmcBEoZgjhWN
zMoV8UUXHU5QxKrzwlbX8DyoOv3D+yxP3xSwz9kxNta0kldXE5LeW73ByMFEgWCV
4CohRCOtWCGBLjvUtRoj9KaiEXq4JZXrQhoeEvQuWoLOwQLfKyOnZgdGnSq/6EjY
7OuJ174dR1ufbLEwg/WIEjzH5fJdLsfYZG/ppS0cEv1fS41AeU2fcOXrhfzyWveg
CpcQaIqUS005FqbdIzifeG58AvoDVO8wNU4BmD/AVhs+/ZYLTwmvQ40XKXHv1QO/
skl+YmIVwblUr9o22UI8CZ/17rxFb9JJz6OZGjTSj9W4/aGQHbJANHm8URv7Y0sv
Pl0poLIGq3QTVRBEibW8jxsrrOZzmGanqxPG0Pa7wzUMKL/c6zwEcmUJuz0X2sto
OGcG5RVYpuZnDzvlaCSpx8C0QhlKfxNoRwsjxgMO1WRK4EcV6RwZCT6OrW0jnGzN
efcWeaf7lVgyVHjj/P2W07lbL2BSUyU13Udtos9xPA+ZxehG7vAdmoFe6ZQAe6MI
hOnffOLc5r6kt0GTY7mFxsI2H5D6Df+YcAxMIXWZMWLK9tpbvPTST1JVZXp/KJZX
G6tW+05Fu/WiGJCm6sqx9rZu1SvqCDz1MQvv2l7O8Qlg4ZPP+IEO2CO46KrUh9c/
1WvSKn88J3HyiN7PfAZdQHHL9JwEsAuY9u7//MYnDgbD3wmj4vuNAaHBOWko6yC9
/UjFt4HKleG/BSH087RkDeFpH7NhIIEuLzhdmyjxSGKlVbG5OdayPc+a8Fv0lNXW
haWClw++lDlkoKeWIv5ySCVtkS/HX5nJ0m3H4yEJH/IxkOsPYtkPyrR0MdHKs5uG
MvqIDYXPDwNsDqJqRub9kakQQuZL1J06C6aNY/ol0ZKGYR9z7oirgpyjc4xxrnIZ
AHKPXY2DZ/qjQDXXMjzTzt/gUGAteC62rnX2YZF07c34zC+efvwWEJdUeU3IXECe
85IEpCcH56I34mZxWZkLEOubOXIyMCqnOlMXPfOFoZXCFPqKE2a8qb0ikl/FgGuc
BeAO0AY7IL0VVYTCF708mo/k8f6DX5QafETqxuaCi1elrEMd+QLiBfdoYroDeTVC
vFyRMPJ4rogtyS3+hXjgHFCBAGkZ527iXDUzAe/F1LaDVMcpIL8zogzKr2dKFNao
xoumtx9Hjb1tHq6G2EdckRhMc/6B4Wql5vWQs1vy77ilfNzixi9if+JLu4izyhfZ
6wrbpfBUYOYYIkd9s/1RvYv8uw9AMir804xE2LTUv3okyHV3l62YrCY8ffLpwYvt
YaXLJOH7KVZoS5hFcoxPR3xvDBzHGPJAPwjHNBWGthdLqnFzw2uF5+/0Xv78ZXEF
X8eBsrr8JdOr1LRBjeMkedoym+2ITtrtntPXYwgc3C9eV3ZvIRStPh26G4sADQOd
Kjt/yd2RaiqlpLispEiu0TrtSRsYRW3PaaFAtnIxHry0QuhQw/b+6L/k/sDaVJKO
feggolWouzZQkaiFcJeFgwae2WrNORJ1oolO7BVNb0aPg17Gg9tkUYjhoPIO8Rda
KCGjeUip5+YjkL+skgtXKLPKk5DisSIBjR5GeUCCRJLnQYtpYpNxKQghlA2dYH1i
hQXbJtqMDKU3nLpiXc2/renWo5pTGkVIFYQjIkvj+SjgZkq4/uG+XIn/uZkip7ZE
XJNvod5ILJ1oEf5PoArM7wVkii54uUy6vscoOlz8h2AxpvrWtBmJN2MvBW8PSOO0
TdUt4gOLn04XmOH0H6HI511QAjjAOtvyxUWPiI3xkFVRPWL1v4mUcXud3qUUqn3O
HJY0eHiGBabdgt2MuLyuEZesRcgvQMW/CuzPxTIBYNnw6M45TWPIK0kZYVt5d4MF
ub3aCst07idp/ik3Y719i8PhsgpyhP/lRgn3wvmtNqc=
`protect END_PROTECTED
