`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ar5eCn+STIfJqDQR8F6QwcWjnRMMOHU8bR5ca2bSQ9TwnFNqPvLg/DqvG6Q4QIjl
bKcU0XUiF0AVk+cFraMVuDWgLr97ZWZRuNG/GlHztg7XgLm8UVdo8Zcytvw3DbH2
9JyEFmbTtE11D21MdG3ptGx2nnhZg6ZqahSkn21tL75bAyw8Ot9gYIekEOaBMbQb
kQJtYsKsQREMeN8Q+kcxiuQjjNIFMzGzfZbHHFfaMarwYoY8tcYkH0I3/EDPDEmN
rK4wJhke4062QOvp9El9xwc7oszz+OslMElIn0J8KTdsF8OhVUMX22BWfeEGI5+3
nZI12JKrljP5XiFy3kyG9+jIqIRzqtlw/WWELt7mSxsgy4zqdqnLRjDoIo6RTW5I
uu2QVeHLYkP8LqHfFi/wI/NpO/mP/heSZA96Sdi5mjPvQdrVYvQhOdUGIndytEl2
iCcf5Z9OhUzMaNH9O1wCuTpR249abMACmdqNADNFTSj8IErkyqXTxKxqRLQX6vcl
ywg1uthriQTxXrJZf6rubJuJBuE2mv54VM4OsAeVILE=
`protect END_PROTECTED
