`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8m68JEhYXf3LkGMMVg56cUsOcsnm30QnILUpa5tXJg9ktBWaNJmzfP3ySi4hvzjI
56Zejh0h692Xwd42wFwf9UJU0ttv2lTKe0/SB2mewWLH4mvHbYWCp3Qb6fBtG+Qm
S6Izn81+g3b+2yCJqGa9D3irgOGVJMiaxzrQnHu+RICTS76aYd8dWeW3VVXO0ok4
hJVuq7J7QQbCrWBjUsX4Y0cLFwyQ6UGCQOAYYG848D9N7EwNbTpFTSgFMuwxGBSG
VrwolANgfEUpL7UzDYUBupEJFjeRS97E2Gsb5uOEnDzrnF3VRyPI+RNozEDzZTKA
HC+ENCwm6BNxQXjhUaZp5YwM9PbEeARVG92dZbHXvhebz8eeKmMtUyNZsmc8z0UC
ubCgUuQ1jP/e9fGxp5Pet70Ah8nTv1065qAJW51mf7yaWKfs1XsJ/RC6Cv5vUJR5
gYM7UScNOdUKYAY8+4dsVpP0qcdwfpm1J96EewIghQ3NaG7Rg/HeWtfb9iRc6Zok
XfD2ZCeXzL3vBmb0ru//Fas76Ek2yQyG8B8YiI+75WqO0Bv1OtoDo3OKcXF21j4/
Eg6Qe+vbwuIKrBqdyGrpRnDgMosN3o2SfNqCZY5Bh8WbaFia+nlXglhJbPv0pp/P
U68wxNDV8lpWF5vERSQYNG1TJRI0En2ZkQhrMSwCbQ/ENlW0S4Ip+fbh7b+2bKxm
LSPHcgqDZ2pVJt8K+thDvrp2MRL8SZzMrvvLxxInnWj4SH0i2XQrj2iG3lHKIDkG
UfoR17YoefxUqEJVE0Z4/NeaCIi/Veeyv1qwEVM5NjGhYImdWb/epcZ+L7XZ41va
UOXDRr+h0nC2+iMEeyz3lw==
`protect END_PROTECTED
