`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T/n/Vvnd1t7VWFA8bdVYNo46oIHR+gFeYXmnab5qZmlIjPjwwlkUv8ylKqy5IhZi
Em8Tdi4B5mkwJoNKo/2lUhWAc5gbuN+Csd1vHHWjQIHz9AtH9USetKsDfDEPPieF
286hj3njiWvzYf3X85kPDtcPaAOGIerIE5EkGvV/bjM6RiH1gvRUB87YyKUFj+kU
TLigubgcbXF+QlvNO4TVaee+fiSu+ILpPcYh9PUFe0s7QP2daZBGHBQxdJ+uDUiN
fz7OK+KXbf2CJo8Pa7lL9IDNz11jQEJUaIilRMzNylYo6alCocV8mpKpO5toE/QQ
D1IIZVYXbpXsTCbODR+p9Fx1lRpcSlBOd2IU8YE5bKi8naKCLMjJ7tImgE1sLXOJ
eQWSPP403Ba4/j/rNWMaUvBNh4mtNHeQooF8qF3bT4+xiyTxZZGjWu03SW9l8KSk
V5XcjEL5gTvfg6ZLIloR4dji5LN0F6NWaqIHIj4t0e5nkxDynhprX2aPt880IvZ/
3jLOJ9JvMtEweheKonZM8P4okHaGr+P6LrX9hwjunWtO00U8wtUb8MDeM+WgkZLh
nGZb4HlOCGEKl7vRO/eQSXSzKS2OxRBd/9Rz9L8PmXzXL86xzskrnPVCaFl/F02N
FncFKEB/23TyPlUAHblgORP+YKl+naxyH5oCso0TcpUXjrrMDdtxSBfCAyAYPr1C
j7By77tMpE88kBIdW+AdjmrB/RVg9YdPCtALk/0+mV980neIP0FtVAku8jsWXO7x
yggc1rln0H+jotRDnCIxSgKNWKqy56XTwFa+LsXcbcc4WkorTp7E0U7hX/szVW0g
GWvWzOyhVjYf4EgAuBJ11S95fcTpMoHXLWtBMtl6qcVQYzRNeyHfvWMEP5sS34OV
7Ox506a437pk++n8+x8JqQ==
`protect END_PROTECTED
