`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U1sHiecvkDBXT+ei+hEEEWNEbmyuh9XeHwEez3VOG5wWwLEszK03RBsMw7rVe/F/
RhGg5l8wZbkYRf0EwyAnr2P4D2/KDw9AKTElkbuY9j+1xFbG1+PszY4Am4UAz2YZ
neKnM8OAkZPe1SMp8FN092q7/ts+IEhIXzoZkHrDVBym5I6hl28R4wuysp3/4tZB
ujseGd5lqhJ1ShLrLN/mRRP9kNYPr9+5wgV6YRjLF+uyDaz8klMP8LRy0ioX8oY6
WoPGkco45qvkoeHWK1Wt35/oMTCYdzkBnH6vkb35klPZbo02VIcI3r6V/lcSREd2
K1jG1WXa/JgqGhrj8Roc2g3zICq3rw2YMcx4gstJtpLsDZ1pMch6UNQ0FPaEjMlS
`protect END_PROTECTED
