`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z7K6k2X1GKWPLdDGNvzP9zOCHI7Guh3tl80/ma+Pm9P5sN9lIAaX/HgVdU/cq9Eg
dabrZcI8XpgjTw9nNlwEW+7FOq0aruIpchBr6C17NwwONSaNqrh+oGFwGz/DboT2
tw5UXzvElbvFxwn56w6GgTkR0gZxdLAUZSsDtWFa3plajGN6Q/1WezROvLODoAz+
T1FweaioLmPx8haWBqP/L/mLwIERK+f5l1+TueIMq7quxuriMMNAypnYw5FV82L9
PJb7r3U2qtnjU+73hbK7FsuP2lRwIoS5RoxILS0QFXqkUJnNqYZdxAwP6GQm2AUh
apnD78KGrKfuV77RQu0US5y8XDwGJGiXhl9vQ8Us1crVAk59J2MHMzN2SwfM55Cp
+g9VPsDV+1YbKB3OZ4lTawE6sVNl3gyp4JkUgpn66dBZanO1MTJCUZjJtv7HL9j2
Dh0YvpnNaW/HvUCuc2T0alC8KdAItTD7R6eh/9bwPoFa3ITeCu9Lu3bP0R18Y0zb
X1TTRWTYE7DQS40Lruse6k4JbiMk/H36HmZF82tKIfT/eVI/jTYax/mEjfxGjNB5
nMgbvNMZe1koHHM85A9ksudWGsnUAlsNeq4tP31NqA7utvytq+ul/CZotOl6KJoA
AN8u92ayZeQPtekfIAWJASn/GiQePXZyZZXNOZp5qGdL30wkFeKpkax6/UFbtA4i
L5ugA0Uo7trMqRxYTmfmEIwHpfV4FCksLlKr+VEzKaiaG/PljZybAppra49jiBOS
e0JoXc8b3zyyQghrIPcp5QT7TNXelbbh7ariArXxreT3EK2p6FME8dEvju5fg/TY
pxx2fxC7opcOFvKbsdtQtqzrYJa3Lmm4w9ZiHhSdvf47z2m4Ie6noGWRKxtdaKNJ
ffZRefUyU6gy+rxj/ZVCoHvI6w2LSl9VeOEuTIMbrVL/2nBa4zQBtnoS6RXd7d4t
ZPCckS++bC2BdpnbIXxBNcISQiRImn4VC/JCJlR1cPOSYjxqwEQaoJH/IlKrXkpM
dmTWQH6bwdTyNfOyqAcUZJFBAh6yQiWQW6/eXf786Gmo4RbGsRsx+ORDCv8jNw80
cxZe/c4+R73bH8GFAavw6U83EhYhjqKUQTHzC3YO7MocWeotLoqYwH9IuY0D1qfh
F0J49gYTivxxVpr5dLgaPEEQzvSg9hj0+cJeSANfISND9dRvaN38eK5PJ8fzPu96
tvVXOGnl1OsouZbgl70bSMxDTS20Okvy6C2/bXwFoLrQTltDhif0tZ4ZZnMUoToA
1r1QASbyBuStS7Iy6oWbUDE4DTm+kKjtxCcvKoEEyWuK7s9s805M1r9mVnj+LSAr
Q3M8wwTJ6XQqmxWovQpFgBWARdWd8AvuFS4Vl0Tc/OgIzujSk+hFSdJ93bK0f9zA
1tkRLWDHVIR2x849H88lILJ+7u5s4dJgMyFHkw7eX1NuOWbUoON6PzC4Jwus4ilo
X8da5EDufxjLcBMUnmkybcIt5JV35Uy+DB9rzqQC2sOrbPJGEhPgOdPcUBTGi3FF
61QSBQJVztdT09Y+BkEssdM6Pzt63y1Bd8bO6V0JF94A/4ONCaI/4pgWDHHSk9xZ
X8pPiTwBx9p52O68QgU0Z+Wkyl+BAL2gkOhOOYIqtpjVg0BH+DbE6JpyXrzYmrZl
is2o472Qw/I+qp6tAq00HsG3WF+VqDgE4EVzqVQ3xce8E8WAalKNJZPSZJlDyxca
CET1scWXTOY2Z/sK/e+mQFydfW3wmyocJVWX+tmpTZNuZ2xcEaV91gE+aqNOWxik
sLWrHxK6CXiTAa9ZpW5KJXoEv3P18rUqH/LKtJFt62IeLgcvc5biTZ8XzPeOF6aB
deVM70OeG77AA0Mwrfm8e6OS4LP0u9z5Qz4iX+x5g8/HLxZPEDwsCwK9msFnP7wt
qmUn5hXf7kbzhLXPqkG8ZPSNcoxqdEJQRUBzMmCOXB5QKlQEcK5loQB95fPm94vm
0CaAenI98PeabtAW0JFvAOHy2xaUvPA7MeqntkO7yJyRSYF3oGOK4tPWXiAKqN5/
KSmipoGvH3qLQ06WMmd9lOn2f8mRBN3nY7iYUg20fI4SHOgUYN7lHjrYBwRfFFc8
zlExzRg/SXyECUhq+nZqSQFTFbAsw7Fel2Nj+jo9nsG66Ppem0mMtlGY694C6+7I
krYIZ9fcGo0pUZ9no3Tut9wVqlfpQ09M/LWCTV1T3tGiXgJCkL1UrXh2+zANJZAS
WH0Wh66UtPOXMt5d05PYXWbiTu9EhGcCWnu+Tp9rkuH8ljMURJkpYvA+5vmAC3qo
7XWkq4Bo+vUjpeafUr83TaiAz4HmXNllpXx1TAyOzr7d7PWueTJrM5H0UQl1xZqt
hZK2tCvSV8YPQcAaAObzajWdbyxEK5zqN0wXyj6/WYsGYqwX8uxGK/Jkz0uZBf4f
r6xsITUyYcotY/sJ8/nSdIc3hqFr2BVo3k6g+e2lWAVYRAZRO5GpD1676ifptOT7
zfnfVGlO5SfVzkZcE1uLsR7Jf96Y+wa9kC5Whyri3WEuXqtSjpCVxt+6/ppRfvI7
9WZ6Z+XQ8JWgdrmchJORMUHEavuCvgNadAlQ17KK0T8Nm1apGIsy7X4fK2lBWGoT
gAWnj1m+Gyxmk4xaxhMIICJmP6NkDirZo2X+4tV1lfUQNT8elFFRBL2uBTGyxm+7
ECfk1dDwabMAeukzAPgXGTjoudRcqZLPiGK3fU4DnJCgdE6l+jxfxjCxZdEScU19
mHgB0YdyKclJXut4po/zTaiWYnOggPriAy0kBYWaoSfVwT4iSUGxCyI+frwieOUw
sYLv2kfOCivwr6AG2rp/Yw/UyS9Dj6mfJg2ImePICLwdv1oKwPRiUCAsdXh4wZBn
ZZ4LVpk9Witkqg4QKSX7VYHD7VIGIkwRh8yN7BipKIO9PSMkUSniEgeCKI8c5ohv
LqpmdiuMt1870x3MfXVXzfvLfN3FYmBjL4658RjVuP8QK9NZlJkW+vIZBFw+bm1k
2qWUBLMULtwz0fCnV8exnErEoLkk6DmzuqUYX65g3Yd00Y092U6PFmTSBMdYKHiP
wW9SKjUe2dsHv9eJ3GBaDq3+5eukAVsnmkRzvcZm4fWF52Ns7XqfoCAW/RH6N6u7
7uf0r8Hyis5dl9cQ0BX5yCeHk59ZVGZ/2/HLjHDvHOO8BTcJ8P7gGAGvlV9nWDsW
2GM3Ffr3eRG3T38RjXsTbOkzYBrf9M9Af/B37+NW0ctZGq7lAn2hDoXtOcE01XOs
qh5ARsjzQsV//i8noSqDjY0hkWzGiJcIK8zjLUpmQKBtBQM/NStn6yJEcOP1uFzV
h+wOqcUg+tTyIECBu/Yi4WkKIhrLis76gsA1KQiijGZ8RUWlSvfP6tt/P7Cp3jVs
BifsYdha9i6Bt1DQpYBFZml29Mu+NJSo9V++Q/L+OyA5yjy9yFPk6Snr6qHmAuOT
KW574Ffx1Zyjm/aiuL8vocS+uzU8KY4aUIuo5jBMJhYPW/1VZAQNRaZ6YR9Vl4Of
i0/zIqAENEdsfsUblRc/9FUMO4NOq6ZZymjPsCISP/9q9mWLfH+DSV48EaI/BCvT
dL1vkWjGDifH75kTEvr/qciZu2WLXez9ONgffxj/OK2XjiM2XxEZymjcwzWH9GTt
PS+HC3vRBPXqaCYTBvlzDruw2wiQs99OzdzumrPFI2V3wU+mjgL+tvy2hz87GOAE
uwK8Rwl/SlehjkGjETQ/UxFdvB1j67vEOEjDOLGxbCYonuMtH5iyzQ8slNEGtkmc
leQd7dOa77UkuMYe514eUA==
`protect END_PROTECTED
