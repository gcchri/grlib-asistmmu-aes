`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eaXrc4oemleGRPf9VVxBt3c0xeavYtcOq2VriXUaolaIDDi5v3iAPU1njFLSv09k
cN8Mj4fHQ0kTc7EVj1blIjuHe4fbg0GUloNl1IWzJT8wWaMbwf09PPySzcG3pijk
hWM6bbOivjwf+l0VdB/B/CG43LE7+KBxubOhtjruwgWqpj5kan2/3/wcmeiZSWkU
t3AlwtjO/q+zWuJdyGsdm8V8fLKk8qIrAzq8n4/UXyD1nM2sZazB0Xm8KWbJEC1y
aS8Xoqb3o1vkWViKix+Ywbmaif7GFIBFFn2ojQ77wD2dW+ip14CpXapyzzNRHLPc
wfGuZWGVn9sZLL90vX/KcWJExksPO/VEEXqCSNCP5a73CeB/WEoWFlhCc/VLeo/H
bOv4xk4ZOtbQbGyqvRS/YYUF627DQKX7KVtMep/vhMtYMdkrNsFCGOHMh8HEycAY
qGGB0UlRMiXyDA5DU+CpZediX3BWzviq7n+wy/ZnoLR7hEtMRMMQHxNxWiOMfUDf
uvh4MacYeNj7z5tsrJmBsGyvjVG4VDe6aGRqvAW/i13YjxiOO/ZmG4Y58sFLqllb
jg/EKhUERJhW6WLVr2M+fPqW+l00uXTuFvTdsH7/sVkpkBZzsd37iV7nqcHciuKE
UsuZ1ru/qIwXftUJjTHaGK3Sz750DYd8/ybMLdFUEHwdBMtFMcRx7HRHV1FZshe1
2/V7/E82bWNUOJdmno0IgRueAaQxUYmwy0qFmAqeW1GpCRcm4sqYJFxFnJ+6jeNA
HEOP22k2Ovud8SifhY0KsOzbbEYP5ieduKBAP7IyfLlyXnCz5C84RGib/6dAlm0A
T+Dektm1PE82lmPQ17hu44fao/19h3ZFk3dDsjk/oFacOkcWdgn8vnRgakkBytaN
MAGFrk3viqQVczzZC/1PFoJyMrkxfoMKXlQ4sPnHTrVE4v+Hq1DFE+lIX4bh/2o2
SMzEtJrtp8FXH+bnDsr7dcM+LMtIjCaODNLjoQfccGc3Do89gxARnblMb4eSaoW4
te2y8oUQ9OcbumUGecDeoGtRCCAR7D1fhp1CICU6k1M2Ma/BktYPnGW0L75bXCu6
29Q8SNfRjNQMJMMfw302FwCfOnWewUf4l9CmcG6lrGzw3BtX5qNpNro+AS0Ssvc4
TL33VZBwdiHnejFRBId8MQcHOoIp4RRzUM49K3b+A3jBtQD0VqKX8HE+bQYYgPpS
kPhwhDzwLRXh/G3tPcH4fFOm3E0i6m74IAzHCegUoP99VuxblOd/mVKX/vaKv2So
37A/MI7KMcytLtZlKxoDIsyn0JKO8HfFhahqmzJOvRPogBS2+XGPGBXtUYz4GS2Y
4PUsaQlwBZeo4DSr96L+gNX7Eqz/7vz7ih9HWXYi+eeOfCjzXqsAl5l9difWyLxv
idtD7PdfBhxGsODJj3YDH09FwPCG6ZFd61F8rDlVZYgWp7vp1fKbciLd12O3dgej
OWVMjLqA98graCz6HIMUcpXutvcGhWJmchwMio7ms6AB+rVYUuvMF6WbichmOTcU
hbTNSSh0mf3/HBLcF7w/jtOw5nQOXce5G08XVGLvZiFoDN1G5LPvRc0PwLNP0TDE
yjRckwjjkimSHKmkw86773GtfnZ9Ozx+uT7QD9/frYxXvUYC+6Ct5lTJp4ts4jek
3KmUWmiRgYFfSkrosevGJNJvlKrKLr9na3B1DLvBnsiuOMX/3czqI7dPK0aSufT4
krUp47GpISOV+9+i08X9D48iBHqEvwqNki9ev/wAPV1BhCyDhhTdmF8+a446tuXU
vq7QVdLMws8nSJsfha0RNuYUKG9Biw5mRjFbac27BjKueb7NyyI3X5TPlAKez9/2
BoPHIM6drOe2pCECGadTX6azhv5lOWYM6fLNCDESNi9C/WTxw4255EqSMTAvtQI4
jud3O/zplsnbBZZxd8xJSH4hHlb3bkOg5/RDOfn6YnH/yacy1VD7k0TpEdRHCZ6K
FUSDKyvIl76ojqL6AtVPn4FJ30u9OG+ROHLkliQNbaFvITKvejbpq12LmOXBW+8M
oBK3jSp/Tko/kZBymD4sFr3W5PHvehW6XqfsrJhHyu9jKa/kaH3lDSWt8W6PtPqg
EBVcnI0YNnQPP7Z/SI5MsjWdoILLNYQBBQNlfDQXyFvJdCp3IAS0/6eDXkyXQX80
uI4Ed2NSEqhDBUrNEZ1WabRbemx95ZntCJgrdhPdC7zkMnOxjdMjqvRRpb9uwjJ1
yZbwsCT/emF5GfdTaqSfKIrlsMtBwtsGxYSTIzlLmxrKVCs25fAaJkaWdLEqtlO0
YC+IRtbg9jhgpgzfMiXozA7EmaXaE3yigROdR/KGDxWOcGG5GIq86gO/BWNTnVe2
bqAbzmvoSBu5ZuELpTj2H53GKCxAjFkks6Hqptehk3H3j85dVxMIwN4DZzspqp9L
lqw4SBnJuhfLy9YPR2JqX8+HXb2vWtsQc1ZHKTx7qwVqVDaE2XKVjR2L3uDzeLg3
oaCr3VI+ane/DjNo95wjqUdCKZmjjz0uQ66wypDqbKWHxD3nVyRcPkoo+4retz3H
m9C7h4SN1UXmd6NjHGlB3fWV97kV9PvcYoZ3zeeRUG6kxibWesIQKvE8fnlKjp0C
8FArdoSJDG/We3C9clHMgalGVvHeyX2+U3tUK2b95EGeo/4sgbXdLzUJnWnSxysF
k08HCWfGd+XF9TuNspn+Wmt4NfiDR2LhRrVQCJErkcsods0yvPZuFSlKiC3piO3n
a4d0y54Gw+KxX/RW921LDca8ULGd+AoVX4HXugAaR4P9Ku6syUz1G4wkyf8TVRf4
26XIyfSV+pH7EwtVCNfn7fhFkK0CjIug6xsPcTzN6VhbkH9sI/32/5S3NMwA6Qnz
8YgI1K+/GnNRTMkl5k3XvVg0RNhAuoaXe7Dyl5qbTFBcXypQiXJbYbpEuS7+pYAf
iDVj+0jCczWWRUwydPT+JCwzOsd6VfZdzX55tgD0mPNrCdhhn4aXsJenfx8PuUfP
dZuc2kCqOQbmVINPai4fYxa8sOpw5O/d6S1JN5VXKf0x/W333pd32CrPU9StmqhV
Frx8x0qj0VXWVwuSgW/01KRAfvqnK6SnA2aZnez0EQrhIaAJ+YP1ZSV7X2ilqLXh
6sKHeE9aWHiTaIPn/t/NcJzdECP7XJIQIYtj3BqOlckTnjl71fZLyAM3UYRm7nYf
V1/dVkJPEI7BkCOTu/cOSMmyeJKY8Lzfj5u1BnEL1bRnQwamDe/XYjTXsl45THoc
eDkQHoNwu5C9LAx6Q15DQ3IVtdLW/olqEIS4Bdfsm7VOIy4yFEPVEA7yLWqpAdut
1z5uK/gRUbwbHbF+BXL1+d7srlMt4s8XCjcKAVK8PwLG+i3ZrCL8PvZjo4hlEwUg
BnejjnvmiUunM+6yUGUT/le96ZOR9LyOkSZIqJOXkPaZNzsqwN7Ip6yQJBhtUQk1
+1YjYTqTGotv1mlKeEUuaespyR3p0ksDu8et1rbVGFB4Sg/ekeFWErkSUQvHbhwr
H354FED6dTxaD1BE1gcRtpHBqZkTtiqdoQKAL9ktizXu54V3ekAlOiVHtlAKR0DT
32FfFDMd8c/DCBWxwaIFUgiLx3UxK9x4cBqeEkw3J7mMpNrGLHnfASN532MYf4uq
T1ExqbLDApW/f/v3LoqEvR1sA8Godlsyt9Hh98lsth6xDiRc0u++vlXjOdEWLV8N
lcASpdeGY7HALJ5KcDEiKmTSzLyU3oTOOzCJ93CX8OFehybo8v+dyi6lTGJijEtO
+624JUuQthGlYy5CgejjsMRLmCQbFzDy9dsvXbhSEjMSjXBhCAnkuALojmdTc0Fk
/nkoABuWBAeuDDwX1GQDSKZuF6TNoP1UcRyYD6ypdr3WeY5dJnVSb69CQelmOCmD
Fu7TXzoLIoojhtDjpmq2WVKl1U73VeYzU6OerEMnHbwmEhTakyqdEVD2aDO1ka6J
GzzkNIL1OSwzjrGeCabdFVkbD+0belgUaPkrPLCKkXKRrI7tBClBtT4WVwux/lBq
b7YYTY+SVpenZgK9TflYPlYahZIZofyMK7U7eDaB1XOlOpjPD0ZP2eoKLZ8MbETp
BEvrDT3VW1he6/ul6JMtWSzRzlqRm/PK1H3Pcz8cUqHTanIrg9GjfIx2bRnsMAhV
50CBs5xGkqpE37mh0A8Wh4gUqykrZ8lgF0CeiLTDa5xW9J1XGFOP70e4TLnXt1J3
IpchF9gSlDJjqWsX0CS0Whwqx9S6ALYDbcYi/znqi3GK90uMN9usMGfK3CfTv6HE
tk8qjv1NVc/J077e+3Ct0Dm5+Fr4CLOkRQjtrfN1++F6MCu10mfED+DBxgRJb8df
9dHpk3eL6yHiVBLQlJNgk+ypnPLIhwIrhISTSYN18wnXh7mgk0t0YudVyaYJz04M
zqXA504MfQnZ2fJxWQ5dBHJzc4UnYdcAcI4oLxKRqaXe5ZON+kge4waIaKec/E1p
UDMJR5yFrbuptE7Ve8dEpYNntq7Yak/B8vqBwpi4c5rIMMxyAAkYTVetgUhiZxp2
XCiWDqO9djloPRz4qJMj9FAIIjFxLvyjfIrzAHSbSSXRNSnOa+wbvulvtQxAjjXD
m2HOhBX7pWLVcZDZu24BbZkkmibIXrZVwWtp+QGQ8e0Fut83OqzXhRYEzJaTA75d
4hsoUMGNNnVK4sAruFmHzKkW1Q21rLnxf4mTV2xsZSXi3YRYe9dQevr/EW4eF7d5
YFDftMfR1oMgFg/UCvYb1r0UVvnOOI3DF5UhIRQ+RX+fsq7q/PCk4GZvQ7AnUjuA
8XO+qVyVCrSXWMqy6nF/z9epWsceOfN0Gcwj/gVeM0hIzZQ3CFOfmJ1lwc1Esrh2
xwHD9gwnPxEWuJIjsxSwAX+UwlnR1UkpHVbgd0Q+lwV53hzv+ePj1pSOiDIc0JtY
btA3FKmsKjyfJAlojhYP3JfkZGAjFrUfWQiEQCS2vl/3M/HEJOMaRhlmdLUCcd/W
4ftkli3UUmt0e+C2JUbdtvbQTCm+mkx8JQJ0E7g3whPlpBQ5c9lPZ/GKzhyIVol8
qeKLdk7JYuEQDFGPTGhOH8S48NxmJq3eBeJE250SqCk1IherNER095+nL5j1k19r
4wla7NbervVFMY1mH86GbVqr7O4CiKi6TYzXU/szu40oLJAxMhuPF7tmdN5v9oFX
4H07gAbA1sWLQz2BTNg2lqDLiht73FhM/DKCleZ7+dy1o1j8n0x7jwyNYqa2gNQR
5y46GUwFOGj6WMV9g2PlZnHseHRJhg8+tva63umTn3uDDT1nXgS0k5DixHAb2imc
E28r9Zn5mRxKgzGM1ItJwjewJiOLMVFl11W8uJ4nQ12IzBJ8WsNBdbbpuTRM7hUU
M2IxmaAolZ/9RPNwM+GECFBzdiYh28KizPIhIjK2tB7ZtdK2lnNj/uy+gTNzkBwO
GWkZuezf8Eb5xd/twQLX6E5TYhKoio7JK28Hu8shLTsxkaHelSrW6carMXToAwGE
znwwbR/Iu0CD9nL050UGAqKLrnv3QUCJz0ANGva927JnwRRY13rDJqJQTPKZH/5C
DL+FkIIlN7J700kwyNP0x2bP1xF1DfUk79UoyS1l6LZcqRCkl5/tO3FO2OIWRdNM
3D3Bkjw/GopkwdJMvZVkW8XaQyUxPsX6BFFp4R2j6GwsSA5xC9+zU7KxoOLVGRgp
cINfvOep42SWQQjDq0SragCC98nbOwIMJzml3xXGynzODelU6Hvyo9uesd38rhaO
6DxcB2Wsk/qWyoQhLw65x0S9Me/J2i83b9HITrtt1pfqgE8MFgQWzYflH46rJol9
jY6B/Xdj+bM/1ojQOfn+2K2g8wI9oQiex/YXbhyRN1phOju/10dgxfrIrN5Io0Nv
kS4MUm8tU5PQjbmJ7jNgr1ElEgr8gWxcdtpKzzOFEEPxQOsJ+XTaOQT0If6ysJMU
wdncdyUagm10MEP5lkj9PSZziPv1Y+fMGD5aTd4bGLnhi169hZWHF9/oG5EVDbUL
5VF0p22u8s8c7f94LUiGgbXtiMGZ/MBmXW9XJXlF0C2MK2MiB+X9p0oU4w0+wDOs
uTXWMbTZWLUngTRvv4YGyWiZOJ6eE0jDbxvH0w92xAgNuZBi6n80x3D4xZE3N4/H
PL75470PLjRS04Ndi6wdNs9B+4Cnr+vzquy3tNs2nzfb59WT/17evwdSEmvcT1Iz
Wyq9LYzH6xk+PI0FPceWKGacILVblxxsIYLbZ+obikQnD8qyIjry696rH5EqeRSC
sF8fG9dqL2SpJQxFNthnarc7XU5lOdJjOEaMDH/L40BA26N2JxsH8Q8q5uZbGpQM
JyITgd74hT/s9/AFCQLepQkWzkxLlazxtbyvI2BDazGUtKkD5lBrZADInAyQX8k8
Q51YsNPn3nLZHmCxKrEATe08N8TWyBNhgUbNIXyHMTUKDoqgz26uQOPzeqlNgdvL
YiEYUwimRKECmxFRz1jjmI2gVSb/4iZrSO9xYuxffeDsP6pccOdGO5bnw7K2U6F8
C5KM5thXSOR1g0vNfVp6MNTaeUjN7MyA7gXhXQ55vloFHODy93SKmRmqQbB8I9PV
NSuZWHqPPEyirkweGIHE71l+cVWHh5M5viHltFhIJG0HrRhCVNqq136g/YrYmdF0
Lxx0sHeblwaRl/d78Q03dqtT6BUJd2zBDZ+8Izqd1FCvh7HT98x/kCiqXPx8kve6
xzdS2ZgsG1O1JJF5iIMXclX4MxEAyKQWfTlm0vhLfb4KgFfz0UnMbE/oW/QCWC0m
Uo2IF1tDs0896ia8SKVw6BIMjZ+OQXyIisntK2FmnU8tjJjgYyhMUJQ9wffPErBw
CX/12BHDp4u89tXeJrdR1QAazwY1KxK3BD5/UyzqEwGTZKsP/OEPTQ9Vu0e63ZKp
u4gBhOPf01QgcyRNk384xyk+sEFPHnFBT6gEPgdz1EPvZr/HmxoRouUUlVkCprC7
ayBeM4/utmVTB3Mk6ZVp+JefhKwp7QzsFMsvQYOsJH1ctR5Tw+iguyWRi1J9C7W3
YV42iaSf1D/cbNTAKrn2LvU5MhUedSe4iST5Ap2ckpAqXhVyELGKqVst4IZh9jqa
pRwKMx5gGGTGJv9HqkhUzhQIyYplSnCQOQALAra7KpJwLGSkovY/cuq0qqo5deY8
nhXyrFlBbK1dV+1RW0UrSJJA8hrAf4yI2PEI+YAZA09UgncXPLKnUN3yuot33BYz
/Zowof+1DMceLFhxNxVlo2vN2yJxdv3CWMXPX1IkVB3egatdeBFlqfBzyTy5zLMM
Y7g14uzjUe5Se/ZFPPjAL5K1MATQppyrWDGkhz9lT4fGse17Gyf9bhpdxp6OLMVZ
zzVNy6quadHd9XyNbyTbXqtzpUSceuOjp5I4uezAyn7Wb7owi+aW/x533OTGa1My
vy1JXyIdlfcD0axUDFIW7ewLlVUayr4BvlD4f72P0PKuyDb0h9BrCci+9ZMh8Azu
qAOmTjA3EAeu/1u+uPYiIn48f88BMGc4fatPM0c0260efyaJ4xGVRN+HcHthIkwr
GFUp3gyXPzHhsr4kudp4XgtGaUXXTaYlzjhhCa+JGJodb9p5Z9R4sQIMxWKVTRYk
Uk9YixHgggc3PGyhtw5NqKWVkK4cCHTOg2HFU8bNhJ60woGEQ4JRKpASsSd8+qfM
pgDtGIm9nRlqUks5LJn6T0SBTqOoxngM1cLzUSusVnWsNyoRAD+P/VhDz7d0b3tY
UMcm/EoD07/9FzeFyztiOn1KRv240gS9/kh1TjyzclSMvnu/jmAi2hOxuMyplpJT
LCxenHDvDvmOSoGRvgYj0pF63yAcUW3GVatWlCnzJ+/uCxNIrhZ9ZYrSb4w0hrsN
vsS8zhZqxEORq9RMdTj7aXHFUJA3SrS+Xtn36Z8mEp1CEWMZ6RNpaV7PbvR7OaZJ
TB80acgpOaHoLqZlvg+L38qk7T2CgjwpQMlNhhRsyAAft1xZDdxurIPsRCYoPqdD
hzz2LmAqTc4wCuqdmebyXwU5MnFLvBrfFfLbq33MV8gVF7zcpykLbBkoFJS7DR4/
dZm4FZXd7QLAcpBakMDnvxFYD2Mpl3Ipa4igKWaOhpiuzyccxN0zw+cSUjo9oglE
tEnmYHdWS4G9pRWEqmQACxGazRt3pSIhfPw6kDgKs57mt8npxSeH/iUPpqkJfmlY
a7+f+jhOXf4VTcc4cHd1VUFUTdzBYrwbzpCRdX0d/36X68wlMUCtD+BVFlVOIHN9
/iiHy7nqP8/TwqPODRJVfhJAmCdTmninJsX7W8946hKgN8mywxtjB73KQCFzKDVC
qpzmHf+gFzkFeEVU2xP0dLNQKicGWySZeYZojLjMKwiBXSx45j99Q0TfuXVBx6R2
/7qJJn554eABiZrelAidZfZ7yIsy+Q5hpsLaV0NS/K/i3EtyrilSfspWKV23WP2c
U0g8SrxFdIXzkvsVMTSBQmaPPYrUC5c4aFjqKg79GgMl59GYzNGYRQ6fXIu+k5/C
4sE1JBCXhLfjRYaeuouO5zcIAvHKPi4lfn+hHAwKFBtW4nvw5BA0xbOrgQRCQV/t
BiFAyiytHC3z/SQwoMXRx1B8zugPjmd1Ef4M1rdLK/bg7kLG37/opMFjxDfxNFZw
uH0i8sdXZ/ubDUSRhR3Y3hqiZ6VYvL8CLZ1D4phltsGQ16pfE6MBetnQcLIJ2ZiK
sxQd/qpXN9XZLgiLq8lwEJs7o/ori+gxiw3/4rlrYkP/k0CTdje7VinvIgwfKB8g
x13PjcyX5aZ2kTgYA7LhHT0XzKljqU9fZe2wIt2RY0L1ovxjdX6m8Vw3Q8TANzU8
04xVSNgoTc4CR/+5ojVH6Otl1KkJppU2siqhSpi6iaod62eLv851vdM9eYCD81eZ
o2Q7HRiefEkbf9EmMBDAUCg5aZ+0xtKfEvhyvTEHYwZ2vETvlb15Bis2y4i0eFCO
/TLcAATwJIY+Iet7sSoA1/Ta2Kh2+yrmcdiPc3TveEcmyPTU6GHlNPwajmk7LGEq
TfEVdASRrk1tl6M39tXUXsZN6AnCB4wOVOiXJewBA1C94Efv1iYcXPi/GjDirC26
XeOULd/MiaGC3fxzZW9Wvio1q9HHuAgSS3oAvp1hO/fK4F7YgnrPNndE18HLmHAd
tzLQ9pXusbh4anSnXHtNlb5dWPgBXGinSjrkaYfQ56vOlj1zRPgWCbHYIn5yK7OL
eQokYeluOUJrVYEWi55iKW+A+NcTHOpfE6wuQieVjshc/NIAKaQM/dlV+kd+w5W3
nzrgZ+TY3an1YBHpCHjZGqSWolq3v0QuBoadKNhcijevsg1xiZm045b6bHj1eCrX
O5awBkbBRGAXIPbpiL8ns9gzNrBjlgjDaj+jua/5tmqQu34jKCK37TOjK5B85FNB
UURmJt2UbWNhftHSQaXZ1sygEhb0/P2qkWo9DQ4BYAQrxaHgzo0RH7u1rlBLIVTi
yH7CLRuTlhoMlvI7OglTY6+6Vg3qmu/9iivA4x/HYy+JBr89Ort0YikUoWXLfYvr
Ip8ThTjPr2xqiObtNZ1oYzMriYsdnIPSFmxzzcAAsX4TrTxezwowlZG6DejUymmO
Ar5agnUONlwQ3MpThRUeqmRpQFrb6jNaEs8/0y3kCJT5yIBpkx8XdAOYbUOnVbCo
s66rZoc2KCLX8D18UubJzaeVrc7LGehuhHSYTI2NAymXwIs0oNoYKvEF16hJXcGi
if8aWc2/HBTE3aRjJ3UVey058gLCQ/8lrSv8gC2cnIA4nlOdfPFoMUJ2fYASO0aM
wUQs5PgrCx0J6SLuKkKuAypsAOb8wKkYwAwJ5KC63AdBjdVm7NB5lJEySKdvEBlz
KgZlIvpHcH38V8IhlFf+vR7YE/uMFQxVjSlvnJGu8jFsEWUgO8o3P9nfCdTLtnsF
AXKvwhk9LuVLBEFNB+EN10hy5l4IqX6UpQYl1FHizVLtphzi9OMo2txjNzbcJvJ2
mFaVJwo4AJ74rN6yVZU0BcviU7tPLirLshAK4OhZygtWP92Htip4O3gAhJeOibhd
35jTj7xDBZ/Nesx3LHQgnKfUFv7iQF2lWSQPpD/L4gGWKMKDtZPxmpVuP1l23mXc
2O3TT/NiJi79ZUwpkEhgsFlHH5jzetmvSVpcDPLQCWl6YiDMvdkPT1yAvNv1jOQY
y8JqyDR8J7ck/klWc+29jqcJ6oAGQSefjvAQ3ShQON1hIFt87csp0DRf48zNbPNA
uol94tsQtcboQ0QyZ3EIEJSuyK8ORhNIb4BfN0Tp5uh5IMR7VGOOtWB0hfyTqhQC
UdEnSB9ZWV/b3oIbudGDyQd9Mp8CSgC9GKgHPcKoI/5zMsajYbunx1EUrASfSlQr
32qAyLis67+KciNdAqKcrzeOQgitsgKOIcJQWMd1Y60Pezy/C/vLFdtoldld6NTT
Wtz9LEo+Lpxrx+cTDb8PGhFLmtm+kxHCYZEDATj6iO4iFLUz2ivWmgp6cAfXWCea
PNqAwYGSnK1SeD2h42oGvWdMUp7h5r2JB2zYsn5bIt0e/jWjtQgGGi1DCjvtk9Rt
Uy7WynRQ2nT60QRcFvkpTHRpJcVpZUQtT5Goi8N0XVR1ZV0Vb7tr7iYeWv2muzYe
DyZXjYf3mdBaV5TfrMy+LtKYUtizijQ9yGOcmtlv9+vz8xwWGQjJyEQxR3VUCStE
/cTlt5EemZCJraW8EDeRf1cH1q09wP9i+nuBSYSfjkyJE34txWawaciEAF9jaohU
49SYhUY/XNA7dIl8aeuLAfbrcY4Zh4vW+MB2hHfg08w8ZerZkzdf/hdBHWipeJHO
2v0IIagvpy4Z8e30sR7rsLTZtYhf77lCKzzB/bokGczre9zQyCUGTA1TGeYBBQiq
/UbRbltOUy0MWieVcFaG/QRvn4KggFTTkioe/Npn8f/JAa+CJBVG9yT/ApNP3cuG
8aJAivANK7O1lcDm4OxoMTMsugoNDDCES7EmWY9Uxw7nWn5Jd6r0l/GYicviZIeQ
sfNiCGQiIWbOPnTf/0JJ6w==
`protect END_PROTECTED
