`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4gVh+heLwVIg+eezt9jsLPtb40oV0836sNfwGeg2hmD/f9gv0byswpdE8Ux+iYhb
fDmTMci4eTMges3kvLU8YaoP/UAeyxIpclfJXuAuSzz02hr1kMZurqQV0lkqVyHM
VBmuDtyn1TIqNRKyR4lI6v+kRPV4BJzMmRV4woZeP+iNcDlqvNcj+Y2i8kxqx5oH
RHxYDgVqBusr84AlI+sn57ANltawC9YDxS8NVp5bBss1JBNImLBNw7dlwJi+iymL
voCYrXiEBFF4BwlG2bNN+F3S+rKlN6QC+uSk43x+L5/pntRs7D3klRBhkkR5Uprm
TenfLFocQt92nAkyEEt9RI6G3WizBsC+gNAMm+Hfxh9CGHS5NSQ/x8f8o6ncJuBZ
mV19doNTEnQYrme8jDYYRqQ4dhO2rvM3MvUwTdQtZoI1n5HbWSfjG4kuKYJqS4I+
TjmZ5KTQ44W5ETuxEjY0Yg==
`protect END_PROTECTED
