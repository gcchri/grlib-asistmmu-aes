`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OZlx/y+QD5aARoqIFeVzg8XNMZ4FLZTcysaFM2VYK2p2ZSHh7hdTsEno6kIWhM79
MkajBph96ldGXSB8xeofYExtaDcPk1Y/JDVS97CctDDPGTKVhsC7ozCwUp78JCVF
QLpbdy54s6H7xgSbLIAOGyIZ9esJYUKgFAD7y7jh5mY7icSdppIEYF/+KHW3NzI7
WIYV/K+aM6DCCDYig641k8JrwA2Ty77iDn06rwtYDiItXRwM2irwQ+Vmw3NO5QBK
/w9RhvZivSousvgBHtUz8LXb0qSAM1e/f4/j7x1zG0WhxIaP0IN16nhqRvwlADnm
35U+n/FNNk55DM3Cqn+wUu9J6p2zUiJZlwaw84cK1NvxZe+qGTZKJ9EJyiMocFPw
2GfeM/x33poWCOVPu/EAzeKsnnQF9AzU1j6eMekHuauyfLfFrkjQ+YAFhe9dSghO
ibybdQoRZa2MSEuz1m+YFoAcSb8wJhPwKwIt0WHbHlOBlZNUbjQcWTzEn1/8ykSU
i9Oh6vUmXH+eCFHWvF3m0UYm9y8i9ZwVUZbhOVg1lztsx1pHW9HqqtOQ6cBnv378
bkYRUznICdW/3Bvx41xwn+CgF73f9ye1Gj5lcae6Lx2o6283FNbCDVQIsmrIQxsO
8Z60GsW5RoPZ0SX7e9JxGQ==
`protect END_PROTECTED
