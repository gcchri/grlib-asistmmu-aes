`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KtC+Qdbl2mUC0ebZXGanCUVgdqwa9oQz/wwnwIbjkWnbkral6chMiLgsLxjAKEfY
ArP5Owf7wBgUBaTOc6TG/ZnHti4683M6j0CamcF7zuSRJhZE+yaS1sW93H70qP0v
MsJ6MfBR0Fzj43qtnsv/T1MOs1l6QsPZ3UtpS/fJ9jNSYPnU4eiiaLSbxaeJzjBw
+gxB/mQbWsjjiqOICjBSxXhhS3oQz+BgCjAeoZKv0xQRL/iFMLEPOg4kRuHF1Hno
1PnK3UaQ4tNDGdZ9GqN/vVK+TOhqMOXeqhNFeq45pcv+Ffqwhxfe8aDV/rcZuVVF
BXczQNGH+sU7M8kUYcjne5DHV6F4JYYD03lNitsyFHvRpavx12OuDUKmPku5kIW4
x1iw/DVAlThIeTazrVXdRqctUoNZKaHlHDvhGcG7QwZVAK9adW7RfmYrU0rpv+M2
YkKMGTZZmWPMbps7ySmBr9Dxtzx05GAzmp/JTWfEhX3hCzrp/dXRchsJHhihftDH
`protect END_PROTECTED
