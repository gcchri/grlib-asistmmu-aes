`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b8HqX9vo4+qcigbXF/kM4JgQdTLj7JUQqJfs95LLgcltKw4o971IsvCW2I1aoKiE
dgngjlSNZ8frcLqqjJfeEtrQya8EjLfwSAraC9/DROlupoaMUSTEyd76sK+ODG05
YSqsJToPRtfnGzmtbEY8TgQkIX8dbnQpv9Q6IxB5EnhxBAOrXjADfa+y7lE5MPSd
3QawuN8LhW3fLLOz2flSD6BTZw7y/KwDopfmFY9VfrGwVEJ3QwoKWRv/tciw+Pwt
G9I/emqJsZvYZzD1OR28AOLVwdm9dLtttlCpoaIKv+6g1WvKgIGIelvcmZmfD+xv
EYYKntg+DU9o4xl8SHoIEP5EL8yYJXfGkul3Mm9fNkRQqrH2oYi/FZkzd4c2pWdd
y/FjSBz+N2tUjwpnPNRUb2k2OCddfhKoQwniqRQHaH41uYyrXV3tAmOmk9HWb0Hw
Vwnxw+2bcWDcMOdFMil9OcFUrt+ps+kb9GIEPkKPt5tmALZGBnCusx3ioxqm0eUi
3671aQDr8d4VJjjwzCXArEZ9wJfgEROj+QtDwbbZ9DN3HVsjqkEZQvruorRPE6HU
ivYU+q+qQMiCatOH+LSzTcy3qT0FV/HqaVTqET/jB12Pf8bVG6MjydQ/IDwzUEpB
AhRRmCEJ/HWwLI5L8VxPyAFLkfxWxxwV6Xkx59Sd2wfk7fZh1I47aKcbM+AUr2SG
9i25YBGI0rFyQFf4R1EruqesOk+V5Ye5UvVYa3YRElSO1V+SKolIhjQtgeq9s3qz
UhV4+SQISzPtAwpUrIeKmcTnXZuny01PjZjCyVSJXmMjtbcWqS0BarV1B7ZTWAf3
7f8mTzWsTFFbAtCGr2b2tlM2voL3YNqHLbZQI71f0rEGPms9FN8iqzjld24f8N5x
TCFHxcTV+efiEocv35fCkNnu3aBUFKw9YDaMXFm6G17SCknsCXfwDRoL34ZyOFLS
MC9Yo5ZCzkTqgL7L8RledtfjxVqBhoe+RVQJHhN90F3In9dpSUjafq9h+MZsucr1
Ew9oz2CBUygpWpWWAfx8jPNRpRo6oZqBf8LpuRAaYqTfJT8xBHWH3Ci2+xbIKafP
di/o2YhZvdsgF/QlKoVv3X3SqYBXDMZzZ40iMLqFO1A12Hw70k5vBmLiTZZwfj3T
izFgpLCeJn8EzG9g/fJIGovyDHDASYGL18DIfZ6Fiw+PlVuGiWfs9KLC2JogaSr8
VRNl4TcWx8S8Fruv8m1YwsBNrEcdEH3z0Wbq7zRKHVW/pjV57uNqioo2Kuig2frg
TEuDe2rTjqGmuYtOOoDHl/7Jh46LHaZaEFa0ksBI6l0/I4QfN7Q9n/a9LRfteaVt
CV4Gjkyyad+wztETRTs9vBSM1SfV1SbPtTkuZ6UdkXgiJ3SPKlbarQ2wOv03gD0H
Hvk/9v0ehnkHFW547cC8w+/BK+CLue3cdCWqAg/FTCBaLeBd+3sJWMkhLIQmrL1S
aY55QCWnByuG7IwRbwJr1df9MJvw1wQ2Wpbzj9PH4R9PtskEEn86npfsLbPPycDP
C2tRIIWhiY+Aewmstv85gIuStwjM6wSXLFzKXI7u+RTD8+plj1YX5RobTijwFxsz
hC8wKhclvMi4iBPy5xHPlNlDzWv+oOul3vObOYn3ldQgXG36tfAaF5mVL1o+v3E3
VwkxufPRjFYggRXFO+e7p7YevFM7ZzIuDCpOOyA6kjJJQHBOHtrKApTg9eAGd8YY
I/TuFmL6uka+wQdNBFCSt2PQIY/g4hz4YZ7BdwOyLa/9Inxg/HtSZgEHcDbyW8UV
SvYR7TzxyJD9v7E6PGop4M+GMaIQRRfyx9m1QB0k5z7yoIm+r/luG6oMmNHcx4wi
x8kr7v5CfXQpzIi3jkSgFlazg/kECN6/UpHgT+SKUxfkPLoFsITYDrlZRWDlF8+4
5M7JYXX/g244m2Ha7w/uSJSp3sFRVzq9dzTmgzVmXj6s5iJeDWCQ8m7H3G3YEfA/
iUzQn9no7eb7rZzgzkYdrhvOfIZcANwHaKvFVYFOprNq7cFzVlWUfgqbvUyneoBo
NRD7aaLYgDMr610CUr6tNUO1hH18zBxuQ0Dy3nR8tBqw8slbibPf45hEsVWmm6k6
YPIwlvO0TYSDvJ36+sYiVPA00FPDJLsushggt2glct9VOb2gvGWx6UUPbvQrXmpC
j9FErNaarMBXK7erGvlyoPqccur1QTXSfQAw/FkLBod/juiWYTVP58IjNxFb6PRg
1DFssERr3xl8XorRLozzZQ5WLS6uDpR5GgzYAbVLrUlgwmnp/QYUsWxSIJfIdZuD
8ySketI3O9G4OjRGj3A2b4EsAD5mkrYFoI2fqNzX9liL2wHZFbii2cf0CnjwkAIz
mcMeIpqNcrDTEd22WwHhAfjXEcPyb2lYFPOvXIuio1hhUV++YhZIdAs3KR0h5F+r
D36t/oVpC+iLcUuYKNQDs0LKVUj9dTA16cu/FSFOppKqHax1FAHpnubEMIu1zzLu
iaW2KKAtVmtqQB07RBhFR4HeG296IlsdPf0RHxrq34npZe3X32/p++eeSH5A0SUN
lfR+JT77E4HZrPpB5iEH9lxSeX/Q2c01JvOWJHIqnto3Pjwm5FBa56AGX+Hrf/Le
NwXkIzsagbBR+MvJ3Be0kynaQlK7YOTl9hb1p2vhX2PKJIiNkGCzY9TB8UIaDgnN
F8f5yeziLmciVnA/EKTQe6lxpSdIImpvJ6pb3ygXrNE/mU3Eh4SNTu3kz0XEVpu4
yYKnS4l6abrn2D0FOe7NCkXvjYyA/D/0M1hfcYT5U8A63ZbHvGrMYNJQX4jLtwuF
RNPK1atc3w2icAhowGNnai7H4LoZ6e7/sY8VB2uyvQQ97NwkZVEKLzvFBEIuTEag
coQPpqNv3IXVDDk7h7G8oJankVehyLb2TIQnKNvbErFt5R/OLb1nCjHYdssY4gDp
u70qlJuEsQXhjfYZwD1TGT2ym8FEtVpuNqcXNjEG557oX1EYNUetLEKbBEMv8WC3
Mzm5oS8x0xrXoFii3+pr66A3YT+sjnZDvbpclHhWAzFSYawpxwCHcylDQ9Ir2ib7
IybI1v1Xev+O37wG0UGTkhKut9a4d+ni1CGvU10QEypvXqcp682ZijGSmPCsFmqu
ymxunsDKCAmFIYnI2JhP2nrxaesR/BqzbIpkXXTHyYOnJXQkw599johAB4Sus8Lw
KKoWHVmfjmV9Rb27zrYGnbcYlsrYbZn/FNLzWRwyL8O7ug+zV3Zg3PmO/s3IUkPz
XQbFZ7x/JySVTf07zIAUIbWMp091GD6K4TnYy/StISO9sR5qgMSG6cMggb3gzyRJ
pGXVjdoRzVkLN3ybsyKO5g41CjoS24loxbBCb6po9pyhF+mTeBV0me85Fq0BSRP5
gAjTBi1d6fY7mAAOjjwtGzNJxaY2eGPCjj3l9ZGB/eoGLOfYLBQKgp+Ct7DLvd9+
8RGY4v0tpJoUQasBkDSapAz1y3HBiqKZzltku8gcqZa7jxP+iZW3ZubeBoPkAZGj
gyjQdomMy1o3xL3FaEMS7uPze/NkvpajEsr8xeDekQozii/1mqCz7wPxbyA4lcx0
YQYKr+GLhqi6f1wi6Up5XuypiNoy5No6gqslBsfwtilyS1Buh0c3D2LDw7AT4NC9
8qRk/C7yG4oBHZsK9K2LXhqeivpvVSlxZalhAvhDctAWFP4eezKBXtzl0wH3c2z9
mEbcLsoTAwnJXf8PQiyAOLzBBTEN8N1mcBdM69Uf0xB43hQC+gZwT/bKiePx2ss/
wYFyjOIrbLdtxZX2kNlXAP5xvIdVxBzM83u9mmbtQd9VmioKvW6PCgAZtd1os4G/
n+qk4nCP2sE2euZHW98teU2niQ2xLS3N3pbqmTLz68LG5vbh7hxX6D7cDxjol//1
0ebENw6o1U8295vK3AsVnflhElnFRxsZJhNW+TvabNpzumteVRjEg5GqbFbi+Abr
7ABVIEK+9w/27pdUtFxLM/3GPFpjEqPmpEpYoBXghIigQwQ6jRuCOUTUpy6kUQp2
p0MfybjOnhw52yJfrd/DfYjAKa0j+9wD3c7yJ2jX+BeI+Mv1TI9LjKnF9/qlqvbZ
qCXZGGQ+DJTGawsuLIEonOYjDwJdAiQ2/Tqkgwyl4EbUth6q+3xj/wOlfOwmRzNG
LBbZTwmTeP6VXsr69PupGDAb5kbEqlfOPoYJDtKTx40zhoqLeeadVOZEBDRNcg8C
G+1C/jO8W/bM2LBsOd3PwkxmgaEa+zd/NkGNsCD5Z73/Cas7XIvQIslg7U1f0q+d
8mqIM4xwphB9ddPPm1O8l3QNUw3Chek0nzV99sBDAnpi3UoFcUMR0oQQkeORjE+C
zrhlBjBT1EErZWsNK4GOFmpxYIz9uVFQFQOb/uM2aTNEe0Mhj+ioKd2vsrcWfcTk
tdBbcovfvd2d7Q1rW9ElOs/MBUQG1PQNo1/+IoHiJWjDU5bTvrCWh8U7WqBZQA7P
QoKQmyPRuDiXSt0E1NYiFANApQJ5E4fLU2Sk846K8r68TorZ3NxaL3vojaoZ+5GH
nNQ1WcgbzFdfpyqBt8QuyzeUP2MFJrJRem/ZP2U2VLU4G/kg0N2NjGeNMuevMPRe
3nZqs9mDq0RdQWdr8hcqKAWHiPzI5tSAVHLHtsDOHht2G3rTyP9HjuE4ud+0T2+h
IAmcylrF4jAdVOV7EyCVMellJrImAMMxpzWBDQGiMcv2xWYOVcTICCHej2MJvFvK
4v5IzccvObKbdHyw2R6FV7uYxlkUiZ9D22qD0KkwcPyvCbMcxt1jWJ76zDiFzwMf
AM7/uJY/dtQuK6pNAF5CRBcUk2ZKjHj+srTDbwti9GVJQAd905U4bZMSlmQptQLZ
Lvx+jHvYo5nRkl/ZLrtLjQ16SwTXvDu6X65MjSRjRyVFbLJBAt/Cs117417vBSqv
gPn4FCj25FeWhvJ7b4BuNx+QzmSKFIfpe40SFgTfmMcB0GoVMZV3cpvLuXag1liI
/c29xl49T2wTgFfjnTvs4k7uYzUNGowgCAU3kgSMDgCCo76plLTkHUvtLG13Y2Ga
5JviuBoQ31lldTBcYNFEq0OAHOPKkFSnXy88Zh3uXiPiNe0Qle/PTiuCY4k/uWPS
ewwlO/dF95IzGhpPfrjhl8OkTjaHhaUPRXU54s6BkiZxd2sAvsc0a6GsiO6Hj6Ct
+TMU73vs0wJBNCWjA9+Z/PKLd6MPxb5ng15o5MaH0i0nY3y5uF8V2hgjEQchXmG5
gnlIEI6gwui85ymIYrsQR5OZRuFMUf8A051Ep6GhkHmVB0GR6k77jM5cI+ZPaTgG
nNyzUAadeNpZlBIpraVX3kar/hQLtrtxSn2TWGtA9NNPrWaHnw1DKawUOgirBY1h
ebvJ4wGM9AB0VdfZxyMdT45q6lvmtAoeaOJpR5PS/U9ZBENUuZAFUUGYeNAkTdHi
l7j7mBWzjBM9jWZ17G4berJy5eR01VGMLLtGsui2VpIkXLLaqK1E7nEKW7OzqyQO
Ow2pkKONPygHiE1Xr/Fu3O0/hGwGkcBrIqLgzkZFLQBWmWiDCXgH2GZUtW9Jhsiq
HjJBXVjlNG6FoDDFEzIE/wm2gUrLDOuM/9YqyLQut9BmWXAzpnjMYSqkGWyql7YP
szNtUwezjum8KHWiYPNNs9WTJtX+TTAzwDOJpjgAdPHIjU7wOXzLZH0OCAGrGhXl
m658ht1CqAqP5Ete5LomUqeiAddnKo11hhLH5+xuyj395B8V1oMG0SB8YRJq064n
GsqlKGfEumzRWtS5SBdwSSAhhggWeZmkBPnR/XhuVwNmmKN6WHYV3pxPZ0jH8Fk6
Tl9zDEi1HSBbcKSu7P5yvtzpe7Azs/NX/sMm8TE/ZjGIvBEhDWD1u+YrDXL7N3R5
OdqTaGcteiyvk4CmgszUk97RWGfzKaNUspotxKLOZs6MD9I+QHnhSvEtw7DyjqdA
LCVygFD57trBxYdv0TZOy2S17jeZIagDlNXVKgDwvAjqYnyLeveGwok3/yZArxtX
ngJfE/++vjEJZd5PLyniaPoSyY50+pMUv627igA4Uk0QEf/IktOKaafThl07Z1Tn
QSlpCrU3Q7M+cvkPuzsr4ddsEbQdxl1Zg7tyz4YaD+y7u/F7IJ2+ajR568SwUUvH
0FLOu317B/tOltmDpoc4BglqWfyIitlCvyP49WqKC9RFsmq7A/ILib8MnPsuBx3g
dyAJqSIx6W4A2G6q03HxqOQ4f+jQmpZ5s4wcvm4Q6rYEnB+A8ucvwE4Qc4B6Cj5L
Fhggebjv0vv/8L8RHDkqli/e4kOX3nz9/Z/Ktb3/8dhx3KldsyuawI3kw/DSjGA8
pTuwuEpAm2c3ncprX44z0zc4foyjA4/05+yEm9NtI/slKONs7lJb+oKHwPRfRj8Z
mywDW7fmu2DgAqnjt5Vszvi4Y89+Un8pb7UKRJT7qFgezUeyunQV2cdZyhEFHvIg
GERUI+Il4TXCqW4CELGsUOdEI6DEKlPZbJDTeUzTzYnROdiG+6/I+CF1Pt5bHVdD
3CZQbobfU6wHwxaT+9RgKDl3hCB3pAKx1dUUKKKDfdk8LpUx4a6CpFxbcrmLNPVS
V2HHFSAFWGbmF2dXmkYfcQ92/K/Ibn+6IcVLdc2vtBKjH9cHiwknftezZlzLY0Ze
fR5mS4srqZwzZ+/L1f1odkdW8fLDOCoH4Tp6CYDE0iqW1nB43Z9munCOG4EKRy7A
oLIaxwtsd639xsS8yDgnadXa/8oALGPfe+AAqLPZ/CQK0kMmsgSrU0iqwvUoH1KW
GzOKsCDgZ1xk8UlMhqoEZhMbMeae/QEmBsR936ubTtPxDDvYijytxwkn5hthK09c
anyyAfY8z6AZYad8UFwRWvtodGCDRX3e27w8RlKPOwIZLg7EMyIie8b2r1t2ujP1
RyEvQ5kZ7ZvPMfX+c9AjqkTbmCFmxZIc+OP9Kdm8HKJnCTE5+MAeMgwIgZ7+TLyN
HzEIobitv9bxRN/YT03AAFhAZ+MZQsRev8+N+plQdIvb/K8p/+27xpHf2AdDHfFV
1dcNW4sbDzXg5+RaWKq9eSWv329fgnBjPB1hw2QqLWIP/tThePX/FEtTFKaIncP4
KQ3Dwj3FWYyP5i4lY/BKPSLk2IR95NcKbbRFO9YIc30XlXVZ6P5RLef8GdYTB7dz
YHxkNIoo06g1eXyAd7eR5j/iH3eKW8/RVtF1zfwHBoah8/R+uH0OmH4h+YzAIYNp
cDgYNK+Lc0NljvOMaIf9J6R+dJYR7pMDU4H/Y+EnR5uZqN3I0crS8zhfx2T8UiA3
9042+vseCPvDdfVVXO9X/8pSbZ9VUlr+sMdz5eqnBhDgdekzlwmEAIGrS/ChPbjt
waZM26A9FXhO1GJV/+qMeTh0fZgdzy2TqDK52YzIF8EinoXVjl9J9CEo+cUNmWZ8
u2RWeWSzHyvimJR8BYNW/f7MXH53GaSv//slaHZrZRNcx9FnD7iXVhUAeefn2HBM
zy6NBL4czo2nBx+T3N3OktmxZGS0wNmNi0NmlkLX73t4gBZwWePX31YFZgSOkqbB
HOR382OdD8cmx6Eq6CtBMXWeOFD1CabjFIPUiAoH86T88HdMlp5sRwu6V5N6hZkI
sN8T98cJYKZBVRa/cV8uYGT4Lrj7TkU1zF/6KB+tEOBP0ik1T5bjl5z+apKos7sk
6w3fqiq6xYBMgisZtttLQcjFDqyv4ak3X/KdyLE4vrUmK7G0FYt+lm7RGJuDj+io
9O0wV9dIXBb1PJPslT/79g==
`protect END_PROTECTED
