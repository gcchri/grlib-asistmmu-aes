`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zUy+jFdYmCn9vfuRXeZKML9ejrobw8gqKyU1GJ/DcS5VTStuwM0l+qSlz5jWgmxY
UHA1FpfRdYQ1Ve2SF7zijzM3rVp8UfNtE2MnKFmAlfE66vXnTYvVQ0hf+8mWsJIE
xqo84FKHHKlxdzgTOONA0tDG/tJX/5LFDr3itx0rv61p7tOla9FEwlcq8QSOQFGE
POF8etPQxSgZVZqemnSBl7oR2/XSciW7h5qkbrnII9vmzngf4ZZ1BBAcrbBFL3ko
PH9+jVsDJREPppwaKETzZAhna9/u4Xy9FBfIExOQ8JaQaaTZAD+skUDYmaA/nsCS
+SX2o1blUX8ISoxdOZKJspPdEXJwC3ZCNH2hvUiOscfUira1Uy3wwzKp+5ks2GwH
ctc8fSpNJE1FuJU1Qm6Bu9+j9EvGOXe2sDTLc2FcMwnF4cXCJideTbQ6n4J9Xc1G
+0jvGJFQRabN0U9HWEUeKdN+1updJcn1HJt/auRcYhzXeRcUgjAEcfvvoY1gElgT
1J834PyBfztzFSpoJXhFrPE1IxiHiptuEtiZVVs/W5YkToM8b7dWFHmLVsqPia1f
JHTAlfKHxHLizlRrivwGfAssSXZG3DIxTGn/72ydqyE64QqMHjawLtMeG4Gt2loA
5UA01YQckK30BobwLJB+tS2d4DS+8U2ErtulR095B1903gzuUxGYPJXzT0DbPk5A
Quwk07efxxu3RGMn1qKcaJRe6YWr5UJ40N2dehGH5b3KtlHgzwF6u29rVscywdUv
lZiR6Q7TYMd9S+bNKUeHuNfbDCa9MKP5fxwk1J3MYkaGRtZnnjaBh0ZwgHoDnirK
4sndN825k2JjGsyuugFKHiJI1UcgOM2T3E6oEAH9POinG6Hw5i7WPZazLnDtDxee
dC34KJeCToREuiLnp+9x1RtOsmBRe6sZ/PiX3xfHYWFZcfaj5eJ3g/EkjdgKi7TR
7+nMvbW5OFq1TN2Dj+0xkv09JMueQhHmG8bYGMfRgpy0wGKL83X55jm8bqj6tkj4
J1/3H3uagqY8cLPuzF3q8Kx98mg2KwJmeR7ueEd5Ad7pmGMouSKx3/J49g3sKblp
SDtf99Ip1EE59A2qKgx3sNRHuZ52FKxch1/JvTndh38jrFGReW7Hn7fN7KWzw14c
2qcjIQtOyzTISampzXmR+l+r4HCGtxkaFrVmHIamLwY9/BdP/UqcJ2kRkxRXDN8k
FypWjnXf8m8Ica5hPsz9w4thZhzMTlkFkC57LVbtZq4WIHUkIUO0NNynF0uSAyov
F39/s1iInopl9hI+fbXfRxwXT+oG32SfS/a4rYwkuQLVYEuGeNDC+lpDWiNm4bpT
enZwk9DJ62nobLQyvAT4UFL2hSyrXA68Ev/6KSSdrzOpPAXjtBf7a5c0vHGNWX/L
hhs0Gpjs66Vdw/mkGvXEYVbeWTAs7OgpzOznF7INCV8OOWH2FdtISr2fQ/yr1pmE
b5ok8Q0gj4Dltg1I09H49ECTqxCbIHs4bkL4vMO7DPYWmm8YUQTkbqlrAWnAfCog
RLhzQrrjJ4M3yCtIHn2aPMw6L/zZLarCpPkPc5cfMyM/1NpReaMadrBdz4DaCHPX
MMWqqQaZZm4Bba1DT6rr+UXiUPqBEAw6LjNfT4uOY+oQEtksc2Z66myOJchZ4vbh
MWTNyw8BKKeRU9iIotTmJqvTrtpm3N2Fp1J1rr+A6tX5kAuVyPTTB7ZY3F9sMj9R
oqb9cB6Ec7zay10pgFULsV75dH1g0KW+pNZdsUnZPvYzcuxXdaaSZ0fgifmYTGPo
Uu9UmwNIB7t9t3UcMykPPl6x9md+AUwZtS6RhySu4gfBROHUnmDi0oKXPpZ0VSg0
xcGL+HW7s77j62Wqqu9GVAaYXjCeXs23EJ+qysGR2UpQLwF/Efspwm0WLHX69rwF
t7RshPbkrrG2Yw3GG1glEgHsQecyjOO36UVznKRUmAGheQ7hI00JMwgAA6KHKcmZ
mA/j44qa68JaWwmyBcaRzg0+pTu4IGsIcOqbufBKptbbvA+/HD+oN+YFygxir+Od
Nt6FlwoOqVHN74nV+LcphT2ylMeahDZ2MFmbwVJh05v9js/xiYCU1wRg/QdB/4ro
xMmt3s0IFQ/fkLx1oqcVtBMj/OG3UX2H2kIpNGdM9IYtLF0IfA9M6x4o/a4e1JqZ
flxpU4/CF3RcMkS+i4ISr1p991bsIG9C6wf3KICAJh+A6v0NpLiMdyC0vGKEg8yy
vIHEUSVNrz43VUIH9ibSdOu6aH0yH+AywRDAJ26mfOk/7Jf7GS6ygT+sMkY7dZDB
NQrP1Hu6I7l21nJbXCLKaC1IW4vH5GLTsAFv8Q1iFZXg8JanNqdXR0qKz6rgmzgj
VGBoZ7662LIrxATm8/otzq06j3pHTy5J+uVgsEhYs1qXurG0ZJGwJRTtCTbolRNS
7R1/48/9lYfwCi4M0p3Na7foeKf5XwJfEKVl0swsus7Seo8lDJUeaKny1Fe1I0Xs
hJs9cLFoxhK4xoajj6cj27N1yRsPYXog3fPe09sRdrnDxlKh35I/DHqBCHvW9w1j
b2GW1jo8GOmf+b0yL9aGNhCEMhaToKHAECIOU09px05a1LMBVEglhJLJ/doUj8xR
hXLPpbl8rTd+/LSMTk9bwgBzL6uE3/pvH4kiI5YEGjqw5Y3rFr/9AVthJP0fD9Ok
ajHNipH9cEKaloBxZuY6jDkBsZS1VT2aFjDkY+FcPr9BW6JucOapg0dDkretMwWP
2LuEQv946GWYAumBV3ihAqmui2225AurkOygcoyD2Sew2MyFAv1NOI/MNBW9fX1E
NA7C8Tsc7eK5ZY7JzaMxp8MNhLdwwuUWuz4zgRv8b66jQwDK4X0JRCFUe3ZJ919F
c8aLcP8ZYvwa6oskVKwNExhqoMWrzA8auCd08hcgrYnXR9E5Bz8yjxj5pND3atwx
+NJCDEgQoOj5eeQYmked68+D2kKi0s8WL19UEkupi5rOUyTMoZ0M4vW6cz7r+h2e
msLr+wlbNfZVoPVJyRGaACel3nGcQiMocEojs0YOVh3mK6m5W32YnLUpenvqRXaz
Uiszu5ct3IKhtUbuxNefhn9/PpGvgg6dRLwc8BZPX6ISLh4tJtBcno9Ku64jCkoD
P7Wc+J8xfrriU+ZJYysREv4sTny2Ta0XaNJumSk0VIgT3yeGQDII2ExFQiDPQwg2
KSHAFDelX+gl+Kl9qFo1Y+t3SnXOQwhGW5q57gIAC6pE/GNt1+UCqx8lacVQOebG
K/gcv9ekYotpkrGPFJVznWUEueOZGzGzmIXeuF/gOFwKir4K3R5sEcmPOu45z1Zt
LsQ/GrOhPrFPXyqsTkzB3MLV6YY+qm0AutbwW29SmCGSZnz4MoJx+QbbMvF775Re
EIXVE5KUlIhy7wLup3Wap0fUgijmHgzaS7CP/OV1blLH4gPe7zlKRf18FZU1+agF
Wr2Ntv4mnrfLU7Nhsvz2BiFa4F5zABjWyZWbA9z28SX0o20zzBI8n/IxZa88oJ+7
P5dVI7y0RytJ7peK8dYu6F6pRfT9P/NU596BW2jJWEI/blaLt3MJpjOHMQ0zmErG
y8lVBl/UBkWlP2VxZscRvbo6ARyD66ipHJTJCqL6pu2Vha7CkbX4bXtfZM3gVsW2
GyM0kyFlXpR6rF3vjQnbGPnHIiiviX3NjlxldsiNYcWsltxJvXPq/0aUD60EWeDR
wCvUwuJTc48EutgFV3nEZkgAnwEJzcnyX6JcszuBPNByzuOohl/aqAWz7fWjjKpN
Qp2cqsUiSaG1mnoX4TFDIuZp2zbDcVfsC/zWQkffAxUQooicoFhje3+s7U2Dw9Qg
SDpK1Z5K50khLQ+tIaoMDrjkY+nWmixVLI55/vqrBgVY0p9G8pgYxJkovdOwEopl
NEpBnPT9xYbWndmApBHit9s6UAcD8Np8h2UJSUnzN5IcW7pP5kmPJXlnU2MGcGci
UVG42DAxgNTkOsHK1ZnvGtGnYAuGEoC0cP4Vw0s3/PjgCqZUgviicPIXkx5lP6UE
4wAKJok8iBUVkNKb1T0b1JwaT51IHYiH1F70o2xtavGiBN8yYZADIphyqJoHrNhq
Wi+oQzfznwL/cuewfm0PurEkYPtW5f9qkvrA1F9zCeaGz0SOKCVGKPJClNahKrwu
sTbro4397fEu4OuiNyZ/L/TCGx5XtvfZ3uqJ4U2pLH0HJuwyA1IcgCMMqA9sDJ9P
Xi00M8U+VoFgB7uJgjf62+r/126TfY+yXZsDZ/oyXvSyH9Ckm2sMHh0GM6OT5Jzk
veRCTXtakcmTiGU/rbCsoLC6BmUkAaEeVfuHkFnb12kdLax/p6rnTFxPjW9z5Eyg
81pFExBF39N+qtlYHaTJDqKsdF3iy1dFZYHJPGjmItKeewQ+ko78KfnyepHoNp5l
XqcS7r7pnbsqCD9U0FnH0fGZiDdP7PjoMZ0owBJC4vDNDV2XbgzPBgl/IaaCC5hD
8/zXKPkHzBSd5Mfm8ONeJmb+fB6iTC7mbmMnuTSBDCIchrwPNDaWYRSW+yZkPf3+
MoiA9vAMc1oHvfWacEWzx2kwo+xYV3jKkAmGk3mnFMXePd74uamHxZ/6pqyawdz3
xRkec6PjovQFquXntRNTyKyRH3gsWlbTgMHOOxfReefUXQoEJ4EAM7qqYI8ihvKc
oeSDZsUMF5FVjEC3Ma3e1+JbCvFg+3FCgZYyB2XbXV82jU3eEApKmwHfVAWUDfPk
EKwvG2irhDECq/3l7e9vBn+0LZwi6bGv1dHfOAmnXxI=
`protect END_PROTECTED
