`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wJvZq7DxAEKzw+XQG4N7HJx2uE6PKIQJk+jCWQNHZwvmBICb0xKYvKGV9pOMXLqL
HfAI5wCiU10qNHWNoPqZnvndTpD0vbzwe4tNak62ZMdV6SMyl0FGMrLizbUDB0gD
koh95n5CKo9KgBCqskGFiLoo0ZBnd7wP7P/8SrTDLpxFZ5LxGJUg4COxxpc/MICT
eqeV9SDbIhSSjwQjAo4y1AVtywr/XatgAhiLkTVxnL47V2IvNQUboTmS+gcx6WHb
G6nzzBJEEGckam6UAcHn+j1MZY6lAHVSVnT4uZ9o1R9xg5W9fkVi3erkgO+U8b/z
bYiZt45KX9KOqV6ndvAMT445MiIWY5E4VQatixWSY7OEKyjhoA5rBx4CgjZ681XX
sg6OgdNRWSCg+WAZG8N2iPXI08NCT8/R3zJC2WPIHlJeSYXAY/GJb9S/0kE3KocA
bF/4VxxNz5VYj5HEfQkuKw==
`protect END_PROTECTED
