`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gMqT/kJZtcWcaIYjHAi/jO08iXgocD3hGCgHP0ucYWiz34TaVXRCRWK/3M+ok2TD
lAuePLqu5REP8ZYdOCi7rGiKB5KTBG389EhJp0l2pcq6ne0T5z/3iQgMKXSilP+m
ua8b1PGHV64VZwD2Gist+eeAbzZ9kWUXMchdt8jTsEiBXJinW491nO0ZpQJ/hSiQ
dmrzumc+u1jFP+AmA6AZVpntxKyEzVQW3eYfWRTCJekSJu1+LpyV69sn7bj5NpvY
LEnBvrvsTYVK7vto2Jb7v1wyd0PyhCiTT23+aKjuQwauXspL1q75qPsivM1YJRDC
BVsqqw/WaJsvQJWAGJLTft7bMlNFEW8MEi51Cf+3pvEKllfNygq/shZ9TJtoILFh
Md89hNtKdnEEyupVo0+y7R1XylPxwn4rfXGmNOn4iHpHKtXQqqGE1LcWp9DA7mvY
bWEN4QD8Jh7uIEuzjc32zQ==
`protect END_PROTECTED
