`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wJLw9ycD9nA+0w5qPqfCTMkRDt/Yjmp4pfnfykQDNkTW+wa4Zj05AGFxCCeDLDjc
0YgnEIwNgBNqsKHuuWnCAfdpdH2mkQywIJcVKeaV6wDi1u4pBuocbZ+1xWYUwqoY
SUu/z1HKwFMCB3uH9giIj5ZsKLo58u2nAiZ4sZnn1VJk4hZ+ZQOjwSOZe4rzabZo
To8GbCc8xE293UDuGpp4guIXzzxju2VYZXi6qbZDMBGDgwnD+oUwkQ5eIXJ2olGy
Mq1om7o7TCQR8xbrsLWMIw==
`protect END_PROTECTED
