`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/4NohpfgRrwbWKW0THQpsZqPgiWh5Z8IgLhcAAGZv5eLYp9hmCcLsHqrDc3Pqtd+
b7SJ8i1UfUBDxPn63KCTfDKNDrKCc89T46ed/b2PQP1C/FbVitD8+SPFumffAK6s
cflnJBPSmk+37qM9H0y5ZzkwpnJtDgoTEZ6FCR6RpLYHqIRo89LGdmcCG6tBaXgl
uI17CkJoc3XZHotctky2BVdaKz+yWHthr8avIlFHoa4dXGE2qrRHC/mdBwVvL/vV
1qcVccgk0RZhW9Vp7DFscKZU+6PPN2WQPih0Oxji3PvQ2whDomwL8lTQUnz2RFRl
6XKqEmNrizM0QbU1WN3Ufnxd9rOge4JNTjTtt0kQhaacu3bqjHrgS1QOslyR7DDx
2dwPdfyl3Wb9rbjjWEFSkbYQGX+x36L9K+qeDgxHji79TnUGx1W59hCGypDNSDf+
ffWnWH4Py6hoYU4icPK6/luNVFfazVFvzjgSlAI3wkVpW9nP6naCe6QLvIOcD7L6
JNGz4Gfm2bthI8RlSQ3gIcg4Vc/T5AbS7PNKyh3oC7ykZrFW8e2iAuk9IQmUwkZA
`protect END_PROTECTED
