`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xXnXvTx+p4iwehIjQJO2PT213s82w2ugR9M+W+oudj1EIFfrJzWgEA4jp7C6mqQi
yG4NdNhCJy3JJ/npB8C9zUiDfms2ufsjSl8U13b7rCvoAtg1fy5cdoDRbhK3hwR5
NUYLcf4UKSvB0z5rKEKJIDvXuHuOdUrfWQD4qX22Zf5pzMKXkB5RVYHF0OPI3iEN
0/GjmtzDHX8HhzOfUPHt8Ui2ZVBgQyEQzrIOwY2kOIseHnmFxf2sDDno8L9Qq4x0
BOC3TyWI7rlgNr7a36UX1ZBWhDJSFaNSkQu80DRTvLY8TJOAYbzPFLLSJC9so6u8
Wreu+GPE5CJhfB7ty3M6v/wC4DCpYxb/PyEdBrxY0C1B8owqxTF6uXuEJo9MGxNQ
R0b+sNS8pCj0l3OZXGrel3vmIZjWlA8GuIru8pi50x/kD2f6BzZdTBc9GTtNBfjT
7AW+06R3U96wxoj/6+QFAMYX6gc2HU6rypQ2FTPmTLXuu94QRUnogrieoxjos9Zv
Jej82y35NsisIWGSD8n1ocLQ7ozls4qFtEkcnHNeIbRUIBEQ4cwro05RfquJPLQm
3PKdQOfmqxXjtUHp4aoMLyY1rmuwsdrZ4wZKGo70PgGu+GYLOpgKTmmd+h/CvOpK
ENcdT+5bdEaVdIeqEogz01qqWehyxdQyA/pioGnVuzpi/IZYJkon8yafv6jorhm5
i5ADcN7D3hjikzNcGbkwW2bv7ULYznpxMxtqyzIw6Nda0D9seja2ZvROKZ7jIA5+
bw+DOZidHjhVQyL8rArg1ygDgxmciYxSsLTjvV7i2BujHXjdrVqP0c+Gn1A9fnbw
VDjWPvhBepD7XoG0cHad5QYORa9xt4SYvtGBgbI2rOZQH3axb+2hpqDE+fJ7RZUV
9k4CGDXxg2764XzUM0MibA+iksfmtDHD+xuFy2vGzQ4=
`protect END_PROTECTED
