`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
irprDuiOyF4tKvSp/iop8kKcK0alAux5MYAq48pxStyvDRsG/UIPMXBek9qjFaAm
mOrJOoFqo/g99QWpwRXlEwvCWRrfT/Gaj2wmakWjErJdS0GdJIapAhg1cuj+j4Du
wCZbqjEhbazq69xrxDlxjp0M93BCzHGg8bW5qJToYJIYfMr/PNA1oZJEUv7PPtTj
PNG4PiEJjo/0sjJ1r5mnloYc0tJVq9vJfC5i+Lwm0qhWgEEF0wTXDSXFREw3D7NL
dzRZYEwGaXwATAGSg6gdS9+XCL1sKGvlOSWP15A5gwT+ynEP08T10ar4E2WbMLLJ
WNxTQbAfIMijUGSo3upYck92AJJ+8d6XqOvuNOM7dwTZzwfiwCI7T5Jz1MPn9zyE
cNZOrIPiwKqQ+XaLqGKRHtRoytrwaPp20kUeoj1PvJEZuoIIuQM/AJ5JsGCj7HSk
uWg8jolUy+RU9Nx9SD9aIR70CAipdfEHjuuus0spQ7ROwSDm4qfAdl8pxE3+pil5
eO633ClIZ+GmeHHq+QwsY98fpT8XqhT3UbnVrKxD6aKb7Aypq9rz8y+Wf50fHXCf
BSXcm7gvFHFZIFA/QUnwAQEZ2vtsyYkGOz1Io/8+yS4kaYxHiCh0ZcQ5X8btiEe3
2e/dLGdVaGs1ntwncVw9exZKCvT3Upr8MxrsvgfbqQgrwcDdegDEBZlbGJ4LkKlj
lPHCes393CbpC11lUmbYQYpZFY+YfFqTRYbym5GuhHWxFDQ68NZp+gKwvMRCvX+s
cPz/8cqaT9OfLQf0r5+myZaz7dd1Vb1Kew+Z7tY9V34xBSQUAMo4cbniMl4QdOyF
RXpBKeI48C9iXiWdtsEqt4QjnGvz1J4cPBlC1DNl2e3Pi2UG11iVfmmbtK5J0Loc
`protect END_PROTECTED
