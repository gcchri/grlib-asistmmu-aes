`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qE73ILPE8EYLChIqyOV63mjbr6N/+y7DRIyn6m30M6Xjpe/c2Kxx6FtVh9a6ug32
CPlh0pTtm1Jh3z2UG9rgLflqzxibHBnLBry5PTAlKp7gEytTP6LSut5bc4bj21FN
w7/AgKyBpb7LQYiR2KnBgMEsWcV6tvdX94jttj+RCRbThQupl82GkLJKYQR7ApIO
YCOAqdrOkgr3hlBWRvoyx58YH6otLmjcZeHc2c9VGEsYL2GF+wyb/ttAZtA6feZu
GNMqYI31mwzC9G+vzC93W3do9aia6U93yeB26x/9H7c5v2xJbayHB0j9vm90uFuT
Y3KMilzMgNdvZ5T6uTvQsDeqcgKfCEcOdb+7BNd/QiOCcW/+djn8hRwwvytf4rOg
zdwC8Vu5YWYFwiiSHXyMDA==
`protect END_PROTECTED
