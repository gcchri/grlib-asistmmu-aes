`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jSHDs89E67UNY1tLwqjBWl5YZjRQEeJfqMosKzOW1466uBAxN60Wzzk/icijxXlV
blFn4PfpMr8inRwqgM/qapEohzTKUEtao8k9pco28prH4RMtm8nedEC6T957iy+i
mG5wVAqr4ni1tPTyvs63U1s+1uAW3oBDoPINVKtibHQeALhbe2s/2frlGpXQzSMA
Q4Jr9ZNdo4LtQ9kpd8o6wSSKzGzspChwOb3fA87nJA2JUiddoeukcDgaSvnK4+DR
og3NdbsqrBzAB6fuFPnVCjRw6Uc0cv6eQvpny4ClWG4bnbG4wnxhNug72qvxHPD3
EZVItjRWb4sUSvO3IOJw51rr6Rn6kUaRHX9t25sWKk5x49etclABCuXKYyZIcJQ6
W2wPEG+3BSedkBIRZRr/ALpBfYePNI/gASlIJ9yNTGJqQtKoKH/GfRJJOia8GLXt
u0m34b+mfn1Qpa02YUpTCy12OIpR7T/AlijFI6WHkdc2PnreGkC0amsiyxnMy7yt
mIagdt5WErtOO4rJuzCeJ2ITg+1XsYak8laO/I+s0fobsOVoDjhIRVwqV5mMWY8A
XuI9otD1p2XSAEfobIrMnltSRIgOjpyAMC7Ustq2wjgfEUQZGNnD8jWCnxpeZQix
qlPbG5q73debuEEbrDUCLAbPtZttRXD0+c0859dI02E9uKR+PzJ23qogbehr8oKP
1LE3FrJkl09Nm8kmoN7hqmVUAg8/W8T4xDbDOHBHgELhTEgkm5P/AUTQG0qKUjQI
EmmZNZ9WNWFyr/xqYYpYf14q2oZZB1j1WDLyX6L0U4iqAy/L5HOyfqNKl9bl/NfY
+ni7fl3AYiRkr7JEM/vk65bL7zNTD/MAM23gyHXEbj7ViLr0H0YyznbHEMfvU5+p
FJQP01G4JlbFNkRbKqprHdvl1rExxo9RUHe6k5E1YZf7Vo6NawOGvFRUqlBb0+nz
EH97XY9f6UW75PntyH5EVDg6zR/eWo5e5q1Vf4dwxmIY88xJvFlnLMU4Z9AT8UUK
Tx9hdEci+H7a6vAI88ICbT7396Tu/jnOYm3SV4ro2zbbOyPT+23FogfiOnBHqYqK
i61wSTTFVIi6/X4EwtkEuOZu5Qpo3Pkni4iu2Ul6VPoto1eDVyaP+JMHf12I0d2x
PzwAkiMu1mngl/qftR2k2uY1K7LkyQ2K68sjyLH0waE/wlDXF3HXTpMakNlKyxWs
/CqiYaRm3G2wAN1F59aOJeh8vJl8dx9tLiZDoDZ6G+5f+TzO7RsUAB2bgOxJbLSc
mn4taH1BERrhW2BIclPw+TnN0DAWJ1CeimagScaHzX5Z7BduSrj8euq+FULzMaKQ
r6PNp/Ay1nXQ2SzNkogPKtYOUbD//nmbTW3juZSng1ZOogiSe0/22fvAhPL8nJJn
J3uXxbDnnJcTt/ChtGJ32mQ7UWnPPgKnzJxsGt1jHk8dfb1gOjonVwkM3QMyWazg
4Btha+zR93q6cQa8Uejgat9cQGWitsGIJcE4cZOqLcVYy/A6xXgIvIHHdim7ft0M
LRNF9zUsTJr+afWE8I2EoXHFsNrYfivCcHKtSIcdm4VimWtQa/AZsBiYPlCXXgh3
drB4zUzw77wJJVKV2Nhgq1KHCbDzVB01R2nU9R8cvgve/77HyH5EATlHGxUugynF
dVvXDY1ySHY0IQ4pU0aMBwaQm4jNPqAyLGZojRxJ3WC5cpvmjvkqMcMzAV49KXQ4
TVpwK8tUOn7s/sxW/7on7STmxViRW51Z5F3MwWnRiD2FWlOtSgmGzZBzB8gKnHK+
TWgPt3Z8rSgjPz9+TO+A731ZkcFC7dlFRlFjthizevBAxmPv+rNfEO1ODOLwTFDA
/9CSamAbuS9e8FPoBBrkmD7OusV9E63bZOLyyWZ8zOfuy9zGwmPQov1jjgClZoRH
jelfNOQBbQTJh27kaPyLYmurIDbb7Uba4hJWScwPdA6NFDXBbISlZguV4BkrqEuE
OBQ10m2kFgwi7orNF4VM04/pBDQVY0QgER9uFmm3Y9NtoMaS/uht0IaU6S6ya8Wn
tkC9FG5doHkoLB/WSYv85dMdCmZxvhLZj/LxT7FiOlE13iNaTBI3lavyxcV2cBUB
JZG3BNDYGU2kwnmX3dz+BNaDFdQ9Uusa0zUjOU4e6ecFTaxRo5R5xPJTwnxafKy2
bsL1uH9MwfxW02rYHshcLrFgPCsFhrMFASwGr8cUuOxxFzAH1elvGuxTFuSxO/DX
RT5U0BwOeKw5uuU+RdwFnyGeePuTf+TPoeLo4zmMmtkQ+zPGOz2+fj8Qx3Fn4Rsd
vBMxM+ywl2MhLQaiXgHg+N1lcuGoTuGAUP/fbQRopffxVUnsvh3JPkWlWl2k4c6D
61pjxmcOd5xJUuvMsNNE8jW/CRnqYbuVM1wR3qBfML4qNjZFjHPMVJHw3JtgIrcy
xY7ubXxQRYac0x4zLonaiQet3WUrtDl6AWqzsxPWQDo4UmNg7jMhwRlYMpiiJ4mU
yOJZ9Fd338j5yZxjWM3QWRQ9t5nLT7GRt2MRWvz5Mz0RIAkX8E9ReqY6YB8Krzey
TYeebz5B2jggG1Z9GXVzoG6noBNQPuuQN5CUeDQ+pwRi7MfXbXkkPmBv7nFUxTc6
a4bw8qgpIlRgYvvzuzHU3wycYNl4ZPqT1gKN3N7kK1H7F9QAURWyRvvtF8v5VPJq
ajChjFX9+sDWdG69MVwKHKM6ho/uLeHQNhKZRDGxh5BjDLtr/wOl6qvcGWIjG+HF
xNU1uWvWqvHyExyBfAmTJx1RzNSXIyDigDQ9dQLSvKquCU2afUoOTMtS7iRJ0xN8
ae+zQUGYdW/lgzWb7bzWfpP1NTgZshQFeUjJO+CnFLqUqRKfCqUx2+eZEYAw6ipJ
vKwMm3+/tqvrGs8ChIj/PTl5cpm7xVa5vAq94KD6LRfUtX14KXQx0Q9wq4sfFz0T
tD43dmhbARJ/FFPDz9SFI/3/9iDjdg3sv9SkALG3DyuKPZ6zgr0lTlzN/Axtv7rZ
eOH8TExSKWJpXNO0mKVVpf4QWklfaucR+l1GSjX85Pv/HyzKiMCNf20+o0trp4Mw
PiRgjWjrKrzpv8ZzSLmVLnEiVueghMajFOE8WlWZLtEyRURPD7Uc+1vJ19Qw1DTa
lnF8pcWFEnr/xXsz0kNuR0DBWJs5KYglCZgUjJcjkery5ZaUEqF+Ny7HtXPvFHgV
lqlWzy3kL6hi1xppd6yuhRXXUykKLx1DTpQS/qqPANyPhQTlxNlPvGX4W6urz34c
lMBPwvhUW+4QwBynMoC0XX6mv3tOf/gp1RcHdwrFyA8QjJFp9MhQ0R5UYG1RfRRy
XtdzGhnU5HS3n42mnCWthP7O02zaIOlMNnmoA8n38O4n0Lz5RGbUYI4TE8x1rjCS
YRnZXJ67ZFdM79wU+NLNhgg5SCmnGIb0++dwL3u+iORwBt1N1N7lIx7xfhtQFF0s
UQGCi3Pz1YEYcxlSFg33aqVNqoDpQ9fS8UZOUGGCCVX440VPfZGR6+lEcPiixjHb
gzzNJRwIkSkIj1j5laC7b0Q+mkoHFakyGuxK+flG5Uhjeewqtfpa6NozayBvxnfT
hpjOmQpDHfveVBTpRu8s9PNlEoIWeLOR2BwrxJRZzu1d40UpurkqtUjVSML+OJJM
skVkBKSfb1S2OcQb20F7XtM2bBNPK7u0k7c6BeOHyTacHt5sjtI9Nl9VpvuR9NV7
WycCH1HAST6jl+TYCtEVKOAVETluuLXT7kbPbve69Ymb+vScLUFXjiADs4GNk1Um
LzbTBcbCXPtRoatHcCWPD00PI6fO2YM2h+S1y5hfVRfb3PtK7gntVtiWV8IFdkm6
6/1UyiUUbNdxgvli/WTbr/pS9Ft0ixGdQm9Phicp7A/SD9zgwMMXSCvTZzricS6p
YTkheOcvBbnjlzchSuA6YkefMdWbdc4QxT7i6H5MXXxSBg9lD4FpBCStqjUTDYAr
tWsPOHd908mmU15DD7icxZFRqIKadPgRf2Ghga6pcZ8X1hrSDVeD8BW75FjofV5h
byIfCrRA4f+cZ/80VxCtH2BpwLaSgC3Baj7pqjakWHYRd/WbnUKVslbSCW0b8kTA
Hs/TcmjaSFb+812QWZuP0zGddCIz4q020SY4bZ6+++CtrP3dXTiw746G3jy8cBCA
ujKh3053ApEj/59T8ycwVOBrMtjfTZrN+nRvfv+q299DX3FIy8mqIVMZv4cMVcYH
NqpW93OcJ/Low180/+szu5zG1c8ISsOHY2Hh8Nu8WvGASzjlacKmNcVjFDqKQ5Dc
LmUTqaYd7XpDOw//bwsMqNpg6xFG8BdUVfjVy85oLH0eQT2rxI1nmPSfSxT7W6Dx
+6sMkwKSTuP+zI6SUSZM6Twn/3YOabwjGvmC2EZ+4q7Rw84E0CCy4cPj8jo50wvX
9V4AY5j4aIaJjnoZulwCScnV8t4b1DphL16JItMDW/GHiipB6N1PPYrTVry1i9ug
qpC+uOnkuhjr0eRObY9FTj+qHg/E88ecv85mwvgauqBZ5rrcBBMb/GmFQHKYuwXV
mT188l8VwTGe5z0EbnkaaubHLVO9KJBSZdBr6gj1RrAlAKHDB8aDHRuqg4vPF/Be
fe9jheTPo8ad1KmPEBhfjVEvajM02Utw4JwsZYor22sIBYJrCrriQFxkrj9Pe35+
IXADPgx+a1yEC6H00OQPNKTab+AD7NpVoRYYVv2ntVUSrIFctonzmA51UFUXXp8L
hKDKAuyncW6Mkc5aliCif55Fmmwe83PXZqmVATw8OBZfOTEdCY/6pZhDhc+dLNyU
MxdApYcZ+K/ZwkuveJT7iV06YGDCbqC+b6QKVHTUDqPkds4IxfVxgKq9yl1pbH1v
IVFxsFaM/Mnwm5Opwpsgoa8lzH60ZIMkZkluz8Mt7LB/LxctVc4jwY+Qeg+oIzgR
EKoDxmvMHqHX8UcrZkYKG1iPO8OF4pGuIgJzzZK8ENveC0EyXC0wjNxVg7svIvWc
g3lPXJd2Sos/hLpD7xOKnc/MP/U9bLQ04AumnD2cvFmW91u1UydUvlyTj3y7a8k2
/u7sJrcVlSP2WMIuLkeaC3iy2xCngJ2rpG1/oDiDgs83Y5FUWA5tVn4JcE1mqOxM
uFGJo01/oQoaPDvuNKXz96X8sCSXiygm1K425ZiuMerkZAKHZy/GPcAXQcYIFK1g
KOUXxcOwhJ7U/wMd7CqcY4X/CmCCFv2hqkVkxicgWpNyVPN6TdpTNDjsec/MFPpU
rWg4wMikAZYEPWeLMSlIiOMnz6T9pyVbuuZThBxzYpbk0pUuxdRrn88zl8i4jPzJ
Zmk1JGnUjlVd1VBQtmk2aAW76+mUJGNU4WcIDqubtYKq81vZn4d0fBFBcnFz74SA
uibTpbW5hZDs6c+oRQr4A3Tsb20Vt1YRE8ebk9pmMq/NsFSD6lmNc1WF32GTEOEY
f3U6aetSUEOqv6p5+uWrviiMSTpwYj3yXPP7P9ckU6lKa2UX1p3Yr4fjvj4DWyKJ
bc8/qC5O33i3yMOPhyGJjuEfIndJ78dmMJNpUYUrW067MEykrbY+5+JL5qAvZ35W
/fYbXtzErxzFhLlLF19TfjTsl38w7bqUqEC01/j7iik/f4rxTt6Esh/1Ydf4n8ms
aEiHxqGJLA4cJYbRgGTijAeCZ9T+2O05V8WYkOXBnZcn7K9m+QmJlObvk6EPIAfD
OVH0CCr2OUiMGle1fIayUwi/IZTxaUCgSIt95sRL9yiLq1rTCYHbJhgUMJ8Q6iWx
yKPfhE5GSk8axD9ndC1Y6+Vb7WYTFnZKY5CKHnuKmj2YTCjauWYWOREcBXio0xiI
K4afQvgSFBsOBsDnx15U1HOmAye4dl6GU/v47C9AbRnUkVherb4gGXXaBjsq10tU
aJyJcQ2jWiw0pVGMXCk7q61or3GMHpy9EfeFCpf7RWCtttFqWJMQwVuXoeLR9EkG
t4BaYkbc8bRrdeBjYKijSoWu6N0tNKVfEuClRojp6SwgkouraHA/j3jWD+juKQkG
m23zS+rdGD81vRhIIvB835kmFkDZnM8b9fqU1vQLJ92QBqEOeCCjW3GLDZF1yhNX
xK5F6++wImq42fhtctPkBDLpfHxk/PFEgxbVZyvaetiyDdS5nLDgmfjanhUCyddw
CGrIqhMoZPnjv+a1xVnY/WEsMwLdOMDyCgywXNBS8dm4hrTYK/bCpIdJidrdsDDs
PcFH8kViP6YvwZ+EbyC1+3acOyDl8qluxmxmtACKVZ/jzwSX2qxqEedYjH3idU63
NQfWqPhuMNpEhF5zK768YNcR8zKJClqPv5RZW50gQsf/OXUrjEsq3672DoCoJGDJ
+PytLexEU0+ujXulveLfD5SMHkYw3zSf1ri0q3f3VAtcuwf+cLKzYi8UiWZCCJKi
n6Drjg1fCqDtyjsQnXRhJaK1X09v3yQcR+Vj9/kMqCJ6fCufGKXyinilStN0AcyQ
wVdNGqgfyxw/034qVhyKNPAMsFw/0U1qKVKTzMpE8EecjMMQk8DER7GOQMN8ROvC
Tw/SDwSfZfjlKTU6ex31pFW7t8vQM2IGKoTj0eX4iIH7lsXZLj5RYQJB3N54esJJ
tDmzd+r9eZaPALiCMrO+Hv4QK/WIknwKcC1rP06fsQtOVjZDNRcNDlm3hm2AtO+w
bom/V1X9GgevEUtd/LXMi9bWP0xo1+2SXnGd3NY/B6+yY9c89xc+9rOvtr6Rvbp6
69R5SaDxCXX6Ia8s/GZavzl11dG5fpwDvZj8+/e7EmddKpTswWfe01ApmXi8aETT
Px41Ls+bD8EKc8tWy72/3+dcbcrRDkxVJuuDjekI4EmqLPo1tLhXdHxFd+rY7qmJ
I1O69Wp+RM3L8Ok/acoFw0ytt7dPGRoMzewvMpun1XFys0U1J+PSiGFDGqU2b8n3
WrxO6J9blppa6egf1/ym024Ea+T6+VgqL6kB0GWbG0+5k6K+j9fv1tiCSUe0EF1w
9lmxr3RY+co7yPeGVdwKyB656elKV+LCInFFeOcKRTgqTbyT4SXqf3MABbwFUYFu
JydP1Y3jV0iUtxi3ejpCUJ1dgwKRwVzG/xf8gVDaQDuUDy4DfS93IgpCtRKnGe+T
ZNR5OmntVggJo8LcFTDm9kjHVLPWNny2iazCuXTV2ijZQko41YMevPdfi+EvX7ip
U/rdF7vLxa9N0iR5AbpWiBBGbAU0BU90Vebqwcg+cpTc3Yzbgn3s3W+G53apaNOS
SJL6Ny4oMeivIN/K/sxIEYiBGXdz48mTy5YssaQogKXWllp90ip/ylteALFksjX4
ukPmmxyeFIzevjkiTmhoLAGDnVhwWqIOIUOYLS+Jqb5f4pD466DLHK4KgGcHYfCA
TfQYpb4lNoWXIgcxzd4gH//LVj8DtLGe0kx80ANlYkc0/Q2jFkU6FHbdHYaZ0tHD
CjPWWgJWfhIzrOhhYNPa1FopZ2EspP6R29YQzFrsthYZlbh07Dd7O2OWxWCMs2tP
fNudtZOmbw2ieEgCB4KY2ma5uCKg+rZwx1CpwCeV3hF7DL9Tj2W4kSy69d9gDkeT
vqgzyBibpuJ27c4g1l2hKWT4HF2m4SzxGq1/ANhmpsqV5DeRMURURyY+yDzi8BGP
SDtRDC6S74YyGnhNBXST1O0/WZWTQku9Se2ANTkEVuOh9cU6OcA9fzCmHoip3Kg7
rquVs6xo9B9uIQL6VnUm4XxcLTDticjj04M9EuO+N1731eeNY/1rdM7ap3aIM9PE
3OVHxMVmTQjov0J3aLIoHpZhwR7UQwzeRs50Kkpn5wfce+JSvF78YDD1YKFtCXrc
NjmXsONbNp3OkeSCt3V+IPQIG6jYlQUnJ/ygY4y2uI4B78rY2Ikv0OYfE01qtjDT
UpWYrpL1RXoYyyUdSZXr+bxDm4S66pWKUoJbtDUHycfz6Dlq17mWK+Iey87qcWOW
v6O4wHKAVbK45vA1iqPFxhOTnAHs8JIKczsi6n7qiX3d6WRuc3T6pQWINiGnTDjS
DMEY4ZdDL81jVyFlH2stqwmjod7HWRKVwwTbGEs84s4sqNVVwPGS2CCqOiN80qUa
+TrO+4Ve6W3mPaneqjtMhLfWwuy8OFtl/80e79h8z7DgJ4UHyFblp+mHg/FG3Woo
C/nRM0Z9RAUumyADSiBTImrEeN2wLLanDdxYwbh929jVJL2pZFLFnIZhM/K+o0Fm
ei4ZYJWAAicNnIBlS3mcDg5cGVJUIHxosbbCLVrEToYA37dc9w2kRpDNPll7eitS
e/EGcAYrvukEMhgDES0xXhqplatWyVbXGIHSk51cY/THvkpeNkMlzupeLwCEsbh2
BMDmVITwFObIZ8O27nHAYNOdHvxdK9li6ugEViIlkkXnRejTgWbPO6GI1/bAfiWF
V0bk8N5ghJmNeAA9JG+pf2IhdmUMZNjj4knnit2mb4/ZJLFGaQ8s2ma99zovzd10
KP/JRPGJb9v3NXQ83m9YRBfVKsQg4wLRs9zjwq/NaXmXlvKUCK9HJFWQq9m6HP7/
+zgXd9wBRI4PRbFXBIrrS/F5xHx9V0dcQhcucMbf8BFqt+SoDev/6owwjjCFpcir
mkcljzDZMbbjw8lbvtbPYZE23JMlz2szsfnrHBN7V1hkmadj+pKWsPesG0IjwpTa
WzK0OwLA7q6SUw0R8kAUtFEOaPXQX9OFjqEDpFyRRpECQYwrIJURrkG1146DMiuE
2oP1aWSU8Kcj6/3qLIzVIS7Ni7PF4lYA6qd0fFgrFgW5GTwfINio+/ZbHASGHOt3
Zm9taq/kFi2Sx+bDbYIvH2dhbjcz9QEUccspdW/y5DYJwQu55yAvtLATrrCk9U/l
CyrPSJYDlB6MUtBfffzYEjel+b0Ywg118vEZE1p6Tfuwunkzo9tSiwQezsRYdIFs
qBegFUFzMiamLBUoqhWTcnQmT9mA9OByiHBhQ6ZAvdhan7T7B+3ECEVkoGStPnG5
LZ4vztKNW+cJyEp7Z8EIDpwKBBTvSlEYSbHj3G2FOswme2pOJqfjXV9d1ARC3Bzx
pQ2INy7WtzutpjbYCmmFCa8MlE2HZJ1NEwsvKB3E9vYHB+SPUqgj23rUDNhLwyJq
OTk4jWcoyMF4DYoxQfZynYu1ytGFs78apPVZMU6gky22gmY+Vd4f6wujW4qGBvDE
HHt8E4PPTLVvaDFrpbd//b3vCs8kYQU6PoF3vfW78/NP78WvZ7spQfY+vXDKy4Zc
zjJxrfHYy+/Re/eXh7s9Tuk5pVdqsc1d+mTisp7VBACq3Lgvj5OjekDK5WNqf0t0
dNwS2JyqK7isA06MOjOG9MvvEiRSB4FtbZsTnDYcl7c3v+UwPdP7578IcBHwq72p
aVRNRcXD7wfatGF1/ybF39M6hDIec+KHbURvsKjKDK7+7rYJfmEauN47cqoCALg5
sOS9AJRkSvSzgXFlTRe/nWApO2tuFvBMZmcurcvQigDpMdNRBhyx17peVDApY65o
F1EQJWliRaNka6ZIzZMsnlozHNm423jFHTKEmQsAc0lEAlnqxBJG5Dhr2APJ8xtF
mJ9Wz7JsVslD45/XRsrwCfBrCDUR8fVCO+WsVUzii91dQG3ucnAjYJcQwiIKFkfR
FTKoy8IsP9Z1lGdQUycg7jjlvyNwAbzqU3cv8GU8p6fwmTTCKCBmECLNj9vN7kvh
kLYWwMnDlWet+bmkKh+thMUEw+V+HdGSUdgg06cl5FDT+EKPG4Wt/wJ1WHuPhiCH
QFCJCQrUnVKzhw/4iHW8KueroIXncvGAz5EZfEoC5gLSXT3Iv5NDlsLKjuDs/Ahg
gLi3Yz0hi3ucW0Y342MBNW3bhwsqilv50SxbU8eVoJexNN2b8SzKbozJbX805NEO
B4q8btrCOTEERblloGtrbhZWgrGIWIBV18uYd0VW+1OkWPhRwJEBNbf09kPmMgU/
9QyDRnyJ3fCfnvRN2xd5FipPzgN5+llc3isERoxnyCSAVfwBqffdwXvYjwQlnnWO
Gyiyt6E7qXHcjLtFSxUE1ao6Ok2bASeUQeiuLo8RwXXCh4nehv0LvxVJGNkqKBrS
JuzyEHsLGuonKfBdHoGTnb44OYW3UVNb4VydOMGlBsnvl9DqxLvkNturrxml3BMa
DhLoqo6a5dGAXO3OUtvDG0ucq/vwkiHPSFlluLYdQsCsNfEApN1IrAi+W5c3ZZiH
0RzRwR4+wWoYQtHa0GgTn3RUN35Cz+s2vcKhrJF77rtt4gMNKirtDdvm9FazsiFZ
psZXnWL0bvEoIVP+zhPFsP5eME69WdZ9XsIsj0xQaxBSd8xVXRLaqbdGMjIQAUmZ
rQIkKRdUomElfNR13hQa6o8TSyHwZ/eX1d/ebiQ4EMXrOp1Q8Npru38ZYSFJ2gXU
l2YWfU9RSJnsAjvtU9qx0jG4E2ZcR8+UgP2BbrOAm5L7YjK0eFTqqnb08/G3Ys3V
1nbjwWGMg3+UWJ2hwwUWzfwpcaDdR/bFkOIAspWkltCgCmXxQS2D3id8REkK21QX
p9CY1LMs9t9/KOvuXL3YvP7NZiphnVSVcsAM1Na5HgJWMYs1Govp0bJOPi02nVeL
2SONEFRKYG8mET2kC5QpPqZAUMZBh6NKCLL3SfLdHkXE664k2vjzCi85TBBxO9Qc
BCSGWcH2MBQhawBj8HLW65SIkiGTb5P3RIUftxHsXuMhtkkXZMz5+I2suXW30/b/
oXs1S+bNY+vVjDojjymT4m+oykfydc/y8T6CEN1W4zlFsEYHLViZyAvJ+glhWHa6
/nE0kvc34KWxH6iFhKD4/IDw33tcSku/MykI/Sb2wmqaWjjJKusNUTJSV6u1+lWT
KMcmzmEbignU3tlfM0nPp+SyRFLWDntySG1jM2FGUaPf97EruklA3wbEUfjjopaL
maYiEynfTXWS754pod47Uh+HJtLNmTLkfR97KdXIp7PRb50rNhiBH+Gmmfmukhdf
C4go2GJdnRwSPl99C1htSST93FPClXf2Dp23OAqYxitGcJYxd2jvUGiEhJ8HUPmz
bXprglIcJcs6ayKUEjUU6Qu5NLjhKXWZ/C18nLt6dlBkCeY2x3Jya9Ic0bqZI5xt
JMQDd3yyS3s01PVsSeATl7shVSjiue488Ukq1qLkzxemYe/HplxyizdE5Ck8UqKi
QwzpDe5ADdNN611HhUKA7k2Spa1y+WGgL/7hLUdHYKZyPT6Yh+UkEc6s7tIU+pTE
dbd0l3ij90n3Bgnsm9gdtdwmNM1C+vWDJoDi0KuG4jBs67XIVYuVHIu9Fm4rQiXv
Emux63rB/tKZG7dzpJLU5UYpgXwR1rehS8fhxHhHrVn6azo/uAzdhmlsW99W3Pgu
KEUVUdUNeGrXUjWLgOYyt/7YRFbiXLzq1G7VDr4ePtAYecpDRHhyOvgtCJ2XvbsS
KTS4w4i+81cqGWgTfb82tmx9WoRYB26iMKIksA8aK7LE0JO5mxnynJyggQ87CY0W
No1NI7C7nR15l4djsuTG36fmtKLqHY4CXX56DNv5stmEE7+uH0GL2PocBjMCjNBe
njGN2MY36b23EtfVS/rzW67ifB3y2VVFyJrgx3AwYBKFpWzI+fXJliiOQPtA5jED
NmersMr9v9/RHOEf5L/uIJmfuem1/Gwz30yXiPqvtIrZav8nnm/IoLvHVxndNGT1
hhj2VL+9owQv9yqUI5K9kAakSpfbHnzPAAy06J4riFCXmjn3bQDWlYxoYoibC9U5
HnN5Kg6UpPWfs4qj0rTi9uxxYMutDpPJJo0hPNk9Sk1Brft4BsYJy5tnekomREdL
JJ2R2nAJlcNFXikIPjuiyLtsfkEa+LqZ4lsQPUVBA6Lu/HOrnap5kv7dCTXgDGCb
/vZlwhi9NzLn308pcLxuhfFHqqck0v3auV1T/33jy/W0Tb2TuwwrXRXtI3FM1a2a
2DAmWET6d8m7wbLfad9U1emQUvH0TR/IexkwwyzFkLNVYKuaMQMeoFEMTShI4J4D
XARuM1vXjWF/uTgvBc7mcYKe/2VBk5+gWw0idpjIbg7gQ0/NZx4aoLSS4tf9vepL
SUWSSs4IGyl7EHfXcG53Ew46w4gxl7dK6OZjOiCyvV+LpgGXdh/cyllDAlR6tfgl
QJyzk5F9Y3mIuzoOrFoonkH68XLd0es5rZFuybVWoLpTWdYk8/YVb/WtNAzL4tEo
14ekIdtJxwN7jSxFytBLwbPnhs3dZXbwpwhm/So2sEe2qYyZgzBAHmtXZ+Re02Kj
Ddbys37fbE6vluwkYPqVgHzok38ncYmHKwEP+Sgt5ltYkhteheg34PKgk8p3bcsL
O6RzMt9ouiRCfgP+FnvIJwdR5BzXq4kNEMBSgr+xtFYPT4M+5Brq5R44bOxp8dKY
PfWOpSO8H7yAAjb0eML0PzKLPe1Zcz+eB+0mIF4LV7TXIWewBQ6/uxFbYp7REo2W
XNd5bItYHSGFvecgUsaf7oO/HZDrfM8Y4Uzy+BGmiOpPya2CPxT7LyTsUVNczi+L
PLo4F2vwoQva0/zuIuV2QqCFU5ss7o6qgozdKp1t8jmg3HkjsmSL6fL1IDtn89+H
vPVOIOpdPvjnPDK70iSC1kswKyZqBZNwpjCgDWDl7k6YIr36Dyb4q2KLVnHnKjT7
NlW97m1qW9rbY66EKTJFSkMk5u9PO4f84N3e21/EXCokaIM5OYY63KOJtZVohXh6
A9bA7dvciyRiA4tQ0UiwN9qArREcZqjrFL6U7yrQZ/yJxsQaxCbCQqlBDRSZ+FeE
fQ5Aa6QwJ6TYyAIM0kFrPtlEWlZc6LCX5pa2Nk8id0PHAThHwcP84MGt2KT9a2QE
qdXgjwLLXHYL1+L9QXyRugbkzz7dIE3HZDHfBX2x2LLv+4dscJWZPKq71JFN2Q2x
6RL3ZP5T3rhhHbNkEYGeaOASk4rbS9NxJngYaUde90V94OZDmcwCM0eFYi4D9Xla
lxiD085ikl2GoMqdN53TpfALITDvevtZGOMb3hE4cS7hQsnch6A+1lQOSXHrx8YI
1QSbw6aOrgg3Q/vfmqtFvrDLupInrsELjNALAZCnTNJZct1lOAzxFI6K6JOPEueV
SDUkRV25C3k/cjT3O87mDKz1dodZo+cmUM1qrRTLdSevCIArUtGhmBZAKxVt1H07
QIS5B7beAc/vCNEQrn7NYZQ3M3JUdIDy8nX5q5ACKYVU/SuRrN6ONtsCKdo4izJN
QojbKyC/wfzxdnsN8M5osacN46mJU0oeFpvWov0Ja50ILu7Sq0nKIg4wNYjMX2wI
avWwUHV2gy4ZhMkz2t50IyKRQrzdo3onLM39hQdezsm1V2trY7LWgOoI02XzVN1w
jDCqLLmDblcr5lzQS+ULmuYSHHLYY9XjYNuCEa19sLIntH9xTFurNxqwkXN2g2bv
nu727nQ+U9Mq9inE6Ql/UehehyuhBScYOc3RjFRHBW5Yamd33uWQ1wq31wF7ZYN0
qMtffD4hgqa8fKOdB8x4ieUu4ZfAiIxEGUmcIlYRjfhoZqJBmAcEgXg926YYqeOl
A8ILbGCsNHsa6jiekLcwDR4b+Ao22WJfDA/DIIPzvSpllTwABPaZlIHpdustKYou
D9OtAG/kOYqVI6LcY7omLgV3CJ5CmCtx796EeQofBWi1eCt+VIY90UDABqUnS+06
2q1D3Sp0Q+47LGhU+bLSNcodBYRM6kueOqKi7dhtTqt0tepQpOvBqpfueZw2tJsq
j044DRHgvRKcP0mGvmYBCK+896QqDIJMCv9StG7yLrglYFdzoq2fYP1flGYZbIZp
Ny5ZIZtxO1kFDlOAouqjqXNFCsY0v61myG9NKt7KtdSGM2SRGBR9Ko+5/oVYdQCS
P3AoNj598Qp+MZEok2XoyOmp39Ixvx5CgeQ7L+AdenaASLOYM9KerHFprlmYz2gs
hzXyoReYKc5Kztr9h8Uh8FFekjgnRVF9UchXzH9YpGiTORgNDPjAT1cuZUIHKGV9
hK0PAyeaxiHv2H3N4Kbscaub6fOQ/oJUgbygWi+kLF+oM3o+xA7JsjeLMnuHWbTu
KyWFSFF00QK1cLpGbSUoWQetpsElp8YknyAMmfZeMq11Xa6SfgJPauTqBoyAY97t
SHyDyi6xJQ1SpSYP7+1teJtBpH3SQCwVHLZcH2LD3TUBi2u+01paed+g/thAWdu2
9ZELghTUfxtm6SeeYfSFyk0q06gJxg6S7OIW6RrTdIzkjYZdGhpMuEqlz37PKCpc
f3Q73TRuL2obi5RiiQ4L3FHOTxaaE+8nSWUQVool0Tv5FUfFcHnOFsfhIzwFz6YG
QTPiOF1XEj0tOybS2ZP4RtHZwKCIqwuxgnN0BbqgsV/S2XJ1+WBpNxaB1EPetDOX
AkYpXAIW22EWIlV54suRdEG8Z/CYzoiIWf/JPcetK+MQSGm7aWK1czhVkBIPUdhb
0v50pLYstk0uofJ5KScSoeAjdYeSOfAc+9j69m6JSMBTXd7Rm+Cy0joPq+B6chkm
MLm3gVxm/EsBfRT9XZW5gQlxvnT+mf2D/DeOnZX49BfHFbCNrrWmS7bsx6fcYSgo
uZdiGBxcOtQQesyB8nWs8rvUeP473YF0ED5D1GSSLpc9Y/Vq0OgCBI/Rs61kOjgr
6e/3nDzrvLZEUw5Apk/snmdcbOVZi6jVzE8b8UecHKYmCOXpmangZ0nJH+reMTwe
uiwTJ/bCkwbxRIns9Kz7zZSycgTIUOWFFyHx8PQe+6aaRGZE/brmeHKFHwDlDefd
GCXbLoFjsfsHmLK6q0PJZ9SKQ662rn2sRfnklQixdf8zQkEpzPQtzQxJ/YfHoh5X
cxyLt3ixaLvT9kj20JJUmx4qh2W7z/g3CyR52a3s3ETjn44WZ84kO9YdCA8tATSb
QtPqYkQF+aujVWkELHSj591sOQ+28jfgpBdUOWKHRporq8ALRgLuT3Mw0WMdPNE4
RUEq8xLzSEY5anK6McCWwA38Pj2LWLFetG2furh05kofsw3Nuchbdh7Dhw90BmPi
LqDbWp4KKK4i6K+bscVp6OrLWoR1porC/0xEdM3FcCDCz9Ye0c3U8Yn/7/DYRQLf
sy3tzo9IXMbhop3E7sq5xmeRj6ExkvElfnOLg/peLcT3xYADGhRqm6q+iXGVFmGZ
lrQ+zSHzP5gDGBrhAGSw3KKY/Zb+vAlo/7nDIUJ9083obLzGZei6NDlhTrqxG76b
+4BjUVYRWq1sqjRTrvyK7vl3gTbgvou7PjJLj6lf7aog2Ot2Zeb6/VdcBU7cP/RC
WxLNUowOwY1BCFlIhCOoK6q2TQXI2PG8DcsKffCjyHvv17eBBBosPfaxEiHPo5Vd
HDhbvFoSSR9M7VZDrfeFtOuGE2Kwov03Woh2SrfPD0MbIwXGSqeuekCqTbTwAgNs
SINP8JzuxZiX7A/44y1W0JL07ohN8pqMjJb/BaEGi0ZJ/iGL0Ll/EdQOJG9xol/5
j6mhLf7S8BXXzsWldA6rBZKzk4857s8DwJIIN5jD5qLwYpSG+V18EytYUbZlW0QA
CvUimw6btSQs1Pora9XlAY3wGKIV4ssW/0VTusLoP3qVCOBBoYuHfZb8vKq4Vfim
I5PG1SaV1MMVCRcI5+nIgORlYhm4wf7p5AeAWHxNzVsxkkXqAGMYHFsiFa/b6TYr
pLg+4prFmZGIAFH3QVaCkVcUbTCrQ1UanoLe9O1UPoGEAozhpJzIlHKmGsA/NyNj
WdBhgEyEJk1T6u25OGn6wW4mhpalx4+Jqq6AkLPhyRAu9reIbM1fOsNmF1yk5n0r
tibJ7TAkjF+R8hvJnfmKEdfoEMrGQ5FUOEcdo7qcyOIrE//zhEniPlB2yt1vRiqR
NcFC9CoDv/VRj2tQBl2DFYHKNn6fI0so/vnn+yLA2LK1q/O93roTG4Y8u58oqJbm
tgwv2AiZdOI3+ROBSAQEh1UcdNPZGj30zGmMEpeOZ4xklrRtIY9ClBPG7lSIgUS1
Gg+5+m/ewuJu1Q+WWTbe5mJN4UJEs5ksLkXE7zRx6z+UAcvZY0DQD810COfrx/80
PQ3gLjWnFC+/JAH/G07zy3VKTIcAZVhviPuNsjSgWzqIAS1ICRkTh4ZjBOOpakL3
1qyXFqB+TahtgAR4fRQdtlA9BXZhNgcU87uW02+YNAdr3STxowyZT8YHUbfCI2MZ
QH8xtnHiwlHLOG6mkRKxBq8eFFjRIpV1NSfBtscE3ZLPGJRNk7MI5J6NMeLKcE6X
ZE02HsfQepcLlDJUK4PA1Pg0FliCYgL3oa4r2mN8sxabIgZ4ieIIFAOQje44XWcE
NKoC6AnLVj6WBmru6ui8VKcJup4Yra5/3wf2pA16aFlrKXFseG8J47VBepqZuB/P
8O41FylnPPU9gWVtkSofGGCrY3o919NxbrapgUXCJ7XeTtV7OcM9z9D8LQJkRkaZ
p1bYFufKfg1efwALyVYz0HgH5IFJ4z4urwtivI1i6gLNowGDPt+4ONhYM3E0ckpl
1hA0y6p84qx5NlT+8cJwmPIk2Pn5BxF5lcRF0Xew2iuiqXw7LSEvlAtgN4F6TsbF
Dlvm8ucmvJUJ+i0EGtx78TyANbvDdrOZfrQ66kfObtq4e3nJSs6NEVwagyOo8wK/
5KaEWVhEjMtbAxV1d5QNhwnO8TMsXCb/G9MWfe0+Z9RqmCIA/PQq96WSPIzwNVH7
XmQ5LHeVvkB8FbntsJM+00/O3xj2roxlDSFXLo8YJpbFdnpZ+g/pzw+zSlMxV0gg
5GkjP4I3Yngi0uGP71Kj7sKxlV1gnkk4xIn4xFGnySqqI7HdhDAEE3D+jYFWZhWg
0SRctyDzJxmn7Sg3vE/SjnJTHFwAnFmcbsz213WrUIsfqK39cQY5KkqBFnomqwnK
Rvl2oEKeDGjBHrXDbBzv8lWiWDQOoqJhzXwaIeDNwLLgxu3p13WBLxfHDFWWqOYs
RrFiDHx/ABDT4awXl1RAxwa0hdq7jZC/Yntb7mWd6o+OQ747ndzf3L/arQmYNn5e
0q3An4MB8NiQ2hSze9SlnlMxFkfz2kvGVuv4jjIvlXEJgAHVbb9kkUc89Xtw1M07
XrRV6mhRA03sUN8e5BAR4Q+5xR1WHI6l1lR0leTjPz/ZFYFpjTVUCX8KjdtTbhKc
xrRUPtuyHyUVsV/5VLzv+tqsqgcEi289F7zpEMxTLRRgMiZU3+RrXp9Vx0cgkzTF
vBK4RcJUx+ADfAUBJZpC0K421MztR962y7UlPSJvFLRBCEAowZy50iGueVj8dpfP
cKKYFKso5dewHe/XG8u2WiewPs/KGhcHmz4/WKc5Sk6huuC5fK8go04oRUpKdgJG
6x2L29fARwRGpUz2vVaF1OJ/4aDaWiX9yxw5iDsrArn9muxkDOeoadAxS36B6m5b
pEVBx5QheNUnkXHnmCXhKr3AIe2+3MoJ7A5Ncf/6nVzbTeaISFJqNtFsXoqYmyec
pdLywiwMPGE6f8lvzBh51gV3jX4Szl9+lA2TuZ53lJoyvleFmR2jNZzb92WxLfjP
MQBkCp2CoKeOmmMBMEE4G4L7lCCRZmpIlBM1DelzMtwzIt4AoMLkeJHJJMHEEJbf
BlCYPwRvIFoDbDpdSdkFUZn/HK1gI6fzOccJRe7ElysNxCA6FI6R21CxHedkNJQt
l1y/3mx4PAajbvlvCXlxrdPMzVD4fDlSbAEMlrBCTFejJtSWvRFn5qcdTPDzj+0T
chvxfYh+ZYRvVBnb5uvvM/qJQ1tTXhxg/NuQIgHIfHGrB2J549T9H55Mivjn8RLO
ze8U1x+/Dsg9OoUN1igYpS5+GfpWyeWrMJ9R+r4QQZxAHpoDWckwV/18F7g5m5jy
Dmv3rd/zjRIiJcq49s43Ll+3bqQaJBZBB1EDZupcahwz0p7Sdc/yju3zrxCJqC/q
0mN/Xtw0T57wXjCw8HdiZ7W0cfie1+JE7Varzb2IvkA0lxqFOJmnI4288bvqrCpr
DakWUHtFA2JH+E7wIpO8lIoqfVB3ZwfIgpKwRd5wyoFr7dlZ6ei7wU+AwTze3Aw4
mCdR0S9cYJ5fpdbqVEe/XJ7OgZDSJagu1ELj2zItLVpHo+tG1p4sDD/erAvV0cfm
RkEcuCBzBEUZX7IBeRtr9abzr2ICUZ3XvOoxbCFtw346ntSZcSgse52YnCLENxo+
FxU0rCyJa0We4lYQQXi1kiZOiuWpWACDgYL4uphMP+BfnRd/X1xUGaOrLWh7LGKK
c+CBsatLUT2Da0uxfPSP242VyaGiKU9mBzg7bhliFQwrZStLn7EiCa+GLiCywu+o
sDf4iyJ54ql93v9XiceL1HCSdDwN1dLsgJw7zaYw7eZTyIDGt3KXCPJ0vOc2+LYz
2EpvlJLFQMuuOwXEzhYHYKCwP6BN9qw7I17uvi3cU5WK7z1W4x/mZUAWVW8i/x0q
+5pKYIbqn24SLy9FiiuRIB93ZmxcjIVmQZfsSoUFmPL2rZj7iOp4SaRhCLBI78W9
YfPx72P/wR1YLJBC0svj39Z3w32AHCQFe6ytgQ5sGKuh9pzVwJX6UEueswFGkRiG
VbNtzx1fMcix/EfTNTj6GKUAOWQnZzmY0pnCeYIBdodHICRPNwnLjYn2x7wOb0b0
L8vU8A+YmHkb9VAvHkMLFurANpIjndVlS1eBhR0aNWjV1DAkNILyzx5qmMzba4BY
K9NUAOoCgpfeE+PIuopaO0Pj1uw/J/VyCdY2OolCKoRwxWMP0Xr9IlRJtOO+jxcL
8T/GlvbAB6wfWE1ShEfzT+Hp8sz56BTdisbHDPfz4ECLSaD6uMjKE3CIGQTXpJ9+
baR9vGE9Y8gQcINoI8n+zypeutafmjq4AlUXpyKqBuG9uUwF2tv55hnmBZZOLIBo
NcHBknI8+2OQ0tQ7UqEkcH9Afi6QzEc21WvH+OSmOxYyuCkiHIM63+tgnJqBv8fN
DUoh85KU/5bqKExuxR+p7VqqRmgy12r1g9PSWH3aKMbT+DstVkNq0zOx60nvcHNu
ou13NWjoeJtt5hC091c6+M8qfSrsurpK0wKfha2HpgfCJgweFgcXSLjy1xeTsXLZ
gvJLMT2O70TlIOlq6FFDuYvtHdualtN7iuHKVSJ5gnD9uLg8EpbZ7+b5nRhzD0b8
e1FlGP7wFnSX4PFphf+zb0JUcbnUnWq1hoDVcHJTugzIeqX9xOHpN2xjBvbwJptc
jjrtn3deMEDnJ/EN2bE8kOZHHE7y2sh94/6+fVeT2ZGSC85T4EPImzxgM+MugxSe
yR5hyI4MBiwhW1L8Fa2cDtlRHl/06Ms3dYf0UvHC5ofiCDZ0rFxBojwW+vEzktRx
rDh6O+FLd1Qs8aDe/Tm4GSKj0+P8XdfzN826zJH2KDsL0+bxMNlW8LICDr/otBTn
5zaG+cQ8Xfjrq5KZ+5rgjbOl0u7nyA0DMTTY1PJ1l9sISPQxH6R2FjrpQctmhD4a
HheO1jokK8B6LeYXZgcP0WcqOKHHdvVcIqw1WOaoPcFMzv/sMTyIOE9GxBlf9aS+
Wu18gGZ0H38xqc0qtvCUEfCkLZWGw8LvM2UNRcRASqzgmeeWFVV9+9XkTX3zkVB9
vOArYxBXvVxytF4B8TzIgTO+sINRfzR0+HYbRViVDRpmVqmIwp/0QOriCyPxe3l5
4MEX4WKKFQI4O7iMkeomZwTD9tWGiJOzscR0rmH3Y65NAs8XLEoez0km+p0Qly0e
cSKFyNvZgj4iF3omea7Rg03dM+z1LLRWwzvF1vDjwxxj7sLa8Bx8oxu/N+qPU3jG
5yUm9vqE0LLzseRNXhOJPk/1sZH0DeQG7QEMMsk2L1ugr5YbOFIcgM42UpIi5h6l
BwieON/L7Zg59+TSoqfwjfFwOkqtKLhaP1jJsHBqg8Vyww2toXHk7Z+aLb/eObik
yrMlfPH90oZp0tJhd2EZw6ynKPwnAc6ns0JNQ5vVpxr/5SaixteA7rGG8U0ZCUjm
rTn1EyDdE174aX2vaGK/DYyk8j9xjBuwy5dcZIyAMMLOo6J35I2Km8t+68VITr9R
3P4uOfXwMe2CMyZXiTBVCEVT2okbEnEe2Sa4N9Y2MhQohwl4gvfVl9b9/KZBkk1x
6GsIQcdr3GyTJD1zFfFfScPNzfIJK+1Np3pyfiZmx5LuMN8inf9+FMY3hZ99bMO9
kpAbHW1hb7UUSAjbBjSx1cidbp+WNiLqdUaxnffbhWkzQif1z9cmPHStRzcMUKF3
H/arbBrHL8O6hLD9qJ4kzlhuB4izS3g4X7hAwcsxnjDScdKVMq0SKd0TZ9tAKdhy
NnqeVMm6jyGe88GRG7xbL7CuVFWd6zyrwsfDKlWOtjP6+de0Fn53NnSh2difBULs
I0NCQMSicpkLvPplYXFolwDm+aVlBi3zbqWOdM9Se4NOIy+wZq/he77nxlnNmHOQ
Unu5MAoXajzZzwlAO4ekbT91gWFP/a3WioWo6FB/C09Y6tfIPeWi1B2kfESZAmb/
xPyd1dLJF8ydo0QFWG89V9MZscPWlJ57B2R11iHYa1EfJUZK1j1ERZUOTEbVTwaU
T8x061aycKLqcKoPHd8QZt3ZFWsf85fu0ZGGeSjfdcT///dd5WD0NU3CIWCwUqrY
hgzQbX6MJhkA8Nn4G3ULFjAuFXhCFcVyR9TRzEZwDrNZtuQvR7TNdOS37pbyR275
onEzagk4pZZRkSbTdGy7ytB5VZaA60AeXlANM+xuik1jupeqvkTBCvDZpg0yx/2I
zpX1VXzLZN69xwvXkQB8lTQzIObMUEVBxtQHnCz3Na99hpFQWdfIf0PKka+ZGtyf
V/gtif13wBkpckjf6g3Jdh4XfcvWhBxRr08zqRPfgXRSy6JnT3cvqVOmUYCHh6W3
uxMBFKcfQVauyDtjxjLkz9TfrJo6/Gpm3x2cTgfMycfTFT08XNb/JnHifpSmyYBd
grSOGrZdzy3Drh/J7iGPhfiPjVsRF2iFscH+WsdassZLYVRMgLQvd0q2gQWjHVF7
BM+DnsNoCqPVgnimDcPsmjr1mX8Q0IC2tGEPkLQdx1ZisjvoNKukzcE2YtGWy3f6
QTLd4nma2oh9s7TOD3gPk6xewH8HiEHcSoz2sj2slE/ilq48gFYVGottm50A83C6
G46A2Dd4r3vlStphbVFWGmx8EhjTsmBj91f+fsX0bQA4YSQSPkXzos8Wbq2htnFX
MzEYIFt/35iwlV5COUNmPxN+auDH3jlW3jEoKA1bJQA7VL3YAOqQr1ZMeOOHQuZo
d6w40H8rTwvbTooOoewkjduW4z1sqWlrv0JRRWV19v7GAUx9ALlFWpTZeuWYiMIi
/DEzptVfanMe3UpCLJm9CR4QHqxBao910Sa1hsmTu3UmP0VJJ5K9rAJ7ApkdKtVc
iX/HoA7ojhlSjD8Ixw42HlicVZbCBc45jm+peJKNdwbZrzeVGN/k/Lk6SuruNM+w
LrhKQ5yG6X5DhEHesowvvrIpxS8NeettP+qJsW12/CqOfH2UV0smssfgqS2fb3hC
14nNF6SUKvvHVTPphozvnw2O7f9kZ/y0wlmElWX5nH4N9WfBzKvOOaIhSCAET8yN
obKBdiqNoRztuacXEtkph6JrrOaMdD6vzDMarALVJKZkIlUwCnyHKvDTM1wUIFzg
Qhe92jYQq6Y4gdhS8XOwWFad+XSA1QOruP7exuFOX0WV9iSVCPmC5TxA7OP3QDgc
pbtwfSkXqY8X0cEiJ5Kto5S4zSjuR757a4mzFvhf3TiSywgGXSoysE6Sswa0sBLs
hSJbJBlDGWvehs6f6uOUXQMYQg6mQjjCo3cfFFr9qIAgcWqF2fAuDoexKB+isd9E
7hq66EWGZLSZCE5D6IXPS3YQLPyJh+jMMWg7Q1tKnVG4MimZHaNceyh39vxN4Mh/
47rGM0iVl/LRsM7zwiHJp4nXahOBXZx1kqSGO3AnA70qZd+Jgyrm+pg0Fxl/7QZW
xIEMZouPtM86gktQCk7rzGcLqDWgUZg2WpyyKVtTEP67bICRKSuMOrPxRnbuF1qs
RoipYEI6TDkbMTt161PSA1fECt56SJIdAXqyLHEhn3c4C4ukhtAWdko1iEjtw+Lb
wk+Y7AJVGfxZzsRx9QkMETdRjmUSnOvSgqzFi4RYGYZz98XHq5VMFwSp+gOqyq8Z
OsxM+7eeC40GK5eEnxMUkZFVJZgXq0UfcWRTEe5ZjL09WywZF3pJMbymW0Kc0zAu
3bE0k70BTRZVTdi65IZdgLow1K2wu5CAQVfE3SX6A8NACUg6oWgkl2hxuO0AlGxJ
9hSwjLK3w4kp2iDien/AK6Qr7mjEHIKsCre8wbN7FyfntuKLyRqgTnOW1TaLAl0i
W6qovQvEvprZ9bzlBlSlpQuWwVm1QMkw9zjR7q7W4TqqTqt6Y43nhNqnvYa6L6ln
38e4D3IsBmO6xtQ/huN7V/PT0jLCFJbBmtfLnYQ9f6uZ2TwUGFansof5iigXNaoS
anMsaoDnF6VS3X5T9qvh71GlNV7DcPqc2djVuD7yf3XSuc1nGa293YgQMHiHdxpH
gcg3cXfaxfGsaPgg2VaIuedFV6Lc1gg79GWVm4WAPua2X0UB74mrKTOFY7+poXk4
hJAe5/Qfxq5yp3n0HRpruEn9ENrBKn6+1fpCVnqlslFeoUEEWqkp0ovpYsr0SRGb
Xed4BNCW0b2firEk4xc4s4CmfScyQLTxF817Hyq7BJNBnqC9ecOrFYA1daoTQwQT
kXm4Uj/mpuluRlH7CFpSI2inZ+mmFrK+K90NlhXCPdWCGCi+FNlAfK4bUx2dRN4D
rGplYWZMPomCWTwi3xopWSjD9F8otro51kQfliaNFu72ZpXdDSCvlSI45tT+55vv
fTbS7wjyxV1d3pJFfuLkLx+SeUwBNBrpULkPfC5KS1UWom42drQ7BlX3selhGH/r
aqpUIu569QYgCmwOsj+WNVOtzqXwnn/Mibe0w6UyIdCGJKUn7L8ltYzB26/b76B3
Ht2OJs6yfwelEUp/hkjydZR+O7k6BcrRv3Xych05U2ad/NPna6rcGePy49SgDsdx
+HmcYLc1t1DHcVcO7dCkFvRoJqfGxEiifiJght16m4WsrR/J0FzJxFtEKVw6WNS9
cR2JNn5/aAbzQZmCkIJeROGJAapTTurkzAkndUOZ2vMs3/vWDxb9I47TPvH0jAYz
M06VLqUUBub8cQkCT/C/YEVr0R2Zr7Xav82zpVmg0VM4TbS1K2O7YenAhpQSPFER
KWk9gIti+MTcX7TOr+9U5iSPh3iz9g3jTT6e7Rt2qLhOGb292BGtbf4HorKMwfVn
WEBJ9X/04H9O3SxvQwni0nlKVMF9JUONp6lCYqpmf21xLy0sACMA0se4NTHEWLkv
vIzzlalcE6hLjMYMAxfWsfb7utJfAoCu/hTd8pHM8lx1OGZpxTQDynk8d8nPekXx
kPwDwemdtpChttKKGlJTd/90FD+NlQuaPQIWo11gkb6ZCp7ZZswYlkw3ZVB2ld5O
VmcjCZ8aYqVDrf2E1BsJyxBq0KCCxEB3G1REictoi3giHRgvP6caV85gf+JiO751
qdsttLiGZ0PyLnIXLxOsv/By4UTA560+9UHq2n7yKW0a3M8zweMmfhwirY3uAbN2
F+Sc0uiuPdVUGGKBU68EAmQvl8gGi7Rbjo76EKJ8EbLmen+x5vaMUZCUJ0Q+/AJV
Z2jA7TPrMDkxLQY4beP8Bo46Pnc2ZZ8XsQOAP9xU/LCfnpyyMM+6vNgOJZwZU/uQ
K82Ai533dOTGPdpB49b1Df6iS3PKQaYrVZmFs4oxMf8x1tgGMfVgj3KNHoMvNb1Y
vNMBj9JNmGtKhvZAj4DcFV8iReMKNOTovSmhmlQKjfGHkIp7xWLc/3KIZrDZjyzW
wKUcu3PogbLyKJq6H1wMnjhYItvlELRYUFEIzhLZjJXn5+gbpWhwoRqGTEhjmPY1
u9okz6VBtdRa/mDsf5qs09jZuJ13gIYQxckmYhlRbtFyfoOPwxben00M14AjmwIc
MuPE6q5T2hmH0exPUAZOWsrzUVDRtixDxGC3WZhw4Tf8IOQy2FyyP5Ty1E7p+Ucn
Qi4ylmt5aTLsFuCeGTaayn4dx6v9dSNOhssQ5n2efn52oXwhygu5rwQCX9fo5aNL
bnwgRSucAT+Bpuf0nTJeO1kzj2UJ4jmQt4ywXPB6h5nCXZSCmy0Uc3Z2PvINwKaT
6FAVh2AanstQEBAcQm9ufjl945MJYqAnbsnqrYxvds8/j9hdJWDtXSHTom7jTvEA
DST/7e4lS2iq0cohNpBu2Gm3eDh/JvMBk4Wt0VAlGx7IWIQWJvsBUh5s6A+wvPMf
JFUDdX4Z+3acahGcRtTR2EfRkZMJJawZYxdTdi5lxjFpx+OlKcGsFQjoSunNXJZt
YaQH0x3yQtqbzWr6qGk80a1g0uKFNrvv+C1yiIpPHlDvcQhSuFZDxtqMWRLW4gRe
47Y0gmCkyWtuI8jNG4RfjU/UyjHqqU+pJ26TlSNSfKPjtUzodzotVEsRysC+T8On
xx8tStXDMbmYccnub8ELpvCD+M7QW1iknTZVRwTRFcpOg/uJqs4mDIIamubjHQC2
1fgGh5OZHSJy6S5QZ0eA3Dn2z1GeZotIlyb4MxkF6KaiVAmsCI8eFrvVynSx1kN4
ehorueZOk6K3KGLZ9OJbURI2coFdbJ8u8W/GZnIZrpCN6v/Bfygt0ji7axCgezG9
tByvZDuzJos3PHCVrghxGX2jYPwWGGscUzyrlBK4+LdX7Ca57FzmiHdY1/BwKZyN
brRvT4pKzeeix/id3hFyS4LiGzRPSA0S/aNcMc1s8jeGYlJWWtTy+zH8DrZsEN/D
5n0qmiLs37BHwUM+H2Udfc16lSm6QTWoQ1m4OxDR3oIe2VhyoF1OpkQNIaeMKi8K
wWgU1RXGWfLJkCJk54pkI8UAfkWZHE54h4bKUKRD7oVXiowhwu/O2bTuv0J+Dkyx
wYOeT7XCz7SXPFQdivdi8QsPgaRx73Le+w/rUfPV7y2qH95e0OII5P7wRxV2QteJ
BNVIvANs9pofUzS3gxjyVotuNtn8FoxvKf7anezfi73XlzwUYc1KMrtsNCKhSGIs
fD98/4t3+pXuXQNFizmVD7d2y2Si5pYZ9FwyiOSaq20P7UmN8vtzdC+rtbpf/j67
+fpTbGdF61uzj5kGfDKmjUXiaDFl7cjVCw+znTE48znAKkJ5RMiptpMQ6bkT7ZwC
opSZ2Z6KVTkRyAfxS0YDz1Zl2mM8DJy6LVK7enNJ0Dx6KQKOfZc/W2xdirQNBds9
DL/EI5dIUfm7PmYYRq8K8HgdTlx2QkIs1ZVZd4Cjp4tcoWNnRUYsBBOezdV3rRaG
nO4cK6mFEX2XZXrOHQaEIWEN2usIbjoRPduDSZGDAyZYMOlWMtMHSh0Cabqkj/Qh
O1OPRB+1HXvEeqwGK4oLuxwv+kjbl3194b/cwi1BcaA5b+v1ZqfTyjZ9A15pt1M7
4UXjYrOjJ7EXkKE5YOGUv9mncMx6KniBS2s5VVbrmR9VqWRoxgnLr+yZARCl+jMg
+DLaebQLxHkHDCmY+VZp7D9EbLYrvUVRg7z6sVUb6wtZZchunkd79i9AVnrl39Mx
xDpnHMwzRMn91q9Pz62ecWod30MJgzdTMvhl7N8/oBByP0soMmeTXoNSumJKOK+q
1Ov6TAvFxgaiYVnc5p0zG/r0drxcbNNV4ibTREXTRFAf2SlOYKinLF5OOWVPEV3O
wHluhDpkStOORacO4rshWls+XUlqNhe27VwiltpJmHk983Czily2Hb67/5qJE5ty
aQU/RCOvOdin6PV6xbB+gnzgRnJIOD2Pf7mWrZIr5e+fXi7+V9mKzgeSlpli3a9u
pe8FUjwAQ3/uPKzRp4ORjk6rMQqWZ6a1h/uRXaZM9T63rHMFL/FQXs/BBllvuk5p
iq4wd+KlhgX4g8V5ffMlZ49TyoHbVOeHDY6AebEYr/CKRoqSBv2lEXxYQvHngugS
hAx7fYbGQ6r3p1HiQkvRqjtTlk/oI12Y6BwI1cknnGwNEbxBhkGVy8rl520wstSi
H+7tB9VHiqp9hWJxBNWVXFG14p3GPw2WNXqsLWYNxYO7wDKsT1zgStTGNSmXWEek
GUOwHHA/PTuTwlfRDHm8TxWulG8J1lQsuZb03jAqGUQpiAQ8g2MbA0UP8dcKJXmo
/pFj85afUEWokAyX++DHKeBiQ73280BvXhvTnhpnrAsBsHYuWf8/SIJ64VZRR0TX
I5H5OCNT4QuKjRRpNImGX2XgVsfVT7c/Yw/AOH2g45Wx8rYpTOJncxoECirN2MNs
ES1JxMvTB4vy37QhP4UxxBzV6IDU28c5fdzVtAWEt0mU2AHRteztraVyztIvG/2c
GZ2UG10LZG3FmUV+J/JgC8/9TXhTOCM3cjEdhd4IA0lDCoCHHY9dPYfGkn7FAJ2O
1KCSCsvzmgPl50CrIjPmUpCA5LpwWhAi0Gso1pMeB3xu7MO9CJgAOThQaLzO/+6p
YyTnQzExNRQH+G1IfgtDmUs0tmRtwTgciTB1MwleNihR7/fX7PMhA0IrU9OAj7/E
pi+AFwcHqfHWzfrYvh3P6JmOzvtA1ODOAE0xasdwGHT3I7pWtFadwM3jktACW2H5
Yz/fHxdy5S1p0FrWfMgdeROC5kOx2YBnZuBaG5k6EXM4A8zTc2FM6w7vOkJxzHvo
vqoveegEvA+hP+7EZUzXl7rdeJ/QlrV+/c/ZPoXzT2D1xmSuuAtF32aTivo/msSB
vvw0hDMV3RiBuLUWN7JvhMMr/ZYHG7yzz80Uc0aL7fyay5CBMToOtn4E0AVn4NsN
ChSwQND359CrVc8TxLhOVqcv2RIya+N0bxjlGYetDvScyzrKmShIPs5e4zis08dT
Gwe2g33LIYvQWyk3QmMiTBvZh598e2P0Nsgore3eziWZC8Q7ZYxGSD8LsC51OPfR
JxsiU8mrBLA7e3vOPGUADPCKRlislSoth/kE2xfFZMtydoMxyGeZ6GvMikEj2bri
WEGO2mUebFiw1ZcUHppmPROjd4mxDDqi0fjOIVx7noqi2SEHJd2XZq8zA2EXLDH7
RNlELUELzwe+oc9q3OoX6ANgUVHgZyMzKROG8TXcVhnSFkWk8+bE1tsTp43RX0mT
/1UHZqPjmnHxiT7MlpBOzyZ3IBg1TFBMd7OUDrilbjDQhjajRwxEEsnN65baTJLw
WVahNpEUrSkirT3j9yoDS5jeMFgmJG4NdODuhlIK6vi0tia25fgjbisFEJ3oEktG
nj7BROz97MSE1RTyVBdtXi1pzj/DbUmIg2gEDe07ZuXvHEbhDSbp1SUPPCL3bNab
traVZwrfqDK8OD/zsOybCVzHJaIjkSn0y/Fao/v9akwVfo/8Mqf/n795+96BrXRO
tz0EcF63b5mfRFFXJsLij96FNx5OV4S8vqTLLrh4h4j7aDowjeXtNaytrFejqIc2
maGp3VeoI8AuW78wqFpfivjJuvnYWTlriNUHkZIu1BGFI/MFEurQRmb7p8ojsuXA
lmMq8ZPs4NSizwVZ3QCneyrKT+IoLpHNOf2bIfrZCz5A9qbvzIK4q0ByqfuC5h+I
RDxmh8Tm5lLtiGISjR6GiQiiQzcbDHcR9eiTRQq6VURY40yRpGnVRJFKMOF08c68
xRGW86EF01VzSvLSp/fvpQhF0clTyfSLYVUB1zlAzl5pG9c0WQgdX06NAYgjvB2b
BSy4hRU+FSVbCbqKdYWSCtiI6d9W3eeC2tANSWBR1h1wbqa1og92bQNV4pC1FYYF
dotAXpcxaJwMmIeCtE9gT3L4gVw5qPRfb3N2ZHNJT8qi5G1IT8K1mi3fTqxsYx5n
hLkgwnHdV11/KX3TFH6hDjy+2FHJWB0erxn+7K70eb7KYM+FwDGQpx9uPisaFH9i
FsUwg99rLp2zH5jMem7PBv5vt227PbcxI5Kf1smczSx9f1FIn3pnN1UobaBtmUgt
bdu7Vcd+kaDkcQuOIxmWnIG8MMkubdDJK5kuTFjMGYv+EVq9eQZ9EF0W3a2yLm1o
cfEdqFqC7g1baoIenwxWLdw/Ht570mxlxjgDui1t9XVsipvVIOgbGWqD9Ws+Me2w
cFGhOK3iV03yE/zKyZePUwrpnq0GjfqIKU+OAq1xhK/PeXATHc+PuP11fbQwDXtj
NP4z0dR5CbA6o6rjWlks+CYW1+JBzuEcHUxWvbHY9V6wRS50RApc9q2Gb9tC5sYI
28UTOEXSsxU7074snoF3YzT4q/Ac4d0e8+KhnUh/ysJBxts1+PMG1X1iU0zWobPy
piq8R+SbNgIo5zNNG4GkUpTK5byxeMA+u7Cpn0vt0vcc3g6Bg9SV81PlO7y+foBA
fEU02d0aspzmEzCmzdf+G9P8LE3VWoAwf/fMYw5ohAWl8QGqMX2Vx6SzP4+94mwh
BUNMCh3UaV0mRj7rCRBqzEbuwf0Puce9r27qEWNdOSH9P2Bi11Fz7LyjtWqvMC2D
XC1ihV7uWVvBJS/8oW+KJFCAiARePXclJLhzv3L2pABWVeMshRPAx34d/ACrfX1V
U0j8dWK7VvjMnY6dZtbSbPfWRJ7UspgAji385/aguCaWQapI/rgLtLIWYU9Zz6wO
gdh3Uw9HcmE08J5VWXs9XaMLINq29AYCObRslaFTcWKEexwv2030ZT2luhB4QBJv
uHY2Urnxa7oDDS5b7in4Ah1wI4LZoMdA9xyb4zHwnefakjDzE3hVfUePSL99yTHD
bvqxPbpP6xlkzKlMfxGmklAE7srhdCCt338UbFDYBIgwDORtTIwuBH4PWwmESkjk
lueV2QYd6DHOFxujZyOqTQMO78svZ5UW59+21mwnbmhc+idGnFOx6A8MXc8ySMAh
8i+HW/AiJamFbs9crsCn0yp9pMU1rMByX7q9p8vICYFKukXnh8Xgru3JxVsNjXYG
8KFNNIBkaFepvC/N3oKAkl6fz2MgUB7Z1kaVk9+C2tMg8hRKo0LoM0H9alQGuvYY
Hi43NYQdG1XddW8aeuWBCM2Q1d0o7OqttKwl+klk4ZS5w/vFSsj7TyK2dzeWwlh2
VPSMCg7runurnZtgH9SITlt3KyQQbIaidQeYpXPLvK8Mmmoni7za5Xpb54IKQb6E
TlGzYepE9bGiEBjLlBmX6qrr/jq7MSj5EfUe44rlaq07nVkKisFmgDIr4biIZLtT
X4GSFcAPHVZq5uMsyLJj/Ddb7LT4jJvrvYDMyO5H4lFv4QdVvwJm5GzkwFY9E9XJ
JgLT0Xp5B6RPxsCizN44IJySf7Mrk/4VbPmXmEjb9DCXpHQAB7oJoX8YGPpMrbJb
3xtULrka4ul+WgXy8awErUQbYTwh6+mM8CArf1nLPe7y/KxmdNegJlNJksnBe6l8
FvMf7SeUdM/W1/oTrpLdXPtvwZodwN6/u/NxWxhN79xzm/BAbbLyfOwzcNvcVrZU
/wJStZNbHHK6P0Wta5mQLhinBOAarx/QrAnLo7uG71HKfnOvVY3AZf58/bEhju9s
/pGDxXdODCoEcCarInqTsH4Maw9LtYGjjmlpVMZEDhuKakTcYBRPH+2Dw3EpL3il
LuywHsvYA3atVF2sDPX3NitCuGXXCdpfMRQWrNsGb5t7UW1d0ZPxECfGFpfTGTEV
s+EMY/4l+LWavvgRdAwt4b5qU84znM7b3A3YXfyKVThDXXrdYd9F1cAtHsybcyh+
FpkYDSA/Vik3fa+VuX5GholYF45HjzqAurWEw2vU/MOpXiMMmoylTIXVHIow0lSl
TYpFgK0imT44+YPs6WKcRaZT8oVZ9+0X66vRkEAMRzRRtX34LVWtVAHKyFgLKOMG
YM/41NsKto9WpICp5qIRvoRz2zXifmxlvbcvGb7UY6xaMNURCvvz7caMtb4BvfbN
mG1yiZttkDlBPu7jCIN/QiYDw9AzBYdI+h9zmK4gWTFEzN05dglmCjejSAMy3fhw
Ja90S0XmjOw4GODT2FeN+13+Nseicz84DKGOJMEm1t/bdKaaXBSLXKsBJWY8GMj6
YJo73ouzgb37k8ig8mxDpnrtxUApcwPh06Ne4keyZSAD8TdV05825xxgoTNWufCN
QWxAG8m3jiJN+QMOlRwtF96RPDbyoEfxEEEpZ2ixpMjh99lsAbbb4+y6C/up2OsA
Lpfy1CNoTRqhWP1p2PPSxp3KgKNmIJzZnaPOGTb2HCTbGkR2W+tACzyz1boafT+4
uRjkpMQ6A4LlVbjP1mp++bNzBcI7i1wo0cMHsitIFucmek+G4Gn3KN6qYt59iQWW
ngxvB4hla8O0VGu7nOeGmCPmwEMNElkIEgo65xKcqJbqM5EUwBlknaP8x1Ix0uNT
WJ/pXRbxzdCt3HG1nEL48egy7uOuoF+DyFl1IqH+s4fOmoOgYsF9h2iugItggD//
hWAObLvhUiAM8GXply6S7cuXq5989oO2aN9Xsz7x0F5z4ELOZzqelLkAnrhBSR2W
2t/pYiDGq3g1snsy+c69AQAZNFxbdvoPSi7rThEdyZrRpR4lbnTXUPOpNHcon3zq
kx0MVGTADF36mqilnRYSYB1MbX65V6UShJdf7Xwh7dlIkTARww5+MJrOjDZYSv7D
Uih/CbXlwM3w5fT83QoSYip93ecLXLAzNp8EI/HFLEuGLVzUktXl3+koGVSAYSyb
c4fyQCF7k0XWm9WGmfvHJDz9STq8rUIzB7vnEcSIWwYqnKsUvg+GL5PYSIpqdJHj
kZrc4fhXX3vbcMla5QGA8pKz4NbQ8jkVtqJRGMAHRaJ7uk2nnSl3+/v03h7DaDAt
7pvi4DibD6NIHXTUUFO2BXyXb3PMX7eZa75s1ihdCtzQaT786b9RLH0BCzsd36e0
3WHThnCLtDmfysawVMFqvTDEwkwoR7ZW+McsM0shjCzdMirlKrpZ/lZfFO6u/Krm
qtsdhjW4JJvR1q4y8eYNFP1/465dvRcUlBVDjiFLKw8XEbDKihuQYJJcFgI6290Z
aZwihVOI7/sW+lxs7LFKzwTlDXE1PGuuqJxRgBOiNNO2oKJw6oAY9hpo1qtbNjZD
p+jNVDoKaaoXwhakUt6Nm5pzruhYFhFk4hBhOK/9nnJeXWv8ciGUW0TFZBjpXIal
+Wh9pg5CQJ5QqqCBMDdbJA2NOV8fQ021Ujt6iouF4SCINkp+gXQEcGcWvftvEfqN
YAbacrym+9zCm5VTR9dkHiBnO/s2lly3qHcajcjjMYYHo6oKEbx9UXy1oYtHN7ct
XqLoQnp3vJKwsBh7G0cb2BykmnT/Yng3WK+5FCqsqN0Fjlv16t/7d5UxlVYOC1ER
4RLEIlOX6uBS5/2sd8zx1BSCA2x75ozmbkLqA2zoKZsfM20VVvCK2GBFmXYROpz1
GsynYqi0z6asC0mJNiZeEilt2wj/L6xs2BiQdQCTDbysAgRLwIFHYIsQtwoNKPtX
L5s5gak8oDekp0ydh7awjj6TINkdiYS6QmsOA+XA37LIavlKBcibJnkEQiabww1I
bM1l04WNUZMmOsaiE6WXI1uE+9muBN8Qn+NW/cVLALd6OYiO5mqii/NlaR2obGFJ
LF/urSN11F8rDsG163IDphW7HNEV5ax1QHn8hbAwGizas2uI9Vlm691rEVpac5OI
r/NOlMoyd68W4TSe/7yKn5qW+JYrb27xPJZcFjAPLVS+xsXCr+S1aZfgW8iYYVze
YxAbsBCAQGA67NnQUCbwERxafrhpX/kPPOOnm4VzDZ/uV0eCPTeVRwFp4sNBFz9K
UkN2fZxoMURVznZ8COrUDHbg70TsyhizGsNmBqbM8JIhFg48oEaqICftLAQEDJBm
h6I7vdhEK+WzcfpY+nGApuYuqejyHbDnqM9Wwo8C9QQaAzvomTlPawknkZm7jsrV
BbrZ/RJGvKz3Q9CNSUu7Y1DPMevT56WAvlYFzqpZn1BCALvnmsvcGhYDxG3gFPb+
+HFpmy6NCXyGectzIR0kXHagWYdwiFZYyJ71OVYuKO8Jre3nc1GPQm5qwoprQgK7
P11DKN7VuhbMClA7/g/yYmFn8wLaHgoAkjCyXfsCJMTYZet2QhyhC6KooUiCpmwO
U2RBa68aLOzQFHzRipEj8rif5l3+MgMJJ6gv/M/+BvHsTbhQtv9/S2wE2uIqA6TH
8AF6NUEgxqnZAubKVBAZfDjHCtU0dvRP4woJ8Glc4pat4AncE1PhnOQMnxbFyphR
8fm08WqwEhtYP9I5+SnIOF/KRMdC8LN92D4mrhEF5fCYtNOUpZK9Mj0JOSNfFK8k
bt3yXnPCmk5hmVtvRnZJGuJ3we8uZ7CKWcJmEcaUkiuyh+62fjFidnBR5rjNo5qC
UwIcfQGwpiTjT2yOddV7yQS6kRMRgTfcvj38kUJcRiaP28y53aFg4g6UUlLkHUn6
FKFlnar+JnmyM953a4sfBWk6s/+V+sKvSeZeKUsNywhqYSsk23NWMg8y3GN9pgmN
opn3eKLhYAHGYuupdiZKc41Jy3NQREXevkLMUSVq3vCdmk0xE7kSo2k8Ew0KrrRu
KDNTxN8w0y2mbiaZDGiBVSNjutyF2GdUCmOuFz0sjKk10wPpKC2kIdR9Wn53mr5P
4/7dbyStuNP+p7trnW527bsUz1B17K+OHkJQ14eBrD9Iipeab4Z73tYPf0ABs1SA
D15WlSa4+pNc8cb7SkpJziJH6nZyl7YthiRz4RIDxIEkPqVGZoQ9T43Xt35n+8uG
lmqP8Nx3ruo/fus2xbcmzoc7X50OKKaLp1zVdvxruOqguzF5sjwdL6zhJLThK3xS
0wy/0FHCHGC2cbAvSTxK7xfxQH6NIqDW3ddny6EZekPAALPBHu85M7XGds7U6998
Spcgszw/dD0drV+p5oJE4MRQ1vPaDgYT3HQhwzNxDq7C3i5N+1A5y5qlSQoUkUag
jKJjpXTecyKY/QuNkhYFBHjiE00m1Fm0WYiQc8hR/pw0E0FyFgSdTdfK7s3OoM/R
QP8uGtMa90gdISYkmM0q64yZ1R1BC6bu1Qtsc3VpdmBUxOstpNvHjAWRwNNuQwlv
Y6zCi6nDMc2elstZYYqesNwj415nVsMNSGI8/SRMYzMBrw4krmLK8inqH5ydDW5W
ycvszz+ioz7L/+EVq+kC7lIast+YnRKMzR854Q4FJPGj0xtLVBkmpwk6/gfn1EYm
LkrwFPdHgj1To80Ud6/qloWbAAQfWGuljHUbbFjFhNV6t9jUiL9LwjeV5s0/KoXN
f5z3XQKJPvvxxPEyu3gqTNH2EJ5sNsPVEcDq7czhcsQLPz/cjDge80Mz3b9zLdJW
a/C6KKKSDyVeWmjkGBTtoeK4eIezEeS6ZHBAAG/dynyT9++zGdybH4tqUVnJ8+6k
tMWdRbLduScnknp6NW02GrM172b15EgGL0VukEKeoMVvOB+GELr998eWZ9YLrg8X
4wCUE4xoUGAZsxR6mTqOgN9TMsLgB7nhtKvhlhZVSotB8GG4BTkZ4VSd/d/3VBdr
FTHntkVKIryEbAfnYBZzk5FxFJuspuMWZtQfe9rgW+v6noU2DBxD+vFTuqHyW+yU
xEIRMzr+WLxLYnA4xgMDPJ0LklBHo8ocl5bfWvAHA42wSnJgAHH9oYnPULqq+kUG
WSLdSonjV0Sck3ksTdVtkjaqNN88ky/iZouVmJPq/t3iCrnSehQg3GvcvflaGXg0
L6r0qVctMNVPrc/EJHVVuSggGjKWdpDk1I5Wriw+mkdmBDtd3uv3ruJUJisHZztc
XgksSvNmNogsLxTW4i1SOinScR/+Q6PhbXa8hXLtD2q2ad83YxCH7GvYr/SzEHTM
0VjMAWPAeJFqBiLg78ZQuHvw6iWFCz7RtiWo/VqKK3bSY63VcVIgPYjOscn/MJBE
mEuN+MioarHO1kn4K4LWBKGLdYmC4wzxFUFomDHTJjLc4pq2seR+VEMkZC/+UrFM
2JzaWUsuuWtSrV34ylnR3ySppvyVIYqOy2qyRS7l1esBcUVoi32aYDd8CiZF0l4x
U4Y2gGpmIIPbDDDAHgfRRfqDPOlDb4Gz8odK8xo0hE+b9BffeBBdzN6bqjUbKPSe
6vbSTklpnvaMW1SnQ15kt5orpmeJLlzmrX/4G4z+MyZhOIn1zzDGgHVdxJHZw/2X
Lksn5vbkSSz4DJcV2WKtxw7yB/fhhAJknVHxouYXULPKDVQ0rm2T8t5SnhCpokB+
dgsfC7F7mO7S35zELsz/7g9cckDioQso5SRT1y9owhaZ1XQ1VTAFGfmt5NcZ0wJP
bqRxPKI27oaqXxANQ+7Q8u95vSyHO9aiBqXAEKcn3kd+YLt9Q7DXxHeZhqtX7O6V
XvIM1t8nWt6tRl0mQsODPRvWF/cO2PpTwVpYgoRV9sBKP4iU5hEoJjwPRCbAeNws
ptRTxLuIJCvf7lin2utDxygc6iTL6Lb6xxPqVMSyQQvuFxabH43sAfweNzvBBz6I
tBUCzDuvw2F014MOuUp9r4wCE/ZjCxjNs7Qc9XBLn0hr+cpaAlziIgiQIp8FFkWS
BblSycbEur2XuKLchG/F8wv/GS2fe+uRdetPBjC7LLBQrD8lyCNQ7ihRrDqNuu5R
0JoQRbZaSYQvCdm5NQUWeeD/5ApOsnO9nulgAuFLEkXSrl23YsrltB3itPgxAQBt
8WCaFAVv+E/tBsjOYpXZEZ5rZvpsIS3fJJ9/RaZPJO9mXXmGE5NrZP96NCKqgRCt
HQJl42VipqNza4wvqPOwVujIACZf/NRoM4SgypCRfPAtpJZ+JHQf4A0uwFoYKM0e
TlGDWm3UwUswGLacpfzOCM6IkdYevkExc1AhhsDMxmvNGB86sATObop+7K5xNRVK
X1Gk++9RupkhYxxoCcXgBERAmEc2WWNkYt7KqK6PIYqa+haNH4tebluP0II+DcV/
x9lNgkvMM5wwPjoaiV6mIx7xCw1Mj2Fk0rJeGCI+eW7pBf5zQeSo1fAx7KQur6df
vXI1euDFPSRYSYyIgT2fLZ8GhO+ZNzx1AFth2+FDaJEgNRiYtPBymCD3DFQ6b48w
I9iAzlKu0lmPLnSjzbi+Xl1TLIzAwTKYRlUdj8FTddflv2Z/qlhky69T7QjTNUxQ
G1VNYMFQ2RRxdQCz1+8wNMwPec7QTxUP14xUrUQaPLIXFITn9XAORmmI623+aAGW
w6MTTsqAtPbJDxV0wGssZQZZjaU/0RPfFSBhWmY5rvd84zwIUvAMpg7cnRrYagjS
fS018qWygKAObcLNv1aGeMDSk/GPjd+iRWh0tZRMhdpKcYc9gDWOjwP+/7vyMU+q
1s0cy33+qTyWyHK29MpkpK80FeFcNrEp8HZAMH4OxJJrPBXICk6SVpDmsd4+FjHj
luo3V2U+zDD54+EIuwk3BP+TzHIG8frfyJWJZbiREAPqyy3rgYgvCWj61maFb0Os
HV9NVAXapW7Pvo6DKS3HymVzPrWtUxvg3l/E7808e9XRvLKCcMPoC56mMceI7vCR
SUrSTqNYa4BgcQ7C+aQFsgXV3acd5wid7OaUG+8OijhDuWNnLqN+TaQXp1Mpud0E
85m9sGICR0J060SjeOXQ0OF7AwNGyNzbAX5XfJs1eqTtgP9n34dHx8oL6irLCrON
H5EPTMTWJt4FvnU0JtgI1dC8zqW78oiorZucqFxqUGeH/si2ldQdV/5sMZVfAkAF
t5dq28W4b19MjhrAS2lPQhkscI2I6TnZW1qFDoX85GPjqPw3UzbVZmmhkGa4UON+
rpF94z42CNu5I78oY0DrLXMt1vejwh8r6KQuMLU2cMIDlb5sBlM2peU48MK622Wn
tLlppQ36CfuqVwv7ad/9psSwpqS0doEA6vHASlhpmb9VfH5zBBLcTdfp5hY8BeRm
+RWNfrSFHMacfyIz+eDCjK4O4xqYcsTpth68wC7qD31NbNw99l+6YHV/MxKEaRc0
3xBH/HXfF96MfsE+6grv78AjVp/Zf0Zc2+rr9JMwt27WWf21Pqyuo84jqivmUu22
5jW2+1VpgG8P85Ao+ni21b66WGkBgt5f17sxkhs5bQUZHwRRnfuf+49I+QWzfqLc
+AJL9JMDIl0tIULl0ByndFo+MPYxRc5QqWqERL/TVJscAFRCgwkIiq5UKEThw0MW
GcgUsJBLNq/5Y7lyZEGs9Bm8wn9ykg/Zwl6xCzSTAixOAXzUhKZ1Pef+KOV4nTyh
XuHl+amCqdS5/03ITxYVTI8sYcR+EEUD9qHY4jaGQptiC2OkJcHQLUUQbMY6UP5k
qHKz+svYaddbthjYZfCtYtvda79XkG76XFSBYrC29wsbTcDxlQvRUrAHPYqpIsGy
1z5vDuiijZyWMHkbTu05eC9XbLsN2isFw+hijfODLulny9XVcSnvPJ6wv0KRjJSF
waD67DgGsper7X8Ign0/e/++X7YMAYDzzlwiGvquMX3UzU8CcfY8+qOEyVaZ4Bp+
WZ/1zS1DcQlgYeGMbWes04PuZqSjC0V3v3VCizo8FrseICe8+eLoRhyRj5QVODBN
vtGes+XR8tQqDHUmlYyScGkpPCkTJjMPF0PXfuj2WRiczNqm6FcYNEXqiDRcuPn5
Quzamw4+rS65l0shWwYhjC460r6Pq03eQmBsAh4ZGg9v+E2OXiDIoE6HdhxeZgMS
FeZuvMuia9Nel+epkhZMgX3RcYGhpU4UPSZaj0hTc2cJZesd65SUvbXAOO+g767C
HE59vl2WmQjWD4n+EE+VXK+i4F0pgrYo2bScfL6izu5YobBh+mhEnyAUV/SZc5BD
Psj+eQph45J/wcO6oeBLIBDbXWjvOU2a6M0ryrZnHg+qwK7otZbu5ykh0fmvTMzM
olMHtKTR1it9NmQibMc3sE5OPNRjcdj21iKQXPbbj2mS84KDotlmwoVdopGvVfRD
Kh1U7Whp8jNROdIFyptETou8AV9W8kZTiauRgp8jffPLsjYf0GfO1SZTc59rpAPm
eZf1+Cm8yD9XE9WDesq8D8vbn7XMYGfldjEO1bE9aXa4UOWWeFOmovUXEQvASj6x
pRTXAl7//KsQaCICCM0ruQQzOc3JqSphg3ee1+ulklMbeL47M73yCszyOLO48xfK
AHdF5ULLpaVgoTtsdqYyWMvrdUO0cEAvfoPo9g5ITv6AAqyUo/cMcmVwfJdCSEkF
6TWghPKg3CUy1pxvgcjs9/QOHlwuiTuVPBG4yZgVd+Zblv38pyfd7N2OXwSjh29B
jJOyviwoAFX6fYQ1NX9I7PSkD1Q5JA2M5tMOtLMJplFoPsP9igrK15gLEv7Z81Kh
lPkrqxomnCXxPjYyFkAJ/G1rMwdojpwNrEIYN+DRTVgAsFnTovIkcoTRrkxsb+4n
Yzi3Ws6eNnkpoO2WUUmbjA2BjSNHUCbhKPfxkBXZ7LKQQeXWkCohZM5ikozHUD0J
lPxPFdUFp+uw3Ps64/Q3mt6kiTIfsgx5lOoy486+p3OTIKl5UWFnWHiWoXUOz54m
R4m3EkJ+Tbl9uk8wR1fmVB8ggHihdp2J88sXe/pyVD0SX/qNiwb6QHIW0lg26Z9M
2OMNd2gSeHa+I2UK5qwUoe4ea5wRt9D9dFsovE2WbbBVIu+yXeODcu+wc/qbwUlg
wLKQKzVk/ScSrzkziCAq1Nzlvuan/RoZ0wlo2fpfU3pRRlmzPcu4o0PjFzGvvwSi
D+VyYnlmhhqbYLNMqvzLpGWrtDo3Fk1nTKo391Ilv3627wHPxQr0nT/euHw8mndF
y+66pd3+aTHazGbMI4tSR68fhGEiE+Oc9u1i6IYcYKd+NuFZZfdeN1A/Zbk5AzFZ
qlP2YH3t4uhvkb9gQYWjcTO25KVkX7BT2PqoKKDb9QruOakoAmSY/mo2EiWoSnz+
Q8wgZgDCjLiAE8eKakUI9gmAXFDZFUyNkXFiY2zA66xTwE4sGnLUUqPuoNZj5EIg
8H54h/VsGXj6Qm57TO+5SdenwhZeEfyvWMY8PN14RZGWlf4ecwiprT9UeV3RiSkM
TdjcAm8s/b1Dc//3lEg/x7f7l2owDm89ytwaJ9QkCejG+Go9ZTtX3gRwRsXxsfvB
G5kXoTe1UPNtDIuGBiIsgooGULeBBgN8cHjnPG7Of9Xsly7d7oTuVXz2Oq/oI9j/
req619+i+tRh9fDrVB62xRBfSXCAI23/yKXZ2Q5bfDOoEiLoHImmwnBiHryIAVd5
P5GuvZ4lh+u8cdBP7MDv6q9TB9rN4cjLdgZtsab0jaS3u6EpvsuFq0QSWk/vHCK7
5bok/NP/gq60NDy7IGN22zHk1xjrEVtcOGeeYLvy/7Px4f7wrrbyLJocsQFmdlSa
sCEtY5/2kaxsHhEurZBXlU3u845SQNm1jYM44rYsZxxl8SSCBJfbALbhRqVDBI5H
KVb3JUzyjL0rq5hqQWQjXNfNzTDdYxyD5Lol3TXUuetZPcUZ255Db3iMLqUvKFvg
6pAxB//fq8uuQeR4EnWx7GaNGsj6f5GieVgu1VwHzOaFLCciNPphjDadErG/oRed
/MZ9R08pJtLjlXnjN10KIyqdlxSBg9M9kp4Vq311sBjnBeb44Lr742O7x7WMV8//
323LYf8TH9tHE3eCAkCZedvtssll3xcFWC6/M+nfaaASYWLBdAwD/UT9qm12iRbx
jpEbW4+3Hx0BK/TYk5AoTD8sWHCrcC0iD5yIWSMeWElAr0CrF3GsLqPsrhQv5bHh
ijnN3RDT+0xoB3I9MuwziCuXgcdOvLGKD4IcZ5IUChAxRUF8u8WPOG5lkVga3Zr5
/i8XAOSZgBSzUFv5Vo3DjycFwnBlXbpN327emYvOIxhKjq28fVy7850h2+WIP/JJ
PW5TMVNoV4DkUX7FENWAS40GNi9mManNgbK+85+wGNmsRyiFfhZj5VgnDqPcs9X3
7G0j0iBdJ4PLMPB08ppbU4PFRK9vEZzuCK0cgxXHy6LmF1w+g7YRK+Yn6tn/tNx9
IyRtPTLB4i/sD2aL/rUr2M3r1gH2SPLFrPf1HfEX6VFbFeWhPJ4klfSPTEIt6meI
LZ5Qao2g7tqOO2tqJ2XszmZQ0PYc6QRBKc+KDVQE0PgthYlPov0mr5I+2YTZiaFw
XheYbhA1/YNCTmX96/cvKzXKi1RISlUppFc35jf/TZ1Ec5e31G5vcfeOB2xlCMZI
OK1wAO13fAAyEPAlNsi9neC2bHnyWzY3IaZzupnBBIrr3Mm5AiQk+vreH9dNfkGH
ifnJ5Pp+sni84Nx+qCVnjeYjD+Uc6iFa6Ax0bZAzg2UXxqDBkLrNMMIKl+IRbIp4
RkBv4xBpyk88Zwo3k5h5Bf32WKfJsCZYy8Bk3I0mNCg6bsn18pmFNuOWVf/EFb33
xtx332o1FydWGvJRlLNp9TxLikTHa//KvBssZfZY/iq5saL2Pv+4L2Eg8A5NwlHf
FNl7fmOUecuCoZ6KFce/qbya4mA4eYM/LPZC31PxJd7aZVxt+Y6HDHOYgWQribWY
KLq+ykinilts+JyfbKN+09+cUYcTn75IQZiO+fzWoRyWfWUGddsPOQfIkvYPItkm
ECA62xGQGkZOKNcKmRVCeo4zN7iME6IbmT3FahwGnSvZnxtW7yUKQrqxEVjRnZ0J
cN1TmQdLB+A2vYVnvSSshCljyZi1RdcImpHDNysfiWdLy4qosGKlP+MUYzxax6gj
h2GSRyWuwsBto37Ggh7i7bdFoT2skEb++EiYO0y+55hDMtbkfKcSM0No6YkoRTM/
hwG/J77ZCjuapR6NVMlz1bEduMRN/HvYDdd3C5xhvUlZ6jZ+imF90hnxTTxtzQz6
Evvv0nDUIok95lgxrod5DTVtuEq02Mtk7luY4YBGrohIM/WGKuq21vED2f65kgNG
+uXKxMJZRMVeu+DWFPp3c2A/pdYVDjuYTN8PEvX1og8u0qfIfWNWWpF6jwnSMwPJ
/tRdgkue3MmlTcHvh0gOSxmofOCuSlETNQNNGM5KgXmWHuiV7fxOJUSBN+cChMMM
JFqo1ATw6q6xnIcaUtCrzO0kKDVsAhSDJAfL5jjYIqSgITAM2zPReJfumY/Zp3gG
N+IYlr6uBJ1e96kmQEX+MwDMpXJdOCGnIYhnMdJsvrYKz7kCUzqaDUwyxUAGFjK/
fqRQzEya0Fi9RtYv1+n9if/wBYQS9/uOoR/zE2Bbs8ke7SAQGQqFgiWRa6t2h+NZ
DuMwHWfxO8Do7QDZASiL5KaZXZGEjrXjaYKCSQ4WfF3H6mdAnadBnI03IIbkCzb4
gnC/8WmvOxCQ1ya/P4VH5L3MkfCD3AOpdPk/AdinAgibZ4V34O3BEAKUez+l16+A
0qRpRmtfIQ8YZLcUATHwPSewKnX0jS8M5nIMyPcTjExbCjZk3EumSriVapGBtdFi
0LXF1toJ9zKA8EulBagMcJGT18hPM6NNvVer0YMN7+s/1+OqJjeBf7VhN2Yilhw7
OnEUdPaAXoMbZP2F26nSTNe7WoI8U5KhOXbrhEKFUQIs6ttZx1r0QxoKKhRsWG9D
//CmnI6lTVq4WYjMmHqBc+xlzIa9AhaE69m+DSh6Oqbo8Mqz8T1DOE9yA/G5JRzd
/a5BYv3vgsNQ4/WlLrqWvvweMFG1MfROgcrisCmOS+dFo5/EGTxmMXnrkTH8gnKj
5a1F1eU6JTdu2OUypGx7jQU8YF+C5SECa+CbqmNgw9yPRVlUC8Z/o9JDjBveP6mv
/PhY+oyHgeTFle3zcHOGudoOD5a/Zk5yyXbFjALG+Lkv945iLn7VBPr2wYV6wdwY
DQVIKLwbvP2dbPWmJMxPCKAHp0ZZ1JbV8iuB6qUIGuAvkCVmk77jlJ8t9rlPOP5C
CkkSJHUfzNM7o6mLQLt7AAiK4FFsmlSvCgQhcxvG1Ixwn7ZC1p69LkOWWhRKwleF
pniRxqxJNrHfpRuzigFTGunmNNU7n+trcZfFsDROwixGKuWQIAxeXx8S25bZL7ob
AS1e5OSDs/W8nYK9schmPHV7CHjtTDxIJT4r3eW4ov4dbSNeywq2Kvl0GBcjccW4
fu5ppsBarJ6PvqX/Yu0b1dfc6j5utdzFS9BV7pJdx62F8eTs1jLTuLpjoREIdUxk
Oe1O/WU3XWdciiwuf1ZSiEivVwXFV2svvv5IuN3W5HJ2hR3869Encvm8WLH/eoQN
pAckLeOUn2hIusP5/M8HeCiuQ34hpuHf8xHW6BJ0ti6NXbdTma7u6OG9GHPAISVS
JhEubebdeqEMXBv+xQxDtMe+RqJgQsiVE4p9JqUoEZabsazC/LLH2TW06yQ6+1/S
FOhBaUTPKj90JsAg0SXGFoOev+sCrqS6yYqvohY2sTbbw0X8YLLPZOuevb8Qq9tU
2xeJJ4VRCC08JcRd208UDo5wUwnWowXGaV9fuedt/0LAE1dYAPODR4fQr/OD7/FD
yEJxvbJn/pDWh9tMFgnTQxJntkwewOytCADcZ8OK3Lq7o46vHM64WRlMqkE1dyXF
5b5R/Zc3f16yE0aq2n2w1uCLNqZqATQEHCstOXyEqx0ClRwvVNbxwYHK6iGEDfer
4KtrebB6We+85vi63aaxTKsHf/l3JaYkZAUwCBlh9RHihRL8Y0CZSwl5vndr02TZ
M9fG1GoVO+g9OInpb0rbJUaZKGfpo0ViuW993pD39fDDjB7+k3BsXQXCJGC5uzul
4OCpzhHvprQeQSU8V6o5F2EjJG9owxS2Br3bQjRco2wzA1MZmdUPpDPnVck2a2I6
5UB16Z+RcgKZxzYmyVnFe4u6ZGDi4FmYrkSfWJAF0e4YsGOXFval6KEtmsI2KmkK
g+0D3POTweR592qiX43Gfdfe9Lwj7jWEKXo9D1at6DJwWIgX0Tq5ZwfG7o6Ty85S
VBq8GrE5GfIg/8ve5G+Lnzvu+e4N2h1MMZKL8/tb1ZNXdHi4zOtRPTJSSugIIfNP
hjBIhVLC5sxLZf5M3KXkmYLfqqXylgpP9Qevpn8gjqzReXR0QBg1ePx/wpovzPdf
1nsaXRsGhhaJvCmZcgyt/VkdnLuUWjapXZ3PiZdTRoGsAoy1LQwCYqdDu5dkxxIW
9QQIX79ARzfPx9OjwQt9iaLqFp2wee9rW9NKiv/MDdMLNMmnS+u7ATDWDFtHcwCr
p3TBoomXmy93jddQ7s9RXANVjWlBjk4vN9RHYaNi3h+VT/xS959dnc03Fndaauww
vsdjkhRzLYH6OuoYxH51ydhzIQfSmfBt5GjdPifqZm4CQD9wcplNZ8npmpCkrRpl
MEHoXKArWaTLnTUqplWim9Ls67Gz6GelAL7TAutjALrhZ513QZs2Rb/9rf/9X9DZ
gku8HsfhnD0uhiKNfukrH2QDEQeH2vifEleIfTZXe+Tu31/faFtCQTKu14RCJjOd
Gw1d4Sk1CXPewi0osuYzsy7/xLQyn8kOU9C6oBOUheT+Yh8VHTpmEkGvqCoSMLYd
cNmxN39eXofvam3Bba4yaklKafH7nvflHBpoyE2gdnLXE0sHM5gGIdnYVlSnOsvJ
esZgIxj2tUDa3KUkVCMDM6H7rn+0IaWs6rrmAyPZVWmuiTUsMRwdHmnj72GYoS6F
/sppNf4S4S1quOLTsFFIei3pkUwPzomumAk4tLYPsYliGOQvfnpma+AnTdoFAqxU
yh6q8vT2wcTT/7RloeHyzAiWLy3Ml5VCvMZKqPMv37LDQYl0CFa11mXgVSo0/S5A
Q6bgK4uSt0ea3J7szIINMq5Jfz8pmC4FAqJfAwqaJc1ZzyKPO52GGB3Xl++kE0BV
iHz0zkQsxUQoieIlwWDWI04kBCdlRPFTt5q5i+uHMtJa4r9OYPuJrHsw4Ij2dmpu
z+4oPSgJdlVLhQRiWjWsk7jNBij3qrIK3l7fG8Z1ZYEUJn/o0y1HCDKq883rKhxw
Hs2mjbsSSag8B0tLoMMYOTeH+LHUme35IHgY4oPrQWmLhTeUOuDQgJTjoMQl2sKB
DKC1wbwwsO0KMnymGXiavOYWx+U7kQNhF6Awv4YQMBHxG3iTudE/TYHB/4ZqjAsq
qEj2t8QnXMM3r5xq/RVhU3QncudGKV2fklOr039+MKAkbqFy0M2p4A3HSZbLuiyp
mpUk3Cgsz17NLhPsvOZehDRYeR+I7dz8CirK6GtlyZXawGog4Y0hWHyX++WKx6fk
HLF9MkH/M9BarYWN6/OQz6ju+1TBdJ+wPMZ0oHO3RvTlh8FgsN5KaEWUpU6+JAV8
pEjAewnwlBS7stsNHslGYbtfNiGPUFoKwHPC1lGd8TT9QIl+cYl51SE1lWLWkb7W
EBFQatzfo3gHOsUY41E8mptXcC7KOrEyOYJaPtmBofQQ4i77/H1pZuFyT6yl9RZR
ctC9P0kfufPSYYFtNN5jxVKx2eFITakWuY1bRRhHuKJtzBtGZAh6Csgn32dzX0ME
9lfeavbiRaMt6/iSuhhN3kQpnANufxFctl/+BNTqD9lFabljaCpi+OY6XOwjPuOL
o6qMfawOr7RyovN5EKvL8Vl6bo3saPxJxmqk1WA6WCoLiB9IuKT99mZhnf5q0d4U
TM0ekPM+TCp5b2neoMsUxyl48QLCX1a3mi8P8eTGwGSWSGkGDQVQpOOjsDxTZ4Hu
IVf/l6pCtafRk89/qXKJuESPTrCXf24jO1Usl3jMvyIXxs5uuDWioUqZmFxV066d
vO5TYd20BKNPtxJLcgqMwZm8bogFHmsMy4NBWICa+5zW5FWSX0Ep7uwu5JXLHzJh
Nv73jJiahTzLi/T7uimNT6VrQIP95Q8SUp1MB/pfWe4X/gRi6af79zp4ZcyckUZU
hoqRgG8BiNzS0dcxqKCEx+pG1+Fergw/D5GRa2gI6kIkS9JNJdiLYsYvwHKF+Zhh
KKVT+LgRvdedPilH2Y0SJxe6xcU7vi1z1ACHtXzWZo0akO757FK6+rJ3vaJvfdAB
VQ0wmxWWclrtpDVRrIq8DRhCwXk+pDA+faA/wENuvKkFkAezDOqzlG5hMfaF4evf
vYNM7Bj+lo2LOg6yTH9RPKpPsjkLpNKHh79bqx+RAhaETQZvxsa92E9fnSClbh4u
+cnOwjNxX1aA0gUqdtT4Hys6gFcrvcMBoCkP41kMkQX/6v4pP3utdbdUMEb5S0P5
D1BG2RiAgFkqjpKoJKFNH9OmfcBbIj8NlugHaLRknt0kqJXVBZHRJC4LrzzYOLOI
tI5YHj1ibYz3ZyWUy8YeqyR+wzkdM6aUD+Q5OkfzJn5jKHCn2hZuntCljM5EUvUl
ONVsAbOgeLq7ybAFcQ08CBt6ePaxC2jOXDQEvYqCbjIM2f/jr48yIivQG2DwgD2F
FXxLoINF0yCHy0wJMHnCviEagb+0xL9RGvyBlzRP0pvxmRf+ZNC/tpKKRw4+0rN9
HinY/pF28BVxEwQuPZLs5SHEvlH908BOJV8GaAQ+4JSZYKlIVYjL2pOoJga77nlk
YUTxNhQbSEYjRO8CPjEW4UZR1ELfX459hDx5vNZGdSw1U9FtUsw0ZfDi4BzNc+CT
GCFXv89RSu6bbTFOEEW8MNAlYCD9XA9GaKmma2MZGQ5nPZ0Ncnv+CBs1ePj9JsbM
92QOOt+7tzILeE/qXCai2OqgMR0JUKII4zqFmwwWvzl07oonWex/f7tRiZOFBDOF
IGge34DrRsOCfeei4yK7zA1bZuuGOphE5vl2Z555vZ9CEKGsgMCCdLXNTrLc0IiK
O2butKdlefpTFxgz6cdmfH573ULu5/PrsG4eKmIq70+it36LiKP9y/DSsJj0hpl6
6W48BvKxcD5Ru1G0b1iwUG1DUe7YhUR+6BTgSJu+HWGnI+Ha3hGmjERIaariZUu/
pa4DN4e86v3RVm7GV9Kr3sr8r3JaK50kuxe8kfhaPRkejzlXrdi6L8bLHrOUz4SG
0AhwIrIqgUZtOJXf7kl4R67AQWaGrkJUz4CetAozEH0EhtFgDI6wFxkpGp3CzTaN
RcQhJp0FFOoMjx2/qC3qeTyzLEohRlH184XOyO88CAyAibJXHPP+D3I0srH6mI4A
EZrlB8xHH9Ssq7a3TqInP1ymxWv61dC/xZP4UAN75E5wfPEcIDop5t+/bKkFcPd0
EhGX/4zhP7rFT1InlC9CpE+ZuATxGg2i2rxVJdenm6OD4NAbJNxr+IzDpl5XeQov
wnVtn8qVGYsPbmOKANt7MS90qng/S//aRa3i/kmB0re9u2C5vd3SgmZ1xceBIqPF
z5uHVPSBbdhxpy/nF+mHXcFgaiffuutOAL0TAE1pl+rMKjyKI3ynbClL0GuOFXWb
Sk3v7z0DbCRJ087o5urPyyLib+L/cHBNKc8ARTlAwIrEI//qmdbgsa2zALopxckj
oSMuzt4gPp11IfpbDo4RM7WbH1PJo8ScpABfL9LbWjOiDjmGZ2Ed1rqpy0Cim8to
LwejDVozjJejVraMARidRqzPhGPJ8poJpMQQ0sUeW6Os7Bxk75LqZJC47dr0T5wf
pLEK3yd8XbA/MFNffZ2cqcNW1dfc2CWjmdFho3t8Z2Sm/OJTwvC3BWRVaAiS4KZ5
O6xaCUuOUDWzp7JttD4Zs3QI9CbQrZCbBwJFe/MBV/U9Wnw2LBpZBmpG0sje6oGp
cCv/dPrujCz7tjJl/ahwweov09anVgLdc3Aj+DA5mKlGrpSTUjzctyWmatPvX91d
QrUAaWr20xTvZG4LHcmyMxy+mZTz5UoUpvv8vID5b/FU5gAGlgMPUrlRO6TuHk8n
ChzsZw5QurVbn9m9zF4MuQNl7XUa9cn3rmdvf+F0Vfa38VhJAmRTG1clQaeBPbH4
XzWDKHWTHUWlLA5Uu46hFp9jCdSod2B11ujSwo1drQmUD56OtXnf6PNfrExPVJf1
vyn7YKgpvZHqr8gqsFWdyvhUR7NJWb4c0a8iHrIJB3vjX+qfQAjnrv24CHe44PLN
HzXD9sVKoJ3kFlFZe+nq7tJQKcqIN2TAIu0q4ewZLVvrH4pFKUMrGSaP7KInr8VS
E5Pyf0SN5gympUEpRfx4xqc2t4JFV2ByMnL/1JtKADV01eYXTrskQ5Z1UODurlb6
N1uIx/DX9pKQd9mYlsZ5r/K7pfJndQZkiPvXENt7cLNG0KirG1auX/zyMT4sodPA
HS0FA1feppboJ/UBuJbpEufKaTlQmevwNvrNeaDD2Re6bnQyP96M27ILgqyalUPP
FiIa8KXE6UAI4jcb6HgARn/MEEPffm5R8W/9myj80fhei9wK5GKKqOrWWgKbX2sY
EBq5w1mnjxYR/6RkJA9ZdkFxkbzaJTXdOmivA16pbhCAM9JYVYqTyEBSGXGj32G/
0aoR276FLPrLFC3PEOOFvxnEDhsm5fx1KTtN08DcRMZgbfY6NAAgPvf8rX6fMevV
R53LCJzX9O0wVx0RG2GARMrPda5+8x/mLLsCELVDiONBCeGERT8If75wevKxo3YA
8bnwF09/c5OH0Q0RcRWlPpNynMrVGutMRM4DLRY2IxfMSYRPiSe89+k2tHuiDtU5
LN/NsePkmHNBHNupevFKc1o7wEQCH+1/3S91aR9nGLGA0hiquAsW7z38Eqa3jnM8
EYM3cglw+TIYzHVJAvsboj9Ek2JazQ8XvTEwZKLc/m7UR+cbnDHKVUadKXKNvnyb
iz23CrgxY3X+X6lJkRVugpyzrb2jlaVyGYIkI7iQSc7b2zLJ189LF/HjlljtWiuC
7XD9fjk/dGtjMsulJEgxlHMHvBbxSOzCx+b9284bBVCYLdZQxvp+O6eZf6PeCDFo
VT63D8wnWaSUVyQaVeRVvLLaj1ksG7g6GCMr7lHmrV+62Lkfip6x7dtEnTDPaxqZ
oazWbGY3Bt16xQqrnNKEziC1/7UOOKOVVNlSy7ckVdZyOqmRjIgVeI5TW45QoUEZ
QaEbBjiooqgJuDMuJWS0BH8ezNKk52Es0zQnk2pMRAWWAhPQ/n7q5Z+Z2UGCdX3G
zIFrgDfaTTcweUkZh4Bl362svHoZrDC2o9wjMI9icxWXpZxTNzCu9errCLytm//v
GQaU7D1VuT/CAd/MQVp5YookPc5aYV8tN9BNzjjMDZ8CqiZWhs8EzYBScy/RiAa3
i0hkWF4OzCpKRSkTy85uUOrPG9LngnJcz50WnUkCv5uKElzyExoc1PMFTRy4vM3n
550YQiaKwPkcFx85dousG4qLV9LLZD9wNAI91/BAebJd8ZHIYHGyyUauKC5Rjmbx
HPxJYdTjlzGNwKUBU1QsQ0r1DBn0H71S2lZWO/CnZQi/ogxnNnUx7DAUvSv6Kw1r
coqxMi99iAaRkRPdL4Fds+UX3O08y4lAJyhzKCRWaDdP3KZtLb7mBUThff7LZW+s
rKEsLAuL5XgQIjRot8HItItgJ5MHhja11wnjosr3fXyxGUKVT9zg9MbZtEOAfhFQ
dfEz+FLyf/ZNO/ytotRoncnWFIymF5fJ42M/Mh+G9o0flVo1RmmQQ2keubrBMYvD
2EL3Tz57Tc6d8iu5OnSd37B6XfhisyFlCO26o0rbz69vCn0L+IlF82KcB1aazVmr
7/8qkNM7GrfoJwrCYWU2L8kz/D8Y1JyHMwi1fMM/o1fZ3DmW5gT+MDR2z35RmwA3
L0tL6YWdwoCduWRxV3N4Vtxgr4NZ5qebkgo7acH/CKWJdCp7//jF/b4XKF5VEifH
g9CxDkHiL3PJVc6qzDrXcdAYghG5l2ucpbqQV4SvUgxhq2NJuxmc79jBlWCOKcUK
95GdfmeUwXaPivoFHvQeRoX87xv/FwcuPqhYYOa2fa/9U9WiwukvutLqo0k32/dr
riRRg4zQGoC4aXWxdF0eOra7TbLioiRRvg3kxaRrnlD3jdAU0z1t0SILfO9F2DJi
1mK2gsVA/IO+nsfcqNuWaWzX9Z2cGXYyvHErviXN19tLyCH9GtYS6wkry9QsP8QG
wekj2cmaVMSq+ytrvt2fDziy/Q+8XitXMxB8eJgoggJoHWPeG2TuOtxDF6dPxCLn
bFzexoONCoznG6js7m41iuXirZRoqdGbb69rz75Ccd8KGfxaiSfV94CdGM1vPe2u
7bWGXh94K8eMjQ3GWNvvNHJAoHbVjCbR8TmJjtfIsKtrn+mgExZuaaKO42p/uDtG
8E8uh1HQ0RyaKdv0ddk+O6PNKBY/C8H8hns5dkDg5vhSCkbLyPW9bbArag5fUnMw
nV3G5qhtf2qjARlWcFAHcYyTN0bjahw3utSHEFoS6G7PgdZ0D6yOSG1olQCHWrVZ
jxwgg3Hudn3P0PTd1s+MXajVPRzUaeSKTmXjVVcMRpKdrszmZSJ2bM7h/j//TEwO
pxwCKeORpo99Hi38UQxL6OGla/tjavnBs0URz5pcLcdxtRILl/PUc+rFYlCt04wf
BB7FDflDv833tvj5lww6XdS89ay9cgkZdzi8TV5P4t/qxR51xvhXVBddibuhT1UA
ucjaEn7zFz0VVI+qQo011BBdYS3G1Q9c2IFWzqCOGct2X+wKI19MM9LIISKTH1oy
eKYY4cR0qFqkc7BhhbDS0I2PfW7Ap98ysWcngsg+gt1uNd5Ac2MUDW3LZUyTv/tX
UrGLxgz+mWur/YyzJ+ZilqkIRslP1auLv5JO5CSKmcrnzTLNAPEreixc1PWhNaey
YD8Soogf3/vWXOm9V5KN1fcz4Q5lfWyDqtD/iQTF9nPWHwHCint9jfsyJBNaGCvT
FNVwQ0wjmZq+gL2zFtnWRBFNXMX5rOIhKGRBp/yL5x8UimyqA/Qc3proX8egHxH6
rGQmWKxI5FOPcWTuseao3DnEq6ME64x7QwhYHv+nBcas69e7sA/GrIsxoPvdsURM
hBqkiXAeiKgXjcT77CmGJJy1th1Y9/G7grBei2mpHgD1Gqu+/ANpJnGFKoIJmVsx
/0OQ2awabCKAKQcCPS+xlLJFMiQaazvM9/GzuzXCATdhh1l9tsuew5Ssji9VYmCa
OvyUJR5mpmyv3HYP++/rtf8DfZOuAIdywyhytkkROYupErvrtfQR4ZXcsI1ATf/o
e19UsdjT6ZOy1o6Gb4cpcfaoUz6LelnTpaQZ1K6GO2u0W0QybeZFsca0JzdCM2QN
T5mmlCrvrICDJFSId5HsX7bfBbwYgcq8brPtzKxS1/wceBJ3zrXoSvXCVe3JvNHx
QkUIg7nJ0jcTCi8eXsNv3ra83RHjilaAsx+7Prpdsm9aVH9cF9/neNFqFGMjGmnL
6m6E2mAUXOatz2YycrNvG4fYcfOewDKR9KPMSQ+yzDZ1hkvEkNT8Psx+NHENpcG3
H7L+0boFEi0heiNnofWGt3esRwx3HZavgWPoTSRCI8qxWA5P3JHFHVzf9sJ5jf4S
CIXNxrJFhkQlavpqQ9h4iiQuZGwpUbqc2t03jDehP8qbru3WSOHJyXF0WOJ+dWMf
y2yqRU2dFdPdjSoIxRjOp9KdDAcvfWmQyJo3d1LElWGIwVnjZsP4vR/OLQrGRsX4
IHrPQ0sMmsF0iFnzCYdmFhKZq8Ny29K00GdbtHJ/Pa3C3ri8RZQBy4KCoXiDfuEC
SjpUFW6gB8a//OOo8C4HTVBsdmkzEmE6bEO+lz6qIurGkTf+y1oSPwWntgVc0nJz
jdY9Lc3yztXIVKTG+G0PtUqff/+BIH3HnIuyNmH0yvzc+vN+NDlWlG52+oFJ2HoG
Na/1hfj8v+PbYxE3q0QwD7PqCI9fFXMq/tlniHdyqeVx02MFklaDO+0d0w+9SI5E
twiMv31YcBQ+PDirUH14Qqc9ZbItW6hxLAKbJPSVGxPXZrNhlU/ioUyjdGU0WeAy
Hb4OML2KUe6t+c7fmBr/TCHJwLIgRffm3L2z7NLN/hkGxe7CnzlLWwbeINUAO8dc
PSQXSotWg+9QXKQdIzvUa4OqF6suLbeAt0O+nQZQNg9L6ExPhdKRlE5l0lkq1n60
ZohG4ATpaumIrI5BeXriTHG5r24DZbvFgLYQV+h1dwCWmR/jUNwIxLB9LUwOJe8k
UpTO9CLOIINWRpSEouhBkhvrMIZ37C2F8nLIsB57F321RBC/Rw9SJUzXtyBfZTwu
UM9Nj7Vq4p6rq5n/GCueZ49y5v3QNntpKM8+ql1iqJpnAJg/4j2oC3UvlHU5ZqhB
0sTj0vlEmpC9/h1re5mXlhfFST2ci19g4a+KSNsHAbh6PfZomAKOihFWvBMTOk5w
+Uez7OB7fMOHohv/o2KcLxndcScOl1oNQnmRD3ex+gQX1fGcduBLqeDVgNFQSwRi
EWIB5QcNXnI6vRiqIlSiJU51gaY7AZsUGOtNjdivO1t4wyl4NlWHz6cN6+KLK372
arMqu41yx46nGrKwTtW45yLnp7cJ4np87uQrUFX78DgzS6QfLWx7oFtqZKUV86s2
YKS9hhnrTDdrv68Sh+qAba5REy9mqAStb8LmqLOEezoeAj8GjZHMZEnTgCyvrHVN
x3ik803FSA6OGXyp5K3T4eAxrKSlmfW/iCjlm7BCK7lBZDHGPDL1kuyOenLVG4H9
JoeDmHkY/+khpcsMiRNsMdxzwowdl6pHeNa2GH7xyvkC59KxTm4hMrbgckXQXevW
UknjplkaH3fVUAczaZ4bhXlBxtYeySFX+tla4gJmPjxMQD4rE69YlfrrWHxkBEh8
2TfakEb+pvKn6qRKx4p4f5suBLJXf8jsiVaEO/H+mCbQVEd2JzpwVUDZEnFYCZCA
eO6OLe0S3AEcIvX89UldQ/cq46KABt1aeWbYGxHg9v8uigRmYEy2Qr2nLG0MpDpo
Gv9PZg8uy4oJknkfSPM+f9QQL+bWQOuEeV8BY1+ZojsywgmqgvkUc2QlPoj40PLF
XYN9/78otBBbaQs/Kv0tz4g6hQz9pYS21tggq8+cAaDUkwPQXR17R2WphWisA3X3
Y2bupMm35ozOMbAnOkRYF9+k8r/U6eLYLtv3J8j7ETFKcRKAaIj6qbwYc9gF+9pC
Bx/RPJoRIOQaYDIds31mZLMaT0f8srzHpWEfGBWNhW8WSSQEHGkr/TzlC5/rIVPX
dM+0YAj82N1dgwMRLjCp0/brQqleesVN/9luy1rgN9redqIrLF9CjpfanczI6ZXh
JJag2py3mWBXOU3D2wJEpzR+Wc/M/0fCa9jWXDKO6Vw8/G/aG90sZhyJqSad+VXP
K8J2yJNAQEqKGDqAgVgugVmm4/k/QFdXXzpLBfp22iBWeaSLRk2F6BeSQBaRWVeo
ZxKo8bSSv2BYTf7+KiKlemKmo/jHwDZfjlUU/rXL3gh9jaNQ//eiuwAeF3LjKkTN
XqqElCIpO7pDZxLjUgmJKDdSSEFsFaNLoNeAIGXZqOJR6P6MsE38lsAykRhuCQUv
SXCtuN3seSo5an3zXTCPNWkmgqMJ70epeAzU/23jQxN6Ute9buBWgGlkGWwKwgtC
+1g8AYCIBPSUsoovaMyl+UitOX6BGdX4gdI2yTpHl4HOSk/4Sbs5SCxI0MBIcq6w
0SZvcNWtBzRbOfvcntjK2obrWf5utElhyoN90pteHroCdhdDJKFVOt+Cgfs2wStP
Lflk9iShBra+9KZeYBGlFf7ZXGu9ub41sPQiFHkZoYKevp77vrU9fsXgtrRH9zib
AtfZytrsInwQMzBctnj0g915bwgb+c5iP1J85Wr/7O0efzBjMjS4ESuSGiJH0poS
a6xUsbN/SW8qVd6kwhtGpnjdAZzCTZvDOpNln+VyKdTwwPwrzPdawNfNMmZOy3HA
OrPbLNE+lWHh4SWzfWoD4XghTCsusgJDAv7HFr1NcVEmrLX8I8qEREylPxg7uW+5
yxrmfuHRe9/CAHHD56pghrzGuFV+JxUxJmc80Wkpc9xNWgmBiM0qQqwKaI7m8a6m
BSR0HSKpRtIByZzOFgHTA0r6Bpr84hyrt4pgQ88/GzNZSGPXkuHgv7FbSluFffFP
f2m5Ojlox86Jo8HP4JqBwnoZPqhPWbsoFqhcBhZGuE6SBTsH7djcQpSKAKWJcnwS
mlGdHTgQW7Hmfx4JQOTWD386Dv1ktQ6712a3kg6MkvhRhMF6GDB5N6HBC9MWiA9G
efJvFVBgLOGBX1fLBHKUXs2qSFnz+oiCIqsW4tb1ZLdsnU87xHUAa1yuL4WE7d4i
oU+fXxWfMDNt/brSPJ6T+zGMtEo7yE5gcEaCNC0U0NGkJqLw8CfaaHD7j0ub7kld
omit6f+BIB3Inpyr6eXMW1+VaPzAKCc1n8NNWzGR1S8tor2PMXvk2U5Pk8GIkJxf
kA1DsNa18vYcoMjaaw93HYaMdUPyQSuLJohSMrmbzY1At/NdYAcpXyhZMlOjEOSO
EpmWp4FioaaIR8LEv0NzHzYmbwzzMJ0bQeARII8v4rrOhAJAMHyR3ObkVxWxE7JR
PksfP8j8A9drp551voM8qqOJv4O6i1EETo7+JHOJUn1LifNeuiJA5GIntkamzbWE
ZH56XF2vM2t7zL2L3wPeTYCqsK+YYuLdwNrThYCJjuo5aCzITJ4dgUI+FeVOyRhR
TlfwKYP//Xeyl+Lw0Owh6MDgBua+B1WLUv4xfzjYqKzD9kQ/G4Tx5w8lOcSMzehS
Te/rQXmhrdBPflDA2zNuW8CLD0IjS6LEGVnfHR7Ang8MMRC/D0pTWzjASSx4RPx8
i9FUjg0nU5NFgaMoIpYM8iCGXc3zPO7myTKO7yNZ3bWdMKIQJlaEB/OyERro1i79
vZ48zTN56eN4GkFvegM9VgR1w0KUjLjwQb2d17TDezQ+QsXBOrGswpjWLS5pshGA
H3Iyeg80/EsmH3FijXSMs4hLeJcIeAjrpHrrWr0z5zDHZmoYBvnLahz99oqgrn84
SVQtK2Mdd9ImsKsBIeLEMUr1F2qcpZTk8y4+uFXltvayZAkoYQIdhTm1MKlPmXNQ
BapQWEo6cJ+GWr313iDrPQYVVOzWx4nXgdKQ+3FeMN8FCeCqHur2HyVUvsC1g88x
/KjaqPXUdgfOWkcsIZdTbOk/BGxn71AN08ySi8O8l9lGWnVZduMKmhiBlTwkb8hQ
5gEwZMsCd0OedaTUzlQS6MCSl/iXdnst+kGzCvqUPZyKpa4LuvHsmovxd92Ezvpm
SsHLSpavS5N/eFvVHeMuIqTxOPhz0/YIGY7TIxTFIQVv0Hz0dGSMrd2vQcgg0zzs
ugCIKnSuOF/mq1nd+YJwi+LJb2/tHtCD9albjlEz3SpR4tnUkuhnXtPjO6YZFwuF
ieZK3wx52xt1TpcYRueBril+h7vKtCEcznLrnuCqo5XzURtHS146Ag2N7NGFh2oe
oVRPzSdPMIfYfFMAmFYR5KhOJUlxyZv9Ih/lb8N9co+46FnxJOzn2r/rP5LtiN0L
uiZxleVINlFCp4sC4XzxImsrL3aT0goMA2zYHjY8WEeUgsNc1FN0cvYTGHcHVl0c
dNQUgJNGyG/TF16eHZOeqxJoQzMrXeHp58pbbMOkBql4UNEMDi7Stl1XMn2Ywkgd
q/ZvcDTjJi2TDLVOG6/hxLMPok+8GNLAWOJO3bVEC1HV2qZkIpOadb1fTMW9t3P2
3UL7UCvuTvJPyCSaM2cweIynyGg+O5hyQCLN4TxZGawNIx9yoo3h7Nx5aUHD0P4h
Ync3dqiATAr+ZHQkyXwpzI0w8y52ZIolCKh3VBa/zuLbfaFVW/vZNiVOhsvYISZV
PswPBN/lm/1vSZGYLZIWljPlngzDLUkKCm/w4a5W5a241vnOuBxv9DKkdFeOiQoT
7b/PBo31oQxHTOaHoRV7Ag2X22n+0Sa8To+1veBTGQXKoYTgiZUKGFseuh9afDqp
3Fdi7gpQZOKxdlqhhCtaxJLXRmsLqlcU2EyXXMv7IVi9DxZDoAeepVDuyFB1JSaP
umBVxthZRqxFxg2ann6rN71/wfl7KugVbO/KYhM3+gz9d3OqD03g2q3V1Vhy1Hb6
cCSne5RniTANSoZU4QeBB1RvjB9Y7yc9iNssLTAcQ2yiYr4RvTAXG0qqc9VYN610
/Jx+ODg0vtgayXFzObuMRFxtcgnF/57wkg4i21vVUO+LSMZYIINAY24LJRb1JjsA
XjhwucwIbAH3cIaGtVrTjv8RAjbQGCXjXP7AAdESToktRH7iLv5cCvYiFI5i9xB+
YzuFOMAGlRyEPLbRKk12A0T/oJMrhPXKCNsL3XPj2tgK8MemDz4SqlEKRfTx2hyJ
HtCNMXafmh+ikesne3u4S/UgjcxorKMkngSH2RJ4p1qLtzzbVQKlvuqN704ELN0n
GmAMdItItAWtiUk9AisRJLC3FVOzjDV8DvP5pM4ZfyPWp+U1tDXTcswUfzvHc0Vr
CSdzIrB2rhe6fbU8on6RCBetRy+6eS7jaxDdpU6vQTfXmMpelcQNsUNxkYeChh/z
5Jat+r1MTNxpf8rzLXWlQyLC1PIh68pETaDBQbUpZ0tkXZH73M+SpF8w8SaQIhTJ
t46qmhezxqwstFVg3ZyzKLTSdPsbcYpfC6MluAEOHuMB2lELOXTU1x/TVbvlROcu
LobD8ceHGb+we39VRqRmtBnZs92wNl9ek/5lHpDWtBNlMVOg46YOLpv+tFcJa/Ck
3L/lvT+Rl5HMwyAY4W0fd6Xtq8HCLuzr+u2Ueaf8XnqtWOh9BB89jaJIX+1yugT+
CM/vUH2Wo6lwiJv9+cgvz/IN/NRwM0v0LIT/JnNc53FJ6rqD1fOZ9E8+gFvXAakQ
hzYZ3sbGZ7Mtwxda9/1ww3E8ey9Hx3oKY64A4lygXVaXDJBSnEBu2w4sNIcbE+ni
NN5RHcHaaL34o1IxoZSN5M9pSI4jEbxUvS2Dc3y/SDtgfH4cfhl64AO6DWKYHYkw
yEpPZTF+bCYElcKxHkzVkfXslzcSjQs/+vIe74uHQpv51HS3zwCLWfGM7i1kAHLD
p8Ix5/jRRjz/6a3fzFqDbfXpAgXEVOBIczlZxx9Ahyx9LY/pesUIrJvKQ6ah3gJU
UU/gTz5GG/t76J+KdnYuCIZEl1j40URwtAaNFBgbS/9nnaupHTAq2Dtk1oi6JBMS
OPYEcNTECR/CrYwmLGR5ToF8aBuoabhFBVFYBQbnAQD64iW0K+bd214gUPeIB8Oc
PkUjRow9NNqQvK8CnFF3rm3lheR2h0U2Pib4eQDzGis+7B1Ghl69IyoO6U1a7/XC
UeNzvnXSCT1hRQ16HBCZomyFrP4JfndQDTFADpAFFpMkMcXYlKVFneN33vrkuHEC
X/AvBDS2YAvi1HlmunrcUqO1Adl97YiJ/R+R4RXxEtBCSmcNNbbNd4sUzuA3M5G+
fRuBugq2YORsxDkMxtZA/k043/YzD6nmkQE+baRWmw48f5U7N3WzBCmBbxAcfldZ
a+j9L88YuVD71ZSY8lBXNofNgGHkQiTSnCRBI7MZi/yNcpqXndyqL8RW8TrhMDO3
zExoVKXPQ+2Li6yNF6uGYuR/+Fx3vj0c+7CdBgnv7F0UEoiW0wSZml7SJBxiIzUr
sE0hbG1j6qlxUbiCSJMgooq3BZvOwJbt/VgqLwG/dm/mfhmqZWZAdH1v1d1fOhww
t1YMDgxP9h2krmc1WSqk4+uQDlJBvtwgFS+eZ5ZYLDB286KxkR4USIOtV9F0HvJO
c2Iu+aSKpDqc16vdHeFSBGPLW6HHNiZJTrIJOPY8dv+P9rq7PTmcFvp+vvhL/bZz
fkRog/BL9CkIIIcTpHNMI0fM+6Bwye24john3lCj0h1eoK9KNvH9DAnS6dEocAMl
TGZvdr6EP+d0Ov8qnvHsiLXXqB3pIIjafk4AAwAcVvVNFYwlIBrxpXO1GVdgFTr1
f2uZu4Z7haxkP15/OwOjZuIE8gkUVDwPupZ/0xIkmlR8iShVUoo6r4xaK8YNvtWt
5MU3uM8bfiUUtQaSUvNcD8gOK8UiLdaQdBQjiHPziBrIJGjoaxYWafbb5efZAGkm
Bro+dKCtxPtW7QxaTxr+rnVK+Y1MjmUPRsNkUmKybSfLvPam+gIiZJTKIvQmgzma
IjD1wQwerVDceyM8YD22LtWbsrzpCpYMH3G3FbiUv8wzFw+FpPCKNJ5oSXAYTmik
0TUjbN0SvxBDNC0zYapMcxMkh9q8As43kvK+ox9HFTEH3yMQpYTjdFX+Md0gxqPy
3pzdBOoAYVYHCVgTLNLGtJJy7CXDB+QmdKq6iXn1coITic6c0G01M5tzZ1UBp3Ac
ENDx08M3OO6iz6dTdPuBXIzeEgw6dYhg6gW55st3umdmW+wGQ3R+SbUe4E6ygUgs
H308si2bR57v9UDNAqAHF9i3bwyQOF8k5Tmf2UZIKkqLtMz43xcaYvfmoFvklL9Z
UkFoIleDNhTPHXI6Kl3dBVCZ20W1rsrl6Yq+BeZc5Z/+ofUZseIMhpDC/x6Lioue
tBKW3Evr4sf4r9iBovZz+FFFyBqxtE5PC2l5DxA4efuhMKpaEP+hF3zI1DfSedY7
MiPEwIxc6YAxsZKnieOpW4HtbnyZZNFfUnkUPoaNagOyQwreVfrAj4UW7gq5naDL
w185lD34y0zyKCOILbYfZj9qWVRXdTyrTXDDgVBqKTEpuV6CssHTOxLxFJi6uyNe
zn7XLf6qtyMj33iL1ItT9WjRfxPqqaevEdU5RcISYf6gvS7OQpBuoZsXhkGudvRG
epHHr3AV6S9cukitlpsA/8cbBUh7C4SGpgxapCIttSftR8ZhxnE3Zc2D8DqUg2d3
jpU1pUWKFwQTxgTv6MBTNHt77ExzjCD89x9TnjoJqzQv75M3cSTQQq5beVnd4vjw
`protect END_PROTECTED
