`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZRPcb9bhQI8b8ERgLpKJZr3dMck9nPLT8+KxamqMU7qytmlvt8uq1msWNJ7Ni84Z
OxkjSVudVenfJ1VPxEsz9Y/0ThnGMIkM34i7KlHrrHtVEoDydofVvmxYaikrT78Z
aTUx13nG0T9h0ndTRprvMvdsfyetqrthfKmC07vK7Cotc6ENn727xGr+pZDQK9bY
bZ2QOk5H9to7SEAEXwKK3YTAdE3TxjocwRcqg9EaIfZuetcc0XupjpkLsnEY1DhZ
ZgxqkQXoHCQlKMgKb5SEwmVDNQcqsxXwu+RxN+Vut6Ydympj5jGHzf5ghyYXN4GC
pxV+DAO/7lfzpbJzEyAFGuALY86QzEvL2/F+8SjuwooWqCWuUeJE89cVb60iHshI
Uo6e81a9PSceOzaQ2fVUnMlTcUW+2gKepyRjacoZvok=
`protect END_PROTECTED
