`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dHq22haVhmY5HuLRHff/OGwOGZd9xnxy/fnC1FtQLoJJFntkrR75BUNwC6gotXQ1
144X+xeZ0nD2ci44zYmukjIRuZa/3M1zcFQOmseibztqJR+gyHoZ6am95bcamZ5K
/GdgBzfmHMs5ginTyFfIKTcNG34dLYvbiAGZYzGrm6N9+fT3ivIW27flRdaHvZLn
/xdhq/SMYS1r8luOmGzRJpv9bDPxTwamQuOW1UhchrJiKilAXLijb6BMi8p2ZlKu
P9iGd/lIlMDMbQBfn/iBOLxGqPutEuDgpOIWheGKSgUIHBqG8x42mVRhLbzMr1uR
6c38SbbOEtSuJRVOW906Jzm/t++w7nqU86q5d+OGQ9PjvuVSFLunFK/6SUWOqLDr
`protect END_PROTECTED
