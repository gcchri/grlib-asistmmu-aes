`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iDqRmj+JByTI1IbXudSSiNPwQNMmcmcK2qIeFPE1moJiELa2U8YLSpRfz4mGzpuT
GcvqwAB+ebvqjxU2+imbXczXsmwwTr7MgrEwoOnwl3pw8NuLfNeJCqkvXhye2b/u
DTJXNAG6PHq5jR/iAhT0qGTb9hR0xvZTOvFEFGPqr6W8vauo/tpzz6GIAeb3GvHQ
77b0LzJOCoKjCCSmZ0FJMyFX9EQEH7Aqq6QRt/cSXuU9GCIp7GDWnWIxrkul279p
re5gk2c0NUhKw8xYJixl8zo1A8Duu4M8CZ8TeGqK1zmHMZJn86ii+XXsKrSI0gQx
iu++z3EUjKizZ/+vVz9uMsOZzwGdgNi1v4E1GzqWntmxqcozRDvhJWo5wTfEjRIL
h+Xqc/uzGDLEBOf04DC3ChDlZdGihef+HRse7qwY/QGNdUW1WEmcYNRkuheaeUBr
TljVVnGLoiDS8EWl83uDGNQxDKeuUey7C0pWVOX4vs5mz9Zks8TgagySDW6UBcCO
pLUffJzCGjkqnv+nS6KG1alhOvGzYkSdUSundiOU7vkOP1MXhAGtc13NNoMvCsrz
9P4/TXrF6WPnteMBBzqpfa6m164/Nv6tq76IinrBz70vBm8oEqgoiLEF8Iyv4tjE
Qq+aVcMqJ1gT1U+QTAMhT00X893ddgis8y1+YxkIYUz37Ag0znmxsLaf5y71T8p7
/suc0CrGoz1AvJvThZDJLriR/aRpI7C+BWHGyV8tKiOuySTBrllE9noHOvxhSR+F
CqAEFgOSUHiLsvYoSU/7I3k+FmyxXAiInr7Y8GrFeWnDLF0es1tk3yPchMe1Kp/o
bhg5It/1GgNhqTiMNl6Iu26SvlZoksPKe6Kev5qa5PBtYO6acJzmc40+1xGAynrz
`protect END_PROTECTED
