`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eLh21du1rc/b7Qfb2QVEoYNJJTtQcTgLLfpqwPOXG5V9SaR1YMwCJ4sSq5YC9QjV
pEQq/8Qz9y/CSDeBaj+WLBCvh5Ywn8L4mU4KmPn8Rcd2i87VrcR9tt7NEDp1JKgQ
O9CfhMBx/xnsjh0WeNCHfCaezLIMAn+RrTDlvlCB9HobDmQkwg3lWGx6+k+BESRt
I1eMdFaThzO4PhWm9LK97lo7KFPdcvSpwK9+8+zMrSUG5H2/K3vvMaHYk3+MHsZV
gvM9Bu+c7OlIxguSRgra18HBXPQCnWjLQRrbiTnKuvMPVJSpK+0AAggtrDA+BLIH
SHGRWK6SkexBJpitAGSzR4F5a28PI1i0FJ/5QBViX9XK/Qa6Ns+0DLuEnrkdRV6V
be/5y6G4ybHTRIhleS/0DU6ZRZG5wlwBb/joj7k0726p3quVkIMI4tvLNkrER7BE
zprIc/fOky9DG6OVWOBaVvdv8YAyOgovDWHzVjMvAgg=
`protect END_PROTECTED
