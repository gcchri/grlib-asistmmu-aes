`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8rcxGMq9MkYHqIhVSXc1DKHZu5WaDlBBRQsYcc0BkNhLyPIQVbRaFCog6ExHKIMW
5mMLeAXeMuYYJbQn6+qqLqKCbJVagDDToXGtNAToMeygJC1eVLEiJI35oAHvGxnL
Yplf0goSYSQgQm1gfnFEx6vcc2ZDLPe/kVnk70oT/FWx6wd4EY+Nu8uGG/eBjWDD
/uMdfYy4DxSTGJUz9oesKMCFnYmIpf08/aYYQJZi2rz5AderehM2zF2dPmUlsXZ+
6ebiUDQQrpspPpVZSmqn0XI+iwYFHBkecfbUZE8poBTU35FCIxSB8T9w5MRxq2sK
`protect END_PROTECTED
