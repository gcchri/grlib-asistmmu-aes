`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fRJVK+KC3kzUCD0mopGxfYiYdoNni9E6to2OWHJiqjKLRs3b1Jl/Aa7Mk6YTRhUY
o3Vt/6N6/t+POzrY2REnazsqOsiEBWVyOJOHGwUxNpc+2bISLLY2ymRLiJJld6J7
9fcse7l7baBvQvvAeSewj5+l53tt6EerlT2zYtXrpz70zgFeu7u3U/amUfONZMTA
36ea4NErJu7iABGj6eTzRYKlIJgrhiZ55lnrYQZOXBH50KCf1PvXCMExnRhSeGUy
i9ZgJS2N3qGknRZAmyOyuArXP5Gq0HdpEgkXlxzUtthJn157ryRBBuHPA1T9J3OX
YT+9KQzXj1SLe757b+1D9E43qGtDfbA2EpIDaA7DQ+DpzRjL2RN2AkYsUAg3E58E
6tC/xGPRQKCOKUaZ67pPJ0cG/fqjwNs9ekwlPAOQ0/9mZvCbU86PLq6jEyIZHB4r
VwQHZrMuYRvUTAj5S1v8NpLYgFMU5OMTtsuSbsX0XH3b1FrpZWTaDhEnNGjHgy4v
fPyzHC8hFLiJnca42VwZzwfcUT70MSyOegXBciFoYgtr57V/h20AQ2/SkRsiVn92
yyloqvIxBOdziBsmWApVR8ojqvWY/NiKsrdcXGmxSmueokTbEEYFF4I6/StAVLib
2UK6nJjGrGflPzrVlSZmt1ll6gWyt9vMObpLUsfGgbugfuA8eDUIwej17b1bhRCW
qoEmV2xufOFY9iLaukfH3P1r/isgsxJOAN9K1MIUjzDe8XtVlw99mAS/pTdJtuao
Bovgvg6J7ZQLoa1CJQHMl4nHPpOkE2YsFRGDznqdN0MwQ1juV9YfhXHs36vfA+Z4
CiTTWDLkufwjK7Enxud4BvxZT8fHcE47kqKI84pUVzPEeidYUHD/qKImiZNgJKXy
xEdQhR5muycSsniSCZ/KoPIgd+3yw9rpVmfnOHXb/rZGBWa+w3+B1SK/pIzZ/0dH
sZN3jfKw27lqS3f+YUcj2fCrzQIy7VLAIAJFJ81+mcWQoEYLrx4U4hIgMYDuFN7v
4aBZfl6vAkUh/V3kuVI1/Yv6N0p60cxfyDdHOqBPTCPBKEXdHhji0aKj/LadQc42
G9KuPOfNMq/2olBPmYjiheK0P/xMD5skgyILa0MWWzZdSjbEo/Q7Gs5u0PWuWfGH
J8fisUlFdpd4wlW1rILUCFJ4zcVQSctIVt4r1zC4la9FgtKBKChHkbgmiFqnNvpl
QsDcDXBMgTSOokv3hcNDZAx24F10W1BJZzCe4zjLS6MigNLv1F1QlHIUhnNpCM9T
Ln2XQq7sPjaGUjUZvWdMOuxlvCN85MYKVJz+u3AAP5pLi+mNJG43Cuy38ghB56gj
5+5gIFMghNyCWY1him2FQtIOFjRcC+Bd8P4gjbIV2fjo+ip4UOW7ylTlq9wdu5oL
g2KPdo9ER82qUAeFNTeKNTZ9nLBdQXYNJLtSS8m4TTqszOoDPXhYIFQHPubE9xzg
tOAHiA5CSCct6wSx4kbdmRmCQA1mnE82aOkIb3wgBs1+jLiK2Q8MxtFYfXVB/0HF
3mUWOrzMsuwdLxZXOD2+hlsh0BQr3+ayj7Ymgp0D91b/sYD19oBldw6RfGywud8m
8W0I8tybp2o72qMNlqVVw7ilOmrzfF4VpffLJl/VvJ3BAMdEixaWUPRxNVt7eZrD
8vQACD9RWtjuqXkhKcjCemzf8ntoNMkmrJwyr1V5B1ZZHkfgl/aWAhZp1BDWuWWX
swKBrDZGlbHKOozp65ljZ0IDEAQ36I8JGko/MU+uyeE4hME6GCfmg7iQdKW+Eqa4
zmB85bKTp4q/+EVhW4/xGtNREhaNPGNINSB72EWbSbB0dKfwZzdfb6Klc4DpZwE1
bH8dNIjfqUz+xL/hu3km04AjmHGTzXeDC1zFpuWpUi27q72pK6QWaOma2iIG4Lir
dNBOdbljwMpEvUbUiNPkoC5XW2+6cXnvcTyEUQ89HPaNISvJChs8fE2oyBXCpfJB
+UE2rZhRASJJP2f4Fly5ham114Z3Xe95SMFaxJ1dRLEQYy2+PU6r+M/q5wRYCeZo
nU3NGHkIU+99EgXif4oxcQDR4WPmBWjjgyTREDgVig7UX5fa2JNqcDSt4+dOdQ+v
8gh6zjF5FFSN9oGfqBsMiqELD2kdUhPsuekD0OkDj9RRD66h0SZS6cg4GhSSpkK/
kxsqYBIIf7Mk35yNZtSKxM3/4a2t/Rr66knKcbyHHT1pAZyIaJHfg5RpMjnRh0vt
n1W9a+Q0ghCSk1STraXSBf8Ore84rAcQMBXYhaAuLktB15RMG0fsjWt7yR13/AN6
3cIr6+LiV27IQ8meHRjDTgApWQrInijHUGnAfOiD9uvB6MzwH5bzDB78PiMBaE+b
+gfN5nA5rZktsYxYPq0kKYUx3tCEyg2Kz3dPPJ+bXMj2i02cpFrrfugOufqLApIf
uBvY5BDIcu+K17mUIh1SzdrM8y6V/YAmgM4jmb5wQiAnxhal8HOTQTbcHYr0tHYP
YW6QPhT1ow0NpIAvgykVXqDSQ2hBijRnBjiaZN8LrgTOTlcJ41Ehhc82NfT5mNHZ
2yMuJ4w2JL6lCoU4UuAhSGpPxvTfZQ2ffQbPntXmX1AOUNTsxsS2tMe38gX9bFr/
vTtjNfweqe8BaEYSW2MAUDAAXMa+o3AL24AgbNR6Ca1pEb1s0RXHb9WTt8w9cCc7
UAD2wMOYtVaSDz89rtR8ZW5+K6P4gprAzzEM4X1V4J2dIdriX2bN1I8yM6C1CnJv
v/bRg9AVWshyRzoVxZIpzhlAJWxTcvEdbDekmmKKZIRqce4wxKmHLDBbcyjBOlNY
IRemmDWiIDL3IJrlya2Jz6EC3I8gA0hvwNg6ZbIBqsWWdUWejIfO9jVx8UWwdjw9
Zpt2539pzxXg2a/jwK59IPxshCZ963t1MJ1PAetGdhsMWlHGc2p49HXmRjwOZqlm
Rzbz+zXyxYmdeMuakmsCfyCO5nXHj46xH6bnfF3hUotnWMoKCIgs0sgXYmvtuB35
c1LBbbBtTWhwKNV9PCDqU+9mjGI5lAE7icGHOUMTJeixubAiS7nCmFodDIikbSOP
9YoDaMiy4CePbksaGX8zRulL0RvzHcZWYwO0jFN8cfDKk6od0gMy0U0VfgPG0r0r
nzFqPusgmPRBRxhyhQP+kZzYLQiH3U1l/CV3MzqrGJAJQq7LV0LeYCDKpepc/+VL
++qt7gRSy3HxO4FqfNdpLct528Lm5gC67Rm3OTC9lmC4ymEXCkLzjBjpOPxO9LAe
bDzQEQKrR6MedBRyuVab8CLSl+rzsTvk2sm1kSQ0/5K9uXiNt1aJd6xPLjGzP76i
JzNGt040K0hJWIN6BixyPNZFqAADFisKTSOHVyeQgA+UYbwsChUsJpiXvt10xP2h
yl53uraV/l+hhuMMIkgXrNImf0A2bquU5OW+mWQ3gXI95yAEzBAf74HprHDtR+T6
wSGzPGOpRdpdY6EtvHh9/hk/jFP+BGvb9bTdX0yORbo+mle8VVZwGpUP7KuIX6bw
GEhlEwsTHKlY6ISA77qKOVScA+3clj0zdjLg8gJZkbOD729GAaWo2wovTVsnplZQ
YmOfDxkRQW3bTPb1Ac9Vz4gA0hmXgR8TxaQx0CUXgJzFE/bOrfp5eqaTQ+A1K8De
gtlCI6yu8pnkI4Xr0Dvx0jvU46l/bCJW3fEMmQGb4SUcj1g4xJT+rknWnuXz+cI5
6nOK+BaF4nyA5hyAMWTNa+CZ6uPMlNYTlNSdhVCBIUJdMq6SCmvAz8V0tKPwHUEJ
rjaJp5ldHuZOdQaflrX7ZB+BgXOFZl+EBE0it15u3mq7DrviANOJbIkmvENiQMM0
hsIlWVA9MDGONMWdgPZWbm3kKJciEu3VvIqzufMQkMIy4Assy7ZUWxzCLv3QznR+
u/S9oyHNF9PD+ML/rRem1tfGXvI2ecIDIRM227osp9qFPx7mTZm2G7VUoKEzSX+W
UYqKj6WQFtKIAw1HIH/RWt897VqeEUxYLirPsf+N8WGZoKm3lXSN5ugqmjVULTkU
1Qx+KMfIbB9D8lbMWLzbTI7y8UZF1PZpVacC2/bP/aHDMGDmQlPQeQoMw2hL8wP5
06UM2X8sYfoUemLaELBEpae0Osfb0HFNv0kqHuV4iCBwFJVfFtu/RR8r6mmWcRN9
9bfRs/W1L/hpoAUY8gUgS+MHQAGMAlVqXo6j6B7HxkJ8pvfM0PzOPaBfxXlkaUgN
gy4pwISPB1mviQEBJuXAjKFSNepMiE1i2l0ovXbTrKFWaQbR4ApIz5bnOZU8coeu
wnUe8wCDJOQ1WYtCd1Xg2vdF1o6oqZ2WhgaoLMCTwvxAxpkKRhbCXSOttlVx6+Iw
8fFKVPFzzYEk0igD62oqg759C5+id/mvDN3fpi7wS4xSIqgfUt77SjGtyV8w4muH
uopECnv0rfx0S7HArugRxhIyaJUoWVRKZzqRi0aIJqrThoMhwpAQKtQ6pLVyeZvR
+X8kkZDEY2CDl4/gSF7rnOKzJjvqOvlFjeQ7l9Yq33OuCiGbxA16EgNLeRYiKhcz
ub3cvR1/3UMYcXNnom52M84KRwSxEmvD9oEjcZZUeXwk7hmX/rdE3JOnB89vlRTf
6pGsWTw6/L+mxv1D9XVi4R4DjXXrE1oQoPsEkY1g1Y6GtVoS3M4w4oy44A4B7wLU
2eOXrTpUL82afPFw9NuA26sTI0fPbqAeiUkWFDjO7CSdcVuOxjqKCAKgvnbWBr+d
qxf7OOitF25337cFydsqfKjwBSwyYngROAMrYqrsB+KaOl56qmOPC5yHc3WtEJd5
9fzfwGEOvXBZZz6sgIuS/qLdJ2tyMwdAu2Obgw+Pe3h2/hSp3TF/dhJUT6uMd6ks
rIM34LR9T2U28OXdqOlr+7aSG9voyg5EV4zV24XIMqZqrrPdJYJbgcHENHSSakFa
0i8Zxejo84o7L3+bEMYHmwZF1E5wKZM2nTc/eN3xqRpXbYEt/y93LZ6/UtPaUMf4
iNvEnEdPQWhqwG3TppsBrg4qCFBxSSPJ+NSWRWmFh6GDpcEBqRYq4FFz/yAelVly
t2cHWarWIOR4yj1pWQy7DjUd2t5cnRGV121Z1SdWIThZy9TlMya/w8smgO6sbU4r
fvV0n97LAJrPeUithu+b9BN+l0t+NEf3yNyVyRyNSDllULE6BGTZVOCKctiYxfEP
AClMi7qxikb27W+10NXoWE5oWcJLLfZVAP2O8jplku9T14gz7cH+2074s9IwaWwE
UhaciNVISI8na6Yc2fzeJdvvyizprwOxSx5Hh3Dhb7iBqc9JQUHSanmzmur6l+DM
H5Nrme+dIRtXgnErIdbAbI38fM+15OpYiK3WQW0bilVc6nMC87vjaEPZIpPG2IYR
j5IrLqXa1B3QQjsykysa5IUNkfzKNhvJL/e5JnPvXLcHoC9OXyP6zL7hAc3zDHX4
LXoRpcwEFxXa3SNB4wv9IucW0ZP4+V2/THopPE9WzG4AhmP2O4BKuQ02vCtW3Y6t
5v5CM+6loR27vgTYrJ9eosRR2o2gfzDFxqPsv1ifycMoP+rwhJ1UqyPQwn+vofDD
y0G+K1ng0oeRJLviPpNAyxip/C+OKGIFLJdNuWfdA9/TT75U7r+R56iAYdKVOaJt
PdDFfE42Ea51Zz2blcBv5ZJEyydxzHFKIJjL0wWQCdikRIVqmffSJqG/c9fKtHmV
mjg1IVSFIqNpuzPkZ/5HeZiUn7Cw56/heKjC13H/kqvx47JAFdFSAbb2rS2RNs6/
2Y51bQ2xPCq5jdraQBzGMuuSZuhee+S3FGpWBCEyhj/k2N54OGxioefUzgsxoUYT
Yk+J/MHetlGM1BUGx9koRju7l8QcWXZ3eBFObqXm9TQ13Md0lu7sQlmUrWV4BrBl
Uw7ZtPuwqEzvqVnqobHzvfqTJhY4dItFuqDcwXbtj9FJArN+90axTj/+w1CRv82h
O7tivp8WyMg3VqHNZYyrPziaDMxspQnzl8t+AmrJknANWSbsMOX6eMGA49omFlP8
IdxPSUXtm1p0WyDmGpZ7uqBFE3FgPGH0sxznn/2U5eH6FUFSMRmqGO7aRR6wSVoy
0ukiVwfSclG/mxYsiIlJJqYe2Uok0Tqfn7p5x8MqKE5wqqg60CH1nC4QexPaZhDF
Qy8jtAfVREz4qZ/ac1jtttNDFZYxAqOln4TN6qD7jwFq3+tsjB8TmBFiZZEY+aJh
71qf6dskGItB5Y0/IpyusbL11KjzuPAOxUpNXaD10P2Sdtv2/onwveSe30vqKbTb
ibiXsbVEVjv9IH6PwvyA7Z6Ji6d76oo4QVZyCpJqwcx4DHBu3a5ss0rUS3Ne4INV
Ff299hjlfy+69Ml1ZQKGrLcIojCyyDN/7XIkRDCB3sgwD+Q0mR49U/0ajQ7rf+UH
TtncJtB5+UboRHavW6D+EsUiTAHPT6urJMiKHAtp6PaoMschNBTW1YOJ8N6esMBR
Z3IdZz+NhkkydsR3ZWJdZ7HP5X2lNWVzkI0XV4REk0o9yVB/N3iuC+/R8gAMTwMV
+PnSGWXisOmxv6rAxUdtk2Xinsx81HLeHzuHnUJ9JSJHR/M4b6ZqJUco3h+kIDVH
dKu5iLIJP4ndQ/79uGa+OfPOSqpCeioK/q5xko62T2yrDvORYwTWtyVjLbP2t3WX
DUFKEVTKY1k7BwEGPdkRUi/KnI6+TX/qyOJwOzhJDrIXHm+F2wIOUyP1dlY2A1X+
/WEnFZf5e/To9+jcKyGYf/iOMxKEv9gtr2qFXUjoMD5WOLke1nAqWLcRgGCQwMo8
vjueyyNGAKVNHFwJrMnCFbPfjrX41xV/V2QLuibiTNSJAMaVa1UDdhRG0hVpqT46
5goBTkYHH00jmoJs6wMgBPwGzdJBOcL+tYdCuydg+NRwiOJ8pMVaaI+c3wHXWCsS
wyVIIS58WoGrWHfcQWDWXaa2e77UxjKtQ+mYVABndhm6oxioUmhpN9GdZndGaPZE
dzLzYvNrUAAXqA2aWdSEWzBhW9NwzGUS5svr/5uZGxxiJ4nuu65bYd7quX9NvwBj
IE/1GRZqi9n1PhoIQm+Je5Uruz+Xu9VL43Kc5EaSC5zGcxtqJL1jRb0hxZfwaQL0
zzvMn+IUxkH1pu47ONNW/sjO3874/1FoQbRIne+yeAkz91jFaGv08rZgTt/sz9k+
pWnbDP+cE08RtNoydVb4/dUHw4WS+lxEUkrhTmUO0ouGF24J2YKGAYzfv+oUjIVt
J0XDiV4feeKRD4NCLsNnJObvoGKMGpg9MCd6nITF3z1zIpra6Mf6GPL9DY2XIhGa
efwjQO0OZNwMGyt3Rty+PSDXTDcXSXoLQfFAwA9oPQQ0mbxCYH884hr76a3U76l8
QSf4P69E8hXgpjpA1qM+1HdfhpGm3gPpqRY82Q/oIvooAIAYQggPvzCz5bBDuk68
J8wg6MMQm9wvcvC6VuznydEhvG9eBFn1e/Vy+ZfQRnzR9b6kxPTYWyfdCr1Op3Hg
7jl7Du9Q/6efheeoofRkGTYkZxCHGsB5BfTaMkF+a+Yyhw6YTEtspeyO3jjGkoJX
gJgXXi9HOUvH4cdCeeaxiyr9eV9S5qme7EFrG9fUJnOwR5NyhJ6kLj/dtmWlf/wp
5NpYd8TD8EF2CQg16gqzCZ2EUoHTUUGQe/s60NUrWfcCBduJT0coQWnGQuYHWuaR
e6u+Lj9rAe6asNTZi+Mtv+7YM+qML/EDWLMPw+q8doFANbTvJ+tgygoOpWyPLuSE
TqjlIgCCPCpGQgZMt87w5j4YXu+GUM+hENYsVyMtOUzQZ1V3pOmH7D9xuFtwu0ui
BCvoRnybFgFASdgLSn4brNw3RdvJ6fAGx9r1m4VBjq0v6+bcAZEmzmwjZ0mkjLdl
AYDP7bb8YYnCSn02gGwTzFLzsrIw1RBTlSEluYdrLpyf3oD+EWrn/lFCBaBgL2j6
JWc13CcXCjuF+tKwcPXg6CAKSeaScOj9lbGLDKbAsODHx1sMWlwxSnbaAdGfmAGF
TTJalAvLCOujPEpHvbDsbQSXkojEnCU28Wbfj8xYmUWiAj7zrSafmeaR6h6v+f7O
kiX5KmufrTMsI8ztPeLxDIpLup1AQGTJPiMa5Q6wHHV9yZupYGO3EKSRew++AFrL
S/X5Emy5LbpgvOsvWBb5D5GDBmyvDj3MORYGCdFusKDoi4muCDRgtSO2C350n46r
Z/c1kf/w3GxZA0aZjs3JQG+oG6nlmyUDJy9YqXXCgovcNHcVHU7HGIXF+vTWP6nP
oMUxmrdfGHlCnPaQSuc0eODkOMaXK26nxxt1V/e8Wmpn7ne0Em8WClUYd9vV87HC
SDvsWP7BSIk5Eq2kuQm6BkwIjE1RggnvyEPpMXV1xGyiXlHFG8/UdgS0DOGDbQ/c
mkMjw4IcialL8klUv1oC+H6zOBOnB0lPWpEp7ui4Tmz7/lkP0KOj9ZCF0p/71x6E
655q3s2O+csQdMDPeKxXT/JLiKfGyk3VAe5RvF+YIiqq+DNrwaH0+6FHmqoi10Dc
t2Iz7kRrJnMvp6I7eAww5iTwJ1LN6MYwWPAtZeeFcenjWxpqJpCHEoE+3ldm6ZLL
OO0N0hv8DKm0+OWQB+IX3DJYC7gFZa7hOazmQn/Gr0WadQUGrjf6ggvCjAx/M6KC
UxtRQaL2nr6V1vqIg53jRp/5+VC7q7Z+5VRW43VHPgjDZbYdXfoYXwBAg5N/7tT4
D8zqfWkcXF5jHOxoM5aGgcYUGjYOJ3Gr8eM4EctpC6VQwpnsfroMbR7w+4+E5TYF
ET/UICsRT24/+hU+59G+IGcw4N94kNiSRIRBtiVq7fS5yVofofAqx5zr5EU15pXp
VyWcGfPM0MLi7SicRUeRIR/QLPwsjVgMQxkX/0SDQkNQO/AIcjIw32MQ6epbceHN
qHTDzZXjo8s+SAcRWe51vFWaeUlxhHd1ZJ3LAPpjtqNQgWbNq4R4ICAkjKXe4VId
ACgIO3dHmhCGwGjw2lNidyacZeT3TVzDB+x522r33IylPrV3yihpzuG/EaL7Ipih
lmuVj8h2jXbd7V7MAq8VohRiAxyatJ3Ww13rinv/KdxerRYj4nP5vKiUoIgiJXbF
rmz/qu+duOl5fRl7CBKyZTBbgLE8IXTm+30qWoKyRJXwAiA/kqHBfzYMh7V/3lzx
q5CrQwqrE/aJTh8X0o0vB6wKEpjgQhUDPwXLTJTtjd2Rweq5gFFNSHRYBb0VqDpY
44VrRGpxpFKwuowFlnD25mHaZAHPLrxP82KHRcRxUe0w4wr5NqmisWhvE4eKTRCQ
VH4AM9v2e9H3Lc9kuf27c+KEXCi+369Iquwb95cUB7y9fRvE9b2JdVRcbink04l+
+hM+k48+Dxmhh0F5iYT66kUp0UX5ayiAGLOSHYrtyQPsJ+rvjBHDTj0KaSwXSAq6
Gn8hLjDMdZ8jhMY7qhQxbCppdjtLd9cbJupEwOVvTTRfR3dVdSVaqRbp7eQ3j6Nt
xrwmr+aSgxTqHHpyxoU+Qy8KkZZrp9Xe9yYXtcjFhEV6jY4FWu9t6JJZdwq6S1oD
qroBpegUzwJov51dYToni5qz6fZ1TLTaByOQ7kPDyh0W1+3AHmlUnoGo6SMWjebW
dHICinkM4fh8vywPqf5fI3YSb/kYVDmuLwiJenvS6s9tmj8hy1xXzjYjOLx7JTO5
Clhd2gVz/jZoNglcriZx17lWc3fDPZAbL8O/29+Kmw8FtV6uL1RLPTTndQ+Ul/IE
pErEHY0eVL6a2p+oXFE5NiOVYnaZ4KvtYSdAev3yMenV8CPMOVjiHx+ONW/LRjMp
jpS1Xs1ZhrJE0AVJjabdJuLrfbRf925e6eclws7wtUTa3tPpZoWslvF0fpAeEjPO
g+ml31WXdC+BWmP9/zD3SW4JQZitLEy/E2g0RVLQyTQFwmDjHPtnMTqhnvN/NcHz
qGmyf0A6O7eNWLhNS+HlKnSLJTFcF78KLkqLIznzkofF6oNvy/qdw1WWE9ympagM
og7YgfSRWU0UHMY0S8EI1A6kMMYYI6v4TL2eeqUQSxIAP/8Fiiy3xGourhIhdrkU
625HRLsdJJ+Z68rrEjvSto71vCuznzegdcSNmlU28TkEjqJWf5kADghNbvMssUZp
IWTUcWnurIsTbXVudIklyVHJ0kUvg6xu4g+JHrpMpMWiBvn5ReaaTo0wIIgGBnGi
GBNth/DiKsdmcEI/F4kx1LFxHVp7vLqqDmxBA0m/W9Aq5aHBW1LYrrvKTneD9M0X
KN1eJQsV0bQ7/NS6Hca+NXeMQ1QjJdGdr7ZZU9kM/MYQ0eY/5qw+dbUzqwtF948K
cSl73JYIvX+XB4a3KS/xwzLUuKmcoEaiZeVUo4KQetvsH4Zff9bNkFRz/5mCUrn3
tAndnc+zMMjT1d22X2JGHOqx/L1gaXt0NAjbcIeLamPM6bVPeYyGmVM2yNArava/
GQdf8GjBsUbB4vIlkKLubkz94O5nDCyS+miAhDYX8mxZWkhn01p1lSzVJQUvNbtR
ZkD7sMfD/rS9Q9drM9VKE9BQ12YkK9Rmlk6duIlelGbCx2nnC7Cnniw/tcrNNEdG
SKSYcsCGnuJzceGtk4Qqof3kxyRslf8VEXVvy91PwpCt72Tg91Js8Qz1R3iS7xWg
DEN7WyLe2NmYiFW4hr2xv2ds37rXPLABFDfj9OnVaS1etf4gioIQpZF1sB+SVIph
PVGsFJKrWJ/tyeR+9Ao2hAfKlDeYpmwRzxeicIFH9SqGGWLK2ZfQ1emC6Ysa7yV8
00Ot7+b8UjHhoxyiTQFUeTWuTaS7pEXTBIy0hP18hsM6hlnnH9c2IGYP4c4YVCxo
SdfPyLq2Yhgo/NYx4Zbae/sAgOdI5V5NrmSIodLi2GbFKR2BcksUtsFNcY/gWTY2
A12dSlyIvvi38caK1ppOhblwqr5XknqimMZ0zypcAKi++W03i/b1Ht3N3MeOEXB6
mqgh9NYFSsRr3vS9TmEtG/dpFzbDPcpdU6tUAzQ6NwZnvnYcs/syFWByIJfbSO1/
1gUJip62Dq8BbENU8MhI5Qs/JalxE0LqDhhpnHxmKcYKnQyn1eTDlwn8IG5VPP3I
KYZvpJ+CndQtvSqNUOOAXh20X0+kRrTfErM2bO3PzfsdmSbM9mYUYNuC1ayHlgww
tLzw7bw/3X4ItpAhqSwn5/b/dDrDSiomqyAc9BwISpNk/dbOvy5W5knWGoBqihsw
kw6/x0igjmt2+nCAMQ4PQQZyhGb4M2K0HJ/Q0zya0bQ1CzegLyPI7mNUakV2oCxU
v0Hh8GNN44zau8Ih5GP4m0/2RpirmR1ZlhldgU2Z8MmxN9YWVM18SB+rfYoADDd3
dXgdCwmJ5NZSDF+cTD9HZgV9TF2eNLpRkwIldFBS7v6bTnbWypwA/mKwYMmrJsUj
n9Je0B+4ZPVFsWPqvYTCbiZN1YnfaQJQSj0CN7LHoeTW7dzijXpCBecBDyTP5Sg4
0h0Ufisngzf7GT+hAcOqr/xRy/uaxqdv8tBrl9rPxfm0DmfQDC9l6VDzUT8kNuDT
X8wV0s6sD4hptDw/TYobGWfv9zTlw1YB5pUY/yEtSlR5Adim/wLn9sPSF+iFtKa+
q66LGbfWOaRt/ABJWmY5ij9dV26+ptlJpjtEMTEo8Dgvuoc1QPkdkUUCpCsvArtH
Yn9lZCQq72x2P7wBKPrakV9fEsIsRomIDqIppAqzTzcFNtXTivkyNYHc7ysjqXB+
dK7Akkbhka4XjC+afgDvPSvt2Srt5hLRq/P2M0bBG6EdQ9VvcqlpXYIL8Y1HqnzT
yDACoK2NVjQqRNGndiVQnGANJvTalmih0m5019Hemwo3voDJa1X39A1SNxvWkSIp
VJZqAUFlfxS73Hzr86zou+jMuotsV7X8REPCSiSMd2C6Caj0rM3cZHa9IPqTBVpx
RVb7SRZkkIfg7hQOcP6IxpcPYF/NDlFEIsaUXQVL+rsJNn/IUTfRagCgfYpA09gl
P4b+HTzxFBhrv63jKbTqm6hqVy6KM2dgMqvwSWw0zgGzaIVeB//aW9DfJw3xMCN8
06esjaLeBMZIafghfdaQMegXjGiS93a+3ZlPZ/XmQ5LUtIFKYgcyO6BQ3YQTcNgC
165qRtrc8dgFojo+EDu66gNVOd0KgyxkLgmS8YsCgfX+hdwHHO7YPx/18ITR49g4
dN1AKGCJVE1/CaKdbxIWj1Za5F8F8zj97WcliPAqEPOHYJSsj1kBYNH5AMuETqF7
AN5VCWH5oHlXohmeUU9nTCbVsABLlzEqi1s/ABpyfv85S0bABk09ruXiBg3LVHAK
EIVWJifF9/Ka/RJHV2A+CHTGbz/qDRj2hPJPFFNRxrO4PTdVMzJQRRQYX3uqKkFv
lmJei/4JlB6eDC2ix3Zls7pBaEwIT0ms3+6sEen3fF0iDI3bFm8PgO8u9fNTKos0
+r+QLr0cbEBZbAfNnYPz/kqCzEAicZ8LT77edN+P+rbXhGx2BTMx5yM3bBwkOTL+
ceXME+47w/FM0QsInXwvI+2Jwk/Wx1TCX0h9Qz32c6rJwqlO72I+EX8UvtAicgfY
1iN6YBEPAYnEOuy7AHTkK00I3jhXqJ5D0ag5if/zo8xvH6M1xnKwnJTj4SJV76dp
QFe4KtXpIpcTIQAQ0Jo6uf1X54A/RO1V2XdufCUcZLrRBU8sc+r+dusOSZedLHCf
PwLeug30O71vddhjFEpcMjk1L777ra/SyCd6L8AkFPSqhjABPXQYOB9bylGncdFG
ECjMgm2zXUpswuyGsoOGraJfv4y/henhep7VQS7LLamcFgIGYeHzqMlqfkzBHCDi
PU82fhxlHEPTF2UVBgCm6oOpBazLgt4d5sSWahaVtzNqDCW7CX8jXm9vSbBLvU7X
ZsBAecOhhdOseJR9/HSfxLc84h8hy9FvTBNhSjbeg3YtFrgxohli62h2+nuzmNDZ
YOwxA8VLU0O/ZtfOBMxxXo5pfn1R5L0BjpoI3K+LZIDuXocjNDuWastdgpcxxSS1
bc8XXWSanx5VUClmBuW+kewI5AN3Ywu+zPHVwuV4Vx6vivsHectPG6yEVkLL5Y0I
bmtKFt2Fmlpm699rD0e1NotxxO4kl832MWvmsZ3fIXf3+DsTxVGZoEC4I4ogE5CZ
lWsS9mQRU0C7Wa+lYXwWtAocN1069TcMYDizc5hvhiijLdDnM6pQIMGPd2KOUtPW
KE1Di1J3+Wgk7c3GnzSIsauAQAGyI9Sw+fvgOvRdab5fAGEdn1EH3lacbOyAFRIO
Os9iHpu7LS04KBvGjyPB2a3U2p24h2ds1/dNu9Z5ZDpyPlt9/4WKX/cXPXe5DIzE
b1SWzEdRGd3/9VIuRTAmEQehGUkfIoTmQEyX3VuRImiKJshVH621CNXlLA5MHvhG
P5Bfe89x2OHPwYPjW4QEEaNBa7tqkEPUPoX/zWZMpPyKOuxsJ9K1TOv5E7SrIJ0S
ZUj2gk5DMSQ/hZ9g/M53Ij2HWJTutd30ASZWJxbGCgy9naYB6Q0oMzBAeKhklHry
ApDHkL21vk/uvR3AL354pJeyzKdKWAMPHEK8oPgyNC/BO1ixUPp23kSWTjx2fIdC
nBMUdL0mTsXSegdDhsnF9qd+za9UqpJ9G//6vn3aAqbsT2gAtilkZq7803E1LZnF
qAWTTQzY9WDj1IgGEb/RP47MmDArV8aJ91b4qi37txxx6Ja4K3k7DDnVlSNCKWVp
J3/DXRJgCfw5BZ/oqd45RHpc5Phz9imUYZrUenMspTlQ/IUhpIDDqlkMFcSgm6K4
kb23kh/TH+h98kkSHxwRW0xrvGCWZiisSKe45V4f13cP1zhELa1hf1tG0G3nwCiV
zu27ykqH56J675Hkf+adG/cljH9y5EhjUxUt+uxI7lt561y65wF+YHePUa4azmZ3
RSGAE5uViVvIJwrWEBb5Qp52WVOXYZ+SKMJgWe7BLfpDi5EsTKhzFrDpa8cGR/AZ
g+fda+OMBqvaB1+SFhLugAtx1RCOJfEY5YWpKsP6vfCaXVQvquimyOvZ72nSOvA/
AIKBuT4u2RqHuXjUL3NDLkwK1EcuWTu3ConFWt/xQwjzBlwBSU6/8waGsxD/nCWW
kdP4QxFxNe7G0R+Il3mR2ivulZ8/LlHgr9iWHCUnbk10NszwVe6Q7EX8+uVUjClg
mNiimH0VDpCLyYv97TZnZ2UuC0945N89cj+gLQAnpXeJx+f6uGYK38OxXb40573l
n7bWJF3CZwa2dHk3eT2Ow5yE0x8wCVvTMNX76LjRekqAiiKtgYrsbp53D6yTgcQs
N8ZB2UNb9pSF3T+C1/vuSvKApLtJeuzgVeJzcHChWZCDQhqkRmiJrN33CBQz2xv0
i9Xf2X5JT20T+ygCZ2gGz6ziBBfNOub3DcFsnbDX9IWhzaUr7r/20qNc+iTNMJnH
Vag3GZFTLMC4DWfF4WPpZ4fYhzQRbg3m53NX6oTCKdwcwIiDOTeJv/LAmc4LyrJS
j8gvQs8xu+pRW5RWv51KRhRt20N+JZDbeX4WPVwu9aOxnMG9DbWRbwP5DFvn0sR9
P5DlpaKAtgVzlJUDqgdxZxNCIeVMP02okN8XLgMYJQuu22VCT6xa2WIFrKNkoMux
brhxp8Gs8sOI8ESs5WzH21j2AmVXohdXwPMd76QaAqpWzT8sRgObTZPeVT8VLrXA
dkWsL9LlXCZ7dI1sTZ+tchIAVlOET6I9mzenzqYgC9AqbFRnGMWAVdbl91HYBdTu
8zXagWBHZPU+6WVLicIjo37BLWED8uWKFY6Jaw+yFGEkvK0jMLyS9lCkYQzr3gzr
38hIihfsfPvZixwWX5SBZzpo+w8L8mdluZGZHymNlSHY0Pe4ogG+8lNc7VQUKqNW
EUqhLy4xoo8uSWQ2cY+utVPIoOw+1Fz26hILXwHj5DSFg5nBJfJlJTbO3agsHqUh
GBaPXP4yb3C7usiFvn0Z7O+0WSWgD6ZnZ39v2eerXM9EVzZfIwvFg4nAgnOlvWUi
q1X+XTpenqyW63Mf68zGrf1QVg0Rx7Rnf3mstV837vCzJKVsroHvffQ315jsFXlH
chlAKoS3nA/XG0nxGLc47RrTHmDOiF+MwNpcPt2qOUN7IrUDifRyuvsjRy2bgLS/
EUDGjiaN6pra8QzVG6wwEbdDUeDTC0/YKCcNRSr/YiZB5Pyyl6EDc+NBxJMKwy1y
mPZ0JXblItbNUtZSLFlh+ki0blAGcu/iC5+RcTZaiOFZKq0q2cxH4hIi9UO5jks9
E4GOBQNluBknZmvqkjh3CY8VxQi95B4icVc6QJLUtX2Wq/VjHquyrVh0I5cMDka3
axs7YSYBVgfgmjCE8tvrByMXKu2fkITJaegtCn1CZm9fX1KaYMi/UQPHHt0UWTX1
qacGhvGTX9AOw/2ISKmDbHrVZ4j9/qqetUTIsC8T3EwPqfJIeSGZTh0eNH261x3i
AG8BwuxIShP1rnJxe0jv4NI8LU/Ec0f0vA5wfcpUPxz/obfR8c5eIwK/bTdLMxt7
Ba1oA3qDruDPxvxc0X+uYo9r/5XD8IJhCGGJZkEu5iIufjv+/WAReV0OQsRhnYcZ
JjSIPm7LoCyLvIW+jVR8cZsBOPCw73axJyg8sSgr9k7g0vN9nj4U7QAIvfZMpu6M
cE4zdyg8L2buYzrUedwa/rwQ+XZS+d+XWFnLSwjOqR/b0yCPM9/NPv9eDZOlytMf
E8h0ExwtLS+6waEJ7lhqgXEUTUaWxxMMO68+1Wgxoi5B3fJ7mnOP3AuyWHJx9+yX
s15xHsFy89KgIeqOFEmIPldiM6FEmVWiiHUh5z7bWD71Y1wtekipRtFNs5LQ8Y/h
YQixL1aOA0FM16ueo6f81gGvBy4UTrVdbZMTzzSSFvO6YeAEK/D9MveasPGk/GcK
ebHvQ9V1l5LwcVYKb7qTnS6ZGT0znqc3dZ76mMHh1WrGbHUl5fztSFPQX+5+a5jN
6dIVOr8T9iFczadQnA2T3gDP8+KRQLirfbR1+ZioEY+vg3GxCguQwPs+5mQTERSk
2tstaVRASEG1K/0q+iJpZKY7J2VXqGd0NrNslK5UtU31i60Bms+1ET0iNmaFULDP
YaJlNIqCIJT5hgdBPfq2bJAk2Nfq+gmn0dxdoN5JSa6j6e10ok3me+qTLUrhYV/0
gPp5HFtQRoZokC1mejHFoZRs1F/OpsT6NYFEa1lDH5zQ0NW/TZ1xm3IfMfUAqGh5
mj8Yz0xfXhwBKnTBFPgQEL2/Vwc9kIQB6OlZUV6ngSiE/J2jWgdZ+LOys1zu1rVO
M8M6/sJ/MU50pzBMCDBaYy12KOZdxxBj8hlzxPeiyIZhKQvpT1Yq/kbMGkggiHoD
vBKLt7JvOK67+XZCoZM1PA1ZCajgNgA4A1H2N9/U1hQDcV4nTBlNsoJj3hZygOkM
Dvg9gQm5NsNlbznGLrdV3cezWjDKCw6/cHu3tU18Y7x8u/rs1o5cm2it533KwddQ
M/V1wb2Pe06VNIh6tsTiL/vpaTvVFLMdZ0/MNHWs7GwTFX9Wqp1U2nm9gHQrgbJh
QncO0RstMj16r1CaIiXsQ2GE25ZE1GEFfnsCWUGt53z1bzaS19ap/cLMmRWQJ1ZO
4vU5XNkkDcI1Tz8zRAACRo9lkJMGVEDJ70aZ/VhYaWcP4sZrXwawbANcf2/Fi0qp
oH4OWoiFZ0E2Pq7quHNK8D88h2+NoClkgW64dINfYOIPbgzBRUw6dVtpFpQx5iRy
C6eJGCnVjqsDshyI/BeQOdcQtKpHxAGRQwmHEBi6w+WpdW3lugAYd+68gGYTFtss
BaBFC31XNfjaXy07VHhZnR+tNLx7rbdfyh7v2+CD5cIoC/+Ps+py9oznf4TRUhCc
1OXo178KcOGw8batMl/TSX6GVSgiit2taed302ol1rwots7dglJVz7yJETUmNosc
PRwLwWnTPmWVdezu//iCL3e+sFBF9L4mvy5g5PQ2h1IZIIMIcJmjd9la9VxyG2M3
rRW2rwXsQZm+tXvnd03Zmg3cJ5IPPmdlDPQCUEaJFrwijH18BY5eTTncM3c6IUQ4
3OPkKomX0OhfIFZDPLqEsEa7o0YFVOtE8baoI6XbnmtIhXjhsgDsx7GJaFNoU4bP
6HTANEJxWuQ4BK4gm1B80kTAQuLiH+iPAmQfMpYqbY7wEjXQmh1Vcu/khO5yzI58
i9U9Qelr1YSOtOnBn1lR2RINnoZo/I06vePQVggejFctTVW/Hws8momOdp0eHwga
Favi+PvBTnEIQFhYjuVunAk3uJ6c5izFY96es7Yo+T6Gb8rGi02AKPSvg2SHa6GK
TlpwPhIQ17+DaAmF0ZblOpsiG6I3OoXoDDAIC1YztMlDbpToylfpdq1McnJXfM9C
3N5kyXsFStUqwJUZH69IMoI6J7Hvd+PPS1do5xwoQiEJvcXz7PLpZt8ZDokCrMuo
K31rYq7efn0qQmcpM06Qjve2j4eQE8vOCgXiV3m7saI8SnUvBZTomx1haCu1kYBu
yvqUqAKGDewqEI6GJFeDES2TozAbPWcaP4wXTohpPA/7uxbWT3GMYWRcfx4pBJta
0IQLfhh054LVSn7ep3ho05Bo21eRXoA9xX611BeJUMCFUKQ2fz0uRhNJKLq4aB3l
Dg5NZPHosxsRNMleks/qj8HcHhSvb/utjCUHwLKObY018/ZWz6rS0nQcmC8lotkW
yMAFc10x6MQslPdxT6WdeMTFM06HHp2Oek1FULPRf99ukjdgq/RWgj6HnHYwHYat
LfjViZE9W9YKRbdhY0j+offPuHc3af4BSl46S+XUuEX8/Rg+Upsecj7Qk3uXG1Zq
IikgL7z43C4d4x7wa5BHNDVnfF+Lem/Uw7Y7W36svJvVpa9K2UpCeVoGZtYR5kE8
LKJTL0EejdogRGCf6S4rwxMafGUjgXg8G68yLHO0Hh2dcFZPObfnhOWqXe9a2lhX
dvrIKhICRQrtkPYR6fBsj6hcWZLgcDj61tH7WcVe1oTK/BIv1uACnC/3fZDbpp3e
NOfXSxK3KWDA3ZQZ9DE4hTMgZSda5uTS378fZY/MXx1Pa7T2dtxk+AE7GNd9JjaV
nYV4aJ3H3Z9XNNZXbCYCVBOMRfAHSuLwVD5X2Y0kooP05pkCdereNyWaiPfno3ja
kqkyHLjOYcO3AQs0b9KBKoS5tCSaK2itTIkHMe+5YRUNR5OwpimDng1S0ttcMEjJ
83L1Y1o99sshBp4FlvTJ9OKYvlr+xq31232Nt4k+9FA6Sv+29B+Jmsus6bW04F8l
iACa5v5dWnveUNpdXP0TwmoT4KA7bS/7OTshGal7SSbIV1ivjmoWt8hHapDAy9qY
WwwfIyL2lS4hD8a0stQoFWkVmM9x0D+DGZBdzAIETtueIpCkTYbS1fpdq79zaaXp
yPMfPzYUj91+y+ATYYtK0zPfACC71ofW4OX2JAaULZKmOHFD0TOLdfQYRq/p4gG9
v30upG/UKh3++x2PuyfgaevzM7AcvoLcNy6ZtNYwRxlPg2V72z/ClGuTf6iazLam
Zr2Pgl8bWMMJzDNZoOU8MbRttLXXMMvh59reIJURnjmq4Mau3dl92h1OMlN7JamT
ffkivagUBxAG8xcLcmHH3l1uAVuFY/nB94APe5Aw8vI1Gpv2zFM3t9Wc6u2gfqkv
11HszzNxpeEdudNz18rKKOszzVhreNYoeDdEkqCiUILblaejpPNLE92O/h+KG1cV
FvfC4pytOuzELin8LYUU+u9bgkzTXXJcrV6xdU+TqYen+qvxpfVmTbICIW4WJAYt
YfqQakHyM2PE04Tzc/7z5ZfiFvb2vzP5EdKQRC5WuioV8G6i/vQnAFZXHNTqfEoa
IaoQbwiytBVsObCSgFs0fzbN76comw+OfxzATE1ayyiUOnO1XRcGspl8izkzLqOm
jwppBXYMh588R4PBFcgipyU6W491HO7fkNDIqFfTPG+qHCRXE7AA9zbXC+o1SAJA
bKUx4Yobfl/2ZUVB/KRobkQhas1IAvPvBvrCazS18Sljg/FC+vdREKN+QvED/i/e
WxtYVzQRlZ+5ZxiMhtD7yq4EMIj/VDA5gOc+8FjfiL90MCggBhH++3whHOBjDOzl
JuCmFAeOEN1iz1qhkB/BBWb2RQ/+Pg5Wc6vmT6tzY+nEkj+12VbIqIzPrVZe07o0
59qQQyeL1+lln/rCNZjQevj33jfcRlZZrI69vBzZ3O3YlHOHcCWYFcAYe3v7eEa4
Vj6aUYS1n9h4BhimpqDOUH56/q1NP1k+XEIWkkSdRa9rX7MVPZ/YZF6T3sxt5wGa
3pyjQ8eEn7iUICY3K+wkrj4SiCfWD9mEcGqD3+WgMjjVjFCWSgF4OsZ71eoucGL+
kAuPjv5TRrIoPZKBO6oEYOi+E5010i2Pa9MrR3vTJPYmAjx/W4rVig4rV31XdJpA
7MhE6KIyaO3J1ZrGkPpKwdcCcsPmrXkUfwF7nAJqN3boyjS2hPOjglk4jQfHHI1z
8hvrp7OxPyKKpJiCnZBUDqq029tF1sRt9ASgy1MO7lLQysI1UExAwoOTwA58t3qi
mil0F6EkKCwz/YHMWdGxbx61hFHD7c8BgontjXDxNgFePX1tg4ZFfQ1ZVf9/J1CG
WjZ2L7iw6FIYd3lNHY0P6pZ+eFFziR7fJbwi9GroxL9MI5v5xXy1TqptsALdaVC9
biIAIZS5MIHG5bgwxDpY608ObhHOk3BlMn6FuUgU5oNhhIxxulZxKVI2X0PinXma
YRKc0z+ZQHWLJzCkveESVpxhlrOQ5L83Ni8+6EhQaQKBDsaVxTmzsqERwmQrFb6q
b7TmP/lqDW/Fva+LRD6xAV5ZteUMPDIX4knS3fE/QS2gFUcAg65TNDqNsQmCyJrR
VGHRiXeON//ZpJpWNYaDPPWrlQylBwznqwwRRIKefgPV4MdWHYAWCHd3JvdKvQQb
dv6s+4FXCM97KupOvFTnk1aNteGO1bFkz9qyzBHP2b4/vI1KOfnk7i9Z2XopaVRC
QnczUd89GzZz7kKVGgIERkciiAL0dBEpivVBAWlWCcgGmkM8M3xEYd9Zt1NTWbms
Bp+ZbFl3SYv+WaVqI48uJSKfbDrOJEg8Qrdnuccr+M7iVlFx1WQsUwo5t3b7yYwE
1MGcT4Ajl0Js681MzbJBeYwo3clOXxQ0cNNJJFmsWhT3waDXYOMCCDqA22v2ozqz
tbp8mJGqtrTB8turFnlN1mqmJkLMs+UEOCFNMIc/vZXb1+mfKudcJFP6qDSZCkeq
UYtbE47sV3FhNwNOwMQM4eOFC6sxOXgxHeNR5JympetNJv7GzImxTAatBOtIxNrZ
e0IMnho9A4hTzaOK8Jpw0pAX3rkQvGXQAJ/tyO3Zu7RSpeOamQUYYWs2uniWgmYt
OAkMvdmgdvJhvLTL5SYwvd+mMVW7hL9DA0FQsju3y6xPQmYbY0RgC2beqW8nvyiC
c8g5vFjsBhivEjuxsMg913uFY31aDRPGP/Snnf9r1SAafYovo65aXWCArHx3Zvim
tSV6kFyPq3xcrx9Uw8OkPOZiFq+zd2t+OmHM+nq/Mj/aTnLlwjx6cs0vSl5A2AcI
SL8V6dbF9lZ6TD0mKF8rUThi7Lz7u4LTICEgZ4w3ZD/by+H3UiRGnhNfo+BXBEUA
ioQqA61PUoOP+xkdnlD5YxixdRkResDoblDa/IqeIwGhDt9XzULnYhbbwmd3ZC5Y
/9B8v6o0Jb3d7sKFQdoPNdzqgWIwulsLyzw8cbZ4wXTTuwSuNl0lxBnZxAdVn0z4
zplc88/iJys+PWD0JITk5Oe9GVH6+8HLKA64+Po2qKrY8TNSUo1UUYVOXb4dzjWK
CbuQalyixPM06M+sf9UbV24ve2zYUcoiF8ioU/QN/qtNfoRyih2VzuJstGbxN1WB
0ZcalWs5j9QJwBC5Lm8AnnuXnJuz0v6+IaABSW9oIBW12EFtuhmzzK6EWUNKptLA
9yfaVUSkSTNyI05hDCEO/tPg8sEXPb13yotdFKesR/A8t2rYK+zAoCYjTylKhROL
vT+VfhL11NqJ9i1bnu10f3MvA7+rDyJEU7FjsIo0Qyn2gr99iqbftpbR+V7orMXv
9hhe59xT3dfpeFvLopf4/zAAglwqIMU6QZZew/ql+/yEfO41Yozyb9VkFWspWj22
ZwTXjTs9VqGCpDyP2mCng0zOvVC9Vie4eTF/SbrkRBvgsubsRR9lEqYKvgRNzp9Q
aCCJaXKzdTVCuGSXEWxJIWzmXSeKPjvtdLjoYCdZs5yalEwWXDFfENGEC/VUosyj
g0VN/cihT6JfTby5Ka4IuvfEHlSHkx8uo6e0b41q+dmFxEYXNDsG8G9NDoC84K4l
WYt1wSnNjR4EKqYcHRINKoOqFfJIp/R8ZsV+sp47VHi91c72yv4tVywLlYbl6vFt
8ORJ2DVz8zA5aycMiVAXl/9STdWNTJwjDzRGbYAl70iUlBlpgAOj+sQZSM40oChk
+VyaOhOWK1rwWfARUOctFIpbhfkvSuCv6T3D33Ud/nZmy2/isfhR8mtxJSN4k2OU
WKaBzinw1IAenw1b6vGw0qjqUW6EIbuW5mQKb1LwewWJZF6hgTg/L6XoeTuAwJgg
5c87jjRJ1JdAfkoKwmnmXOrY2Lq3WwPOwbHP6S6WwaiUc7EUkbGsXEJa4GKlovnb
h7H5dArVVIkmKFPF527Mv0FTVrMHFtyP0vVOJKF5stduSe+7QUEgd9fpQqEFjXXe
Zx+9QmOc56PmaQ0ZhQ7UC8Fwkkbp5kZ/DcRpAvakyB3IT8hOCRwvekbpKUYcpiQh
OS1K111s4Ww/x/vnBG32SlFL2MoYWuD2m2vPVbNiLStXHn4uD1QszzojfVfmO0Md
dlrHZ/d8IimnW/71aN/s2Nd2Y6/HPXTHGerxgS90Rj3QGZUbnaXRjKQcgfbgF+Yw
E7Y88RMWho/fYYOyhC7fs6F7NqoCFamG7qaSMafwqICrei9kSWA3mEw181pXCNcI
Ca2GSo5MqYKDNxKBJgs5yEgKE2OJfqFgV4QiS9HiPG5Ex5NYRVoS7C3odRFWCm47
tOIZTA2rcSh9QKbZ9/FnCEHZe0JW/ChChJ0dtlxo8lKx88voUxxIRSohn4EWT3bA
OV/3cErMNZMLfgAsSBI92ixT/OvpudKWhiNYhSVQ3FnRJ0SOn7op8hhuNsAmFhql
vFYzvcffUtSvb9IEKT3aAnDAKQiJ7sdNav8fAuNMsnIbrzzQJkxLvKZcbPtWki5m
/u/PCh40WJQtf5LfsdM32Xy/heokh0awGbPhSl1KCUiM2eviLqD42AERk5MDYpWi
aPS4bV5MMo7tb7B6c4LuLgJ2i55upO5Iv9b24KiX1LkLLz15Z7QAzVW0C1eAMu8Y
/BpPwAhHq29elZLnNP9YQGVTfzcwnqjPYba9//M3df1ylyjqapwjDHxJzPvg5GI0
VEUwdqzKf/YjrZGqxB7Ka3Z6/OEigwfy+p0JGPjfJ8MQAsVrzmCkm9xQqc+yAV0c
r3XgooLlXjqFoHaWnxRgrm8yafHCA2R23zmfUrnKcbwWTHoC7tKvxEPs/Ca6UUTH
q+g7dtyTW2buwYqVo67v4zPe7ta7bvy2RD2aZzpRejIRXYgM8eCqr5Rouk8nDTC5
WxxsFVXxNNW8SOz4x7j9qhMgMyMTmktt3Ap6vHcUxNN28ndqJccCw1A9TDhRo9ZR
f4zucDTlBXGA5Xo3Xi947B+TDaYsMz++VTaob65IqV8aNBzkNhxsDB/SAMQGb3JW
gZepEXoivmMyyUEpogJkPWkAnIfq34T/LCk6N1MUVGhFNG9TaMfW6ZnBgmJ8xvVW
jIawsVcVPCvICy9+PhYYk+TIh9pp6vxfIUB+atnljmYmwGfM4x4OxFPG+6wN1Yme
IUYuKGzHkKibTi4kAM5q88qrdvth3bugplxuEfgi0cqu9BvQKZIs1Rx7TdUR+CmC
DOZSlzbmUaOctE5GwLx84vnXw6IPnOmVprYuZ7iA7CDry5XsmHrGLowW3nSd64yv
au9eFt2rFjWHqIeyqcugCsaRkYfX1DpIfKdFm8t+NlCm0lvJOnUY/zcHOHl9G73A
oj/mhU2ksD6iytaOhUaekufjREVTs6/XtJQyQshdYykcN+RX7SAzum7TNLIBwMuC
MuWf1xjGbaRV1UWBPo75yn7wqHWMbMAbing1P9eZdpZTQ2r2IcPeOQi3/Fe2hpyB
NNBIWKVbB76uA314Qoqs0nLB90f9jsb/bKYMZvuIxU0973wbO93phqhU9WRIVvEx
w2nvv7izn4RIbCzchrzQSL/8y/tEWJTf7J8Ku3iAcjXx4oHy1ucYFo2FPFMyqeVr
i4MKcdjPtM5CCH1EA0PcoPpaCMvItJ/HNoRwA5al/L8eo3qUvvbJnMdc1oqsCiOi
wWPcbf0w5kJwKCOJ7ZtYpaZupCrTWRHNmzuXmElS1Dxq+0iGXPG+L3EaDytFZL8L
OpCPLdyMqHfsNDB2+blRQH9pN/RZytORf5WJCIrZe3dXBdNtHJttcQllFsx1rW6j
5y7D9NUbKE5koVS16vpbGEYD0YhNoxc2DUAoqE8pI0pYdXerQ9IvhOkLqwNiTIjx
AFxzJOoeQyeOMc+ThTLhuBekiZpdse5F3PUzc+F1UByTrlEvmhzz9D5zZwIbR01M
fsD6sehxAdCsz/WedBxOyKmHeW/gSUzXUawyYBhC+7uUff5pfcPx1CrNOTyXo8dg
ptk7wSXTSfC7PWrV7xCwzJXcgwavyVDNBb8kpLmd8wh7Tkk2PT5dw46a/uQHulm+
0jpzy37aqkqaxkNGmy9RuVqPecgbbd2JcU5tqwyNbp5cd3OtaZGuAhBH/0aMYykH
ijfxrTcwEj/3dAbZMUIwfGrnvJCRuaWu9M78/U9T/B21JRchMisYHx2YdZx4uRy9
0BoMLPqrHFSGytyYCqKq/rlu/VcfShCbzCOv3C9GWguMkIFX2PTgw7iiq97BXmKs
HovcKkT0JR6ePqfyPXYLpSqtyp806lQm+IthUw9QiQfnMcDDyMHP9cMhWM5Gi0kJ
Q8i6tn7b7TrKHsNBeaTOcx6hkwX1xm61031FlggYVk8vAr6ZTXK9WwjtONzeTVqV
CgfFngf00EMjWhA0cZ8lZsZrA6ntelxexMp1JVqRvDn8vRvfeoJvDtLwHbA3VOmw
uyBUeZ5wOl6bWNfOR59tpFCfgUOlJcqdQDMbPEn18wynYueEWyVGsajTgA/vFbdq
S4nSm+hIypIATpVeFTR0C7izCjRNGTUDze+nP8gvfvr+/gAHxNiKSUTyieJl/dyX
l8Rt/27z2omfv9aQwfrTGPURUFRLn7e4dm0SroxNVfN7RUbL5DxiyWJiSAxSwzbx
P0fq9iGiP+WbpLHxPLDMuWCFXbnxXphbZtbcNJtLuaFXsFUX7HJ2eO/TWQ7MwS/s
4cZ1JXxqUfHo3IfzBUYuyFIXuKVCEBQyZErZzj4Nc4YC1x5ezJR3O815OklrUT1m
WhNuAgBqo6FwQRcDEa4iLE4ZQVEPiTozIgOGwRCqg7pnfe5F9yYFWi2VAR0RH8Az
ls6ICJacAnM2v337bRb2UFKZkZh+hUYrFL5dE+h5AxX5IG6C/R2FThPHYJnCvKqV
mUOGlEWd6Fy0bn+vlsgosO3GPKaasyvprEafjkejSROkbFBjm2RSsELNJcreqVa4
VFt2DNpCh8eqW0PoKPZ/rfChEBN7HYumgAlorBXPTPLonqw88A9JfxQho//flp3H
PaDe5TIoQTMuwm7orM0bCilzF8Jb7hHaNdftR1HGT8jZVNDE51h52I2CI3z4PkI5
ES6389mkWQTRt9g/z99LT+mgwm2gWgJTwjFDDidb/yk0yJOBE0jW7o0o/U5yBEU1
9pSmUNjNOwVfhSNt9JI2Pm2jVph4gG9zimOyzLu5lHJYXO3575CiuPEIYxaYgV/Y
3yKNTtMkHyznbprl7jGcG8O+yI+UXIcwRP37RBjHJlGVL7TvMm9IQ/3s7UBTuHON
LnP52SnC8FtVUlIdSva8vef39oo88mjC9VWAj85uvdb5QuaDOPx8SB4qhFuJ/ZUR
MDvTRv5365rXRMLoHFoL9BKZ+Fi44dzNydsBHrzrR7cYY6xLHM4DhlLzIbM30jg+
KssG969M5O3rAFTuHl1bY5K2Ao+qYkR4rVE4KT7UByXvFXKfoZdmS8nLx2H5A4Z7
q8tHxL4dKv5Ia2MDOSpcwRvfy0+v02j1MbaRjW9fAuORdzCLEuchvtmoQAhLlFCl
n+ZJ2NEc6Itd41Em3i5CLE2LbMrwUS6yvBEy4adO35FcWsxh08dgPbT1rnWv58uu
D6T18CflwikqdvODmXtj5m81NTxRrnolEkv51hOs36aBM350ebXzll1wWllbVjIS
IoGQdhAcImOU+X1IM1qebVOBl2KUPOD1M9X7vc73ozXQotMMuHojDZvNxBmk2C07
BwMCzZ1Cn2twaMsJehXAQxZtFXI15u9lz9Sl9aY/wGmvGPbFUQkzK0msNQFCqPpr
g0u8ENG6Paplnbxd03myQ4A4AkrC9/I44XgRxxB49vLFgxGJqlWhnFwPAmLiIRSS
Y8Npm0TBIdseJkv9fnm6+Xbn/py9LKd5tLp1nAzhSp5/giTjf0I3XIWV0tsmweda
HFNxm+eJKtE6iQ0MbG9mXDMWKU6WBwPv1yG8hSw50ALDDdadHwn+0CI9nRY9bPev
kL9O6i4GlzDuo8ho83tDEChn8nD4UnAwxzcwlJsOZa4i1zvr8Iq3534yRvPPzycS
Lx3Ssjv7KvLCDvTfbg/HiEnmbxW9wu4UZ2JSt5Y3bTSeAytm5/GIrRn+p2vgkiMG
i2J1NZamqaT10JpWvD78EdmEHFByZsc4V1JHx41iQnqZxEFWyhvO0olgKNDGgr+T
IAncTgGrqZfx4VX1VK+WkpqYfQq3N9jWG+uW9HnLFpdieJ2ZJO0HNd09moRCfPCk
5hx94WpjuyVrwga/K/HjmCxvPAIoGSovqv3/SeqxKH+biQSZZ99UgMUHo6kvLX9a
vfziE+cJHgTJmVfVCcpwKvGGDLRtk4tx/4/dJUOrxMX3W2UBJxpqYVdMz4H1YDaP
3MLn09WB6t8oQLgxIFM8OBRqYmLm5F+szIEIA4RcO27c5kfe73eFglV1dTDNXIXy
PZ7lGk/C/vty7vUk80iVjbUCKCZXPKOexEi+WpoP28CAjNMyOh4uVyon9OUZJ+x9
lUwwHO+2wTIOd3XygTpp/ak6DlO9jGaN7TfTVwDg5NAbNXSqOp8aYN2lYl/y0FxY
28yT7bfWRj/Or5o64TiSBf2sa065n5ryv8jhTH9FDyl9Oq21PIoQ+DsGvWNTBwTu
6YzQBD8aV88zC/ZrCLLGmIaxXzvX3gT48x5HIdsl6E5Ckh/eBi5JNENh6vs7E9pj
YBzK5nBJbQ6OtXApgUOXK8Z6qvHjnH72RCxoayrxx0/m81ACV+UNx2LttSslTzwf
WF9jvaKu705ci2d3fCdg+n53WYrYUY7z5Z5/911pu//y0D4Mgwg00QmEFlNNirD/
Bc3bAk3VpbIgP1W2WcH3FNKcGmEhsIZk5RKG1mM+CEz8nEGY/bXlNmoC0JMzEA+n
YY3SP3bfU5AbGx4HvJK0L0J9Jz9bjEkmiu2DPsHX0xBHpTvQJahJ9ox09fa86Pd0
cck67sktOmXr2tPop0lJ1wVzvXn4GxO8/rbhSaU9OpCTGft9QWGatMcWogmG1/H8
LZNFX1A/Ns3U1pJmJzvkienLkp2ltYsOnxVev6JML1p4degXOiKz5ssgLBj8c7/s
mwy2FZNQtzClIYuLDJRoBRf4E9ikE/4TRewbcpecum1yiSo7gNOmwFoGfu/udK5A
caCuMPPiohE6sFr0QWEfQhMJXeDa1GHz6Q8ogje9cxGO8exEiZkAG0s2jyaP1C8U
PKqxcHN3hrj0leZMsKZxfSYXJBoR+LEjTf+10Xmju+bC/6T9B0zHqVidATOksx1+
R+bpweO0k5ns2/EITZg7xD7m1mrNkkzn6UtF/uVvlWeNH/mEDpF1c/oxtfWFoGwE
bWg4Bn0dPg1WEASbaQVERomVkFJK+f6HU+01LgHaxFcwFB3XNgHMaskM1fBpBAZ8
K1FY4j86joFX6xivzyJZPuXI+XKtRgzxOAUAAhy5w+7EB6rjBiBXZrFsBwT4OZKz
2+ME0FkexHY7f+f2KoDmpabgpNko2tWJ13rF/6Z+lEpOdSjICsBcsf8XE9p2XF7H
h90MQg9RAHOcNG5QRJOYU/OdC77B8v1GhEsVo5baJyPCy1UeeoiECsh3s2sq02qs
MKYltOQ4PVAnMrrfMmPF5L64lnCcBfgyXAAguOOtGnBsj4s443CLN6qkwqaVC6xW
WpD5evPbIIhApTYdltWdM4Cr2DYxJlSM0D7i0INCOm36RdIOqiWg0lTuzyRHP8v3
n332ElNaNVvtm86Dzd/Zb2G8zpC4MT5Erie+zXmZwbKbnh9AXSUezAtXbClW1T7x
Hv+6jzBceqxIDzscubYsxS3itVVnTweIbeG42wy/uHfmgwtpPvKR9XpgHUiN5XdW
FnQin1kOz/Q0BEm7otjGcCwaJE6JUx6YTFqiAEqjzaaDXQmuvdqtEAOrHVWiAOau
D1WlIQcxSInY4KfxBNp6ynMuVEI5igwoIR8lC+xWp0usMR1K68uBtyInAj546lf3
YMP23Bpn5ihiGvqX7ZDPHfv7i3CQds+GaDP5u/0x/pPLTHgmQQRGBO7+ylW/9bOA
uRs+c1XinWOmqDOl+35mW8IfovIlDkiInVtuFoE1KF/UyqM1tBAsRV8eMOdU9+Up
rvxRMAcjnJAhB5QH6IPF088/FginxBNk6Ip94aFeKzFfjKefpqznCj+cTG+WPSs9
gPJxUMpTP30w5+VdLl1u+b8azjhNXnvnWTZYOfwVsziDJidiyhtV0024x+OkGPTl
LaN2dDHr5jUQ3Hdq9TpgaeeuK4wcxpfSmgjV0fVxqACvJGc40y9teR+XrbR0FDn6
XCM5uZpcNIhXCaFXhayfC6xe6749NcqRFlruqVL+ysl7GSB9hbTAkjL/wis/9BPU
h53sULso0s3rop+MLSMsg4G/r/p125NB0NG7MHBm6LF6hy8IgYLewoEiNUCwwDRZ
FYvLOdGNz4k60ldbSxF7Pu4v03qs5w9JpL/9udrPfUOZhKrasgRktUKBOfSoWXAd
uzNjzAbPZHbqIy+7L2W9Yqm7GhdwxGyq/vZM4bLMazczweOqy8+CuDCHgqQvgHio
saIflQWS/Sb0+2mQ6ceRuzwCON15D6LDx6gls0fw+zEA594sqRvHuTXg82TedeUx
i8Dw9JLOOdcIA2MkvuoBPN56U/EosSg+r2/KAClxUrNyjF3YdMGhUvwa33ZeJrpK
OBnW2niPTTjxG1AA8v/PhatOQ/e+jd/xa8IwcPxGS8KOn5kjBFUHlPNb6uxOamal
NqEpqPbb0gmc9ByS4wcR5hAAkyzdKcgvoT7EQQL2nGp2X2Fx9uz5eHM8MhfzsyoU
MGRy9kOV5Fla6mODmMxMlBXRj2gGsfL7bzF2STQaHa4oL15HEU7fNVNQFm8bGRJO
5oWR4lBh+s8P+KhesoCiXVXKozt+lh0bdtblZ7S/4tbtxYr2ZEqP28NwLy2SydUx
lN8TdKHV2znTSPdIBddA7lO3YOBbjKEqYvr+AbbbAiKexaaPlFutyQjn1xmxAvsw
PUbZEBmhvCYcy65rxdb4nVRGurHwabAqQv1FbGthv0+kylOS6HT5wzsI4T8x0YX1
PIulrcUOG47+8dCGmNyWjB3CQ66tnsQXcTDsb6DMdxvVSpFPmOe3Ny86I9btLjH/
oSGUOvol/2OXgOW+FInkAe9MrZ0g0rK9TqwZBj5LAnPdR8A4Exx24dBv4ua5t37V
M8zbHOWgb5PwC4DQvDv9e4MPS+ijgb2+hASCnm+c85KgZ1YB8Mvfu9V0FX0nZcsL
PJiGrnaWXDuNtyiKANOvohESgQX6Pb4rXnRRJ1VXsxn5eEceZecTtohtII3gZqVG
iVEozkYKYCaYbFhtpt4+PhcRZUCIcIIbueQO3PxXYmipdqTkZtDXdIe1pcB5QAUZ
XfVgigX6wTs07kSepsSYxhOWfFwoeJlWGd0L9ea/Op8BcINibO6meYL4ySKj/uiJ
w+Y5KxdOCHgxgax0mdVK6kH3p3vhlj5+s9b0C1C4xUP0HuFka5ys+z0mc1MgKZZD
2g785JLPc9N/JQNM5Pbi7UrHFsq5t2WISAzWPucklcmZetJRYwCES41Zc1zZy6DY
0KDAfuJcy2bWv6QPfcwojv614Gm06MAQxp5wMb5554M58zDJhwNZS40i3gmnrH93
Hy7Y2rtu4G77KSwNnTb7LkNqHnxtCA9IUYLiu3En8C5DDCkOZRndf21XfyEJkq4V
+2J0MHvs3EhBaCYWu+u9VLF0wkEr3r63d78PkNHn/l4+4Rw3quwUMqe5yDi8Uved
452YNvxInTcTz6XUm7slIT7YGiClp0J83UMYYTeLvzVN38MuCZqjFB20lvcu8/62
DkXVBcHx4lveiGKwHxqTIBT38Q1xSSrvoniZkuIAGlrlXDe9KOhUPg3JfymRSov7
uqpjYPu4vA+ISQg4RUaio4hbuv/h1BsbiD/DuEHtoMDq/cG51vcd2yhKSLyzG/Tq
74bKMJu13RHkgxwDoM2WRQI00gFddP/umpazdfSM8PyRoaIkInckYAJCL/01jGBu
iePqSzInuTsPq/hZdROHWQtgQaagSLEdbCQXaRagwTgai9EFubYQdeyX8CnOAyHR
/VgsXHu3+0KybOojwlTxaNPzanxediMDdddsQbJECrWGYsccmJGuK2S343FbD6A4
+HFRCuEu3zpt64chzEoF4ajzfbtqVzmzJNHVmBCXJwDN4c/eTLVX9KFuDwAYjD1k
0vQQEz1c58MRto66XOG6dlhYVcF17K19DwSuoxAQvZn9y/3sv0zOIUWe9Sq1+1us
CWrdZLJPkiUGtOdAJXQZMMjwa0DEtlkT2GOIk9j0KAzoyC1g6GG1svO/bP4upgZb
THeI0cJRpBqrNC8FJ7o4rCjcOzG9kzdCGpi60Htz87kf2Zm/VCqAUVvczIqLr1xw
/COeD9UvPIY379khjB9rSByXVeOmNIgzYayb88cvY7w9Xs+qHDZcVUhjMyOCbRix
YroElAdfvkxtIHqEDXkLM5AJp4e8YsbRjGqOAXDZB0gl5OeAJoglYqA8PzglljkY
IwKjrp+LFdx9hO9LIWbA3DGvn140ra7Gi2gHfzW6BAP2ANKpGPJfsOGJQToRYoC+
XgQHLeWrP+PA8y/JhN1gAvUN+Hr2Wd2LFoKHd0E4jURA7aw+cf2htSNLBGrwyHuK
DPlvVG1mEnvPc4TuoKBg7ilymyFUBmMEa1/OyDx+/yEWf+N+IPxGYI3tdbMc+QB5
5ctqWaHlVi3IJhjlVCWlZVqHHzi/3G51FGWTAQiFJpTmFs/Szq8QPU6z+YSeBmAh
hnJ7qqkNRuHScsVqRppnqnizsxJs7PcvR8yxW415RPv2FTlkm1PeQdjbDGccHXDT
r9YjhtAcQ5YYrS4kDhAC9K7SFu6DM4iLJdSm72QijOEQlfSUhjMH1GtZuGoUWs+o
S1Fqumr8h2XBBP+4EMuxS98EUGXovBVI0XfnoagQ1vQ5Kj1mZr4NZAo/UkbXc3cX
LEsxLt0IQi4NDNKimJge7mAZzDRPRE4+rOpGXPesmxc23YNKssqTOgNq1nWfWYNI
TyIgBaz0BecuwkOXXMf4MSHuTD7BGzUV6Ay78l8ooYtRVB4WQVQiBAW8/byP5kzp
QdN6P7L0O4CnZKH4EO18PGzSL4gD3+RSbJuQfTeSxqdw8nFBpOdtb/3rESL46ff2
WtCijaZpZNAyLCSO0dcgJVhmuXkCBoRB/X0aa1sn/rsW7A3NmwEZd/2gYxEs4NP1
i3Dq9JncgKeZ2fXWE0H3JQl+gyNGIVVtODLw9z5uO1DWQ18Ic2ehxoiTXczfIJ/h
S2IANEP/RAl7wA+f4F0u2knLnvYRUAH60TEe14RXzVWmVVwvK+kNUVnKPy91BXfW
pwF5ZjIUNoud0deCoCy7v+q5/2aVL+1vjDTgF/NEWxI/UaGysX1Sg8+hUZGzV0jc
/w5Acm1VyrjGjuNsM/AmqEWIGhx9ucxDxiCOI7hek2e6+hau2NUJHnvUwd14KQ5F
Cva7gW/Ioj5jGMEXCY2Bt30YGwothXqQwFjc+hAEyaQOqcbXGHd7RRLh0eBmjzJS
oUQ6kCZokt4PkEWmYo/LPbsNwQXKaf8vPb4VVjm1kR+NTU1a0I3btr1ee1BBznt0
QquWQYxkq10v6n8QgFa5hGc1Yrr2fuot2eHlYo/79asPnhOJBvwpQad6BOQRkSxA
f3RzO5ZOZu63hM/+IYmNeJgumEYSRa5x2i+3YmkcGFUJnjzpppNyC/I29sYmiwCs
Bfei9WmTTRjEGBCoGQBlcPSING4hMBymP/+3zg7DIejPccbeKeWgJAhZugzeo68w
YVZgxYlFmxwVDI1qPoNZ0eQXAwHCHw3uqzGPrJC3TXlbiteQ2Lk8KsiIrc1UnUGu
hFYey71aDlEKjZdMw2R48ISHhcGTuwMFLOOhrln1+fZiDyZ2/9B3jifJZXXJi2FP
UC24aBWinIHypyIoAXuSl7IdHUlbkeEZIp156PuQwvXl32NcbLUQv03TZo4g996P
yGbr9bwp1ORcloC/dZGG0iX96nMD1312mHVvw+4hiHf1pG95wvN3rB4Xxoskylbt
BpKIxNpwsXrV4GDWgfprY85Kf5BfFF0Zh920rfAhcbHCueh5TcIeLkoX5xftIiEQ
2kNEZe6OeuR2EnlqOkAUmQ8Vl33T4yUrXm2JvZC2tGKh9/7EOfYwB6QbaHYyNlZC
JgW3MdmUBd9Y63yTJNVazN8aoVnpxF3jY/6/3TI6GjdyKK2S5C1yh2u1sspzEETd
qavRxCFV75uD6EKTFlneR2qx6TtlaseLBvhyPXLcFQmhW9jsw1IEY0XbErt/r4eE
S8FXp9QjTmrG8CF5/Ei8dFG7Wjqj8prbz5dcVXmwMeOy2PySdPLlVyafxaDw/leZ
ghUyhmiSNaXg/Usua3lpezlp5Wg8LRn3av4aaLJiaJf14qSeBDHY1UxwPgm585aw
6abKSmTmG2JI0mJGGpuX6MICIGyzLtJ1HkoPy+Qmc2OqM0OLXLAABnYQh97CtwvG
Xd9ul5AiTO5flQEOPQ9wVQs/mITfbqCK2IImKXxL4IEdu0LIv+LoZC0Nz52Ihe9e
j6yabpvDbJzeclszv1HbKejI1iFWsBTs5cg4+1zrZ95GvliT1e85NevGPMNnCzlS
gb0KGawilBvCxRfLihebkaw2dSLpEA8JN1ggVXkGXvMx/1/YayakIlVUOqsnBW6Y
HZNPFvPPAuvMYjf7pyGkXyx0HfT2/KAX291KgnuZxZXxwPnnTn0HlbgvW1YhdAHg
3/P7MXC5NCg8uW/bHmiGDz/8LKB9HS3CyvaDu376rljlpUWw73WabIZpN+DQE+2S
LzDE8cZpyfHa47APnRKf6st3J8UEq0EX3pmWTnnMIq+FqWPwL77fkA73m1wlncyT
YdyjQCJdSkPLAtwmHZ4vUMTIGAsAMoprbyHKJUfZb2coY4ntkXYUiszPvUUcgTJp
9HpLJb5EdxC3LabnOHdY6inQkpz2zrsgcz+pCC3Y41sLl3ZJL2zS6f6Jct0pr1Cz
AVkryHMgKy3BvoPTJFEwnO2F90rA00+VhxXCDBswbZCb+yOTrXjiqkChloe2ceEA
APaEXFgk77qS20jOZZw1ugeODEicgbKZ9ROQ1fVMkNg6k21hZ0kDC2lDELHZ9d+N
eMIUYUZL0bKX1yZVAtvnE7QlAi36pVy4mRstO0ogvzte00PDc5RBOb3txUWizUfP
MgUVfH1hqRsE4Vg7g27YiX/P4uYvD5aowcXYJYADv584rKNMme9BFr/ZAYdXtEzq
HXcq2m0dAr0Jee9936WpFtCBd6sv+r++S02eFO5EbcgJf3fSYCMejOHUPbTMVdPx
fcUn60D9zYydoz1DMtHLAjuWsjj404hVaC0HrhjkS756LQRLOV1Y8Z6P18lx1b2O
WE4uweWZYvmzRdRcEDnKN0l/CEN9/Ox+HOT3F8HVHi9Twg/x8JLfmYa+RUF8+xfd
6SWJc2rxdswLkeZnoMpolk+bPki6EGOdxQl0cqjZkpp7IOMLFwVWh9u6CM7nGiOM
dbzf19VkVofCzxwV9oN0RB+n1TlD+JY3ICy4VphmF4iQLFKux3VAObkKVsuZT6fM
r4Tag2RiMxxGjW9Dmgp/WIS/7widRVQVUzskfE//M2KOMwkQoWgSqz2EsBox8pVd
Ih/zzMVqw0YV0LTk0yaFLCgBt4PGT3nSmh1qv3mQcvbJNO7ZmXIAfPy7P3zje+p6
Fro3w9JPbQhGu4kq3U1t637eCN76rAoSDC0KaGsYYlxuQ0lwmYLVwcE1OFktwisS
t8WEDqoW6BEz+JSH7wtCWWmrnY7TJdfcTJdUzshHtxF5cfdY7WSTP5ktQyV+4qA/
5xAYnhb0Z2rRm4Bhbw0PTLaP8mrgjcNHm+N19x9lTB32j8aY/hgEe42BIbTPj+Qq
FtTUZHa7ke3BC/VuXEZRS7nOiOiBL3zZf6pigPOM3mIxmbWnR99V+txIgdxzQYWq
jGCBh0pvfLQGWMw7Ds5dAutBxV/HnYRpNBX/GzIvi4Z3LuCKRvr1zPDeJ4Sj2vJ9
x0RnBn04l48akyxtwARG6sarkxaBCdt18oBtRQ5p4R1BY/dpWoF7YVUexY+3Tb5I
iS+pI4d/2YAXc2sI7oGZcNY27F1FdzVH/fXGEVzpiLjNmN8d50SltEnWEAX/zYMG
o7EJ6RBT5Iz81Ux8elzHHcDd81WtdRYnzeaoU4FjfbSxXSp1HWiXNIcF3PZB4LAP
uE9oGld2aOl/AAm7xybDNuph81/MW9H6acRtDWQPJzcJ+Vzo6xLl7k/FTiNViJaj
xXzz05NCDwFvWBBNIbRujSwBNu8erhLqMDV7wKXUh2f0tRqxR2tSSjEe+rjHHGub
CvAcgXTB2sAaGX2PP4xsOl2C8OEjQzIjjBOghlyPGraKay8kwow/eOII3tG/fUM0
Hep5BzAMtG9su8nPG7CdaIdpZVpyUvMixGQH/pYJHiLFhacZ5IPyD16CuemtumDe
SS04cdqIVTrN8FJUo7h37Q19XDHx5HC/VQI0B02JLzRb/SYNdAq+RQ/I4dQKM92n
Ok9eVyunxqK47r1ImYzyifofqaqyrAH/BiLV7U7I0SCA6TyK7VKo2J0PACUQ2ySK
LMRJ9RB6gPMQpOJDigKuQ6Q3G2nCiVDlfp2p/mt2iD3wNoprDfq83eP9j2rnoA1A
nkOqAsSphBkGVuziCkSaaG40WCqTvF1HrD2oaIcu7u4QdXBfRKWzCTY8d7bIZLgI
BC1LN3bFWhEVZqNKH/Xnjl25N4AA9fEurlQmvMfRI1dL9Q9dHrdqQycRSJsppzB0
NLr7dscbf2cyyrZE3+pRQ407XSZcKMJ8sqFfxZJmUKZkC6uocPNScLPgWyW6dyT5
9b2Ho/Q2Ysbsst+6H+h7uL+cz42OpfKW0++yNwYyKEpAoXw84mzxe6vdZL/u7yQ2
lGJZw9OE75H37VYGG/fJ2Tpy3fbSmQ04LKnzspME9A+DJaujT6OR/dNsQE8QE/60
lqzHfhRxh2bQ8cPExlaFq9p8B5tOKd/ASTaNBqjKR/OpsQpkEGPixdz9FXQNXt0S
mNHnGecGRTdjR2MooeUNqqeP7iC90qX5LZFpIdSPwgMjGjWxq7ezvXQ6P9AE1vL2
i4At2DEMHw4et3KhXcB/Ml0uS2+/TkWpTuvXeNAjjc3H1myD43C4mKb6JIKesHy6
PpvvUPJCujesE1h/HX2n9SnrkuHtp07RuT4ZhLqv9btC+DiA7nuXtrE+JPIBqaVA
64LXdIzlrt5kBtMaHugrA3RKmtWt49knmM405cLH9WO7W2BaLVXeb053TJpWDTJr
bIL70Ynx1reoLk+3+YAdu3wiAVyyYT/nw10kM8A44a/2n2smmutzQIEGpiXUzWp8
FfmCDaVZhhYdI0upHMNTl2IcNCf256DcYZ32+krNtXazy09guhOp7UWfkug5V5to
Y/d8kLyEY0w4+MXOiUoGfiU/EqIS+1PwfamsMiq1oVF9rvlRuDuI3n4i/svc7saq
U4qWudFQ0U7ijc+LUxl3DvADxK73KvIKkoIqkaVkVHyv5lWCti//YO13AuqR354a
4mM1lVkEIr1iUxf5ZMin8NcRnML6id6Shm4RwX++hKvDK9ZnwPrzzDAf70c9h+p6
sX4Aq2l/JNIslQAZq+YRhjUhQsU+9SQOBOBUw8pXBIUauP23co3ZHcoAQ/Sz6zUm
B+2oV773sLLfDxHibdR8zqTWaPRboIBejylSzBF+n+LSf7EzKRlW3g7IsYwgQ0sG
4ao7jnU/sfj9AdHAMHXb3Ut0URg9uBZGJS/p7jFyoGE1NgKKJd2ZfCguVfi2S4Ju
NfM9VtNgqaO4aLHm7ITN2t6R+pAnetsL+uri1czZGLbOSo/5TTKlxsIsBJS0TfDA
vVdmEkZvGj1ka6j1JwA4bi0g95GkHimrr5ogVgm8C0Ah2A6C+R9vtpoyoz7HkG0v
lSk+AHVOmO9Rp74r4rNRHeC+mht2f5f/Xt7qLsDrAJyNRph2H/qepCGBI06DcpDt
xey+Q/Q/0oYolpJ8lUu9HkPkePDveFAYV50O5P1Ut8yR8WG9Kgrr2cMCBiny1OlB
zcnbNuAXve9QsB4lLqeh5tCaIsmnc9fuCOTd9PUDzrE7yPAZSDL/j9vJRFaC2EDG
SJPxuPOkzXLjwwd26YmPKXUd5YiSjqBz1jfhbGRkRzneO7jMJP8bcXZhFpkk4Jdy
je2thFrTzRnCyIQ22mbIc+6I9OtC9As+v/iBLCcXenyGzAH5X3AWu8mUGRLAGE+v
Em8o3vrdxUlcsVow0VAnMl1rjmGUhHpWAHkIEEYF3+RoiQ9j6+jtRVsgzzUaGH4a
O+oka0xi5cc8NGaf1RKQKyTtdxuDFy4wXM8zUadwMUXN/F/I9Cbq9yzsluUg3OnX
fJB+cD4NzwYAt3orO0oXUVa1f3a86Qb9dlvNjUiW+cGlpbuhu/pyBvCs9QXT2xV+
HqrPMhLIZuSlfmH6RMRV3hok2FG2v1RtMcfhKOnwhPbjIigPIhR/Fd3/nXGG5bwZ
SCgQk5MVQXvu5xcrD5mQ1vZM5e+LJpZycpO8h0V8M3jjV+0mDv/hqcOg4Tdlvtfw
Es8CQVb5dPvwlOZtU86m2ISTPeJRjPgk042wcAlWIMllp3/qA7+mApZQGg/ts9NT
x0ZZW4jXvaSWXqfAeRDWpoSlXWSLIIZgMmuyPZ24LhUMjAisHYWpwXxkr9Ko5/Ga
lVdLLq7DeOYJLvqTXfGOEY9p6HmGtKpvTa5KwVlDJ97LJpnHLi1R3QIUu2xWsWia
ARmerAceD7P4qqGh8BTF72jpJ2Tz+89yrs7493ppsiwUwhcd/DkmgylUIOpzA1C0
avjeZyWgtjrZ8AgPWnTcx3Nfy7BL88beYlJ1r01mu7UAr9diazZ/W9BW/OYLRmyg
OoQSqNvEE98nUZnx6nLihqmuEF4cCuBXSoQHpUfQxf47N1xUb89xAeHKpf/Byc5c
iulXVofeEK0kZUWGdneS7hc+I0UNyBzIDqu0wC+Me5/7l/ain1YDQUtnQVSV3XwR
YbZ0SXWcHWS1lEhaqHlEMvCt9g6ksawgt0toH+/5yX+Wq07SrZ4FpPGM0zEIRZzc
fjRKnVYh8BK7IQCLNAk6Fj4kI4rc1F+BhJYInnNvePFUXgivmbUHJvmS+6j/ySb2
RrWrWIOHGTzuM9Kh4+1YypPxYkyrZsV4bjBnqi8+2YpTD+2bD50UG40q5bI9yIK6
LN0mb4ehybeXgORUO7d9uZbTvxvZnHn9LyRsaEJxmjLsRs4eKPKQA+R6tCvzh4MS
R9agTG4Ustip5OaRZxHaS49PAILfxEzLA76udLqljgJaiZttcvsIYe15ruJZyM7r
tv/oixh63+PEQY+IirnnjucBNiPLFVuJIJ1Ltz5SFUapKTvsiWazpGP+XsYHWCun
ZjMbj+8rkgTTzhpzh1fMoW16AUl4KJ2V3goKRpwSX8LKZdEo81puN0BPVkVl4kge
jfMef8ptPHrj8VwNIW7s9RrYeM9lPPt0GyeooefAwIkhOxlhqZ8kXQrQbFSDik7s
Sy+KgIF8lgpxtt3wNbk5XMo8SELyJOx5M64BT82RiqJcCjgNcxwCH82XxWjjVZK6
XlMWKj5h4bgr9Z8VoKdRldo1jR260dPjgys9AF8MvsyDVgCOWtEf7bA+B0QYmWsl
bkzU8tzHSLgaG/sbBwMdD8fUsxAhuy2B43FpBFzxuOUEj9Gvg+KqJ/4Cy1N8zt6e
9MpNx6TvmLLeYVwEgAlIJy+W/gM5UY25G1qqKiG/MiJ+AC3849TEm7k2JeExAkZX
I//bnzVRPDRNbntMfJ91tJWPzIzsgENKzVMS2cEXUt7rTYNvoS5F1hJvGDquEKaX
XRdMEgReCFtsnz0CPhGk0VFjgBK/ffD5gri5ooqrEAQYAZUTY+AR0m25IjvhPPfE
qZ4uXefJtB0TQ3LqyCJYZoeYxum7UANii4P+4rvB0hLISWtRczvfybkeShjurR14
r48tFmSH8TpqWBKwWlaOitxVOM9e4o8mHVMquz7aMulqYX4oLJltUyxhviDNY1kD
noNFLjnJf47hls5tmXYGYp9Yb+v33DNwwX4KzXhf8xsHrDee/QSIVgNq8PInS14Y
ibllbxWgk/ouEs3+jvBhcEOSUaxGp7L0kZ8PpkkXu35ol4FTALmTWQ8wXJXxXjIo
Nh/0g3+awdsodZZCiOMIDFEFEWz3Jup1VlsTjMt1OfArYtTkHMjob8CbiHIc1djj
WYsi26ZVeOW4hRseYQYc6uXpvi67yNTnKG4ihXfYndUQaaJRqyzTsDF7zXib8jkS
GaPYcrchGErJrbvSWkWcpAlh/RJ1Pnmm/HBS58Qf3hPeCcWxSuSWaXY27gIr0nO7
grJVV98P3hVV8rQRJtmjzmZ3eTcpHchDtKG4BX8j7Ro/CsrSs8INhoNS9ALxILpT
9rToPFXec6whkBHcSpaPS2qmwwzauofdDrfM9Zdz8y/IRDuT2Gftga+cljKKUi5i
25rIkNaSwnr7aGopXs5Ymr571Xm1wKz/38FKvdJYIOyP6NFK9xyFRzLYY1NCjCe3
fDXW/aEDThLRevXwbDtDkcB0VYGJDHxC3enbQAgy17Hn8z379D+R+Oq/7x8I9GJr
AwIg35TGg6OiBYUhR8/Tc0QUnCo5f/YZvPwQPLzYng+4vpW16knvf2Z5FPJTvUtj
xMt52ajjB0SOJWPyFCR8gJegyamxlCQT7MkjR2Hyj0XL9sXdu7NZUPSZRfRHq/cg
3o8nyb9Nc7dFSJyvZq8P7Y1/C/8cbh/DignvYUEszR38Kg68Lul8+wQaxB2fqON4
/hzcyygmlXIvVkF81y9axeOD4GDmj2yZJv2XJPjuwsy2FfSHiSQJtlDONoRE5OHz
RK1M0yAHg1TVke3XfpjCaqDKm679At6khyhNj2XZlPd6LwJhAkXkrLGacRV2IGw1
6MD6ND2ND+Z/kSPjDzj2w1KdQ6ak0rzafrBYrpDj3fX+F2zMpzXxudgX+Z0mSARL
KOzdCpKHeVhOTVnWbVDNy8sMjXvHi1II68Wd3VWGkcbHY7W4nAoconcxOn4osDj9
gba59ST/DfecCURvQgweT4dhi5YxUjhWcSfO8yGiOnCKvLfCvfGlpJdgvdu9fWV1
MCcWw2F6bx6hH75v+Huj6eLHiAW57Fk7tLrz2SP+qNtMJRJ7wzSMUgFel4K+ZK6G
2llgX4B/O+r4LigHsLbX2NOo1T+Tq/O1UlCeMcI84i4mo3YJLG0C1ksFwQ2k9QuP
zK7/f7mpLeVUusBYEUz3vhLByM6BYFEiWH0j+NKckTHlWRXPg0v9zfmDFqYVjQPs
hF6tWWgBj/YqWW5HgrnUJgI0PbKkuh21+1Y+QO5BPGtGm/U4aR9RAXeIfPJh2jTA
HMJwNdB6MQnRivAb1L7/ZQK9Zu7xBrb1TV48DUWMxo9VEZl1G0YWH4uPSB73taeW
lh3wWRylE+B+ie9zMkG/Vwgzfdp0eyNxwJCoD3DbWm7Z0WPSf70BQ3wiByWSjBkM
dqi5M2Lgi/6+lQBc1XlN3X/p1i4rA3hMeGZqTS3z2W96HR5X3mbzCxVPnjIrx91P
1CL7bMAwMtx1JhdtxEhZ3PG9MF47DUeLNmXNzO9FO6waOS2rXN4Lr+mR88SrtGEE
f/MM1Y84pG7BmRNZBTg7AqXhQyq+cnVvrSwiu/fmhjVfacaiywn6XmYHr9JKUfbw
M2xAt3qZpFUeeLfGU37CAfGHk6PcUDN/eyHS94RstPcyCL9b0yCu3hkAjxkcfumY
FmL1wUJSVQyVvsuAxqzsVfjDobZBS98nLDVuSNd8//QMzKal22iQGpLSR8fHwa+X
tyF45574H4xXSPEDiMTFxTblgvFiengRpouW+UJCr8MIVJN1MJEawaHFqidBzYN8
oqApW0Ip77GXKta0282w0ITWiHoYwI/gzHSj/upRe5LNwlGRjCUw/j0Q1BqhYKRz
I+9FFWo8AKi9vaIYgaDViDU3IHog/jtHn9SW0YoYRr2DaICaGrgp/u+z02LqiGU2
n/7esy5kNkI2uBRHRLI6fqgrYtfTHHox+wvmbUPAAzL/5FYOf083hrPzjBH/f1vZ
cPSAUL+G5ZFQ7j0SN94mJbk7/TTaw6axgfqU20RMmGoI3fwJENVQcVChyTeIVJ9h
J6sgzhOOrEmLtEGqrrRl19kjMcBcf8StJFaL1BSBP8Ahr548/1SGiSzG9OlMJZZM
s4wdDl15wwfunVW7LzrBVbimKGHPkYPd0l097Md8ejnek27n6WzVydOESSIVjRFG
rinAHe01feTzsIAN4wFXrlm3Drm+71K72kaUV5vYrNg9dy9biKNGwe6rBYUZb15n
5Umh0HGeHVDGQid/0YNZ5sSZvE2pAwp2r3KaQfKVRPriozw+CxwrgOSbaxezsFnz
TW5b/iqiEnmNshZUVrJNnIUAvXjum/xeewWcoA9sDHrUwLgSvyeXlXzwx9wi1HmZ
8GnzFG2wK2VneQs4A7rH8W3QzsmyqAuOtXUAVyIO1zGQtga9XEk6OI2JgTtsbxQl
R+OZqcRwAnB+QITvhRDfSrKlV9h2frZFziKYGmJrAMo1XX1uJEM4+5invb8Pyq59
ZM7foB33NLpA1p7xn52IyHPncHWxfGspQREEdTA27wEWiOXIEcagsKxY2Gl07rty
flDwI7cHGU2xdrhgLNFY/n3pnt/BeGi5F0gkCYXphqC6mFEPSmro3cmgV+P8Rpwc
5vQXVgcaWRLK9yND+aHBOaWkETiNO0M65GFCS9MGsVZwQ2mNeh8H8tkBzJSvDXg/
lDBaeHthVd44qheJWtuNgPPqsj2U48y2EDcoJ61IzZm0eZILqeJrBgtQnanil9zQ
/tw7rvOlAIVFIgpmFoMhgEflzMYNRzZ5iVLHBl5qx8ciCqlwvmnPcGMnQNvZz5+J
U10UQrGb4qbrxJGnR1zUeRpKGUxVlvJzPxANvkSwic+erkRizfnDHDvW9B6GSQFZ
CJfiOQjQaeqYvmFPE2c/9ti0SYB1LaaEg6tyAQh9C2eWWj0PnO8d2x0MAr1QD2Dy
yYEtoQnBIyxZBDyDCYGOeGsGRVCYj9K4HR/teY4RK9+Xd00kdMAjji20W1v9T1rz
iU830ndESfTO+bnRejq+bBMMKJGQcN0fNCmMiQzmy9xPwzt0KHnMRJqFNOwqAUDU
ELUhXRwTTdEqzxh1OUSTN8FWM5OFE13ArTghwKD5MUVZOP7Rf5x1h14MjE02NiIk
5PmItHnhPCaLeWOj6CwgW/i2HKomO54XtD205X+NPxNs0l4AFhg7QEWvqezx3LQV
JzaL3hOFzX9a0xcmIBvRe7NkuYUUA/z8Mnb8aZdOJymEbxkOILajQMc/x1BHpJT1
o8xnzTxowDxkiaEel9NO/mjppsLoeu5wo7t+OV19LBdaGuBzlCd8zTgxb8nZrA7z
IXdjnoYINU2pUAJSngj8jJ2+Z2Mpv/8GDwLvaN1NVf3ilefdvkhanT7K/pUDfpaD
6T2yci5j8ZSY/7e3NuJv6FNl1Lze7RRjqvInhn0oXPJTMrjK+zVwe41F0gV39vwH
YVYMy27opsh4xqG2CY1/UxFXN3Ta43DEljOGlF1SyzXYemi1RT4xFfJbWpS7G3T7
6VGHF/kTyTTERyUlGG9dcbsxy6GK/sQHqItcwv7GpwZghX//zmZLVh6RZSY19C8k
2QmTazWN4PHOLBywTnkxbW1fm4CUBC1fwBeK1n3P9Yevw6ksvArFtGR6o/fRRQJx
lXsrnpkZ79gNEo8pRAOXu1R/L9rssSIeLCdxf3rPxAh4jrhTUcymD8sHMAwEam0Y
E2tlSJYybNoA7t5dmMtzvBpmRgrc8PMRYaL23lHkZOB+55iTVaYSj0m2cOHbsMQu
NGZsbXf3RXjcswtfzTkbC+HHz3tJzfu2pmu8IX2NVBLW58tX28mHLFfQ5pCrBVKl
AbLvM8Y0Kk1GEJ+xZ8dEwmxOrUFE/lbaSEsaxO4m8E1yrpZgr6Gu9UzRgNokmgJ0
xfA3lGhq2C2kgMq45Ybel/R5J6xmHEc57DvD8c+MlV/aNLkqWEm03VhLWk6kdkUK
TD8F9O+rUZ9d/Tkl5esoVORhjXV5S0F0ww3ERElMMKts4aDjYZaTC5SA0DN4T4sA
S03eOoWoW1JXModAo7WosqMYyNm2daBq91F3T3v/4u93BtppyTP/cCMtETenL/yX
RSeG+9tL1beNgUbO9Jxg3OdH8CmNOqoV74eArM6P4LZIEh8b2BpdbNojr7qLf88v
SjThltC957dSKDiK8pKIFAhykxVWVD11mYi5RDbJAP1PWljFyAluF3BvDPT3HtIK
cHazjWJUPdp8MhIg8smKjeYHmfyB+bf2RvbSLlcnTbD5TQCwp4SMEz2Z5rIoM6gO
ogPPIFlJesopf/QBBFIvqZzL719sUzknp9m+nVKeMIaD6N66BquwcYT2U8nOYDSg
NgF9w9XWp4frlsDpM8AO74CNwiKKdJ+/TGoi7UiXscAC2bHW47WxFAPx1y7QLpkr
E5OQ6pBMCRsi2suiUM9SQ4m8S0H0LVqermnfZ0Oz2Nh9VMhI8sUCxUaWwVzLQ3YH
ZdhFvrSlDF2pzQlsERR586CFA+iq78lx4bwsFH5f13rxBKCpPsQtFQQiGea4NK6u
x/aKRe8XaOBh5LFUGuGPKAyK7Ac3QOz/KPB9Rf/I8ujj24NwEJIddehK414FqdIt
dNdnwZo7PEINubIlZaSwF+5z3a7mt21gkl9Is+PiQgl95cpXnPHbqZgZ7jpj4AJq
gJV1vtuO67YnG4L98V46kcB+GpYWRutNUy2F/q+qE/f03+QCm8mNNSrarud9Of0y
o7I9WE/Lg4LqhQo6dccnXn3fBv69+ngng2qx7Pd2GYtOxJbhkPLObdt/97s1+jf4
X4fbW2eC2M9gF5golq0YNjQDK+TkaCp3AsK4aPGFap+X2EkS5aLe7bLLe8E33ojd
H7ZB0Q7yYo08Av7ZJz31IqZz4IkQL5mu6jC5Jib8yJIsGD6hQsmUxpeTBDmpP70M
ywT2rtNu7kOepb5OngB0ijiawIvcHbvCMtoyzqmNcxHeIAO6tDFsPTEh95onqbfQ
YI71BzFqG8vmrOeGVg+0wKVONJLd5ew1zVLwJ3T1X4rNaNcteQ/qfFt2fGEkvCkJ
WFoxGHFC6NRXd6QjC1uXfO5nSJ/QyfFG4WjTWpHg/zAxaxNzhsmZqXxp9TeykIbt
rc+DxKnRwB7b0ZRwdu4Fiwp6j2GyTwsAXqt75hLhtNf4D0Nz0CUT/BsFS6DnL7M6
GmrC6F8RdOsVSP68UQw+ABpiyXnn7I8YaP72vLz14Sx/ZHpia28LdTmstXsTBA/L
goYGsrEQZ4XNKZWBGCdlWJODS3TP5puQbuK2GoSPXjdD83UmfX3Bz9zwt/Y4OCOC
bU8tLp8t7S9MPZmIfJ694gdFaPuJo6+k9CMw4o7fmuWyiog6VMLb/HTKX5wjlksn
b76NEeARhzSeywznJYkw5uSwMQxQuILm4aGhR2o3j7I34FvqY3EMcBTx4qNHhXAI
4HxgAwS8yaQtel3/3Myc6NDzCET7RAZ9OrkG/NdjhfqbMiUylRFLRBpi7k53CV66
BVvmbOox0qWbUCRB7+GxEjBAbSYQGw/MAmROC9SDJ+QeFcOECDtZPFGBPgx8xFNw
ui5AdgxIEvOPyDe+cUK1JeUuSVuDH65o7QEBVymAzubMhCHFdhyPEIgmtjyhTECe
K2RRtMOyNGlVdwZYBxEV91+TnrJGNWwVD3qDhWNwVlFG3X9+qSBHBseHDKgqe/L+
e+WOCB8IzLtOqpi02js2m4w1z22rst0xfkqzWl59Bx/HVFP2mGwb2jq4KsPt4U2/
1J6Kb5opgR3Ymj0eA9y5qVm8QWvfQsQzb9x6LRdWV5uKkq45aXK/KGwm7If5nT/g
RJSafiUtGaUdq7ACQ4i+yl2Fhav3olE0+BS/6DB8qtcEHaZLRYFTbjjR00O6mCl5
X/rQP+bkPBxox8kwuuVRSx6QIOFeIXFlNH9ncVPynsV7Bsm4tss8a6yPfDn6EpVu
OQxWo/TWspzxr6ogNkLZ5+XM7YO/lk0mBo3inMxkDRWwWdDDtJdww8zMASiwJvYu
n8NuCfD66Sxi6yZ28LCLRBag+IFJVMM9eGJfzVujOGI17vrr96a+LGpohx47mKiZ
+RhG7SXUmkr0L3N1r0p1MVSNVJf3xL80bmR2QXZXlcEtL8O6Jxm8JJ/IAYsbZUo5
db/dJOuQPW3iWgDNru7npwli1QgVnjN4yg/yA33UOH5W6UfN5hkrC5V9QWZHXBu2
0ngNq5/lFzAGUjLtbk1+6ljPwOtlVxkiNB/ZfPUG+YyY9AAoEmxJSGA/re6ksyOX
frzJyUzcVude8fVYFftUbbkL/JGbjDTRLroHADl/HzIP34feT7lO2hdmLRfl95m1
/J13e5qG2n6H8ww+oEFVNp3A/WxuIPW53Ez1xMTFFERspB9LMhh7mk4wIIDB5WkJ
8fjfPxiFGGyOyBPpzBsZVd6HaVy+dXUWGryMk7ePV4JKiVBKUdTuBpZ49MwSL2hK
eTRuBXCx+wuWvZ+X2SHISG1jyMw07PROf93ZuaczjjovR4y0jQHi/RDUpVxYq68X
e0vdX7AxoWj/8FZUCHGQ9OkCtx3znZpwVqIkA9lFJn7DWa7j9iTjH1ONWnUq5qDU
EDCrv1VSeSJokFshMxxNaca8Y91gG/BeQRg2iI0ZA+cZm4FUmoSneXzAKFi8k+mr
fzHuytJtdOsLylCSZkd1jr8eHL9IgbxczhoSf0Lx13hEZgLM7myFjFC2hdIPM1z6
9nqZUWMyCITB6+ODugt2Nqdy+5WxmBhhgxm138iFL2RhllJGJklQtTOiwV+E7/u0
RrP2O+YAmQfz1ClBVEx5azx/2jtISIZP6c3JtCFuRZsFbVEXwxXvpQAD09oUCVSg
L0cJiNqCuFkDWAEa+gv/BV00qMLwKnMp3DiWtjscDyulGhaQI4vy0EKjMWLYRCuU
3AlsHScM/vw4NNwve33lKmlCsYMJ1ZpPIJPcqpXaZ/puhg0zDaqPTMpv0ybQ3asO
uKq2UqHBxM+Vbjtg3veuFN+6Sz2EwO9BnTXGMupKweg+0aHbmYZp//QJch+8BtOA
BOcAlJinOITSnDs/drdgJvLOfx/Qviz1xqNPnaEGqU4O+UGue5tjiHhbJkFoq5Dp
ThLyWCkglUPqgaVMxegt9wZfT2wCyrM4wcZUy1g9fDmec7ZJshZ/HNheUqNhMtib
0wlY44Q0x33lXkng0CJqfv/uCq4roByvwG8/03Y2nIA4CO0Z3a/2sDwH7gjqH1X4
okgRJZMRY9914Ldb6Ow39mCKRN5pui/xDJXxE729q+u/bKvs0g/E1LbnONx6JUK7
tywSBqyZYhrufZbWhWGyNEDXZSq3uBQetlQF8Fzi3ojK47+AoGegXDMiH3e0+cK1
bFD1VsGzhNVrJqpWs4L3pfnf29ktT/EbX0sLfPbp0Bb0DzPfsLFvyjREuDTym3UX
h6WQJEh51FiPxwHEcJV3/GQeeH1TAdyY9JbdYyH9Wc1nvQItrw526a9bmO8wy3OL
U/+j5OXHqo9sFhHsZKWGhf9iyE6FJhequgS2TGKjT1AvN/6zemgNRKwZxMQesWsT
RZLl7T8lrKS295Chu6kgUnexH8qjQGRZEee9v/hn+gYeETNQIpd8N+xK9x3g6Seh
pQa3pqrtPZYfrvg8wLWukawbMeo1NV0WHN1bn3BhmXPRBnocIc9r/NyOjsoHsStC
WjCfjxrU4T+SLxgQGJdo/eipGLM3K/hFnGMfqwlJUtGuWK9fQRDYjVAYcjkLJzZW
aCMheZei6cQwNxS4kCfhxeIDOfpDoxh6lJJLCYBxHiOKi8xMydLe0Qv0UnNmsf1E
3+fBuD1fGgwWYcn7GXn1z9oEOl+HYkKcC2a2Mm18luHHef0OFl/bJx6f1yeRkHzr
qgeojdSmSmxl4V6J6KZgg5oiMglMBxcdYCSZGAY42xCTmkK1cHj6RBcZXz7t8cCI
dkoPzYMdVKJAZqEfH3gHK6yubjDExGrdZX/TntyXTxxt+M7L9eXROx3DlYQwSH3z
JxZ9e0BybHbFKvtCMV79QTdimssEqr8MQAWfaNvAINTgwFhrKacTB86sMfXE9I6l
fuhmERtD/Ny/gWV1w/zCtLFPIimTXb5wn65Gov+7coU3MnfUyd7xCz4QVdQy38Jp
9aGxa5VaNhhL8TLTUU1JNOKzsnhRnBn+hFkGbwGYn0UNZEzs8JEZLyduf0rO0Cyk
IRPsi/jKBPG+5Ff5ZwGOmeVAyn6k2l/DxP8zDy7GCsg4s95e+Oz9gOm2pSMnif3M
VssxQMdaoXSOex9CBKXsHQ/87tem17zB5LC9gU8YE8y73jaK4fhGRpf15HFfcO5B
eIxmnVdoB6TNmsPiCxgBypQuDDc2He7FqhUW9+OZ8QO0yhseo/FUKw+hgC5THXik
igJv2WZSpL0f0yxlinUx3DljR8scG8mB1E1WxSARu7f6a4tnR9+OmPDOQt8yo1dU
GtLqOU+UW8V6ZQXSOFjWUxAue9VYJ2kt/pSU2grq32QAyD2Q0umjg3KLGwCDLdKi
nh56SU+Of7JXgjCeYIlIRF86mbMWoH/RWRP+l8sEtTT0HYknNH3EKG37hjk1ud0T
52ScKZ9Zg3+UMkxFMq7fiBHn3EwyHWQAsi0BRLKL78s65IybawNf4bvP8oKuaTxC
WUIV9wtaoxXGlXqkZOkALGUbG0qASA+zh90bMfIdJ8dL2LMCrcHhYsSnnKR3r1bS
DnxjmVR7P7AYbx2gZNeZVR/M7ca6lLZSK5eglBr2TiNBHxVd39i8L3Y5Fad8Phyl
0x9/38m7wFUtl6iJoUzXB+PKMPFG9bUQ5oxNiH7HBaFKSfodO9gw/MKGFwRKhx/4
iPRsRGSL+sA7OfzcqibrEg4rJvJmSB1xMhUxEpn8mEpkVLe94yhxQ+9Tc+Z/uhIK
8XP1uwknL0wB8TvmWWfexJDTCI/uimroelOnlzqlrf0WE67j51Wu58EuK1HK3not
eqtBP/OI1vOEJWCVwosb2gSLRLuOr1z8FSn8iG57l6FQCcJwgPXYhhulhLvtxBJ3
aHoiY63H02dxWHH9qKSbcYMDQkyskEeZMpSSJSHj8IsX6PIouCFPuCNengNHWXUX
8eDTXSRbaffD5OzTXxHGWxkh4+Ngxv2mGhThn+J4/IDm44SKgk792i/jUIuG+zQe
cx96XBqVgQrY4pIUNWoPcHg2BkumUuT+jtOzZV/nOttnKsIUBOsW8YoS8fwW1pCI
Ug/d+aJGerEo7QPrLvmSVnq3y82kxxuX1RReNC5DwgT1zuhe4jfL3g61YsJCFkOT
t6nUYCYYB8T0YQc+NewDn9tQB2RyrYhuNb8DkvL5y41Dx51W0jWD0lCFFprqz76N
HZgFJ8l6wnnLpjw8arYg44BTt/xwJrRTwxAdlN5qJeC12lcIHW/tCeilIYVRWGfx
tfmxXV3mUxv75u7xDzhX8XB0WSc0vBXJeF1c4EtJmiBHbBioV6PP4frJNkX4Ijqn
d/mESp4BoZdk5bVjzbPcK5MQvxlRF1EdSTjYsYbBgQ6rZvdMiE8LQRo2NhLJlb8B
kLTSePuqhOC/68MLU6iCsFhP812XFaTG055a6kfqYsPbQSr7ef3F2KC5C1WHv3m4
6++61cugmz2lkGGnIHMuAxUyYG0pQWgQPMEA8pTUUgEn1+YfBUjcKqhNrPywToSd
dfzaVqIwaAPKnggRFX74XckxvSkSewdZVQyfeXrzjjYxAEQNO+Sau614LT/Yy0af
ghOc58XllyB5jMSmskvfMm+hs46SUPJnQh55hZTRC8U5VSLTZOiV5QdypDMStkz6
PWiAs6qOzv6urB0X96cHN5Z06381H4GFWlTFidz1nDuAXAAW1QH0LfvERu7K5/C5
qiBlMxI29Zb2Jv0nkTszhcPf+G9kiRKbiw8yfEZn7JtflmvT2BOx0gH84pOiKuUs
e1ilpx/QcBWXLmRH+GiyoVpR0uqmHllpLkHKlsin42mjobWaZKPPCXUgg2UPZ05z
/PKIXY98WFiwQs1gtIZhUodJpvg1EjMOVYM5VB2eZH0sA5YnDkLTcYkaD5+UrL4F
/MEw6/s2DYn+iTIVktrYMk5te3U2gr40DBV45kG/Pu9aOnlrZRdgvXAmjQNBG+bw
2LBqJmzlKdYIFTrxWIGlOvvm1ORmFd0fwGejVHmAZViLkpcfsQXzzbnE7jkpi/qH
azgcBvbfWOEmbr2tLrUwVDWuzxsBK/BKhedlNMsh7o7IUTqzJXx/Cv9vKX+Jtfsx
AgZgX6weeN7/E+NkRbmW0EJRf4XJRF/35BOheBfd8GzuiSsESLxJlegmxIVQwWa0
dGkjMFGMD8WR5wTJibH0dtlZLu+8uuiqQb8ZLbG8kXqOZEAev6VIsyhCxc53O6g9
q68AxAGScnTsGVbFrGK+IucQz8MFs2NDyD9tK1ELX0qOJ33cQcWv4rJvaE8+sbjm
P6R0C7S+z6AlqvIeta+5Sq9r26mbdsIqoL5RH/FN2QbPruO4I+E+q+gya8m8VeDG
Qp/ZlnymgLCfxvzDfBvuZyUqu3IGJwgUuSAfnXw4QU2Jh5HVprttI+vL3SKZMgHq
O+tbsG//VnAKCYlIZpbYd3PiWitGTSuar1D4yecpI/70BcDqMUaQRyvaKB8GBSQ7
tqvS77wX4SfjE5O1yd/lAau2wvHMKYABzA0LM/QUiOQ6xHnRW/afv4i6ji/JfHn2
rUSCa3W5fcl8JU3JvxPOaxsFObfWt/QiBT4T8qGKFEbqNtlKHr57AGFj+tM71yT/
j/+/OrPqE4qkuzfxL7aBTnM4c2nsR4ZoI9II9oyZl9NyhQiIqJ96XFbPjyNuayMz
pbWpPk0h+PH6HJ4avnnMDncJ/QuYq0kSul1uYiqQxXswvg3qbKSRg24ZONfQhR2T
S6PK4tndMRFNbsoNpOyoEXevEtIenqBpKNl5vjNz8s5BEPUt7sR5gXhrVWlrIonq
htRg8oDZBjfULTe7R2zjgj3WSktYEhxAodz1gdGY8u2HcP0U5vWCdiwKGUaxhd1x
g6rABHwppaSi3lvAByRnsF2AmMqk4Gmmr+4N7Rh0AgID+DFjLHD0Q06oGR0w8EyU
RRpJNdS5+h20gjspxg405T3ymJt7y6f/nxO5pa5YfJHPOaDdlQ1OdWqAP2IavHW9
1NF+eVzEWJ5RuBkMwKIds4zj36l/YIbU19QOy54ItWCJtCkQnVfhPue21XS3Dqzm
7cbSt/RaWQHb7iWv6ZxAcrUKv3mtiD2aqLvPx8FtQlmQvandWqjB9SmjKA47rfc4
JrMuGrRtanB9e3P4Lk2THG88uXduTG0KtTmcegcbHEeQ/McVDJyObiSGqZGliEOe
Rj+uLteN5QNM0ifE4ZTq8XrWAQNZ2WzBl+iova6Pgmt4Anlyez8OwoRHFMbb8Sbr
+47OlZB0TImoimZ0pi6onwQjjxAh0LA8fLdxBaFzIV+ASBRb50IC6sdEteaVd253
G0p2sCJbQGOBdYuacOfIgnPQtuwL2vOHFeJXNUdqHL0szQAtZalWPaHh6Yj6yWh8
ptQcZNcChb/ooxilBF/fC0Yx4VFlTC9ZC0UQY8IarUUEQDtdjRTqStw2rTXK3zbY
NIQfNyrLY8GoW4nPCSVR1jOD3+9tv4ohWRFVPB/KTaW2tMyvPvdGp73ivrN3IsBF
w2YLopWRnRFx5DOG2YITruIrE8jXMWu78EaBIGgoWCo4o5GerdA0MyZyhFCsnCTd
+lMXdg5bG3znR/C1a1Xct1csjGslqTnhgFSxUAYr3hCWL7TCC1vo6iGi2tGRcdj3
DJSM4HOMW3iwzS3BeSzaEAHSoww01wwn+7tQKPJMSU1bSGjSkL4sb6fZJFWGH4te
xbxxEkVJdOTas/490nxa+OMjvhLbC1rHQaxkLXnnyVu5In288xrrAUHaqNFG5uhK
kypkWpoFl82JjtGYDQ/SzGBLX6HgJoxYhh4TmLmsvtF4F0GdDBZmz69GPNfjuiRg
EXtdDGZ0IfdTyfw+0AUKuY2awpsYSBi1e+TAw/iFOLDgNgzS8ADiaVWE3SX1sMDu
UhAO3SEXTjocI41CD/Z03kfPvFG1qzm+XKPlP3C3pggIdctddeMPArr2rvLjJgT4
3Y9N+fOc0XDUneu6t6H0G2wKbY3fIfE2Rzx5Slg95ZA+1Aw4DtzOLJbmCy68Dip2
BgyLFPbvUBxAi9Gi3IbwgwpxqA6ZitYIRzt/0oMAswcqmXeKv1M78GFbg1EvE2fH
5XacKpDDk+NqCnVboAsnHD6nCuNi3Xaf/xZklz0+B5IsC0Ichlq7yZ8WICIf6bpz
sgvq7ypR7qhlV1hYvMk3hMaa//Jl9KpF5mus8/ECImPv3oUfLJvshNSZNr6vfr0M
OSkNiFoC40AJoRZY/ZTxFyO0UauGmJJtKw2PziTF0E1om6IsuAdZcLdGqRaJeKnd
pJhFT3Ggk/PJ3Dg0G3mOGmYI8gLX886G/YQjwY5azegosxtTqXhu68ijAtLlkQgV
oMQ2WRuG3XLHzttBazPGm6K3MiyCXHutav21jlibhAN7MEYbreutFW2LShvOJ6MZ
N8yAVAarLHDq8okXrXFrc38GykP7XMv/h3tEQEUmOwl+gRIb1hWMcNAJijEpYrk7
aCEOQLV36FF653m9E+/jzt+TO8wlS3RxZ4b5KivlsgyYpWBTzRw+JdEZ/BLUU1n3
RQ38HPYKwxwxTks2Hi741SeM488KTUXlvXHH+2Eu20QyYzkwd1Gi8DNqo5V7gn3i
ti82SopKQUY5CaW4q9DMWgzUb8haencWbOoDgVv1g33sMrQ9Pa9T5k0P7iZ6WJfW
yh0h7B5OPDaAwYLz7UxjDlbC/xUYhNzs/R7P4zdEF2PDl3jI7zRq2u1fPyxX/Hdb
6CnjO6MEHbkUBMITvdLMwzKEi1hqB9d5PYYKCMyBP+HKQytmIZbsgMEy6g1yHaza
cqUkrlP4eOEIYiVuYuinTXYKdlah8p9XMH3bAfnrXiD0MkIUjqBOpHyn6E4lvT/+
8qsgCHfXyDyiLxSLpAbHUyKTCCwbuOSnWX4fcJsiyzxmQN/eXT9jbJCr8zB9iXDX
fcZQiHWYS5/N2Ke46/zqO8jLtla7ZVuvPbW8c83K2i4AmtHZRryIzwAzmiyYF6Pi
oMO6JOZwB9bhGbwrRn1rtOsXXedDxZ3riGq3zlRnsLkA37AYwLChVkW8kvR0p8lU
1E2MHD3GV/xA25ToZ1PPP6b9UPBQWOgnmICESbx9huT3DzZwgJj/WxrDSIVgqPeP
ZME76ycLc7Eq/Fhv69BcpJ5pb0wSL8EKGsdf7rC50d0qtJyk3eQ/atMZwvr04lgN
TiIOZU2T+TqIBfO7lEL4JujDDmfD+VCEFaAEg9pd5I86WIR94WRrH8BZ2bkLq37Y
o3VFLaFyYHnj/3s3fMSyknWxYx0bEeMeXnpLOjXtF3RAOZTAeZ82NbPUZ335KRBe
TMyaaRZBjnDw6ZtOwGyTSIRmGW36y/74fJlJHM4ABCv/L3KejCcG14SPQ7ygD9pN
QYZ6B3sQBqW7oNJGL88kz9CMm18MoNXYzL46thD2o/hqK5Th6gnYQ1u64/UjFQnd
HmKLl16ZVHXTPMfO3N5SVXKocSrQ33PrWKNRACBOr/NRxAcLJ/HF2+L/sWeEswtJ
6lafvSvlGx/UYRErnHrqzFSBt0lVEU6Lk3yLzRZq+bLbUgSXC62L2D72za8QqPwt
OpDYIB8sVrp0HUPBJ6fQDpP4o651iDmudqRaFFhXSI1mkSyeBm2Rv0Szp/a3RD4U
WZD2dvsffCShEqfsN1S8fddPaYespUXE+60/V/RmnfO38KvGyplVcTYO4+ewgKen
RC+qUP9gHnk3paG0iMHmIP7cztY0VKcJlSDfhlk+DVNRO0JMwEhS6qyn8FK/+o//
dsDa92NTJ/Zb7/YAltdHSF35YAL6NWzdwnnx1eou1plyHwwsVyy+xynxKw8Q059+
ngDKIuILlaQzCE/4yBr4zx0TyCAMHaHa8Y3GqT6Ec5D+Bk14PZB3FXwuxc+XHjrU
7aNdHxcvPEeb6a2EOlxeDl+BZT/oQI76OtmvaEA1QgQZl5KZjcm/Hy8l6F2PSmkf
utAlY1y9PCu/zRg/AKQu2yYBflzeUxz5atqQfaPl7RVbTeGcG6zzucC48raQ36xg
vm4Lvnj1p6/tCJn+gAu8YrUi7UwKvIqPlZ4AoCHakKO9uI8Dqzu/+xTxjY9GT8ZS
d78og4+4jg2+QIkjI6fZV70pdFlrwSI8t0VBDa0Pg2/Hz1/z+oGuwilNrmpaRRwY
GY1r4dM4wgSQYSekKv08cZF1Osb7zUBtyC8imDLGGDzZm7EE4iPKwAVqsYL67/eV
QjB3KzecqI/1SG6+4hxVxPztn+zsSMdYNjcVqOWOZVajcwuFd5VZpkNC+vovoj/d
ZXxdpH02LkHWnDxIZnHLGv8eXvkpR291bK3AFvR8eHzUyMQNfFxBPJjkiC99sKgn
eGEIe6UR6MQqCRU5Imosm6HNH/M1qqB+K2DBosGv9VUcxo3Nurg0Q/emqM8y/SxA
HG8VklCn1cwlno9z5YuuHg9tg7+EeN0lWBOEpyX4EwoALhhdQkw5fbKukIeUywNo
nUF3zW8+Vkp9vG1y0SLZtjfticC8QhrdEoUvWiBsXvLIvWfWyKWrTuWpvgmk2SxG
p8PKC8FYLJv0r6jjYP6ipHSLVLDzWAGO63KFPXJPnR+K2HfNFqw7B5rJGLA7UUuO
BlbfweHPPp5tPkeookN1kHjccQzP2Q8IlE9DJGv2A7+h68r81ImZXbprpiQoASqT
sPKjUcwOB1SAyndsW8DyvYmql4JWeYLDsdtWL9vp3naflyuK2ySHiGHykf85IrN6
voLveINT5+qC6UMCTpZo/xKN5N3LxXfomMzb8tS7SvwqVHE8XuFoxH6Esb1sBZwb
5GL6PfhaRB4Bj6E9x+yPqCwKhJEVllXCETaqIVFtRZelyiBg41O5XyqpyS6DtStF
Nzp5N1cRtkxsTCo/mEHIjYQ9wiPN9wK0Ql9A3hY5uC2SZLNPTrfcmcWaUeWGxxIC
heWFy831VIKpAVdxY320+4uXc71p8WGT/ZlG7BnetuirQEf8SUsAqzUyeABPg9zg
+OHXO84eEq78E7mxl8mpvImbcal9MvbtqDoaJSumod1STqsWvIGLPtMQa9UypNK4
dTL5/0A5NC6arcOiSLtFYto9UnFabHGITc0yENYveTZQby6N4xoOYl5XCzjhkUaZ
05KH+KL32NP6oQxgnvayOxGo9yMD2ygpy5sBSQ1eeiArY9KHTb8gVbDWjJm7zA7Y
NadNFzHZHIuBosoDT7J23N4NMFiQH45OX9Pz/FIO6c1ibR5vsLlmebE5nJm2Zrzy
EmvISYpPPMoe9yfhD3jS4FcZxqKNFJyGJ+OsVJXFRaK4gSW/pocz4eOtNrlJUL7/
3brSXxBgTzsHVkWkSwfJjCcmeougN5ACU5YQzlWhXEQF1iZmwuWz5C9MUGX5omja
pFHSpjMB+V9DB/pnYJN4cAXII+DzFbgSzCfTqKOEgjdlgkMQAt/TzjUQcSlJidkZ
tvOo4BzvnIXODA3FTAzBqtR8JV+YuIQDLB8fM+1KX9nQETFSB/gBNo06pHtvXycr
eWI72Wjwa7KLI7/FZBejrPO5k5CA7p/T+2Iiw9bZyczwFk1XU7WxHDGrXpwtYSp0
98QznhEpbJM3Zb/K7rJlM1BC+4QzCGAhPyLpCbUKTm/8mTZITEY1N8eBLy0QTko/
F1eytXYUsqe+xe3LdnPLIcgcc7ZNE3BatjU1n/pEEnUXjPVO8/nUwwOj+LLpy2/0
F8cvujsclCacw+EN9rJ+mdjZFpH25uUEDDgNYx2qW4eHM6aY9nvx3XJVyT3ZTlwZ
iFz+gTHyTipUEWkYE70OPUWb+gccmZTtoKCWhHawgjv+4UKPlNIR4FS1mXzqwK2k
eLcHxEAP5xVkxUIdmRUCnqCpukNz9ZPp2vgSkCjLs5HB0iQCKc8Fbkb/yglAB32S
KHSjM5T2Lmlu7HRMjMdd+pCOJBUYJg0cchZxA5vTz+wsKrhHH1L7XW+F4GMcy/NC
sjjekE3btUjFPGgb6fUNV9eflQdFyhG+SfS4fgw0qqQJHEY4VvIltAoYIA0W+TkL
QeUvCThjTJUoPUxI21fm8qytl32dF0Jq1yDD0f9INVQ4pjjiNGu0GJK4Z3gsa7fl
X9mtezrtHjH4SC0Us2dIIf4XMwEQbMBMDjW24fNruDLdKa+N2i6XGxF1r5Z8feAO
pH1PEXx8D3Ji7CBn0pUqWH9xcStpz5MR3QzorKb5bv3YD5Fmh9ZTpkNsqBWNAreE
c/BAhV2bs8yeRbhPMCNW4/zb17z6PJ1TCRvgZT2w3aRGY0IeoXft5Iqy31ngyy3j
t5ZjtStVia7xjOu9oExSlgVx63nAj2lTkRuR/lQXIyoHMDHk9ENLBigRAztWJhrY
uSUTGUrBVoJc/Y69cBWXfgkFHReePYQrVBlF4kSB722VrUojX4Pkq5LAIyBsaYqm
2/jjdmD1qSUdG0FtwnhYmoYnDDiJchE2matrrafny+VZ3lxWP9erITcubSUPPMRQ
uFhiN/7OCKQTfAVNlzzMqP9VGCxZRgAY8sNTZlgqbAy0WQbkNPKmS9boVWGVgNNw
VgvAd80jazrss8fHRHQvePyObHVaAoECBrH5TOohVJd+Dam7rfy2wEQgHPjjJNjH
eKMbCv/6YPYbaZBeIhsUQNjiebZSQ/GVGGHzHDipUJdHwTJdoXEGRgSOK2doqly/
yhgjUlCpfvPzJ39gPAOoYAUS7lE2AIMJBstPOEniRgxfNNp0gsftqayrMJAIWu7o
HnJfgRTgRcle+NDW2SkT54m1RjT5sHT+h79u4xwum0sZFhVVkolB9/1URWkp54Lh
aMiy8qZ9Wy7waxBUS+TpdGB/lVAgcGKfqiE+oIFU3bqSo/TRncL1bqKtGfIxlF0G
XMGv7KmZBmmk1hNQBogIULKvW7cVbwaLbJ7vb/A55ZeBJ8rJGRriacw5FlIi7yQC
Bp0BnOjvdTfp6FSnXnEX1aefKvOghuzhfGZCqoUemLe3zfjeV7NmAMedo73cOLOa
Ng2WBHc1jXvghgqWYLcojCrLnDPQmomgwvfYv4g4S4JWgg9awEMGcl9UvEzdAhQH
q/AkihMXV2upug5h+YcQhOFcSff/RWDMM3aYhluG8Ft1F8Xmui+Mk5viCAymTRQN
0gXx+SUnuoigGiQBOtDnxEFdTsNL2w30XrNYWb4eN9RvJaOHjXv5c9NA/Tg3DiQs
NnxQU7dxecqUIIJOsHzxM8IGdAlIZzUeY+uDB9WYfJMEp0A161GzQaExKjcaCxPm
RM76d5DW3LeDhZgo9dy28UXVOtECO74r1iH1tZ8ea2f2ucZBmT3L2EuYTbEQcTMR
7u6CYwZiWMSksWRiKQrPAbt/gN6RLPOREia05cKxi/+ug+e/Uo5FvKO6DXEmT4cn
qwQal/SxA99N7p5cl5/koejf7HJtzGtj0J5ClVk79UimA8bIfVszy9hs6/hxLRFV
Y1xtRDWfOn/CuIcXffc0mgXQCIRtjAKiLZY1zW/esAA7UUvwWPydIpEfP8/2JNem
N0dLzxi89TOkouox+mBbNMXJMp3SBMQmZpvUFWLkGi/PCEWOwDuS9lOkEnS/aXLI
tJYIko1Sc/15LtSNitf5C2v0DcqqusA1uL3yzs+lO/aHIenQ9bfBSrtigxDn7ES8
IA2m3sxF+wk9a+6I9OwfXUXvKFsMCkXqa1srKtNQZqflNVONtTAq/RQhzm6v0dfv
ht4sjYN/u+b3QIRgK9/W2Mpe/n4ADAr+dmGi68ugGFoCiBMLv8/U8pV/pepkg0/J
zxK4iWhmKH62T9zQEUaGLrdBq18Ea3xMB1K3faOBc4n/CZYpwlZ36+8g/RFIAkXE
ToVGfO8uyY8TB706Seqr9egtX74nvkDaPaunW5mV64gP9DckBRVUmSJcC2diqCrA
b1NlUj/s7CqFrefDTfPW3VprFGOtIpZEK7/2MN5ckdkCM/BXh+VzeeHCeG9sXB73
2vrILcm013FhSzyWzNNR7IPeR+WWRPN2hW0cRh3dTwWVNs5lkG6eSunHB/OR2W46
pU6KAypK5WNwK1GjTggw92wjmU9IHTrIFvz/eVsFR9AymJCgVvNCPsBVU+Ee6zWV
bkFaHD3MSq073M+3GqmTNr0jH9Ht6vVTID9+8KTIXwnicESrWWFj9+U8xhFTNQDS
FGIIllT0zOUymPIFUCPq7ob5soJ6LFIXVL9Iwa2pBePVdaK4DbL4mqUUxtGdwUXj
ZXyt2QU8rbdM/yG0K8AoZnusE2pQkCjmVylK3YCg1j2XV5HimFeICoRgDbKkYqPy
2w2eA5dyjuu8EK4W5VWQneKUz4laKdjGLzZHaJEm0fx95qL5k7Ha9kHpa0OrxtYt
hM4YDPhE9Q1tMABz+eCCDHrV9HscNFB3uAr4c+rXpBDmzLKHsLOZFKbWLNCEUiRu
6mLLJwTZ0C5po4NkWZJkmiouwRs8uey/rmCMsyJ6aGuu6TFaqfyV+0M4MGUk9VhN
g15ujbZjCng34V4K/edL5FoF5sxjcH2lUUP/zSQrXDo+CbT0QTjvbu4tX6xVu6BN
6jbL0LgXGCX9YIX4vtW7dHiCZxkijhd4wHZJZi2sZ7lByyGH1DQvg6cW0aZh0DSN
K/6RGOnqJg4nLkvKLkuJTxY6ICY1lixdE5Lgy4rDkYHNy7KX91buO2HwmoWDdpr+
F+c12idS1LOpWTN/nBtd7H4Vg/Kpt7pq78BOJ5dmMqq7PRCmHypyySk2p/ZuiOwe
49WLqgVWTZqDOteTz5H0gctNst0lv85/d1BSMykRAbz7CueoMeyJ96cqOGmXdbK2
udWf6GMcWxbQbO7pDW5AxivLNjwjOSRH1fbxzyEjp3JzjCQMPh+dGinbOqM9tmB4
xKb7VPwwhVMTTGBXQrCaA1nCNObTJtSXxWI2yEIwafxeFVrtC1X79erkHC7F0l1V
IXfjwxc/p8R6JAbGqBoqgECkNmn8cbOXzQOpDOmqTKazqS4Vgs3F6HEYo9y2IpWG
ME3elJyexQe6b1QlHt4jgPPeFH23A0vq0yviRK8RSofh8iVfBYo639ZJfYb9wWA8
JFv8bhuJUl1WIYrNB/qAqn3Xv+86Jk1rDRMabRQ2Wk/FulJDAA8MPlgh3KJ/Pu/6
hbZSZOy+cVUtISpJdCM+oEahWDIRKldwKTpe7WrYUzyGapatuH4OhUEnOVGTZ6zY
NQwJe7Kqe0KrGfeoRNsTIOPzEJxoN2vs03wWvOATcHA+DHdC/inPBKeNtLhnv4rE
+mB+pzTH+xG3DyyyKLDtGp5cdocqKEIdh3Vi20T1iuQoy+y7nZfcAOILOq129H8I
8RwST3ZvzdZGKUt3LjwH1Xhdxf+VIFX0BpL97x+yYgFamb8P8QIvRtNYm08DWcRQ
TC/kmhGCFiwMpAXbzfSQ9SWcY3jeSoYPOJ5vOhB2/7uTvdxXH1ec5/z7lat4iijA
pcXGWxWNC+fjgChn01z9ZSFDYBAQKY4d8ASDUFEMaowOoBgYIczTspJJrIX1bCV/
Nt1fWdk9PXoXc7rELWU17qK4cc8olUREA/dCWtdUExTHZ9oEmlPwvKWWQo/UOGUD
eZbJM4B+GTbuElvT5GVKV0VdlKKDZ5qcYcdfgS6u4Mu83gsckiGgDKyxreS0eHma
bFIAZQhtqTHTiHQVX5yDwN5DrkHRaq2FTfvXKtiW/TjK/WIYHoNDf4aaE1v0NYvX
Y/8InhBK8QWDKI8OEy9NW19s4HX8hU4N0tXc2uzrpAHkg61a9F9PYROVUD7VxozX
OhZuG5g9l7DWxA5qsEtFOD8FMvhBI+6U9mVgR4f3a9vqC8dRPYKZbPW+EQaDArGq
tksA31w+4/lCV7E4TbwOhzYXFgKD7KFg+bk8+t1OpaTzNCDgd75kFe4I+Uk8pvmX
h8aRVuyneCYXlvmK5OBVB2nqlsCMySCMEyh8QeTut1TwKE7pXDnCg8zgR3KnCW7P
FhZqguF5b+UvXYo0po7V9LlE/bVb3xlt6NmlwWCZ8wKmwuwNjhdCiSGfcD8RaZld
fhrJ808uOgoUTALCl0BwFYLsWTVAmr9LWVxG2y1fZAydhVZwewqka87PVXG7ZCzi
Ev/RGKzQsOSespMwapF8vV/XZv6uT3xku4T1NpqDZ+vZwglPifKHYcxzlHelLaxP
UyDKA6N1jgkKaobgokC0pZMrvw53uqhmJxQ84vihJYFvIRr1yG8XWoN8C2w5IhWu
mE53FaFFkfampRL1FV88iKCaTsAt8vJubP5ro+G11Wbt/FV2qMiW3xZJgNlhQLxl
D5zpZdDpUxAk3egEenlf+aA7zR/Rr1+HIJlXT5agy+XF3xk6+ApgNa2R7V2PpWOo
h73iCDinXe7sXsdmyXpcwHG+GRZIJrvjRxRm46K6NZJQ1IQA0c0eqPQ4oOa/S1H/
XXLxThe7QHPjCJ2wCcIOEaBaPXWWc7EgTpjcn0OVjSwISSH8AKqxOMylr3RTiKzF
DPbp+Womtas3Ak0Yy6qXCbYQSbHeHMwuR7uirG1KwRhCNUWUCD0MzMFe9VfViBZ/
9WQ/4EAdqK3an1y0gzE8ZC5YGbJe0OyQwWuYO/hLqjaWQ3Psf6SMd8tHwR2kRJV5
cD6X/IDES+/fWhzW7x1UdVQLCHKScHI7E6w2Mlz+iBzZ0pH6xXca66gfAnjk5A42
F5cBcKJLf9Hvd6SYP18/eelw/n/lU3TvlZ0FCQdQfHQ78nu5adYHcWHApPRQRIpv
I0vB9dj4D4BspvLhdrT+0Ezb5ULvPufGMGE4pUGhuT5eevF1MJfWI7yuoVzFUKeQ
vGHSy6Jtpyc/i7J4zi9RWZ9/A0mESLQ83wjnreYXI4ZI+QFYK6G2f67qr6TsYNXl
wEkxQkYvP6hALgIA482/Ra0KOuB43JeCrhlPSdqXMkHEQaPj93JKEn2xfFalIUVs
e0U7Dk6B3lEhaiX2vlNbkkDrVjf6NjBPT9ctAe1Khu+XXn/5wvZnHiHnJmVq6MKJ
kjoR89DHDXH5lGjCa0JNIpz3eSdCPlnsuH4uzk/ot/8J5KMttfb+GnPnFcY/gGl+
qYxPq/CZa9byKG6ajBRPC0n4HrUDLP/LezA4aQIWypnQvUr+yAxpo92ouPvo/AAc
Vmrg0X9OujEgm23UHdkBa85dY7JXJ414x1/R2E/EnC0TMEIoq6DRhytbIZQ3Uepd
IzyChRcCMxcqfff0sgMp62JHQX+oDRKGy66fFbJ/x6ktAw0Xi9hh2LkTfUG15O9i
spZhb3nK0JIV4XejcpJDODzzrcbz4Ad4+ynusaVv4LWsPB6fbXvcuFgTk+HTXQdT
cuspZtbhaqkh1JHGhPaCDgqDx4eGw0aaE96wq2/oBdc4EX7zJukmZ0y1F7EFgaIW
zBLlMnPc+/1wmXq+VEPm0chBWHQ6+UIFlcRZdy/NxXLzisL4iyKT9pZ5Jh+kZkCc
YSKQ/a5cbCNqcJXtdeG/pDsSJv5x+9D9RXGQIfZ+UuvOaRp9xqwU8ttVndFX+Xcy
mp+mGCUGaNP+5tDmTWPb8Bju8ADnPn6Rq5Td8Gl+JjGL/r/fcy/mKTfYaDzZ2lPN
hZfoS1E/q3jOK5vJ1zC9o9VcfUofZJa/10Z/UHD4ez0iOBbWBEicqh0msBpVdjgg
e9Y4gyw8Pfal2c8p/y2U40aIOYMukkjc19FVtj4A68HUr/tpsbCpycTtphTxHTPK
u6AILnk2C2nxlTV+Qt0Yx3xW5wm8ctN6JVNtVW6i5fwdAZxZYanuy+WW0Qud2NS3
BwNYRezDeubcyCfmFgwO5s8mkVqLjCB1JDQ3wH5AeDL2ZiJdCQ+4QQxtEZ+Qb1G9
4k6AdSewdz5VM8P9NzS51aCph6PvHznaNlFEsuw8aHhIl2RFB/lgLChNgoIf3qAa
ZMR5DRGyJAi8ir3nNaygkiqC8/airAKfDQWyrzk/HWydVE1b7VJWUuj8Ba+pyufc
Va9VyehpUGMRUGttsfVRl6uyWAY4VH0pfPMl389OYEgmtZQvwV7m++n5k9GDBHOx
QY80RRolWouksKp29SHPvowE2g5aWkTYwOcz5UDuLRtGL5OE/ipw8yBtkrXvl1sN
04dJOFhY3sin5mqbOubdWPvV3hkkqCK+HIVdx6Er6vS4dpeYDtZn5ppM/2XaAcGg
TCEnPx8xxxJYnnSC818MJVl/9WIlngAjcPeslLaRXuTicfmeJ1E7s6zrWzyytNfq
J2Pmx6MGXrvETbc7saVcJq/wCmqJwl0ZQXJm7xa7xq8J503106lZNMJkcNDYxmUD
KIFbXAisXwvAoF/ELA1XtCt0/HX+es81Cf+52TkidMY8I5VdF/T01FpNO60bkuTY
FVgzrNzDcXJyLEzJfHdK503YB3ntBsK2YC4aa+4z4qC4LW2LIbcHowK/Z/LGC4FV
y/pms7VtHXXRhkF1hUgbcOISBoOFqpBBklm4qW9MQwlWtn5KrmUHV8Kzkhpu5ctq
cAPmHeeACuwvyDUnp0kUnyKJAtTxx9nojsJGy7HZg+ItovGzpLZoCmaeH9jUXEtZ
avsJv8KbH1ql55ecLtkiaOFX3x2iD0ocLybxxhEXaJkQ2Qz9doUrwfm8I7W/E8AS
b0GuWHgBRsrgK9CF0jiGx3oQ6dcjSBtP2C0tKrdpZvAXFNL+ikBJtigS7El8hDSZ
2MdVbSAs7SS4BJ6XNeDxc5puYqcUpOfhzTJI4i89RPaIKqWXvPV72wSBCvO4hmdg
qHsu8xLx9OK3+W7B2hlozvcAdZ0g9fK/1kVxVGtdF5lg7qOiTqIbAyvcK81/S4EW
LMEWzArBFylBeBTjFjPx2Jx/RE/Pu8cHs4D6igf21gPPCObq08pOI56L86DO5QAK
ytZyVwsx5x0MWdbdZLn7RqTmlYFQZUukmIkn80d/fzXZwadKsWjoyti+N7xg4VFM
iMtE2etDXPVEh8REUa/7aFBAhogdAuFIg+er+PBHfwxqS0XP/TygjB0Jg7k5kSis
lQd1/wxhTUaoZzu5nyttrslhQr93eG6IdcJZWa3m2lTM3Rn1T3Qx9PNRVH0p8O6v
qaoYDLeIVRdfL/vuJq3iEfOgOB8OO3zE+cpfETJceezW5fFDr0zhCDiyp6QPRFAm
rfw67/gquK6n71hlsjTFbMA6znE/nXjU4iFM7Wx172iffSyqsM7LXQdfp9QHl0g7
Ucprpl8ujB2F52DH7CV+YBqZfPTF8Wcohgw9GfE77Q56ygU+1opXfwsW3Bw0Bj5Z
HJBYKwzp6BmMuT2iYSa0Z/Xhit8+BAPpQIJivDnnObogYdXAhBKWejkUmUnKVq8/
FVN5kazKV2og3Q+YoV7HZEauqg45YtqytM7PfZR4FiF4CmQjlm4JBNYFj9ITPkRr
91CRF15gxkA1s9eu5PgcrgicmbvNmid0yUvR4F5PCObZJMqz61N+3j+kc1lkcGp1
5FFrhSC58wsUu1id9rWLEMgfOyILHh3LVWea9sqE01L1xO6N8F8XUKJV9b/xzmdy
nbtiiZLQO2TOZfZYeOsJz/pXiv0CzKbmDl3qlLrwFNfYWsue0NDhgHO9yCNgmrYi
f4720DJFQQ8xmNAJiDm7iEL4GdD9LqzlDEznvicKpLl7uKi8NCNyT6PoEaRnMh/Z
KBliH0WyQUbjm9uM8S0vvzq7ekdwQ+7Tc9rpF5c9bMDLPhf4DmAfy19ZWNKrcsiQ
4CwNyYWWEU35T5K/crgWzfVJiW1Uwc9pttgpftGlskxV8HF8NyTLuqsPKQb2rzCg
eH5wIv9VaHwuz0tTHqrsDbrJKG9/2AEOKxlLiYvh8GBSrFOzJExe6aJk7+7KQWFK
PDNYBLjXqpYZSwbX9s5ugargaXl1fsLneP6U9uO38tHJUML5/ineohRgrojRHOTA
T0N3FKWlM5lg+bJmfj2T/UoIvsyQWp6NaU/txb9OOnxVTBnECNJP9YXnohfbLrSO
AAGCm1a2aDFKx9q1W1SzgeZRJmKtd8nsH6ZO5eH7C7Kqr9g21gexiILekQkLncAF
+kRU2jxxA6rwS/5/ex4EXmqaaJtuM+FChlyWcMl1B/6MQYmSlssMgQtVDtJZQ/Ne
r6msXBBKIZffovAa5d46A2TQxv8LUb5XQI0RGBcpuj59kqlMLN4N+EC8JNBu5wex
9lRlB0vrlfbiVxIbJX6xDiJ5rkxe9iYfvsOmmKVZXWcWgGgcP9eWx651j4Nvt2+S
GngEf07arKICBl5MRef3vmhjnp9bFdOuNiE5Upintp5cX1fNLQeOFLbsFbSRiL82
nyDqgYPk/tc/pqrQ6sgTem0x69+awAsCGdl/BcquTyf1M66AnowRlMtgUdJSIGBR
4YaC2ZGlkLpjwsQmBTn3i9onkKwut4Mnqgvv5F3+VwR6dNQJeoquFvVTUNPMDWO4
B0REOGrMPEF9ullVe7dPcA6iouKreUImkj8b6tHmO1tzkr2lPNgboF6n19vAKvD/
Xjv7cR1JzzqpFt5FaNNbvWNZRHjqBZ1Bmf1nuKoqz5qaGfPOTnps2fjSbyUKlS3s
Uv9OkWUaN8EgC8H2+6UGetsLbcyfL10Nf739MkIY16/iOhfXfkxiHd45pZz6sno9
fJAGDXKWYeWzO/2IZcmzkSEuf7U5yoeAtfxbD8PoJr/leyD/nKWJ2l0vdrLv8Uha
fBjGYAxWRen51idjNcEhSGFvD8b6/tNQd5WVl0Htz9NOX8YhfT3Avighb35KRQ0O
thGMEcwq9eVxyQ/njQtPFHO2EcJ9iEwaMQX6Hr34juBOMF2UB3swqHJ4/why01pS
oDeFpGoIRinzUA1ES2B0NQwjqOlOs5sWcSxay+5KUagmZe8xQ/KZISJeKxXnBk2o
8EGVXCpGZFxXRJez8f5iKWH7xmSHEUOQpT35+ryAfyHXc8zMRTK0HHHm6uMw7Tan
tcKmjxGKBiKwuJfoAgDM7QH+Z0sqd3e61cAa5m+5pECR1rG5LhShWBGiqYrRqvKT
h3RHKPNULUQGE4/voYFPpbuYhS7xLaP8SzAHZpdSiVrUwAqGo9kJ24uUe1HJqsmw
uuXozXlptyM78ljOER8A0/JyDsjtZhWe6/jbHiPuVQD5RqDYgQDZokXvcJ+i1miO
BsRjLy+6ntKbtF1WE1ChFZa4N3Dz8Ew9CW5Sla0JMHxhpdKlR7SGpXZlwXDFzGYy
npba01qrXfzYaNUQ+pdVbEvoz/mNJpUkz2OOyZQz0tmMMgsnAaPMtLzxZOz8rWl9
8sS8CSi7t3tR3IO0U2ZEYtQ5laygN651SIRf/5cMKq5FGc8uARB2DWCKiTxEh7c2
uPWHmsKp9aW+1dhTfJbI59HdIZB7vZ0Kcwc+0Mrg8MflVQN4xA2eRXhV3HBzo8pV
aB+Ebt9L+p8jk0kbOyiu51R/i5B9ky6Pwz81+49G2a14Tq5tooYRwMD7rLmsHOXw
r5nRFlXro7ZaYXDwws+kKwFjq1BTjjs22hAnbvZBXenHM1DasKMkai9YO9lK6HVw
qE1uJV6IEeCjjR5g+Rc5FHGFRDFCGmP8gEbrtsbqCsrM97H+UWUU0q7L2noNvyzF
FZwSpH3nuO7dJmufXOoXHid/rtG2JcPRWM8004bcNb8YeebefKf6miDyFqu5abTD
2a+oDY/rqyHnrj2LA71CV44baMpBPB8RnYMwYFrw0xXjMeNm7pag3XbYnq2n3s3v
t0r3egrKWdvhkg1Jt/K9U/6XdNadrzb86BEI7gKw3HFjhDSsluvh0X9DzKPZWoU6
sxV0LneLejbp9Hc1sXe4+ySmZEIKNATSgDGVNyR2EIxFIu6bOTf2TkvX+thB40PR
ASBMWPLnQsOSGCYvhBGSWAz/2SppPQZsEIs9OHc9Y9rxSPzHoN5U/bVBu/Wie9bg
1t+gAhwSzbsQRBdEAmXhzfD/id6sDwxyx7wsbJ9QNGUqY8y6malWcFlbnUL7akpl
xEIo6/Mk27G38MwdC+HVRAzeE27XDIMlXuR7eRvGU/KpgBNMZPPMuWh1swtMomwi
JaZhlYqtpxH06grBVXq6U/8s+C+t2TvUwOVK6KoE4BE21aqjJu0iOdsCvxP9i9Ox
NieHrtKfOf5zdIkYuxmSlGovm63+aCAqlSzLTZAyEPlqmL0Ua/ufu1+W0lHTFkX2
qDgPtSK3pTLuOBXujqtPMr1+kJGNcV5k0RDGGLRUEfSd658Q+OMnHU7Yl+Wui6aA
ZjolKSqWz8LEiMpXdji9tZ+mSREEpHAXSUgJa50cLG+0ITcmT89dCUTGRLTTtpBw
F+Db59kp3weE4Yb7lM5XqgG/orUuBQxOnoYcoDMJiLEMhKoc9DiA1yZDHbgIrjbu
FyZohmQsf+W6rUKg+hHMQYURr9xfK+rWCMZcAosPBgwe6lFWGZo9NGy5scnuaDk2
2DtGq5zgXG4/sYMIIXUWkdoetwRmjArqaBCY2gWyDbS7m6zNcSEO25vVRzjIecZk
fHl2BhyiWiLsn5+Fnt7nuAJ0UzUBEyR9hap8kCVCBDXoub2xaDXqcfBayplGdD3H
z6+arMMc9XQChE2U+FTXnpuUD+XI8/2tHYOPvo8gIpbl6wkbA75SrlUHJCe5ToLT
Zn2k+TzoIbjYCy5eGcZQN9pFX6Eov3bqLhqr7sHXTZQ3waTxUn2HOfqZjfSOvSrc
R0HoHVP8Ww0eKQfr3jGhSOGzg6kKy8L7Mbp2S0DvxcWvS+zEM7xAmYdqgbcYsNYq
+evRh+8wtY7lYKvszT45MBFNALC+zD9Y5IId3ymmGCnfuILeLeglhm0uv1GV65Cm
EUuevHAocOYCqYhDVtnIjsomWTIBLuTaqYsNJnf4wTpkrxClL3Qi6FWGBbe9ORdK
kkKK18FL2A71CR11ah0N3GK15vgesYEJ58lxiOaiY8XrYrV275MYUNEbSLM1ym3T
SENwOCGfhSdftCEGUhcPgLAO65KNfy14uRxVtaD5mCD4vPw/sZvv6A0qp43gSHpP
ABA62yK1FDCIG8kIIDJqgUwRiLjRyGsn/uBZdIdB75eS8mr7fKJkWfE+e0idSAOj
j5jpqoCpitEDyH7A63gA5q+DSxFWUmIkT+cQwdv/kBNQvnlxl+P2J8eyP4gr0XHX
0dsl/RrMGnK9Pr2O3Xdk/bccCUvZcORMcG3b6xpZBFbO+yH8EVTj+pwj15Whexg/
BKLTnPJgFGooaCofaWQEv2azq+i6fWQdLxqrWOzySfxtPoI0jyiIAJD8c3DUGz2b
sQtaQC3E0icexOBpcx4o+BN5zdng7I15/MTsi/MLmxGn3fAQivK2FsLEBdgw7Mjw
utkZshsaxTw/aXUGRN2WfFgDvizySjE+xrB0tH+SOteOXziNaDaF4Kxqh6oSQ3Nb
4EH+EllFj+ycyyQ+4AUEeIjRB5KXzzUC2F0aVygGA1+gZLXQsdoVptLeeFf5wV8f
l9hsT6DppRbjNzHCHEm5UHDBSAtAWeGiVo7JP3Rj+zytof8MFQ3JSdtLZVR5rOwC
SB09D7ej6UKj0B9lxyqINdLsBEJen7815VGCGBRbXaad8CH3oyFEi/eLtCqgjFnM
e1LBk+S19zXhh1Blu58TiRVGyrz+fCGYwgrlXvLU8q1JiEXh75lfKN+eMoge2Wb8
amMt65vR6cJ2t+lrbxYdHDPtqQWY1v75mlll+Whaq8PrfNSlY9eVGA0UFZ6xH2+Z
yDib3k5T4+ZrqGOz8aqkiZUX0l8vIQXt6jK+FF/2Q7AyjiSwxsT4XcgYnV84IurH
QBN6DGNW86Uzc8tkKQXw2sB6oBzYY0wlAEVOoO0tfzw/Q+3jyc8kwKRuNtbcf/r1
CV0jzSb7RWoFCoY2ebbXZML12OTqEaGJcJECVZ4LXPC0ii+hXqzY8CwflYzYg3ck
KpT7MYO7GY3/823Go7abtyF6QMqUW2KxnauP2V4nhelTUoxdmmuuUMd7XAOhcgLE
p+rDidV8u7WVTQDQC3v3LCMXc1m9zNeB1V4N8Z7T1DSb9BIOzFdQGV160fnILA8R
FnxtrOKPPEEG+do5VN78Uyl4JXkTITVN5cjHlEvXv+8dC8+Stq7MrPqE/2cyZkQp
BtZDzLUZ2sZHp5vZn80moOgXm4D6N1TsD7CCC15xRDiQvFmBedQez9PWaRErdth9
qMPWhTwNHvIrdMi3TzNfJCVBlIvxYsLK73FJfW3f4AjEib9JUXVa/H6YnrZihj3H
JOsWJVDtAPZrmUZS36KJpcYmOaU8FqbSFvsH25QpT53K80UEhEWFtpqbMUb1Ci7C
cJJq/3OzAOBkYNPfwP+U8RzY21L2FiF2pITdqE1PW9WRiQze0cHCwMyZriGMJSm7
rM8KduK8p201vTBkS6nAOf5X/GKUwXCBYI+D3PcPHtr+Zi3hHgnP/D2c3/ki0Ll+
uhEsQX0dmO88z9BMhWVeECpplWOD10IE6nU4yNmzL1F9+/JqKk7vUDzHJnwfl/Kz
tYHYXB/s70wNDNsSNNRutucSM1Nr1gPzHaTTUq7RPknwdEnbn+yyXFoeWluOHFLw
3la08TOx7QfF38ts2V90f96hz6gbDbEHYZrHrn1fW+bfAyU71FQC3ukKxAR6/PkK
wdBDTMH7Od9PybxM3OnvigwlRR1rfUwwk6tzXpjNZ55qn+cAY0M5ROYym3OwPEKo
xK85OdvWKOiZSjnAcgRnTj8ZqI2xPNK3Dg/Wf8F7Fqy5ON5F0dkCOtdRd3Xo3+HR
RhAZcfqU7olbezPqgh31ormDuhpljhaQheg3kUWlsoGpRh6nQ8OmJ+I74O1x11yC
R/of4L5R3daprbEg9yQ4ZQwWWgFImqKpnMbS8YtkOzRgohYrDSl+e58RQW7cvSlb
wInBE8tUzBcXuPSgPgoDb2I7kguprQ6dbL/G8fEMLkaXIA5iE5ZtZ6sStGnnPLD4
5mvydJXUDblG98jpw71P2tjI9XzRdsjZo732MHYfun1dQPUSQXYMj/hejdf1RmkF
IER6XVG/JrIC4YFU4yOX8NRJgCwhJbi49wRLPQnw0x8gyJXmcTBAHpZstqnW4ZKI
HmTVUwuL4q8Ud7AVBWacTINU2W+Ix9CJOdPQh8OH9Wy2iyOQgy2iF7oKEMnKQkgZ
nCsjhackzFV1pS2Hnmnd9pRhxp76ptyafgILvjMjcQf1mKuf2/42mf13F+dAvML6
GgMV1tmz1zJiYLzTtigM8OeCjZQokGVSVfKzyvfmUsFGTLTBbD64ivzJvTFelPII
1CvGtwAsLS82h/Ks/QiwfeW3vCH5TT2E88djIgQjJ/9985tDmHC1bc+E7G7BuRw5
kTew3ZE32ODomlPQSReOjcdi893j6XLqx1LU1ooqtbVF0dgn/BttcIWx8t+jKjT+
8e1cxYzq/AQlQ6thtnySzRmNziWyRFU4ZPuKt2MVlDRmpnqBK/H4nm82J8myIL5K
1xuufdcOuvfK/K/ooxDLmqvDFf3wUIzQ0V/qfKMQr+5cM0LyHeBrYdlFgwBWMMYG
9zG61Gj+LYqw+qnQbsrzkeKeLyaOn3D3y0U4dZPA0svSymN0pTpXW6DmPy908M4A
PK1NCTFnmr1eRnu3fXJIN3cPntndK7G7jiqXoJzhmqfGoN548Yo/fbylumkT/pjR
7QAWDX4rNjXFLntpsj7a7U9VziHILxFSoNpd0p3nOyan8+VcZ1u8lKPW5AFJ7tgS
/hXZNXkjrzr+xnGD761pYsCR4mIyyjhD5L2n5etcBOjpgKX8B4lsTM+BYQQC8J2J
9SjEPeBNQokTvuBaxT+FacLa+d7TqtlkXURyExd3MYvutO4aRsGhzQcY3jdWR2YL
pXIhdoF/YJPRL6l2qI5UbuK0jLFsmJXmLONJ7eu77bZgNQj80AF0oGGmT9zaeKym
DvKWYZXINnEqSn6Uei0YrltZ9+vY/yUDzXk4uR+a+I/q8bp+j0CxHJE277Teyenq
Bjt3PQl1M6205xb5kGkklZGodTMNRZ4s2hV8Tmygaypj8egqtNBFNHoS0ly+43Eu
gorNug0lCDDyAhdmxzmxGqOR4gUDFf/moqg2pnCQ5jaGIi+4wKiU4qewq5puUB2w
6Uw1De/bPk7iZtLkNKV4ADzwua0HOOWxTBx2Tf5yHxDmoSgBZ2treM8UhRxnYZDn
LNw6QtGCKh7kKNemvoFpaXvyYC616gwNehYUNkqmdt474YF2T5pz99hRhvLI+vSx
QgrgUwk1SckbsF0nVrC3Txm9jLJ0XPPHa+5k4uiHGY+fzWtsL0awJ6u7DuZT5Smw
4VALMmfAUn3mh6R5bKv1SsqwR1sCRgTIdBwkov5YZQK9vxzngoxpbbIlqFq15wjG
zSklfUqEODE0G7CfQvQqBLc7gXo60uy767CMLq1zmuEp1TTdYdORPWtxH5lsAiX+
sEFyibS5R228c6P3F32umVy97n00F+4EXXnI0xB2xl95cPIO5wuxhgOvtZABBOEc
4EmvT6V8+HDlYU0I3H1PiTBITOOh7eBHAzpXggNrbq7wctU+YpacQa/q3SXkqctu
3Lzb1EmNOucbX6P4GDi9o8FOHpq/0mfBIKCZ9KqfaIRV4kxt4RaJdkbDcj4PPhJi
oR+NNT3bU08QxnYiw3pcji9j7ymtdDytf4LFeZeIjjd/wS3njDOXeJpWEGEBs+sP
bTqpRHvjz71pDylDDzhq8ZtpwMUN1G4G+cT6nqsZ7YVWLX1qJ2m13f30V9khscbS
x7A7yBAU2kTRG7o0gpNiLhpcY8iCG6xFLTES0tYtfYE/08e3sBeZa+r1j2sWQAzE
654ZtjUyNMxJ8re18D5OYmgCQZHzSiOPaKFRE5DfvMXnwVoc7602Sjscxx0r6Bwk
28w4HjWczScnTvZ8Wjy8ONNLMC1zI3kY59oQjmLMwyuH/XdwNUEWuDt90UMy2I6L
9Zn5ZDOhjsESHv5+CBDK+xMFNTWMBK08i06HcDE0UTTthRDhJEOl4fPKy2DC1vEp
Lwf+JPZOgkoZOyykXUMvwsMMCMCQw+HtG1n5ouOD3Wgo5OjNhHYI2TpO7fr6IolK
QOhRfWBYVBgM7FqHn6BULRV+ZBB7+/8Cit5C9/nYIkzaPfTDryMP90ZXqW+OYAVP
eIKTtWjYljanBe40GrVfprZzhB9yhdiVhr4oFhN6fpgtjyr8S+4N8QiwtMf0Q/KJ
mk/yJ94ZjDj1pLkkQnmuVJ3ZMih8tb6QVVSlmac53JRfeCXHq8LGO8kg2jzCAr0/
Ds3gnreElhq+qYmJqe4mYsvQ0+9TUrWzCq+w19GZHq6omg//NEG8W3P0HMlhYfbK
IKwd5zbPSxgGVmWaIcIEu11QpIXLi7GPCuni5Cy0HhtvgzFuRucaDMdcgX0SX5Ef
AgXo0si662qkgoXNEMnz3o7KXQMHyuxQa/+kkBjp5j3UBqBvfJjIanMYQqUbcexr
zqPRJTsBcoHVodUiqdNu+VB4/T7QYBa+4tJYUX/2owrDf8Vvng1LjK6tzxs3E85o
kYG+pAesyYXAwKKOY9oRQLjpGfz38Ax7tZ56aQaPBp6biUfnICtJd5E6OTjxaeQg
BzvN1fUQBJYbHF1ghfi+Pjkpvp3qjmpwtcY6nMtODViQkvqvwId7U9c3LkTwiCcI
COhTkfgW0XYmzsMeSI9KznCo5pNw7zXvxpO91pH46/gJiqych/KSmR1E28AY4nJa
nVXM/rW8BpJzl3QRQgB784BN/JO/DjXRWqRCyepjUKoOE8AlDewld2wxbBb2SLw8
iJh0HKsNy13DwDJOAQQFoJAQvLfn7oB2UcbQEwMtTZDGrtlJ5YiMYoJhRGwKMbjK
ul8Our4yMTV/oS6491RTdhNIK6CVctcNOq76oiI6o7gDyFGUSHOtIp9jdNS2YQqj
B4wdPD/J2lIb9j5n9h4z+2Laik/2l5U1cH0kgUcGcxPJC83cqH3UgkIe1Zq0d73c
G74LTcBTnJ47VBoJuZd9HXLIQT2YkcYUpLj4mAPZ4E1eeBHQDvELrSHALVBZV+k3
1J9DhJpYJ/5pi2pMaMO9aiZXjiRWvmZ1lftWTGLcyFFmZGmY+vfEa1toSVYA5Tf3
rhThejVhYjt0nD0X0irtW9NgJ/ZT35h+hiTs6WIhz6sU/Pe0daQEI6sWCMRsB+WG
La6JBRJuspeSlMTZuwrWrz0VfMR6t8Jp7JqHYV/hb+lrrqvu6gjxesneYGPulpKB
CO6jvbbh3A1ib7xyNl5E7mViNhvqrK/iz1EoCtdDYGL7npbjKddoHizgdmLDyID+
L8BEN9eldS9WPcUInSQ0x9y6nY7X4EdQomsfOzGHng00PQjiSV/arDCWHaASEU4y
GnS0hUALS1VNuG7lX+pM2hon4KyoOKDRP7uI160DCzGlv/qz9nDs/ieAwd6ket8k
69a3712XZuAFqw+o/tUnt1iENs1yoe4SCNQqQKIxU12p6uDebuE68UjC2HwlnbZr
E+1h4nf/XworHlloT+IOGhjv0MkuO6AMOVRvwhgDVS5yA0oHaaqU4V1UDf98BdJN
xfWjhzD3hTejyB9aFeAwurk8CpcRVS2gyU35FANevkTeTVdA8eVNYrO/iaCHd+8V
XaZMrTOMnXgdXlnpV9vFeeBOqDDHehWVF5P6tZI5JruwoYzHiuO0Lt9zOfRPRKMs
8XZsNoNIjoMUDkh3hwrmdy4OF/VarssRWAvMdEfjr+v/B1Ip27Yv9mpa29J+/uTG
/1dhrz1UVND46wrfeCraXPPuqm493mmYca0OZW4y863vtXIIOX9DwfVcnJ+Ziv6N
YraicNeL54K91vrz/QBOos91Mv+zs5fwmVGGym78ycUtJVPXFadCCSFD/XHMMLba
MdHbInl97IRairNA1ZsCSk9S/NANDyFehIb9jiqLVIz98Frt1SNl96ccV6BTG69H
WE55PeXfg4lXAY7Vnz5UfYR+L8nafmGWFKyMkRPWmTHakvw4oqFiO4sLnJT62j8C
5aa8evPlnDYcF/t4tYYzwmu7VECS/vXE+CpaVcfCYt5xc0wTpI7YfHsUOC8i42Ul
lLrfkTnicFL6QU00UGeWY+cB4Ph07yzRyLbIqrzm0silnvXDIsg1XyAsXcVimFjz
9i2jZI6T5zyEn+ISPmZxK2STIHxYcFS10ABodRC3JOpWVqSoow7cwFhbFH4Wr26z
ujzmMH14T6ah085gwtzk/4AVm6uf0Lw3GvxYXfW5DJSoerioRzY4XhSPCTnjzJdS
iiMU00KHqpQfAlcUh0bwbgKW4Mc7bCoNJNLeW8QbM9dugFz2+fteigqVcdYIoOF5
wJMah9Y+DWGU45DvPJru06jyRGsZKVSVXxloTaIarFX441Gn5FX8edFA0nTdThO9
B5BEn5H7WoVxqKOgVyKroehXz79Pfu0dORbZx/BZkqh7TUIWyQpNz+9K4DGk+Eyo
DyNDgZm5pnKNzEMBwlIl7UEGZSRWXrMYkJYwV6I2qIU28nUCfckypw07HMxJYajH
MJrZjXI4w8jHqsf549q/05eW+QbU28cYRtATdR88YFXw19LyTf5xveqmsqL+lps8
xXH08H1+Tx78bYxrp+cPTGJxUCeccXzxxZabpzpPIsi2DoZjpit0r2tJKy/z6JRV
7wnQaNbE1mC4zzRd475cZwxC0LRq4RBi1sUa6/9nnlNDuLr/MVP6dYi0Q9dcZg2S
VxuKkxtXP4CKl1xX0fJjJDZOQEUIZSFiRTp2v99aaiXq3kevKLqeK+hh/axoHZ/z
NvBETZ4NiTI2VPQNIUAQ2oeMCvuoC4HKxOPrhx9Waix7geIpjRmmx8bxdjfrSDBF
WiTSl4yaMr+ha7pKIv4i8U46R+VPiHCT+CBfWTwyPP2BCEAHwIerAdHuAn4sDw4n
8Jp6JotzLf2sqPjkhlxiDu+wpdI17c4grtq7OzG5X6CBAI3inN571DIfS9uAv1Jn
rjaWnRXucGxpDMeQwIovABi1EGZ4L+5U/UEOIH1ajPwsRe8xd/DkArGhYmG+2Lix
KoIW0qN4uky5t1JDpRq2s4kDE0p2AVbhrg2x4D9P9Zhrvc3YadPMc92ruTWjtdHt
cYVXQqLGgOY0JEkGJlB/6T8Fopm4YRSc4FfI0+sIagx+GXDZ0vG4zhqYtsF3G23Q
YeZbZVeEelcDgDqjEenGewHZqqxUdTJoQoml1WwdMwRAdJShcd0Lmsh+fc0J2AhR
DmdWbtgGWCOouvpvvrW5vFd1McdeaThSIhchvdvthTZhHHMxD/fyvL05n5nTwd8b
t1oqo3WUsQg0wArHlTgEpkoyiuW5UATqDgH8b+LHV2MfqAU0q294yBc/14UgHYGF
7W1cAkiUYcu3PEqoskZ/PZaiN0lp41DLXzsMoU+0kMuMtryfBInSsJfzlWllEx8p
fzJWYWaKhKMW1D2lSeC3doLVkLkfI9+kfxeCjqWXhY/NcPseH1lfvrZkN5sZGI9F
qImMTBGccXsb5yPWLaMDPORgdjqdr1foqBwXbzt+NvhaVbvW93z1ec7QHeZlH2FH
64sa/Bz/dFqRlT3/PxTYlpLWkmW+Le6hBmx0kmf8fXQTINq/zgXCzbMO3nleNFrY
i/2XttJDjIIo0mO9gJPibDp0Bu3kdWl0ZAJFfxsrmUPRAU24dpo1VCLav3ZwWx+6
8guEnndbM//rfssUzMpQ1Ox/gEc4a2cT+pXP/7xd/hm+IYS5ORc2fo5pkw65RFZf
KPE7FQYWnxczocNrOIUykQ7pr6fjq86wwP3r9kFq1N2viyAyG+sekUzz8vxKmJhd
rpLCE+LGBXTC2VhCZgo91uZUznorEHBuQNCl06Y2Hgc5PP3qlrmfj+f77h+t9CJK
g0PJtUyQL1p9QrM3d8ZLq1LVFhJI/JbbbeJQqWBvIz2KrwxH0TK4RSozB8fRUX3U
c4T+J2s10iEc3v0Ph0Bp53RuXCb4Aquk2oili6CDLzm/DaBT48Ap7jFD6klOP/zN
mFHDu4Gnmb5ckj7f7dU3a1YG3EsR/wndznhrQtHFKJWDKoM5AisICP3BuBCC1lGB
McUSZCgXKxxOWeT3+/M7PQ3HoE91jeLLd2sLa8Hyd/jttsWj4InKEItkphI8+2Rs
H+FuWYVP/s+lF1rJPO4RFSoHxefYJqpa7ahC7YzK0HKTbataIGg3qDh4qLHxj/zv
1Euu35RsyzMgQ5qPYVD9sFSh2gGcVPPIVChb3u1WJSB0mris2nDXARLQFsYcq+Jh
2azfCtDGiiHXd5TudvVOn1TRczRqDtj8kfPFd+uVenyPSUuczOE5ZMNt+HtbFQq8
5KbG/YTww6JVVBsKxd6DXlsX5wu0j6afZM7lbLwIRf8TKnFJlcs0W1ucE2oot3HX
8o16xNk9U6PVAq3byn2j8henp03CQ3wM8wXkraAT3+8g2aLjSp4AS679m6pn0MAE
395aJcYgQNVENz06czjUaL67KDk8spMhSSQzKKGCSYb8pkC1iOsKINLLFttKF9/Z
wIr+5MHW6zqS+JebaT8hlg/Ib7ggdLt8eD+t1p51D8MeiHilrn3dRXD/W23ZHho1
ba7pL3xboUd6LgNgRONYaM0V8NefM/yFFx10TF6wHQTONMlF2zE7gdLsT2ZZKeEj
V+8JTCg9xtIxyu9zbMEGBvuoPmeBBxX5fknEAsV83KI2g387eSKAZlIOXU9c4ka+
IcFIBQdBhxzPGQ2XoraZf0Hhdc3YEdCxp4OU9FBaaBBQzpmiW0TAAIqHWj+mCG1o
rkNpzGR+nGx97MCWdNYeecd6X4YNRhFlIqIb8vB1CODeC8oIDzyakExOvBpKjEpi
zIcA9WHMwb+K8xrmagLHbdpG51XD5hjg+xJqwbMdsP9Mu9Kd8odqlUo/odXf2aR7
fD0FpKOtHBMSTTC1mmdw+Ox8GnuBKM9DSUmMm8Ai7oqB9Mu8Gc4pOSFoc2Fc4vYm
DZafiRaQPN6b8KwSbQl4lcykzc5jrEzaCy/Zsc7vlcdreP47dFNui8HaQRJto3QY
eHvKuTqL7+oUSoZwjg26IsAvENZ52LOeKRGntUEZMorSJVsKecpShNpGPRq8iCgQ
R0xqvT3W4Syg3vX1M6v3XqhPsNnXCNT4OGahL3AO1VO1QD/7vXCKM5cCqqSQj5uX
bKkCNoIvpEle5ecyrcKND3jKW5YGZiuuBjBCwZieI5jEpowjuV6BWHb4zYCI7hsI
O3FebYOtPgE0NSoylE5D5ZCSOTpR4sR5/OfbDfFQD9DlOSWY6UfyY+TxVrhh5wBj
AiziwvcYdAlfXHDGxj6Up6xVCydPAHUVBkVMkn4AbyU=
`protect END_PROTECTED
