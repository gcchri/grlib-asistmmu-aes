`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MBWAtBwT5YbuD5I0isuvxRa1bZsfw8nfboRdlDqozENTYrrzVoKF2v1fbWdMQdcg
Yt+0j5krLho0iNSCvEyHK6MMhG6Yj7VJ5zthV0SJo5heOpB3MUBTpDlmult0yyVX
4aCriT9reNn6yeHEbBLi8i+BBiJhZEKk/ALCcUJ78p8+uPhn055x/X+sIoEsvUb6
ln8hrg/s8rdN3ohUXMu9Q/+k+KL7557/GXVF5XXGtRYSd1cnjkIspfo55lRN4+ED
+8AiY4MVaNKiyv/eYPIHh8QbjgNWxNJrsKfa6kS6YffaheYPbaCfO9tf2FL3eN6Y
tBe2xFpzCLXRPndRrROhuM3NwSVD0zlCEWInCf2u24ZlHQYgrFgalyRdLbed0YM2
+USdcRQ8iilKas08k0qLqjG6LLrktGCRuclUzmjXaxL7l2dxieUQkfWE3P3DzHE5
+iyVaL+D7jPNZ4LvTeBfVyP1XHhbyAaCejgDnUUgZDsBsFErR6X3C8JjfWfzft0o
cNvOqh8fyMiwuPOC2X1z+Q==
`protect END_PROTECTED
