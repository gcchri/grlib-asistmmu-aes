`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c6KC3sZsSLSFDXgJyUbLlz3CH3cv+6uOIzvc2celLx/idqRMYGam/BZe3Kq7BKbE
GHWM9ubMq1DaEji8zyKhn9vYAC4fkidV4woMK7hlav2leYkHvnfLJbeRYTmSfV10
mPeIgUfL7XFqg0ouV/VwLg==
`protect END_PROTECTED
