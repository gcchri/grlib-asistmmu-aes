`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dR9Sy69yZzFkdWfe/zknzBVjTKDk4lVtgxthkk+jgqwVV90pu+rTtdgVZnYncWvg
96H/6fAaHV4rEeNzq73aiUS2cs4vXlgR9K5xPWnVl8XAAkQU2n6Wd7hFguvKk805
OV3JfCsSNcE2Z9nTjM+IiT4zT5/rgzXtXii7TmPLYIxnDnSeMV4w52hreaNY5+Ij
uu2DjrMVZCeVXL82yH9KwG38eDwxB97/S1+Og4V7D5EVfgSzMNgLW1Ec+rthgi7c
x87MG1RUOoBG7k9A9d4Ms/nS1hfBF/IrkoSL8ZdJ6B5Je7ASvFtKR7461/77HZ3S
9JayTkpULw+syXVzKyzMtLIK8lAs8OpumMTXL66g45VumLjHBsQrt69nBXqgcfXx
BMPeXKvpdNLByYVWPAWXqMzytFB0fNnQUbaA0TCwQF4NXsijEqGSQAKieil92Zzv
Li1HeRiLoBL5vsdRj9lD+ae7nK0pgHK58Qq4gmIBuxUkXBC7ZZKg1/VwV1l6ZFnV
tD/IQF+JqqlE1bEicHkMivJsCydLX9kqVBMUx/F4s6RTsF8kAXjpEY7xnCQjhOPn
/8fojhIX+uYOxhggW3EWe+38YbFma8w++dcZ7ve2PEV7VmnYaGWeylDgaRJA9ClO
ny0zj7sN2KyyxFclkqjmeg==
`protect END_PROTECTED
