`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
353j9S0eTenhok1uzhEhiDAA90GgiN9agBtARqBnhNlZP5GmeapCRmslrT+J9wMs
CeMZqSVw+A8Zu1IbeCiuXl7M819cWSv9zPy6l6MePBvl3XlaM6ux+6aMgDNAUzQg
fel7AGjGOXnOwRcgNsWgWnuDH4xAFfobleMEB7rFAARUGmIBCErY+/nAtEtnKDwO
8qS+B8J7qQzezh+Upqy3lS2s24uZs+WmFrajxeSId7y0K5c/jF0Z0XxI1UGOs+j+
LWpTvgRKOCs/wYj7n2jlun6r2NlgRb+QO5SkTpUTCllv5n4mnFVvBkL2G1MzbY7o
JTg7NmB5paRxReefbru3KGqNWPUdxzQPAxVaeBCnFFk=
`protect END_PROTECTED
