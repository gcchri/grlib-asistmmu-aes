`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q9AvMqbr9aLTddEVLbUAz8lQ3D0TdlW2dkeiZdo9TRxOa1GUI7RLHhw4glfWsyRo
KNdrqHRw28XhGJd4Rz0qcOirDYO5oa187qWJH3Cjbxy+mwskseVQq5SALDjzqIXV
CEuBpEeDon/uYur7DNn491tDCSKIv//rVcEUSK3nPsS/ZHrxbf995KCkldelHFfu
mY/nKUrxS8CO9NmL6zhlyqx2h9qd9fEYvRe6kGEmy/cfcM7D23KTGyhXoWltiN7O
SzWyKk5UozcqAt8ghInuMdIdebZPb5kbTD64XHo0bVqbC1hpA0Xf5e/VIJFqYXz9
zP3zG+EsKNQAOmkFBxR0b2HO+tzUeWTC0piy7KX7G2WBzY22unjHbdLTZQ+tWtqn
8o3RPiHQZlVOOTC/v6g6uJ8V1ilW3akKal2TGE7wytHaDK3AGQTbUqA86rNWz5Ax
iou+qvyPs3+4ILNpfw3crXaICSFfRSLwixUkyWthO8Wy4QSjSQQ53CohYBXkPB/+
qA8d4x872eiZObYcprubWwLrbtadrldjyxR1rEKE3i8HIhTa1LZSvvJZYImPbPiI
TYRXgF64LpF2gPnwjiwZlDekbhgMaw2uBP2Hyfn49+G4hPZw75pJZ8lM25gvgapf
`protect END_PROTECTED
