`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i89Azs82ekOVROGKFxSjjSuwa4+YMT82ku8dSRe5SuuNTAA259ZMkwkEmlg1Id5k
nRQrhrtThxbUsPf6TUBiUzhFRZEH/eIyhzXEQvYfAaQ2oDup+haia149kHcthr9x
OLcrMbD4v8MrVyyxKz486t+qhXek6OHVyfVEhHZlb1MnyxIolui+1xSsgCJBfnrp
vpGVZkJvHosnrC8C4GCghD1IyyS6Ia98HhAQXU2ATRB7LBgOxTwHuz3hx6C/5UU0
Pr3j7aeSzx1HxRjG+AnmHrn4Ie1bcL+ldBFhQ8oB66y3yk//r4fuUjTcs6SgwjEs
a6tr4EUrKr4XadLdB0seEUWgSfCtp74Z6gLJted2yfvQalOkKOEQNBhMSlD/UyY2
`protect END_PROTECTED
