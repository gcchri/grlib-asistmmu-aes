`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wLdMO2kBQ+1ZZt+Ka7tD7HtoTkjCyuVS8GRL9nNBQwc/yYbSfjL+nIXuwztLjnpY
s/9oIw+euakMxHBidoBjqGZSfBxouo+sWW0vaUry+V2cOsi6mrFVgtXdEl0YOuPE
NoAdq6uLe0WBzcZHy0y+KVx+vOXIUFgczMeDyYUU4dX9dPXB5UM3e+qt0dNWSICQ
pZmwvNJSL/TxuZc7xwwzGczLAb0Gifv+PaUnke7EBtuYy2FvNUepINlgmdbQccGX
0qTpdLmXA5h77oLRP0VVu0RPzVV+M9zQESj9+vlBhpTruXVMOJ2SGAunYeGYdRgn
DrD41aSbxYjeCE8qo4N+wP1uxRKb2cdMVODsiBbSk77m8HCQoHuJ4zLZf8z6WtwH
CwdXJjEU6g1/rGmkWn2IQAYJKnE1/s7qRAwnNyRaOiQUJlpDmY2HUnOmGGW1QZLy
5W+sK/1uMWJOSy0+lWbae5oddKdZRE41qB81qBykaaZ091FIG3zogFX3yOZVYpT6
bKOQARuJOkE2qBq54oiCWw==
`protect END_PROTECTED
