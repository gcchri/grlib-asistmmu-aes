`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GyLSghMoZ3g6E3I3UzvK2QQcvJlYoZzbYASPv7yPeJZ03gnS+ubXMRUOpyeH2DEk
uB9YYZC2zT9fm38j2ZRbFZta8+IzLLs1dj/lmMrLUOjw9Y65H0uBo4JKBg3sVxMV
FExgGYe4xDGZUpbPCN6kEYANQ3rMG5g7HxjeOThRkKb+Jard97YcnQfn9qDFQDsq
G9e1PtCjV6adaZaogJGQR9IZlvWp4aJfLGgZt9QqygT5EIGiC4wq+gRt9UlcZ4fN
424VAbhLEmO4vZ3sQPHkJITJiDhWxAUyWAlT1yRXZXn/vF52EeRN/1sWXD7f97df
+W7E8xoIxwfHtx1I/+Hvx95gCZRQOPbzYEQGin+6LUhsjYhBsdtXpk4s6LnckqRA
ArOB/S9/Suw3IBp24xTCl5lP47wxYgqKSqljwtXmlgmW24UeK6339A5+7NhPCJKt
lRqnvlMLwRSsaVRUPIBZnhYsLm5tu3n92cgUDRRuMfuqnXsk2samIE3SBzVbSe5I
Qg6gNRf2SfOB+AxVznSMv6Cd9UFaNKMToj4/BNvyjaDREQWe2YyyRLZ2p2cKzmIp
JSnkeKCWfEhaKR1HbDXWBgOQEROt9CZMtS8TYlh+GyNH8sU2UIXlpDtAjPXDDGqx
W+5y6Mhms72Rcm0l6Q7aHAOdT1LKDP0QRXeQGLVEHvHro8+wGIAVAdpdqsKptHU/
I5sDhswSDpD07D1a/bpDRA+NNlAtN0s01CkOUA01H1+5MWiMK489hmQUUOBKPAPg
TEFEschY8nUw4DuCw95yKC4/KxJNSDUBfl00NakdzvCSzL+txm5mG7dOnMWKspcn
6/Q42kb36M4Z96bJhk8TyZNKn86fpu8bytwt+l1gJIa7N1jbnGxeMTQ0UVaBWwAL
+2fxpylUd8tVMi1pnpj3EZmPi7OtrNl2Y9Lc9H8OkrL0+AifnXggoWXUByfpPeuk
v9PNxJ8mvqeXi4/5ub4sFT9viPPgl9FjQYzourpMD1xn1eH2XCiSmRVm+b9ZFbiZ
1nQDTj3ehKlCZVKPjyVRv2BASAFNdTryDIyNkhLcM0TlKVJT0Fuv/lWTMJGgszLY
/rO6qCv1tps2FaOmjsLQWxmBELnnBMBm1Z8rsBo9+lVOCApEpnqqmOkPz0RkPVV1
5Gv910DyHl0/QPPyyOZiYUYFt9dQMg2T5/RcbZbulkAKTV8NDsIyIfKncM0XpLAP
LC7csZttWGll8Qx2I5fA8nlXNXwnERe/gowvJQWdftRQG8QHIWB+QrKtsI4ZYt+y
jLxRfTKIkm8MR+4x9hmhdj64L17w07n7BYuHfgLGcKy9IkC6PXnvlRevEGDSQvMz
43UxoC0sOjdCvXueFzqSQL9lo+hH2KohQ7HrAtszbs+kVM2uX400m2Gl2zXa9PDK
ua4ccP0nQHPIv9QNKaw1A4Ts1/25e8yUKjxX+fwfJsCWBTRySunj1YsFCx31jb7p
e49jktbIcfZWUwlRnSF2CU3W3uvkoRildC/CIWaZRvcS5q6+HO2rt+Qkc5NX4fv1
TcUio6j2UmIUX7nRFqliB7958Yl3FwNzQp16mRWvEiy28b+IbYfU/1hsp1jICX/g
/IFl/HRQJ3gGBiwJmL5PmB62CktDX9g3OTyDKo+DbTmzJHaIO3nTcdujfZYxvsbw
M21a5RYMCOxSDO+LZDvp1sW7Gxw1440eg5+zQOSk0B0vQm2HFaDitU3+8GrymCLx
hiAy8tzd773wNd60FC7+HCXfYKHKAOjPqvIrFdtoEWAv6z9XnlYcTJ5OcnvEKUN9
UR61MbS9a+IkSeI80vnciFYg4kxGN7J5BtN+cNleiEGILw/zR3Rsd4PVGMQxMyKO
gwzXX6zKRZR83YxV3XeTTKxmdKFl16akCcOX0/VZiWy7BOhY+RtsSHFFHbIJiEdY
Pbu7mhQ2pIx1pRrlYtLAc3IrIYgbAH+7eSFqHqxhgR47qtIrwP82jdX592YiHiBb
OTBBow8QAvd09cWMWJ/mFIDP8PiZtdLrEH+02Mk9jh+9Jwn3h9bIWPaDBU8U+KCN
F6O6GidRXQwJdO1mU3cSHEOSxMCGEOrDytcePDrCK7A14F64VSuV3NrBhJL0mRtW
bGoBDHK1ENMjXpxrXSATTW11X0tBkFdtPZWSghkyPMlOyfvZ1eLrhvZZHxX5030F
rfIpwchLYUDX4LuriDUg4nAwC8Opi05os4Ct1cR/zLegHWPJy4fWRC28P75x5Eej
JfBBF0ucDvXyNOVvDn0G8jgSJC1NudTjpTWrHlyTWchafA+LxpjYsuM41x5+N8NZ
OIj0XAb9cUvCt2QOII6Q8OBupDA4AaszWOxKAjCMNgqjh195Gr4//LAB5tzekHCd
Bt59VQUlPZk0w8bgIFx898GHHk2ao1AzqhA6pRQZrnnDlHNmeufEKv9KJemNYAy1
maZqW3B4ZI23hmBeji0wkNzD9PxusmDyntAFz1LcHnb8sphexWKXRct9vJOEAJ9a
gss7TRt9VaWfWZjzR1IFwrQtXAibrUPki3LQZ6KxaQPMrMb7nM1U9N2ULIUJPvhm
KdtP44QEN9rIKnsI/dp32tvCKJt6aahyrp+ys6lOo2dzb3Wm5Pujqooya06gJyZz
2v5eyXzeTPtpzglXi9B30lw6iHX7viv4JV0kZa5Lmgazo6+lGikbcpjm+XG2K2+i
wLNFekAwiqfwF93G5IwK2C5BiRhOZ0FUKFExYyhdLNpDopc5ZjZFC7HwGc5sjBRv
Y4MnxRIARap9aCRJJF/XaFAhdT1hCJK7tsaKtNp0anho/rQKKc2kJ2aBbmgtZ8yN
hb6sugGpOLXsPto8xWQIszr0oU07XT+FfvO+PRK45w8lZOsAEbGvKRrDxqQAXZA0
3L7qOXjSNJXCpozd5N6qEP3K33qZ7qy/XEaPu6mbR5echl0kuH4Yb6i//ZqEfWya
RUBM8Gy1ly76o+T6C615Nv64D1MNF3+37V6WLkD3n+U=
`protect END_PROTECTED
