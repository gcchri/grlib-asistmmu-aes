`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ODBvWDuEf4LBO0rw4Ae5hnAyB1o32Xl0fU91wdipgIBRkA91Hfthm8UxucdSn64S
OaZGenbNG+z1EVZ01zT08cY/Nzf6lPLpk7bGn1Qj1Uve/94JpWreamCDGkLS/yqk
YECNn19WdzImIqc+8b4YjN7PW5liGDwJEDReVVmVJsKlGV/nK2HxBZvp+rn+FxCn
68cWksYiacky9g7uttI6Tv8PDdB8kvSwzksL+WI6Ug151THZmMW1CUZx98q7Mvjq
`protect END_PROTECTED
