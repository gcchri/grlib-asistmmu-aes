`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G3QJSxltS/0rx9arIXvhI0xD2nmDB4mPhLDCVgbCKayhhzgS1a8iPWHurqdUt04S
bQtas36CXXyaEcjO5+2HCyPk+FVq6hRsyxadnusGOrXdiPD9O3yN7X1GmJWCIRFz
qvdU1W2tLU+nSMXdUINN8o1hYRBtn2MGQP9gdSyRXHjVXO8GQF1ET/We8R9AiYa+
fzQKDjx/+URsC9whLoc6kiCbN9rebQbd2qpCISO0KeuP6NBPlm4zfkxJ/pcNVzwi
Y1hhlFQabvBqlL/qDPPrQvpKss3XAsdWzOCSduka7to9LhXiufw1pW6Kxojh5LlQ
eGx2AjiNv7k8HsGxpnC9RItNYhxNLW7GVM16fVL2KRvvLbHG57pR50WRFHDIt7kl
WdPIzL1N0qBk08LY5ve0N5uA36PkCvG2scVFnsIMlly+UO1kYeKyBb4ZPpobSNQK
LLS+YAylkbDb37+MfUuFx4tNcSTtX1dXjXlfV/KrKy+ELya391A+PyCgLCx0YUQ2
5WBXC78I+nvpwWSCwFNX6lIPFtLmULUezdB6q3yYyu8Q12vZ/UpUywdl5N4xIo6v
CUj50sFXFsEeEvDReQtVQhrZz17xC9bKc7/eM2ZY8uNnq0uhQS0VwcZErTztaYkd
EYnHoa3XVSl1PHHVWUjvWQ==
`protect END_PROTECTED
