`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/xa7Ty3W0TCBAPA35+kS/VovnItMmjPpg6W6FEIzzjYRplYaWjrxIAbQoQ5ZBT1N
aTYgb3zz5sQ9p3+uUqvnE3B/zAcGaJZl8lwZZ/hK3NMU5j/BmM4CHzuy7CzKaKHX
xCaAVbW50XWx4XvYb9kWZj3oFL7ZUR9FGz86LHWe4rfc+ymfSOcoFMHch1XI7ahE
SvwcISSKUY9jjD5O3Ee/UamtsZaJyQPuCNibyGWkiKjUZJ2gmfm9GNCdBmj837By
asUCT83Cqy7mKRdZmrFJgo/T/DNRfRwcMUof8rqt02Vi2FQSrPG1p2bhb8qwOd0g
uW5CwhXP5Jw32hgLaMGOh5aO7k9NIOailjCOqV/Iccw=
`protect END_PROTECTED
