`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oYfP/UWXxlzoAdR+iYH3oT2J9GDDgEpMYgVeHqMsuvBpYZ00sDSGqD1Pb+zTyv9a
OwXk+2wO4twQYJ9QIEhetke4MSyyj5xdTqEOnk5/sVPGtXphufeeIytLlaZ4Z60k
Rd2OZysKB6huF6HlEE0DaA4xxPqQKS4Ri9h5y9imJwp9ooKrwR7UPZS7QYnvHFee
T/h32kphgP3kqR2RGulhYD5IjXtgAxYRTDHGZdPiln1HC0K7e8VH5S2jzbV4KUo6
/na/sXJnyqKijgW1FU7s/Q==
`protect END_PROTECTED
