`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rITIA2eXPORzCrvbs4Z0k2Kj0o5I/FMI0UsIkugMuEiDqAqk0bEpFAKxuOnGL81G
CBx7tiF9ZWnNAyN1GV2n52/ggCA2CdGcrpoD9SvkGiIQ4/aUBqfRhMtaONedGIOk
U8OdwQM8Q6riTTQVu5S3Z9rdIbeFiK6RPkkK0XaEd/AgSV8xLDDsWmNDFoPqaAMi
KA+O+I0jmucG/Q3U8JvgXJVkLzmtsXosCMuC+Pf6gMZYRbhKTZpQF6f0nFbnDCMv
AF6zW3/FGztQgOVXtyox33J/eP/f03K3mSiu7EAiRTjAiYb1pEyaFoDDyB9Afz6W
5ZxLZQaUjUOf8gqkDdSUb2SvIX0jd/RZrfAi2wuzX/V8QlKGAMm8FjCoh4YlZErH
/2G2EjurWYk4o35Y+8xSu2yq/T9Sj+aVt8o12w7dsx+NRbElzopy7swLgdQpVbid
ELtyTWZa/aohRpTmBD4rnmh+uDqiHT/mowgIsGD23By5gav2xOX5B/PqVqJUHn/J
mUEiX7OeLsABHM+6lcrLEQWl05By6QDFsDSTKcwFl+v6ic1bzW9d2Qt4z4TXgnvA
HlE7IUCb23JY0A6hIOq5lk91SfPGOiXA9BhxlC5tQKkS1kPqAvMj8Jd/Da4QzCab
yGLiMm5ZLXNLRYQFLKX/ycEJ2jsDLQ2HB7b0RDkF8ukVNFCGtxnytcpiRaTAvpLn
J4PhnYuymrBPpbe/9/cZb5S09vKJVy/+uEJYXj0jm/MpxyoqhS0DLNswSQzLFnS0
Y8G/i4UMPxcqnpn8H4gQHlT5LRo2gGXc9k2njiVKUB4ro6no3NY/L9vb+R5ER7lK
1L+gu7ENCKjEt/DO+fIC4wLy+gI/psuvwP6vga7MITobKZLsoCDDIFvrRtu6XVRT
2VAJNScgIFXY4cyP2mBFYblJS9JWAn4dKLCAKlioYeNasMA8As3C1BFf9/PM6c2L
O4X6WVJFqRTjVb0lcaS6pZ0s7V3fpMsoseNlrqmp7Y91m3UvRAksVEEBu+NNdtmN
wPa08n27Z72SwRUsf3jXNorZWOfqPUtHPl3bjI7TvGWWFjktPOCc7HJFrU2+992R
eiNiaVcu+nu9tlU9F4gifDLD6OCqJgEUp4tX6xiOjsMOs9AogsTpfUYyKNWIYQFE
WRK/FBe5aA2caLOpdIOAR9rpGj55TX5oBwN4vxkw/J+XZHYrGo1AgnCs8+Q81PJO
Od3czeA3KKrWT8tuOn+8OUZR30TE481MT+/MkXukSu3LSsuyX2sakLugCgB9C2RV
2ZXuJpU8IbKGxGpxmTLQfQOzWILjSa9Q8ucRUgSBqLXPQNRYcgCEgokRciUQG1br
FcbR1s+4tgBx2cH1YI/sMTVRtptcdgxlpE/ZB+OEWqDoOGrQH7EoIPea8BEqFo4W
uXjpajc3Y5hVyqXGSRHoVjJOs0mvI9FY1j4iTP/lGbvIyYckxScHg+uBqHYq4+30
fTVfkluyU0N3IhX1o7hps5Yufwd2Bds8cDdgwKi/UHYMxKPGlrVMO8h3dzMdHi1O
TeGu+VAz6RJGUdohv7hY+KD3ZxyDzwExaMcmFf2yEji++iD/H+Kl3LRN+9eDl2pp
ZVufKzpuG3FnKnzjLH9g7/p4noSqWIZw30BJ9MzWQmJr26OQkzpQu2GwdHh9nRUf
9E3Nwz8Fsq2Azb7qVvVK/RYvOPdmNQ04ku9ZDnWXQNAKWcHJWadoExwiomj4wGyy
WF0L4r1tDJhseU+KldQW5VAUUlKptB+9EPqetOZqrwgRlbM46o7gRbY7hpzojFi/
zGO7b4wS9vYdKd/0Mg+jUT6BPbQC2Os7Wu+KPsek6JLp00e1aFtX4WIxPIkTuaSE
RPcVLE9N6woyx32THM46Gi2lTi2OWnp5XyJgieJsFdpbRghrEM7GU0hLE4o3Y2b8
cfnqPcsolrNBsWdXklsqMtgHqhFhP6QdAIg6cn9+nVdfTsNUVkt5Sok1++8fSCXN
vbdYhgQOYUlkUppIkufIW3w+nV5XrMcdFuv7LqSpxSzApnF23tKi6tG2ePxkg/EN
YWN4qehr8Lf7/NUoE0JHGa1Dl8H71c0vJKCzabJ/7IGW1xNLCB1hXGm54PQXRDRy
ZwQsqzatiQaiVI+4G6WL8VnjThIQPSzZaOBUPUAP+84pjZBqyTv2MezShlhmc0s3
b3UueKTBO15mlL8EzyyyGnX8QYUjGAXIUW9gWo/33FYEgf0UJJlzlhS/aLSHaxtE
juWr1CkOBloBNhSe0y6TMoIDfoXVf8P9pBF617LRHH+X1eZwuB1DxWoe9Z76xh7t
KEIXrgGRMf/Gn3hW7U+Dg+uVbE2e4oswKFqTK91yRv/CpGOWw9271wEfw1B0GLN+
tvf3cIAWmGI0Rk5yX0EMyDgVrnC/6Yo7mnO8fc2DyqWBgMPOm/Ssv54hxbvWv6Mz
L3BysBsiJlIXJNAUXhKpBkr2ISpcJVRAISmrSEpVFgxigkdRMyxEzNGPIy6oLZiQ
zeqHoqKS9lzyycAeI0ngB4TapjeHLZ8dFCxvHD+hbYW6oOGElqoiOH+te7tZijc+
B6KlyGcYbGLALLfmUHfnILPe2Wi3PtXyhEweEyhQhXhiqETYy38gI8tWBSunKDfr
Vjl5YU6jZh9P/kj9iH//cyeVBRaxW4Cx9ovxpjN4Ej3q76MY+qc0sQEqwRjI8vw5
Ajk1AbCgR8R/JqCBUVnNRMN6DEki7TK9z9NN9oTELxO+nEphtFy/N2lDOnPxp3k/
UQScKk89DLPC6Rq+XNG4jX9XFDUAuubEPpLJuyPUC9tit2yJytEHHYSAlPObWPJm
2wi2ArgEvFgUVxTKn3GS8HDb5V3xY5+ptuQzjGB6QsqUf6ONFVgrlDeESd2NbzQ9
7bPuwlVotOE983kQvOAA5Gq3+adLFhzwV5Uj4O1LQlbhnnvbgEvgDXjoCCTlWsOz
xct7vHt7EhiYho1er+HUZya/JbD4tVsiK1RoqYsaV4rPzBkuRq73l3/sItvpMBM7
8b6cARCfw7h/hW4m1O6CnftpW8BpLROQ9SyC1eBkQHmnsnXgIS22KiqSn5N6zd9n
qaSGqs+rF1JYalg+FVAX7LHXn7F1pnmuQT/PURTBKMYDfdctRiZvKsCP8j+Q6bov
sl5cPqtDu8KH9tWuqjAE+zRxNl3cx0Kx5TBror07k86lPmXYlT8rQ9xIBx6eSZix
yt7oTkyKum9WbNYMPVSrSHUtcREVmDRisESLH6Wi5+B7gLty2que360+mkKz9dJO
mS2bMU1zoweIUS+gMHm3ZdB7X/jqxundpPRP59iQ/5KsLvC6/SektYTia2mm3XIR
RtH8IyOy5YZ6ymwx8Is702obZ3W6ej/lwYX4RUguDe65yfudvzubWchsHxrDITSE
LyNuEh30FQdxphjKr7jNOj2U32zfU0erQ0sodjND36dMIbP/tz6GoMxKeYHd1dM4
+ODsM4hr4gOPKezhobsNx5/aUfMea+YAOpJTLlm7I4TVLxfwdZ6Hivoqeh4dTKzP
qUd2c+EDqT7jW9zDPlYrt06l6yorKcrthwnc5r6IJdE1XxTiGlaaCcXUAw1eDiKe
+9c0Au0M9e8H1GaCn5eROc+mq8rJGl4IylrEJ98HOH80mWuf0nQIbFOij7ue4KLK
zO3Vx6ItGXMs8/03Xjw8sbib0GG2CCAw3IBikpMiDMAQQAAnE9o+lp+RERe3Yo1l
g70V5pqmysE8rAgDpQ+pPzWa6z0Awtlmq9Ge2kFkqv260f0nFyc8r9Ipg7uapwES
Gbhs6gc+1wWzPiZew6EalOHhYOZu2UMlFAZk/0LzYpGQbtAN2J1aLu88CXERDT3e
hVYEbJ4CFp5UxMRmgiZTBticnRp+uffPr3QMuQQdxpg3PiwVeOmq/dnVIbCmp+Ka
8k70bg1XLnOxSDbzlMiPBAyYnr376ggRCECSglbs3qbjN3mZjx74lhGj0xe51Mde
EYCHtidt3J7dlUrhhv5rn9MdErx5g5GPjNcnlLfXuJDj2zZt5aUSoQB81Iy/3M2w
ouUP1PqpkRe07CljYKuxJyHjT/jvRALbD/YuyGjxbweULri22moYZdKgJP79rePF
qVAuFgqzi51VG/SbQyc6KQZNY9aeuZ2hKuHg+iXfLuV5LdhXPizCG3JjPYG6xPYT
4TNdd8RXExvIXpX9lwr3Vb++l7Ut4ZkcMA8OJz2WO7U1KYnBdfOfNHJrssBvdXv0
yh8tSCfYsIlnKCohKBOCYxa40kVjwLc3GfJrQD0qhB1Z9sM7UHkuRzhNEcNAlqfY
n22sUuHPK110TfT7SHWhQfMMPh3xU56N3KvGfcPfjAEdhEEvjvmujBZmvFSE+t9M
ranIdN37ih4aihVzWyECBREp18a0lv4owz6L/t9wPdO3NwdnnFVxbMicVTelWz5P
MqAqXapOVupJYefQtozA5/haD7HFSeLmyT99ejNsbwJj9JJc/fOt6hpXczbf60tC
cRmkRvPOq27PnKGUzNFir1q19Gb7obom262XzTk9/s7Yw5rf0hnz2WtBo8KdR+kQ
KUWN44OoNwlW5ssXtlL6cZVyXgwRqH81lH+Fejirj+Hdr6bCY2rZK5zvCCdm8l5v
mAPc9BLYaIguzAIuRRL5M+3VcjbxpQ9jTI3tVYwkR4V2Eo7t1OfC6vcS69ieNnAB
Wcr8y/vkHpYTpuLWoLMVAMo+G7U3eX0ncQ0ppLua4V0MFoOpUDlixcWHOIINYYuu
pJ9jEbbIIP2asyY3SJYWKUAdMenQOmz+xSvIvCECdPvH6IA2WfIUj9B6YC1jRiVG
Vf2NMafLSjmPokPH3c8CUNQPRzhQS+Akg3Hbr9ibWVjiNESP2GV6WmzKppAFkDaC
I0+8HJVn1XHkbsU6uHyfK3XGu/zbuCiJYljoLXF+PecJoTL9zfyCSemwtRE/8zRb
aoIr83UNwDzfMxm9zg2wNawecs5QWCfOOBLgXWkFragQYfavVtOHJwPbSd3cr3J9
vdD5EQmjjqVJAR2aXpJd79p5Y4JWphx41CWbVUmqGDPjdHZEiGYAR91FoOTh9jtl
GYew/NtOJSEqnLUjOhRVYvCnK32lClWS1OzO7nX3FzltdyDGArdHq9lUMMqrv9gT
cL9H5JyZm1by8EdhN7vq+e4x+5Auq//CRY4Mi8oPtZ3n4NH8Xz+rQaI4K+jWWqHr
xm3VpEW/CwrrYwQfy+nTi0qK+i1aCYjtN7X3keEfoO7cMf0pkJXZ0MQJZWwcCU6h
DQCT8eCGB0HvEiRxCzpGCsYA0v95mcKrfRis1Z9kMZzMjLmXG+nybDz9BDjLFToS
/Z03oDk6VHd6kBrS6WDG0wM4M1cBMhnUxQHO0yJ4rsVf0fymgAzmmnGNWxZQaQ6k
8dIbSCXR/KyREoxxh+jFA+e3hZagmIKbBxfoltUAUeFgyRkRWSl/lZls9N9ruAXe
AKi24jU/C3ZnRWZbo3beVWncPauKy43N5SOBGQKBAgV6PoHZMbGUAFsZnWR6x8Ta
UQK6SClpwa2AcDIEx1hBVJOP7H5L9yjox9YWzsGiOdKCmsbw7RP/MiR5QHIL7ZWB
6YqW9pFj2/mLFHdKZHWLgorSkhGF8Js2EwCToHB3V94L4F6aalsnPlokv1kGbqX3
9TI1Y5TmoXN2z06TQzsLoed97JoaecE0rDBUjJ6qMr1yaUtY8tz5mHfADKZ5tpNP
K9Cxmeju2A8MxZhwZDQtp1YLyy/LEDzN2E/Twh8vmBSmbxO4mptqlDXDEBCI1Zg+
8ziZIt64YJEP3mEW/nejYGUp4mxJIDwOyJWIX6Oq01tZhAjL5a52B14x7SvIwFMn
9OFUQ1ThdgESKObOVGwx1WUxYmtQesOM0Ayu7DssC0bgmyX3+gomtu3prPlOwert
tJ/JAc6Owpc8TOH0zfvO4vm6sVH/2RMmhVN1iMGJhtq+3v+wWvPyXZQfSm98P4/I
ttunHjOsUI67nos6i0eeIMVDut+7tPF2dn5nPyrIlJV+i/ZzmI+67Tp8AlMTXTLE
AJt/SVLkY/LRgLaNsUMQHmOGEQMEpGL+Br4E6HoRe7fiJEwSaPZDCsI9k6bkuSjf
D4OQCDBPuHDfV+wrsFHudId3BVgIv80Zd1G+1zOsv4DpEng78zRkqbMbf01AWj+N
QFJKYcsOeyWfpE5lzNtdQziBMbWVKB9LJ9ul9rL9HZlqmlSTqmeinvIdNqp4JHRQ
vm+UUrZc+6stze0VEUOHJ7FA2/mA7rdMjZuLsYnA+glXUIIMybi2WJcR+RdQqZTv
s7qJZVj+6AH2SxAmSfPNVOVsZfufCQfXQ0GRga/8r9VeXzOMO/zrG1VAqgUOXb+R
TtaKhmLm4GXK4A4eUfNo4H0v+lcIR6gXZ2nlVIqtIcb83tsYXUf17nkMLApTFr6l
HC6RtGDqDJ5c8y5vrZxk5GAzJWcLzLKwOdfLrFrTLKfu1DzThVC90BDV40dt9Oi3
/ezorHNJfDSq01Hr7uOptT+rzv5XUtytPoH2TZC2hL9ybHp7E1LXJVo/D287oyRD
UL/56qLF9j0pbKWbLAybXqPpDqto+hClqPl5EdJWY1m5fPiql5hoGtg9Va2Pugue
Z/s/l/O6y5nQe1RIn4TEmBEq2gZNY9zDYjsFwj0yRMgdc6Tzm1kAqhwKeVboNvDq
bmpz5xj1ROAMR/SQ17zU9cqCwsj61V65fWHp7yVbrh7brdbJ2c0qF5zli4OwTvMy
GVruWVguIabzkZqMu+gE43bJsTsj9CRYiGFN256/12eh21Jb32+7RzsZz4kA2u4/
GP39wcA8CrAt97antFmq319huaYI0RiX3xDtzbS0nfalolqlAlniqHYNBrKsYPwX
CxWWApWiIDSKsdWa37CnNOjfjS68MTWPz0bkybKclpQrJHtbujzB3Af/xW8htpIJ
cJePNbq13kH6Ld9EnOymqdtSjJ9+LhmQYDvE02sWW/SDkEQdfdxi9psQT8re+Prp
1K4NmHP9PZID5Q3ZLpS2O+TTHwpllofudzvQWp0A9+SwcwGe4YZhjlmCjisJIc58
bApjAzDNxuFiT0e9HNSZ2gRcePMPcBY9o9TUHLxbdUA/hAKDz0qrsBHc/zQkMqFQ
rSIGZttZkJt+wNWbzvwqnrZaT2JtmAyTO5KVoUTe9/E+P7UyzMUvRC80l2d8SzDq
6Tmv+WyADHtxx9MZWG26uk8WQNpVogGnUYLBHarilN55OPX95wRImswb5t7uDn4s
MmFQgLB9LWVaYHV6mp5jcU26ZZ6E66DQQ3A3nY9ZfL31+i9QpygMS7mMGUYN3V+I
aGTqQDcQjK0I8NqUHZzcbr0AIPMrhD1CNkgwQdHJuwSBwMbNYV6zJn6cgYh27EeE
Cbc+CtqBZGl4CS3EAParTg/F5mfaYJsG+rXJOd5PeXr1b3cw6d76YhTg583rgVlb
daYdmn8m6G0VtjJNM6X/W+KRtf+Jvi4usHHsBABYeGaCUXRFhs9agabGHvrkLAV2
6WucgoidLhxX5NK/evYXmWwb46/1LzalIIOfc4jlwigjaivnNb9q+CnO1SG3Tvit
LCxh5xWpzuYvKK70fXgaR/znx6RpYFtMspG/xBH5hfr9/yB5unT6OeoXfHA9/4Fs
C+vXiQyYvl4W/e4CpDPvG1ZMAQs+3UV1MN6gutytMLh6exQbSTk59pbYB+JxnBFF
2uNuzdBHVBBlw9LyBYNA5w1QI2Z3GUlUd3NDar6j5E/LXXOUg/3MT983cGsWFgzA
ERYQypk/pMCpOhJMb6mdAlOzyRRPxkuZldnxEbHNkTa2YZrAEp0CpJPoO2ZbRqF7
tjhog5MgBdbh2DQmwoF/Zxkp8zAtUAbtvboZj7W5tjxvo1OgWXsU6kJkPIOLBe/a
BDFXlBavIX1lOz0OdYTlfLJVffe7pIkgxAXIRJa7mNd3oUmeRU/1tf0L/UAeXLF/
gpqAdqdY6dR3mPzemzgKz3SIbAvRiH53Y6btZLXebKWpD0uej6ViCto82vGVwz4M
g3M8jWNnI3klC7z05zwZEwMkRK4ig9bHcr6GuIxQM6MYTTQc00ky2JSVJLRZtFoA
s2jPlCUYaLrBcIVGhKOqnBtsx/0wytP0GvkdIdtUjp2M6XfuctKafQosOcfH/AiT
SplUqM23XIcwRCsN9eSwnrYFd7vnsXPyUcm5lQOb89Bdii2qKX0REeR3+szLGd5C
`protect END_PROTECTED
