`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z5vR9ud0WhWI4rPWrhQXsPeklWDLcdi/B9/FCeC5NSpuT/wnXgGsRFJhYlBXCB3C
XmN1K8zCFRNQCvNd7NL8N5X3q+8mBDoXFCOHloeirBZ0li+C4VgHNx6nWpNBMEZ1
TmWV6ezDX5EWbYAeunSLFUIDVfctf48hv/EjySFWzVfW9hEUWZYVmDkYPa/v8w7X
TeHzIfrJB9k0qMTJqfOEzyNBZjsn21h+n34uzctNCkZOTcHD1ktJDD0JeUC9BVBb
z520iYYY6KAps2IHR8D/t7by8fmx6TUwS/C8U1XvJToKKg1qyCWlOXBiZxGyGxiJ
PxoL8qr7lKPmU/yRKCp2HBDDrDDxVa9bB2le8r4086VGhqM8J1KGr2lwJqZtpWN8
anzO6cpqJPKr811QnVJ9soweDQKgQitvPUYXTb4TLIVFJjFgJvzUZya6ce+5Z147
3SV6uUBlOS/OlFeDT5wpCzRDjo/syDbP9lz21/ZfgKRI9AEfcM3lNsF8G5pPnmB4
ZSiOn9ZwRTuBGhQgdA2RIETu1cYqtlQ+3qd9zGe89461ISfJ3wOG7ojDb88zekqI
wMz5yR/NTOxQRGf1KXsUSqoy9ffByiYtt7LJKzeQR48ycWFffnu4/CWS+PepIYDa
rJw20lH+rcg3m6+7io91TNpphf6zHJfd9FvGGWgpHBV2u1z8KwX/tis9USE1oP64
3W2/M4ueEdgdZyeb3xiThHzlPlO9e3H68xrcmHjszwBl+LsaYqIw2HeXcmGjzah0
a3/W6D7C9ca8nHbdy46e8tOQsNx9PoKsunGx9vdJiGwnyzkkN3D5/KcBzAn/G4Ur
3ukbyqJqBz8jaesRNLJrkw==
`protect END_PROTECTED
