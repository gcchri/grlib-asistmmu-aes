`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w7f06ygxzutZJIwj80YphzyugUwrTMq4osURYN88EuBMFdfifrIE/ZnYz8IZsEol
RFfegz3qftckiJ3rB9MQp/h0n+HBplaY9OvwxZu/+h+Faa04KiKu0ED3uwlW5r2H
XyF1xYoSjMGr2rgjz8pyOnDf2e16DPJm2J2kv7zFs1QjffMUlWKhtaNniki8wXQE
FhUW+WWHqVsSdyFIXU0Zx+YSPe2lW8yWEz1RMB1vVyOkqE/4OYf1qeeoh4aXNJ81
0f+XDdUqeTWGb/GdDt0A4UM2xf7hf8j/WY3KaYph/ZNmW5FVH1iu4xA3nYfHlAdR
Z29pezDAnmB0DIZj5lku5OHnVQEBAmS/3J7dFksWJjEh8eO44pX8LthouzSzwdRf
4beYn5KSgVZplfAbew70gUHO6PtSErL2JtNaVHmQSXg=
`protect END_PROTECTED
