`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3iAPupSvBR8TAfJrCMc+p6WryDFgkwQqTo6GtXZmXWmsRYF753mKE8YVAn9q9TLQ
Bx0n2W7pxNZUymLN5knybZOAGakmBQQiQAH9iGYQ6ahmlu+Gtm4HRWPeenz//cLU
DH4xjNN+wLx8tKXBVJWDY8r5DUpEVVc2j1Lx2WHrd9IikrHNq7ccgq7xOTr2accp
jYwgEbQOj/6QTQs94cuyizf2s3zsFE5IBbPYoC5kqNc/NrGOwqFtAKMJLoWcx6iU
S9b33UD5rK6Sp2MmuP75hP0KyIcSM7xz9TNBhKeKjJfObNAeYd6ArJIVUThieoi7
NbuFEwtf902qNSkP/rpdbfy41vczzvnZKi8GpTDHyiNXbZe5Hc5EK2HPGkOSMgmf
QRfNlsiNPLz4rTtLryu+a798/VWCl4lD4A4OQmn7NAXi44aiuU62Ta/LsEfL5RaE
YgGnhJgjwY1nqA34R1a1GF25O0Ax9tfgsY9iD4l4DEb19n+2zRMCUJ9gXy2RLzc5
X59iKIFDalZWojgDPbDZWfxKY7seOf8R/ukBvFfmHYYfRvn89VNiIgKP3XponKRW
sIBGzlddT3s+A8ceyN2dbw==
`protect END_PROTECTED
