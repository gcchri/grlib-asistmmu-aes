`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w0cEIYfgXvkJXDhi7nOFPf/STQfdamyuSF5ZXNDvTqkcTk/7ecfMNHOuR5ag2Ukv
b70IdWZvIfV4IBXUjWchLYoGprhx9nIWCIukVc9nibSQiCMIyvtyOdlax2NnWkTr
A1WgaoAn3E0mcKNlzI+CCZIt6TC+RP5bqmBSz4b+nUPBbsNfdIML1M89ej92OIPk
F6Kv+6UDk5Bm/T8scuKUT+bG2RKYRM6JO9f9qreD54+28K1HCr+dceRe1WWE7XTb
yDy2OgzrBpoDlL5mJ3sgX9vDqXYtnDZTLeDT/FicSLmMIShtYNkY785ae8wYZbvQ
95PsNe1/6+0BGoYY4qiwSAR2LaFJycbuVapPPwjunUSFCTPv4WYp5KK7ujoLSy6M
2lpnnEg6+DvZPD5VqgHTVqXvFF36MjVqcPjRaqKF4K9dd00V4aJHNebhCTwK+ERB
t2Yi6Gi6oh+/hjo/rI0ELhLdjzxht2DwelaA/dGGtcLKYSjgXP65w49GOpbkp2ib
QJ0EmVx2E+qOiMqkBliSQkGnTualgNHox20rnt4Arl37qQ2+upUsiPuDIRL53lN5
/c2I1RGxNEzcLVxynW4Wy5MNyIBHLKf1IlkTpDK6oZG5JZuZ1bnQw143AJ3YdNiG
ZafZXuLR7Fn1xa8LkZLs47SzRg2qTmwW3q3fQgxNrjsB3HRQvEZT6sdhAc6WeL3V
uYuUUNoTxYd3QUGoEE83L6mFo0buMNJRXO7Ps9HzyHIbMHQ8EQVOmm2FKOu/mn9X
xJ0+Sc7lj66qLBTvwmF26g==
`protect END_PROTECTED
