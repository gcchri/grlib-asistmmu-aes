`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ICaMgDpP0ga9Uy0hcfW5V3oa29XdbQkUojXYMNfUN4rDO0sM5iYOfONwKjkcm15H
nMCYNokzP4TePc7KsLjvNWpVBiw9JO26zry2uO3Mxq/oitGVyLTdGvr+7n7aMSft
I9ETYxKfqyhZ9nZZD31xtFm0n3/y2NkFGIQTt+/9uPzPqHeXNlHonRZ3CeqSW65e
6F5P11jaaLU8syyajERSTPwGdh8dIjCremYWEdip3+A9uiXVfBgRcC0Nbtl1LwcB
cq7EOg9YocXmSBrfRzhSYstkiUVwuNOY5y4Q2C29fsZhCLiZ18L3i0cxo4pLK+9Y
eT7S9X4I5ya0IZB3xaG8YLwMRTrnOj8Gp1E5oTbTV5rf+znJppB/w5g17e9bPx2W
jMYRKlairhzb+uDTVEFV2XfhFcZknJ3P6JPeGyuseyUwOQN4lNmfm4z3ZF5joVsw
G/qaG0F1L506kvv0kL2jvzocEkp2Yr0i1+JVw9hsFhJwDKn87srvQUxETbzSZPGn
Hnkv06wef9u66iDdCMT4J4Sh1nvP3ZOP4yTqJfJU6EdXGB1I4SfMuHSz/tzWFMsx
T+vFjBDSHm+gUNZoQ04yhmilviTsttfU34R5Lnsx5fajyDHUmKJ+Y3v3X/hw6PNJ
dcWbhmz2o44bjNR/X8RftKK/yFSaqPMDuqlPgdv6tUsEuAerD9TtIl9+8w9wj6j7
5q07SI5GjbDqIoAC5yo25Q2rLd+wcH0M6ER6yklg82t9ZWBzWToCNEf6bDFIWTqa
1izfd2w3qt+qHfURQte4+R33AHgTAy6rZkfZ5vnjoXaBTQgJj34IC5cOv66SZedB
kO9NG0wq6VjZvmHN65rnB9bbJJHUca9bdguRQ8sI8LOw0t/kKpd5bhg/OeSmrbuW
yiulzDHumA/cc4/sy+CGy2L+jVUB7n8wN60ohx2b+RGjYFqUa357bGaFHG9uyvdr
duAhpvJLN3ji7c03Otm3QNeb8bw2BDpNKQ+GNkHaachZP7427VKY2h/t5OM2in/w
oIesRtq07TOWbzQ+y14GpA45rf63daxr3pPbiEbJZDmoxc5npVH8I4fXgJdiLidZ
Rq9/ZDHhmnbzBRIEBsKEUx2o/d9Hu6b18MHzCLrFpaR8LxgGhDEnwbwMFo/gvmNr
KHTJA8VoiLngOo8hnKNES+Sq+g7m/K3Ccq9Mlg0GG0QrJ6t1rwSHAKihmqowHhzQ
dI3j4piTJ6LRWFlHZ3ZvAmlUOJImiNHprMA43WUOaiY0mUh7zZP1RYqNUXaMLUEt
gN19J26BuxK0RjbsTKxYMIk2H7sDfpv2YbXwykvy6sc9U3D2Nz7jIFPzJBCbpstA
kDj4QtMm5CpUk+qVUxc16ZFCyDTI2sp757ai82vV1USD4nzpTamnKxHjKcfuImB4
wbPzRQV92qHPXG9O0cufSdhlFDqgA4zGZ+gGwfjOIx7TacUjiYUTvGJSM8JTAEHM
WGa6MVHoATzL+fmmdEobq7sinb1r51O6L7FfLIoa9vTPeziA6/ml1bMXR0qAVe6b
Q586XamBw2QadIr7aDPaE3kOdG6dI3utBeFGp2OdSgxdYB07SsV/pmPdH2k6aDBN
yy77X6Y0VxJM7fkSqT0+LNAzVPbVVoiXHzvpx4SFgUgJHCfGJpg0gTNeJBrrOk57
8vZJz8u0UtRyv9VFgrPmwfvqVtVBv/CQP708Puq8LXq+gUi4t2F1xmLymmHqZI2L
RPYNYTUI/FxOV+66c95t3AtI31cAwMytkzCfaRWhGb3USV3IyvQU+ZV5TjBfSUY2
+CBhhYCoPkvoAHfSYMcBXjsY7pBtBJpmoXQdv9sv0wIaiZla/wnIZST/NdvU+4LB
TT0Izu9yek+P+E/FxJ8w7nGMYy4LyfUrdOTEmNFS4NP5slbLbQGXXD+8agYQ0NoI
RaYRUDDdG+OpxSDUIhmtyw8Uie5Ue9OAtRrEx2nd8ofs1nU7fdBjO4piKnInRzO5
C0uiIfPH/eUb/JEWYFLk8rie3s3uNv+9meFqkRI5sTjqpv9ZqwNrqVGSzV8Kmzhm
CiJpO0Bhvqv0GJS4Wplo7JDDn1vh/yXL4qa2g53XjcXBRyWdHVCGVdaHs+kgbAE+
tsWgu2qaLmRKeXtLMWr/VL6ZcA2Sq8FKPvu2c9oQBL/eT4GV2I47kY0vcpihXcYC
bfu1n3xH/veRHphOz7G2Y/i3mx4NNUEm+QegpFEVEsURHZh1eAZZ74+XQADFib4a
YUlXNcRaTm6upF7MNsYon1bytvlCWlG31Ol6q41+ip5EYEcWeUWRsLbs1uUwmUvi
q5NQKNfoutv76WKmbq6LTb4qwZu6NAw3Gz5hJSc8sMwxhhqOAzKC2bawQcaVOMKI
AnsoxuomZkOVF0/lnBNoUDst93CtJrYZvhxeomjJwsTocoDRZkpWWYsy6kdh36YL
6Vyu+rNoujdP5jYEOXRJgg2EJfwtwKPgcSQe9prAH3hLlGwwFmAOXmZS4mkyhAvD
MS6Oj8sa6LihcRn3XR3FVLWTP9qkbm8jrKtB4Q0n0GqpkKwI3h2OsE6+9h/Ecopv
7sz8fPOQSu59V6Y306kPqO8hIzPBk7BENrhnm326AMpOciOeKzYCjGz+ty3b91gq
lHLp75SU3Bu3JZji7izCzCZroTjEZczz4R3SJZQknlD1/TeFrjTPE0/0euuwjxiC
rZpkhaRk1j6k9ku8AmKoBPApF8gZ7nOZefhKQ33Hg3/7XMaBUQxyy5S9DfmPQMdj
gOjOP00pLpLWuOk6dj/uC3Nqh/LOoAxp1VH1fiImeTO+8DduJCdQ+giPekRVNKXT
BflUOYxBHKu/Q7PLFjIPGW8Zb3NndCPGEhGcRXQ6gKb5U/I26BC5u5tTy7vkDFD2
yhqxkxGoonzCPPry0Nf1pPhTVpsUhRwauD0a7ejK5zIRZBOoehSSvxpg9uLs5FMQ
iCqXqjC2k8VvIuNI38aDl8fu4oQ8nIL4RI646y+LHcFJbt3eywthveiw1IW6sJiw
EG6RoXE0UdsA+v+WDj7o7iPa4nn7/83KnD/6uV3H+GfpBU2QM89XEChV5JxU5oXm
kWkZ8Bpz67QpkJcmVHFW6HrwrYh7hvC+b/FnLwgYwcy8wqajmO3+D54KzD6XkgDF
OKy5WAXyRE6GAk0/EBAehslTJwTdNoug91vlFe3JuePkBNyxzd0aHmHHVU2Z3/BS
KOJNxZVMsK93SMW9L6TuMXI1tosGfwiS6AUy6krL3jcGZmadTNF7YZpeA15YGYw0
LOr+5jxn4GlEzUO1vtfSYlCzXv5wGpN6Shv9s3i77sriBOEOZ7XNnm/UggRoaOow
Dp+NliJmkCQG1gYUE4VUP4H7c79NIu7tNoSUpoN/rJWRw7cToLeLq+Ntoadj3vut
pm8sDh1hEEkAzOLFtNXGFgUViL6Sz4EeVDyDHIOOmqDzmUlb7+Ur+dRB7iAQQgAm
RiOrekbBKJEBUhEA74S32xEgY4tzcZ8cB07RjfxMeSbmEVXu5KMS9dGfrbVtq1Ql
8J1ACUAeQ8xk017xwJmezfLzxxaGT7IVjUl+gqHr9nsHqb1VvgmKZJ3/naVosEVs
uMeBcw21iqsJZyJtf4O3B5Wbd+IlVfTzp+O7XWlrpigHKe6mZcLsknKF2LCYNXsS
iSnzvISn8CFL9gq8xMdH3wsd0nuEgZRQMtVULjvVHuBSTDVirGg5rZm9M3l1LvZ6
qMjuPIkeGdqPO+81FZX9bV0E1Zrlj/Wvn7TJ9Qy07CKCXB0wqe2m/HUfZy1kBGBW
P8O522ZVwGKjhhAhNYdyiBcxfXALG9HmXN5Y8l4CZMp1h/UF/iC2iAR6EW+XVJTf
xXpFFfGE1OYMhwlrfWCghVOhDKH/zMIGeDSkHQuZqE3bZLILeZN+DAMMgFdEM5aA
CeDT+N8Oju/hJY/5HZUU+GNLaaHFQSldoVDmLD0rPz2JaqNxm6fXrC35OxzSibg+
+aQPMUo3A3OF9dNNwYzJLXoRRHJaCrqjrcAFSEdfK9y+dldGN3jBam/P39rerAnF
TTRMx095HzmYr1xTCHiGCkVKCyI8dXAAuGtbpQVzBGxFfTXJ3MOqetjma6pxYMgi
RkJE9ydhs0th2MXRawI1WAJZlzWGJtgawtNT+lqTrMhtaLgT4sIIwAOLVIdd9s1q
FkGwrrXOD1M28yDTpZ6YVWQuczWMRT5FPaTmbJML5phzGK6iYB9TuOCNuHRnCA5u
a19qEIPYVEBilEjV67LPtEgSxVHLzf/OPimWuHhrWV8VPSgI7lZgtYlDpnzSt5yQ
YeZ188tSJ+XW2Pi3WgZs+sGsWqZyniVA6RgzDGyNiPzCGh/iGdAuZ2VGAOFoICwS
HzTobq80M4M1BLrk52oO78/rYOmJVaqiXIRYr1rzbWRk6GH8PUe9jAFP1qNYgdDE
i6vo9dQ1rJ4npXP27np0GsfKl2V+3ncQuFk48tDG69H4XNoUh+2UGU3u2KeXRKsu
i7a1KalFHRQJKPZrv7fTiIoZ+FsB6ze2PKqvSIUETu7r3Jozx6VXI84iDevVsY8e
Dgy9LstqTFc77XZSOMHg7KHIc5ET91kDdxYBqAsGPnqAb8JN36+jd39vB0qsjwbo
AoEEBkpo2Dj/CL0ktt76KFw4FeN8FlvtjTLSADq2RpuVo9IC7+d6IG06EnLRYQAi
Tz3vfCOmzdC92+1LM68gbm2VqPbf2ek2zuLBbFRb4DPbIoVDuuEb6NAn7CNMMHHi
hGuHLCJiwY2UXYw7zXY7RQerNuz/VUR/cyXwtFhc48TVhD1kojNErBsPWSxEYP8z
08uJJpsBmKKhf6b6H0DP8kmk58Lz+eFFI9NGiF73PEZmN4WRWH7u4AvneU86nkS5
tRCbVTQFcw/UpQqViAfizijJ9S7YO7fINyg6SmSP5deRe4vIAsDGapeKDM6uCuM0
iGob0Jbt2iByc14PNdFpjJmV/QGlnFCxVHur2AVI4BRPlI+zmU5SPocglUfh/lMB
qWLchDaZ1xdHM58u0hIH8/Q1hxMh4Q7IsOLG3JIDkBfxvFH/KN4zo2rveP25MOyf
J3JRoBfdYVBfghNb5LcVRhKQqAphN+MaPkNK00MX3wPBviWwQFoY2NGiNN69YIML
4i4AeNCOXeYaGcTs9NHjkoR8fk7GfR9daWnHgDRa4MNAHJOEzBallwMPbU+QcOaK
xYgPbFmw6YTq5kBluYr8rRjqIEg0OAPs5t/BLFOqca2g0T9ZbNqZeNJ449EZCFKi
Zkrw0Ns6aAcw8OWYH1G5MwpvGHvnzEulG5DkSxVQs9EAnz12orwZiqaVDnt1JqJd
ag5azxm1MBqkIcvUV23reFgO3QIoco3HpInTCtHDPFy1HyK9fmfT5FxRBHCOh8xP
Tv4MVywsUBOHHQs1u1ijUDZGN6SGlNVV7LEmlr0o1HOZPhuXwZJhH0e4QskUH8yg
+QejrsG0dTtFgvWu8iCgxbrBjG+MYbYj+nmJGCelqyskAmiQSuQLbnmtQmekf7DK
zSffKX/hy6aCFeFqap81vcDfmVXRKJUXbiovIGlRnPmj15d1z0Mp4cTI4ckLEFro
ii9M3SL2GzNOtTNGpB/1zYpHPgdFJIKavvhskGVzyXw7h+qJDd+ChpM4w6PyPQ92
TiIgDM6s3XGj8w7qCGEk0/9G+vRCGQCecjykZGF1CkNcU5v9W4pADJmMHwpEh5b9
1LlzWokRNFw2i8tfnRWjVbBvyeu06mbstfDwa2GsDFz4wTAQeeLbHZSZTyF7pCL1
x8GpMIXdLfOkKypHrCbjhaBtw7XWIwyb/LrVOxqJxjQlaAzvMSGkx81NnodyyayB
kRMWcw82HV3a2AW/VXhC5aWVO3uu5cBOCU/06Zux4WMpFSL6jDrUNILCWkbzZiY1
jvPxYw56qlic/rhwqRKn2k1LF+Cyi7Chyg6u+aXvd2nqANPwAzlG6aHyB0t0amcy
VrjxuVJS8eNp3AA9MgwucR2xALdfJyiqIeuMNsCTIS0Nb/fEJv7814rysFhNR1V2
Vcc3JhsW1E7URTG9F3OHSmUJKjiVNHbFsc6mqJVyAU+ec1siMkNO33oC2wG2APx5
pyv1mI8mDy8oymB164af+cs8xJIOZMmzaIE2p4LWJlFdPR57AJmzMLgaaTVvirbf
unP6tfw5OZuLc/Qf4ML1V2NrUjoBD5kBkCzEWXEHau2ii1Guq9Uw8/tp2JGTzoQ8
ZDrGoX9BAyp1RiR5bLJXbdE56dVDB/fgp368L0Dh4pRdi5SCX9cBZmKc7ld9Wj4p
AaNPlLRwyBdV20Bm1ShpTvijnax8yENnObgJ8755ccKPD4Zy8Re11CW4JRrEihDW
uQucJSF43xY6/8GlYbK7W06Kax6XLhsBao/ObVU8dQefFcBYjnC2rzqh93OcpDDz
06f7veiUqm1UWTsFQEWO+Qh4i+wWIvo/2xfCNvZDog42HOJZi0cHy091eBjIPEsP
YxRObxhkWRgC35mcFyIi5h41C7NYNFFwbm2LDDSfT23qaK35t9zuADi5xe8tkl4J
xvcR3xJ68E5Q6QxF6C6b0d2VcSkHkLR/8iutIjQOre2sKSZJd7rstazzQQ+XMj/h
0U66a7fzEYg0OcrdWCmgTksAs2P0YReGITHB1cC1c0bZ10D+CilXALxR2AOuALNy
szV4CQP2UYNJhwXHr2QV68v6HfFMWhfrasLB25/V7T0VigOcMJKDqh7xcqaZCrnz
NEeuU8oZZdy/c0z2A8UBus1/tJPzy73D3G6afoCxLsLcPUIVlkA/+gMxuxsGFtAK
91PvvPYwaFtZs8b2eDyYBVQbbYdT8jnFabpv363Pvt9LTVevGC7sWHvVDZARLz80
HpYScNSL6eb6PwNZLxvhwkkO3pOjExCu9ucetOlSu0cbmhO6f1U7jSz29Jfvphan
ddJ4uPUvwIMpWe6cBrGKU0XRVwMlixYi3cjuNUNDOZPTBdZK7uz/WRrCITcK/eIB
kupJGfzPCjuKWuOL4UY1idurfHZPHg1SZb1wePADNSu6snYOqgQXyKG5yX+++BqL
OSIaUJpa9SL70hiKGEYzPS4AIamfRCMoxVRVOGWXsgBDm7xIflE+onT0wjLDwDM7
hOCdUuNZlQl1NlharULS/t4oYcbh9Me2Vib4oUQIDvjRNJBZHZunJ9Vn7Eg3Ig8z
ZjC87HOLko/W3zIiM2gUm6hHWtnm2a/9NjFYa5w7WTBfhBlTiPfjwnhiYzOVitEn
/4vv4u1t9xoxzV0C1Kty/9m1vXgrxLEMgMRUSpQ5Hw7tbUMiDdEi3APTZEnpZ7zA
1kdLrgBNwrg72+bqw2KCvdQk9ekCZXlRgV3aLOB7ufUH0fZLntFDRTursTLSx/D+
cXQGcvLVZ8ArEWscgNgJzIN3ltAiR9QDofo7FtQoXHd3X8zzGLTr0dQrMf0MyGPC
PXEdvkGXr7MUk2CfcahsFo6EMTawLRYOHrJDw5dQveinZMLE9Oi3zp3IyWAObvsv
ONVXXjyzgqONwgZlgXywX0n38bFadFydCN2at8ISoj3e/RIWHhEGashbNFmyodIt
ZiVIebj3HdqY7HB1kr/To1AAUl0bUaBzH60mJ0HsUDJVveNl722UOu6pMLeQNcaN
a/Qyl8gA7qBWVvDc3+PJ/kRGZOTPKzO79B330etoiOvLlBk3ATX0Md8koXSF2VbG
oVrauOqIuz7GXsHPDMqSSZ9X9bLo6lirBqWr+IqaGdeumjfAHH5ReCEONaqDOrcf
6ZwQ3nTCKC1k63p8OXDa53dbrhShPgI7uyzP4ODV8r+5NWN2tTgazJuhACBF0q4A
keozH02NoobQuFEPgPGQFEdVelx79SlbRdDTdTJUZVnm5MnjqQ+XiZ+JvhI7Hiek
F3JKUcTVBb9t7muoKwXJtedi6GTo65LJu6qqBbdaDborNHtngDUdPGV3Bqa3LEwp
poKFILUdpWaXaW86dt6WFDGLfjKfEaY4lHylEwn7Ig+oQ67e6Qu9fvEMKdUMi5mP
baZhnipGUmPsUmdi54FIxRYhNKkokEXobt+SGqadeamMLlgffrxxybD9WJKr1XfQ
3yIuApDM4jnYNV8CdedRNxugh/kjb1Tk9CXiieYvc7NuqNNZv9P7JQRpvraWN1Nb
kqD3VrFJxj8+1So0WUMsz6ReBOs+wOvy3hOaxizpaUXw73Psnx0reWXIRB6TBQml
5qCcQVTll5PhQa4x0b30EAavpF3wm83DljFyu57R8FKkAqKzSGzaB61Vaq4EtPeL
8t9sEN6TNkOHurl4d6HVu7ct1MGLZrENw3kFvtW7DLn6ILCPvq5QJqsVQBmBH0I+
e/0RKy4Dx3mh/HmqsD/XHw5PD+vghMpW8X+Vg8FvjUrDkVyNWLh0HbBRQX7oh+b3
e//INZ3NBZ/aLhCBi//2tiwaqN+vv3M9/dgVfgL1l5PePcgfBZRD40o3piin/Q58
TINuQJqKim97yCwNnRgQlbI13/YdvuTo+76fzpFCLNHZ32IBAe0RJf9bj8hKgh/H
+91tbvCpaxo/DEZ9U0o96yxRgmG3Wuk53VkuxHpxH9054kwrDuQqA2JYEm0VtPUn
Vdvg7fjIYQBhsmSCpFv3Z3U81DfW5+CvQTrRjBYcfaDETXMtoy5S+QCCSQV0d/Et
Z37Vdf1KqrVyCU7r49xoBC9uM6IXMsbH/xK6mn8Nuh2RhRtYcApTJZbHIhsv8L5Y
5TfnOZLuOxhySrXQ/GCW93Zp4GmBRILXHAAzZnlx+PYFcQYDZm2aKBHY3hN1EYGx
pWQXDhXtdY8qk8NU1qt6KLxsdWfPmh0LolLsLgKPoBSuPkS4OQThlJGgtOS3cCrz
tUfQE62JrfxkV5GYzseQRMAJYW+S7KvV19lyCghyDYsPsxhKRzzJrXYKQ4kjVJ0p
3Cp75BW06YcUooHrDUWARLUUev3isp1voVRCVCzTckhkRy12PYGwNIFHw2eECMod
lpGDaW3hzMLne2hA4RDKv4NDBx9+Fe9fb6m9A4jpS+2bFXv7maIHF7PGpY/cscwn
qbSvTMDsjAHmwsJi6SmYOqdVG8H9UJfYBjhWqlWL0upD20Tz8LmM+OxxOBQ1aG7d
pdoH25VslAJTHtsxT2cb/LvewOUoqKHVXkd+ZfbdDP6LYFOQr3r5aD/3s05CJb50
fAxCkBmK+gI4l9bXsWDPSN9YkT9J5UQ26pbuUj5ZEtjHkTguKo6N2LdZykbD0zEe
3Hq8UHEMDssHJ1SFlr70nmwd/SEJscycKunWiTuSuvZOdPDcArN75lL9Xwu8N6eY
6MNYNfjyJmGebr6gaXYG+lffJenuQmfjyRiKNK7WbpbXO93o59UpZCSTh29AFdZm
yIA+BetWc/tOmrAwaHrL1n/WE2FdrEWsxxva7rxo4BBUSIpkq8THT4+ijlzflnk5
XXM7nltAoTcO9iMNg4mlj4wlwRiXS1lALUMvQRgob03Qu4IpjCkZ1/D7ti6Ks1SI
qCG3qbNnSpXtRmxbm+OSYI1g6K8ovzpxhLe9hPXtprlMTe/yPGmUiAV3/Vk0GWuw
XZtoQWpXAfjyxOEdLXguXLPywZOhVW1v6eCHmHuWjlSlF5u97lvejBveYEuSSaqO
KYBqtW169KIaPBQqQme9alEc4mkz7J/OktfQ89i4o6aVMKOefqpaGBMIMR1PRgz6
4q97iqrYCoXC9R3hZLhO1mn6UDk1EaCh4gsJYe8s7JquiEB25z9wl7OBLMnrIv8r
DvHZgKQ10/74QHstfrJ95wAuasNv1qv7Y91gBVJG+WAeDHThnP/zSUlQoGhIDmI5
IOM3jUWPd4VxKSty7Uxg9PubvX8BxeGV4QrYotGM6+7qPCf2Oz9MXioayki/lOFu
+9OGLKnRYrOspDB347D+Y87jeQo8yHMLP+LuCdQVnUzy4z/CAY4JbtxNgYrJfqQn
0kFeVSqxduIRYoBfXYPUx7f/l3gJBPxy123J9HQsKR59mGl2MPONVIDhrOD5YUTZ
opExgWWmObBXEDu0eZWHyK8IN2SAn/k6ThKW+Pe0S/TKL4A/j9LWjgJNRK+lm+M0
Rkv0/MQSKTwchjM9N7wQnNePQ1kXgkuDsa8Yb8+mMVytGcGe0aZMzRKIfFYROyIC
fkbtDj6ljPGoHlw1TSYcxWq3ECQP46NN4pYvy5tMZ692zcNYKNKJkhhyETD0uTR3
nhcbavxiBoLz7xiYzMXV5dxi/drXf8K/nUGh4ldqU3+Qx32Yx/WpLLYje5MIYxDK
Hkv3a9PKQecHc68NrzT5moaxIFO7Qdyop3lIywvJAF1iGnYiFLgahMj83WUJExVs
J0YiO8BoNH87daABNwEknyOe7GdmTmgXhwkHcul1NSn4N+Nhz8CuRnG38hwbbucV
b7jYBQVd84De5guc0w4dVTiz0WPdQgo2x0Hp5LabxxPQb/sQT3lGB1dIpx+Sl+Jo
4gPhTMUPtSNPhWaNlAmqmo4nBPcmFUe0ZiWwIRha7MVP6xZcvvsO8J0boxeyYrPo
iNl9hJAVoEUPo4s1kI2IibYOeGgqmIiS9LW2h53zcbsL3DtMSgTuA6c8eMsRNnUc
mNUi6nwlhDjBo+tepnB/oMBAjJjjmwkV1RknDsmvTvLlv8fwFIJCb+P9+whu0q8C
J7XoAKLN3WIBLQuI0s4Cj7Z15Dbtmq6LaNUKkkOhk2DJQE32w6lvV9F88XliaCFp
iUptJfFXPO1c81rWCD1XPUnrtz6GFT5ssjJwaujhCVilAnIp+r3oOq9OrpqrMDAP
u6HR/HZhJZM2S5bfaV3FlTSsH0hoUPRnItV18ffWZiNw8ml7fqMN23hFrSDL3GgR
Gnkx1+de4VCyvwaymzEsiEtuQs3L3eG9KDfE3ssaU+y1uQS/BtKR0QZSR2rkK/Gv
XWVtsFlqG8Aa3ffAp3sW9B9WXy2WgiRuUAVDRZ87n+tIJwccE1NE0KHZHSC2UMMh
K6EkB7zh6akma+gY2LCsxPmP28m22XThsqN+QRLc28HeyHUN6IemlO/HnwUud7zJ
VFVsWRBaklkOOU2Y5gpUV6MPr9Fw2I4RwXzjoUZM0kwoerAY6ZnGEUaOfhBg+XS1
G8puUm6hNigfoB01qXiGuEzBmk8Yfe6DflHWYWZRp9f1mjA2ihwsItdlW/90vKBm
6VRxoLEzmfK/bzeQN/pvQpWnswuEGWANJHlZodTPjTzqBVwaZi5Cnckq4rcSpPbp
I7XTiWDpx/wR7FupFblIlwoNdExV1Vd7CBsuXqpVXediLXKnxe6v6ocL7lrBrABu
mfCEf21YcDzCsNIDX/XtMko/y/KazLey+z8xEuScy2qDJzduacqNMH0d6QI7KuZh
YDlDxsOtIcFFyISh991bTtK4lnVZoB/DCN2muhyrg+AUi6TOm2Z265yeW14chmtX
9ohw38P5QaaoZNH5pAXvrsPIv0uGWM1BoeZD2n/3mM1DNhTPoLG/L23WKUDvawr9
dRstDKo4FIeMaNyOg3mxH4sY4vW5PNifioVn6zMO3+qdFZWXLJpO7YqsWMqwQEAz
EZabE440+eY/gko5KdL9ICIbOMlQ+NWhPraGMfwHvn2mtsTiZm/AYaeVrj+s1qpP
Yt2igJhTVX4EL1Zs1ZswFm5/KMJvZXr4W/TEWEYokviVd9hSEX7B4ZtrIoQ1Y2t7
uwGeUSQrnz9cv+56GJA0bDTmfcFfFnjenNPMxiRO70AerFKqfuJxiBM2VJ6zIFHF
FU86dDtK11FLlQhyTDEPJR0WXSKgw+u2BaZgMhRJLgvZvt+2Mu4jSg0g/E63u97A
Cquzbp2LRkSOeTIU1QsA8wPyBCsm15fdpVhj0vXa+adlg3d8A338F4vMWDmzGQWx
hEQcAdBn1CXAw2TGt9NyTomymrg65IB66zTGHDeEWCYqBkeFdgPjCEO7flwVzy8z
h4GUrOHxsdsBNI8lCNtQcbYi/Vqa3ATLGAJ7Z90RtL0ZYZUoyWO451FMSN455nha
VYEIRNNPFTh1nb9e+zxeE3LCJf9eXSBix2Wnbu0dQ+U+8jKDNcvV8nOrektY2QLJ
xnNnzEOXsLsUdiM1l4HmMwmrwFiuGwI9R6+PaBKlIxDrNJEHa08sSlSOxgUCJrw4
ZZPHWvoT8quPpgRxG7NFR/CfvwWLveVrwrIkfYZhYiV+rwV7YNmqGbn65Nis7G5H
P82IiuYgFD/81qDFXV5FF+Ghf2wTuVfO+hq29/ojbcl2nvRsbIob5whJ6+lBavuH
yyKhvdFcLcInq0VQvzgx9riaw7cSgDqlo+it9skqPL+JVzS3ShQiK0dXfqqFZdM1
PobVnKrElWpd3wzUZHAm2pOO6bayGOAKbkVJ595JIZC+jRtapKzFjMpUtlVOEuVE
U+BjTYWrXaVv3jrN5CsgUPq21UZfzb3pBontCyCQNtN/h7PDPWVXNWlxcOGFCHqn
vdhHcI8/u4EgqnXx3Z56dYZ1OD0g2qUXNs/okCCdUvXctdPwCwevGUS/73gz1Nqb
yznYRvdFm+W5jxYEwSrCQ8/haArVrWQICUqmnns3kcoi8alYiX9bEFLGvgkBgxo4
au+xc9A8Y0RlvxRdKA/NTzlApQyQA4Hc1rJEOa8/OJeW1BkF7sQ1XJg/cm7j/jen
ZjiT/CyT1W9/JVplfryfZUoFMkGgY4ouf8Uk307NsGP6QGzhx5F4o6AvC63lML+f
eRV9S+/sGM7G+8FfYcKbDz7J75nGt6kcsVMS9CI0DCfKJIUSjlge4LJdML5R+oHP
j0gKtVOmkl1+TWp7k5wA7ux7d02w/Yqrx39E/SKzcbxOK+behJKtyGJPAmEkKf7U
XxITOKFfG9TI7UD/20w3GcngdHPPd4gEhIL+Tokvrp0=
`protect END_PROTECTED
