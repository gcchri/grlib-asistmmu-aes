`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
870t+Tsc2Wzc7uHR6utJiukO41mMPZ7KBymrGV+g5AqLsQjDXFizyGtqzWYfskIp
qfyRCD96Me7wYJonHgbmM2DLsd65FVoUe1qSG1yDMnddlZRtXv5117iKHawbQYp+
M4DVOYJ7rNFdd4+BSLouMIVI26ZSxtLDKh9ECKXRj7xfX5HNvZccvHhB1OCC1GcT
FryGKPbdxQeacgJ9MuDRyLYxHpEGmFcKHndlrdV78N3C62ecLiU0K6ReRettKCNp
`protect END_PROTECTED
