`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+dQW+rI9tfaDb9ls/922b9iBhOvd6I+bQz/MmLzjx8EZfjKWAYyetVX/CvXPqvKD
xTlBm7TXhrwGZtzlS7ceg5L5AuVdeO+eiArvzXLVJUvIRC5mEVD7Ur93wPw8weeQ
Y6y/O35kXmfWpaBqL3dv4lhwh3QoMP1PrdFTMHvKNSLb+qTlveDtWRGRiw8WJGQM
cII6CaJCyXDk3/K/1xVDNi4t8SeLzT8IW3wNNhuGtp6n9Faw2WtCzwL7xLbRKCAZ
KWpSFyONbwo0Zs3vD7ZB/2DnR8xJQScScrheuAtwmb6yY6NkwGVxiS9a8DZqLJ2R
k2w85taTXD+wpfhk1Sr6LLjyZHelatGLplvtn9Y+uGUDeJhUnuwLln/IX1TvbCe0
cded4x5NNa1VB9Gx9mJ+wOOhSK905xbrvMLgAS8XBKkJahR+0vTIN2aoBwMdGfvW
LQ1V9dKDqk2uqpwtFbgDQ+xFzqdXBSu+bj1E9GKsqr0zvRjXLicj3xLn2+l/ApAW
lO2hnnxKRVgNXMn144xECzndaafYV/9VycGGDnVwryY=
`protect END_PROTECTED
