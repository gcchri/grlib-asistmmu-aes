`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OzCplAi02UclzQPCKw+DXMQRhpeTm0/WsPpaT2da3Cik86TnerDvJa3FffTCymWQ
kYe2RpaElR58BQXNd8dLaEn7S+pYfd7v9Gs7Bo27oOCByrUE7w1dDya2/RAMgy8X
vdmdYQJvlROy0D7X+vfmyzOAew4O2BCgs6h5XCqGjCosYwGNgji8IEQ+l9fjbWZk
Zb/Cg0q9npZaFniqMvyGy8ZVIpoLNR2Qg8ieo/tRF02PpIih7vQmBIBwkaRnGp24
PzYMdwHkusNSHjxcVU+UJMVfyHLvOgS1g96hldMaMY0GAj+kd6RdnWthaCAi4Kcj
ZJr/v4v1VnbUd1QM+R/BfKh9yMmf/bwYNhh+GC3aHz6G+Hw7mDZMr3zgH2JS7gZ9
XuOPYFFjpA69bLg9eG1qvHhB04TMlaECVGFr40W03iWxk7s3gpFB4vbE9TjaukUu
6fOoO/zfeWWdx6ct2i2KIgVZZohOVlNt8yEzAm9+5pUL0IFUTTwZ80Dg/fuFAFZq
qzgEmT7RqGQjYd9zYykN7+UwkSOJxXlNg3p8TeMfMHQWNnnqbQsRaTFBAeaeJgnF
awHZPMJierXrFXIErAA8bgf4qO+KsaYyS4zblXAkkxJVuSV10V0eLiuGQlpMHerC
98MtyApuJj9Up/J4zewnxA==
`protect END_PROTECTED
