`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fqM+PhjctaRvI+OGe5oWHQrq0tsI8i5KBgwzdHHE5JvyENTbeaqVS5X6mS1YhkoP
j9xBpmMBCsULqDqSURQQKsgVJPDQ91DezdPH+qgsLcu4ggib07s5CXuH2YAzcwE0
4kb7nYvJn9zHcj8F6EXBfmeAnFDSWTHIQjopDCtNLx89gDp0nBZFBhnE2/iHcaiL
fbVE0XskugAe6FYy5ZmgRp7mvYuSJd3AIJoj61XmFkCwwUmlB5SYOlyeyffsTYLj
pSkfhWRGXZC8mFFFXOfs2ZGQWNKpWTN3l1LzjNLThlMuRaXHtdohKlVMnWTs77Ia
YMtFXeeaYG92Jrvd4TAY1TeyKX6gjoJHvOFb4Uj+4j79ho3F+dOTieefVx98Bpk6
6CGgkmdEK512u6NzoKl6D/OS9m8LrxmWxwVY46imxGEJYt0E2od38JGoOZXq2rmp
lnVdTmyoXjHIx8gzoHyZjdFesWeUNWAFGsREprnTtiw=
`protect END_PROTECTED
