`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VSBcvnXtF4YVgKjFlLyG28kTTJoX4WMBRqXDg2wosTIO6524rvaEBaPlkhYQp455
rynLD82qQTxxKLC2VQ/snHwEvZPUGEnQpLJsE3VxQjBrPp+DPdba94I4HC1odY1O
P1mXTIDTfN9ZOhfmZI+zGZtWMoy/oCzf4PoVJY6H0SJefDqU+6oCFxkH6NtC35nO
5V9CwSxlmnQVxsolPMd8Xv+0QGntENI6P+Gut9d6fW/vuZZuxNCwvf/LChnljxWb
IpTPrwaCx6XVlN7OQIxBvoX9vnDup4EAxtEt9t9N9PyXqznIweEqp3yDRvVmUai9
KEFtIumpG/fDtJ7K3wseirtnfgEIG8sSgm7MrUuGYd3oB3x/eEeuLMzfcQ0ZDMXS
FOUuTqh0yR0Ha5qvAHY/TQrtPpTyAz8hDZtHyP/Wx/sf4GVi6RM8SuklyGtOQsJ1
+7bkxepMbZ49ZI6stdDJH8rDexrTUvnVY3WcQ5FIPWQ=
`protect END_PROTECTED
