`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oCDG2Fjy+91g+GlazKjdobRM5WXFYnupWhjiqgU1/y0lj4WB9UbcnphW1TNUU87U
ZUQBUyVcaInB9bDP2D5Q6ihcbRELBuf/Cr9ZsaGcGrCnIhvEZXWGMBcjgxGhregI
SIewgvEZwaNCvVgLeTOgkX9fQ1Cjx7aE3jr7xrQtLy0RilmDvvpHBUmHCfwicrCn
XlED/6od793V0SKqGdNiIYXBn7A8NgijYCDXkORWHiQZXvpNNrMT6y/BLrTgaJxj
UnB+4ltJsyKZkYueD79FOTz3OsUK2dobOfu3OpLBBzY=
`protect END_PROTECTED
