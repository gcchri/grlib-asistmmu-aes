`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J4mhoZaQmQGUZFLNyKCNwu3DdtBYmi1Kf4syVyabdm1F0nPxBdtfv85kv5Or+LrM
unAtNETBtWQZTYYBbSo3YYBm6AoGm39/14RnVSZxl4ZkCpxGILt8C1aVSqkplGH2
MtDhgSRUK6elVBKMsMUmJ6X02M+h/fqh7SLt1gMDwXSwRCY+eOn9Y2tw1DcR0eCF
Bh9s4Bs6asKYNHIKK4D58gbmwYRj0CzdJKqrHZllzzs0es71wtI+IGxqRlQ2U2YM
+kHSCAIs83BqJi0CyxvZIBmPxsyYQDZdYNzpC2ZkoaLQBV3ovZxWrj2EY2fBh+TJ
xNnlTK49aAH7gfpr3Jh5pXsd0Org1jJwOkL86xsw//lyBmMfHJ+cv836A5uzG9X9
`protect END_PROTECTED
