`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oqxUU+HZEaIfkpa4DyokmzXlIOfNdBdUc9t0Uwt/pwkAgUjeGGwWN4DDfRkadFih
J++PWFEf1ltQG014I+kdtX7QqQGpW2gBZ0e/+f/SERSF6P8FAiyEc5LlEtAaDqmk
fh0X+LCJaaSkMmcD3q7DogTooeAcxz9Y+mcNV1qFNTrU1kTNWKYGo/MoHLF/q/Rw
qdfw+XSJP9gJcQ5mMvgp+jMGZxQKFzR6SH3LYmChi7oZC1GkrJEMk+MpqUl6nmmO
Fz+hJjrhGBEDoAZq50+yPwEtR5XmjnV0oPyb5ALKPE2Z99JZ4YIZ7/pnxHL0K5jh
Hn7jo1Dq8pXeQbfHjE/tni/MFaTC3x5YrYJx+03R+zqFncIQ70D5yBpdkbImScSV
8rdHw3MryIavOB/kU4MHFStTd0HPlS7EsNA1YXc93kz4bLWJhYiJDXJJF8NNOLL4
KrFsIPqMtx8c1Ew+gXJ3K9B9SpHFaa7PoomqJtK8aLyjInu9ajj0+dUgM8QluK25
gJZ1/FadOu31TvgheOQHxkiNkp4l3S51+jbngPiMrUTNwT1bVSKOCHKomc2UmfE4
SriWrXUk+Fahg1h7BpKBdbvmxqZ18AwZ29Nu3fgBEX2/JXCIzlHVnLV8KYyRylDl
FOpMlO9lA+u2hg+cGTsqoAUwJe6ABVlUJfhwNWSP72USvm3fwaYWBtFbVlJTNSXZ
45ygzw+bjPJLwK5js5ZMqt///pMfiGy85Bc4NcaGvnCkbP2QQDRNn2SAZZ4yqZDD
PC6PkgCf+MmY9se/nf7cARO55WwmicKHnkdT1dP85xHUnpCwMe7cKdVc+WFYLySA
srNMDpfgTRIt13VEhrbuYbCWkYw1oadeJbAWLHD6bgJlj968v95A6x+wyQbfCJkH
K88m5LuxQDHqku97I9boMXggpgQzlF8nAYL+2S48mw4DW4xXGs7t2sLVLJKJ6w7O
VYeFeousS+2ABD4iQcktInAnmwuOTNkZjLnzRoYVUt0oZov+N2kChTYj6nG8au/C
6qOOn3KQulmndB4FP7hvUt/dLkfiOfCl3DwgloRCc8QAGGzaDw3DwNiuAl4kBnsr
/+wUdiHdca9FAy8VmYy/5y1ctbSKU9QU5phojFrN7WiioNHKk+dVXbNLqepCQ+FM
46hGHT/kJRdX5a9JRYBD2lAxdVlVBJ3ujl6SwMCZbXwV6e/si53cn7pA+LXnP8WO
xp3SDc2pZMOsN2k8WegMhmIJrHWVjCzodzrJB7z1QB3rt+nHcJ0wcQUuvkZX5xrb
O41+eNvKIIArF1+xTvN9vt+k3jQLW38CAKc6xwlVGTfQP7T1lK/KGEiqt8TV9qY7
cQ41Ozdw1028fG8sTS2S0DqBV0tPyXAimbG62RFSoPanXCTgxgvDHMSAp0si/iS1
ElToi27Bn53tHoqFFLQ9kPRc185y5cFt63a5DfSL78ORkt+20cGnbmQHpFI7iXEh
8yjPPtB8vpxny2Mf3FfwEDury6u+KrXJNAakT7wMELQUFquspRQ2/+WZ7/wlFpug
XGc0iYI9mgUfNuMkvxT5QjtvmEAIC81c+Wg37mmZuhB8/6iFm2c/IorDvJLWJ9Xs
LCz9IQO//dxNLqFszxf5jJWA9G6nk3BQwIhrGiWaPq8pTEPWHi8K57m7dgVQeLvU
ImroOQDtIBCu9ybvX698zapZFgg4rsI6d/loxBlOkYAHKhK4JS4aGWrB+dbx0qLJ
A6uXkKqYxGeNK/3q+bPKIKskM7XynYqYMQfD4JrBRmdpBql6ElpDYd04VI/m7F23
pWS+zoYQH5gaLgT6jGbTcA3cNjh5z0a0f0F9CTdmTsBaT5jyEnHzFbMAPhLPypUV
jeA6MHa3YPEwAuhiVas+c/1Bpl3ozxNed5+FZY/rL+ypATqrNxLZtAYLroJKa6ff
KTFu3GNI5rQvBTgeZ8rnfO0q33sPdSIVUOQNdhFRPrb6GVVl6DxYL5eKM5s9mZaC
NbACJai2akst1udZ4siX7MXTPI5ThBbiiw9EDU2Cb7AnxzgHmzip6hRuDakUz7NV
NLlo2EKCNhZCxoA9hLoQfkjb4+sGZpJvM/kFgqDOdBHipZ139acggJjbamKgZGMN
aoGxSJI4uqT0GWX0Z5J+SrizLe0D1f9T3ejT4u4yWR9bCt4uXkRXoW2KypXH09SX
LZK1lZfE0fPcxuZijEohe/WlKDwBbScwadQc/VYzDYB7XA9+U5WcER8scXnn79LP
BwDbq6udQf0PqOigGhH+ZgOvQuJ2zAFGH1bBm05B3wDgVFAxWK3Rr0w2yBmjL7ms
QjVxiSqlRVkyQGLanSEwH5pig2iSIhce57DocY21NjjMNUHzjS5nZ/dnqFh+RcEa
VT2DfxAlq4JtkUkHCPUi3Q3CCDWQdCdgVpRkIJjVQhO7FNZiwGt7XyLoUxkf59MF
kYxzT0KsaJgQh0YIMGnDhgS0Aol5a5aI+eOFojpmA6NUcdkEbpf85NLlxN0u8ObO
3uUH9wrmQX5As4KGIt1JaxkygJR99qCp+oKK60d5mmGp1pdt1g2TyMEzZXMtTiip
nUkma9/J8GS7U0x9tsHFwj6bgmWlmthwNHKY/OADWVi9NhNDCnk/zv6WWe5L0u+M
Loicc/ttHnGyosTlSmOzsr+k136FlLSifWN0eLixXronng/lWx5qSkdnAve/OrGH
WBWdeTMKwfHTwgc23D2HG/VSNJxFjl2wtBJXMnu5wlc+/S3rkvV0QgxvqHrUy/Nv
5DjAq85EMsFvmZOMlCmVZaEzacCLeQDx3CHiIyjPz1Eq3b+VUYccynPSuMlU2iL+
jcXWItI/ZxCGfvDKyzwJZ/sriGtLFDO8wRaeuLMPa+7Eme8fb/GKGRI4JizPmlGJ
o2NDzjuYI2SOHh5A16EkNwXBW6EtnyVr8Twp15s8k9npSrypEQxjAkeEbQERF+jh
kI+OMFvtIRWaGJBXrFbe/gAvzBggU84x7dBdUx5K6hU=
`protect END_PROTECTED
