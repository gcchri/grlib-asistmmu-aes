`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xC3vXCQJ6GwidNStxahz7AEja4YxivYoFLGx885KsDzxB+A2HU0fFIISvEytC4fw
H9mAN1dIMI937wXRvcvXWi8iO8nVACn7C2bSCe4V5tqT1fyu4OW5dhPiIpJpAnQR
V4K5jll2tH5NEZwEgxiHeiGCgJiancb1imL3yk+g/ddntlYeOjrAJj/WZA77cZ/g
/KdT0xOvQfeeWc+4jNQxwhiK3Q0Id9OJ7m3h+IdWzrjwGMYv3HDgWXlpuVTG219j
VjDA1VZJu4Zb2asykSgX7TAQ7H6VaTSrf3Hh8YQ1ngncZ8LllkKyXSCGrneMoKTe
W5sgkQFtrM4PVBmcqdze2MDPaiITjCdZKG+cG/iDACH2w4lbVwoL1Vtju8G+YGbw
HTMmx5seNCNeYwO+Pq48CJqkdRL2D1tquuwPJ1eVh50=
`protect END_PROTECTED
