`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nteuu8pwUU/qGZ2tT1YmvOSA6277jCG9gNvZOHJjtoH+TpMLiim+s6NtP5kei9En
cEAqAR7aQkPr9LTE5gq8dDHjcJYlj0tizmwOtHOwaU/1QaDnSvUbFL/41g+5ssEi
tS4kILlpcl25tyoqdd/T0fspIuV2jEL/Fsh75AuPFPNItUiB2Mjx19f8Bqc554Gk
VpCaPojFzwrYs/N92ronTGyys0m4XyvBAsNHEErfOYJ6xQn7rkHry+lNXDAyEf1s
J0g85xmJfQ+NtHSv1Hr1xU7Vj1ePNZ8/5jCgtdaHKmAJm0q3SmK0EIwdvsD5gA64
QNuMvXHpxUPkHB9Kr6c3/jtigGi9XkXy4Vo3fTPC+9Jgg7QOWlK5Zrjk8oQo1wUu
awXoqU01876dcvX+T6W1vlt0k2yzBllBI52DUeoXQ+VTTcEqyFXZ+jDBQjQZICtO
uJeDhI1dkzTZhsIimC6RL5en5ri1KG13Zk2KPhHVxFRtV6vJwmC+E9ywnDjiGw2c
eLKmOOlMYTb1FbY40Qv9e89AgkjncMqOtwXQdJZRiuJjnUlW2xaLvmWnB19ebKc0
/gKK0z7yBzSnI5smHQs/+Nxzd6chAZ5U2EcCW/Iwd/cqx95wfJAFOSSfG9ZTOWKQ
yNCc1D8wpGp1/aF8UtP3hfq+8FEUYADh+tCYigV8mNFthSvWE39Ghrfp3krXQwRf
N/un2YGZZfLsQ5/SkkihQ3NfkO2hcHBNYgtIQ3bTJoQ=
`protect END_PROTECTED
