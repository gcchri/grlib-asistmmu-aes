`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+GYMxtAUBxfj0iuaulqprHZCUKFiED3dlc0zmHcXPMk8yfUX0MBhB4pJy7pxblPN
bOaiN/RkT28nZhzz229IO4VWFcLrjpoOvjjrh66VbZxHN6+lKcKHUSDnnF0K72VF
/TWdsvffDmF+h/0ygQYLP1Hehd/wVj/E2nnJbuKEZ/3kZ8GC8MV97q4h9xDuhEvc
GTbcrhsbYumMsOxk3SdACcB6BNWgsWGvTT6ms/xnTJORu4x0K54o1AZ8btmkkTmf
WnfZUE8Qua8sBLM9kwAP3ZC3CvLZM7Z4ntOdkMazTNIQOTU8+yN+5UexkgGhuYL5
tJ1BiuhCYBPN9x+P9Fiqkcr/hS0Ecn3NR4GldtGg0aqR+n+G7ENjbecLpz7wek+K
zQpdvmFlvywn9C+u3mg8gwdFsXbARYsfQ9Cqs1dSziN8cLehcoA9xqRllJ1aj9mL
8RcVWWSjhtm05IaMyFgf30/IdQTeHNWujZ0h604LMPuW7fguTC6try7JtvYW4Vpa
ArBReHfR/WlBSEIpeWnebwJ3LRD8IWUWNZuDE7JnfFobfy6EQ7Eg9TmXxNxc8BwR
3Amu1EMn3x6oTS2u0d63ONBRy7FuAeRKjZ0Po/sGZ7KbwOoGRjA+NO3OLimdUjTj
2muWyPi4SNEfT2gvb4b8OdaJ7isRHpUKORgZW9ZtX5yLuTi1U0yAinm2rIDYrhGM
qvK7IdeTjgdeL35Z+i0sUrGcEP2EyN15TcdRCU0XdLMJGtTgUOhfgdzExFN5LMeG
+eNZsPJxFqvjr5uPU2xbrrjcYdE6AGvuqMr33j6lDmdOiUjTc6qllDFGP4f4/nUl
jcyKw9hC9nCNRe/kN1HNQqx6WWxESkt0SRm8MPE6mZ4sw/FPBM61MQMQYrV1CsH1
MIKRPdnWFnp22NUvnmzxXDjWdFdqkNS35UDHj/CqfZoVDpR8qB4cpQIpYc9qEX4C
HCOZgU0ChF8CQ4Mdzd7LHwCbJeo/krPdks3aQ3rcMUskSgHtzAwzphbd0bolHwh/
8sI40fQVup2rYKKzjJQ/CJ/gCYobnxOC7VA5ENW1aMj7//7e+YiE1CP2Zncy85iO
n0FcpwQW/zuWWFvEb1JKWNPKdBI/yIEgleYhVuPhLBO5oSBfUZFJD3v8RgfpXfHE
p1C8r8h6ABpnRG/cpSguureBX3oJDxHmd/HuXGtSRPzNezbL941EIsf2Ec1rHILm
XxCPzmub2V3JqHeML859Dy7asoU3O8pkfcisCtDuzPZwRyr4Zsno6uQacgJZ7b2H
+x1QxI4ntTS2/9Gv74baOVaJm57bEkiVj1wLzj5Z6/wB6+2n8acmfR2r/J0ONivX
0N8iir4mKGAoNy+77kwMNe6ix7GdwZkIA0CHUwUjF5/mk7pLi75kAtE6nwd19Xng
6S+ZSwj9QBw7ZbVvk3uDrA==
`protect END_PROTECTED
