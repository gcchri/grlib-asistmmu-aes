`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ah/2WtczjMyFB3Mim0ubru+irWBsL8BHEl2IbP7Jzvuw+IZHzTgKVQAjN4S60O2R
9gppcBZzJ5+AfrubgY8BymH6UvfbXTDN1u07i2iDqW3ylK1ifiZPXB+nSg6MtTPd
CaY98XH4plly+2/4rTYzWkqJhD4Y+o9Jg1lVTpInNjE46gM/iFKQNk/poWfUCsp7
RTZsmZfrSAgRBEuCnIeClQR6BrNrd/p5kwmg/XbzV38FezkF9qDlzauAudwe/lfe
mm/ZcT9WyfOo309Jf5e8RA9mfXBEsg9XuIa56WgT5HoN6gZPjSmzPpu0Mp+F86yw
YKTMb+hPFQcQ1uQ4ojXCdufcfVNbuRKuH1gKOALFh2g=
`protect END_PROTECTED
