`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ujmv6PGIRJh7AS5wp9Wdj2d2KWLbc8cc9IV7nRofP1Kb9wS8Pf/X1f9z1mcDvcqB
fjsP1g2vpVzDEz5gR6+NOlm7KS7olAqByl/lCt+F2nopdIE0wsirASXuBThKAbRY
a0qSiWaxQAC1Gwqoi+mBiwylbtpk/5oRXEk95WnKwTGXyTdO2x9w7kwFq0nZKM7v
NMk4Guy8+3weKjBT4dJeof77c3qU7jYYlHdHMUw0H7694uIODUDPbycbLSbPQaMn
Gxm2vaFxp78YQ9VgJrPgafttrZowA6SEypZjv9oB0GniulDvYBKodA+IYDs3nQRV
xVZkR4ihF9PmtRLbYiz1o6imb90IzSOBZEv4WnLS6+2Cc4zncnguvls9HYJxmNzU
Rv6BmTqUefmZkjMfwVfnqAgxwVCTtIEgmkmuFk2rYjUfVT+RFZj5A1+ioM7j5HbA
ZKZgFKokU/1DUiI0mTnDVA==
`protect END_PROTECTED
