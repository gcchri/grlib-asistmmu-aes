`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kdtYTZ+ifwLGGycGJoDVSRFknCzID249zjIr0s6ociIf17JPJ1fpE31HBBOFC2F9
Z5qdRxulFC9kQn8+rmmneLVgHaykl1p9noGnWMs/KROsP4UgCfjerY4QfpFTxZkg
7+VUEYKynl6ueOAM7vy0iSzIGUWIps6T6G6wlt5s+F9xlFx5a7zSSfNBwoeYfni6
/FExewz29ezSbZ8uw6rZUqqJAHQ3LzGytd8UcPTZpOlkgstM7uY03ikBS0O4498o
DCom2uZhN8IFrTn57KLq7Uo6yzGC6lKwj+I6fwJ7YbpeLuoviAn1pn7tgPIpLzOy
pgqWP2G/elf9FhXQSWA7gI0MkVbPbidtP7dUEuDw1NfOpZcWy+/9bk9FhikXHfgo
XLvgqRb/1wkuzyk4Mmn1rNJcI5FwZcaJn9khWEEgrXsBucJ3V+CVM9BRpJMTzujE
Y8w9idD75zYY+hRDT3fxbORQlQnJsZgjYcl+2pVlJubzdQyiy5MkeJY4Y8PXw6D+
brEAU9DNVLaPHjYnqsmOJA==
`protect END_PROTECTED
