`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AqHzYG4VxK50hdokm1xa1ptT7IHUw8N+1WcvA1AtKvdq0nEeqFiQ4BUWM/5GVezX
7YpBjVnsFuKn2mC/7mRxPrmocn3yBc+sHqnCNjcncvOVltK9s1NEzohI2mV8EXzn
NEvNd8xAIaN3ylusLrisZ92x78CvudxZ5gCvyD1Z5cnVSMeGZsWrhE3b/uMlBalW
Z2teUsSAYbNBhQ6sPOWmoKjBUpppQRtXBwiSsvyUs9EX1DzxrUimn8FiDzfLdn/c
82STlpPX3vNjN40dN/dw0g+IwB/GtBT+wxQlIOoDt4dZmyPm/6w9kcsF/27ayxT/
jhIkzPaZF/u3Z9DbHRGQthpFPQo2DJ9DsRqmMxN0Pj7ZOmNoDor5/pJ3p5rXsVIH
/1uAaDl98CuAUJS2SQmnQNl7zmRI2AexUI708RvxojpMC710hAqVt8FJT5+Ppe57
8OQ+Hr8hd+SGnyZjDoCkQVBkmCwQFphqHhsXxABswMGexpZROMRkScdoJCEznm2O
07E/hqzfW9qr8mdpgJ/Xph2+MFGXLBAUnnhpsO5Qxg8QUt01AUEBs697pcMUdvYr
baOQj0sXm86//FO/ACh3AA2+AdpP82ku+XHHMtYxCWQ+cwZdAiCeX7DFOYo2VZjy
vhkBk7meuBksjBWF1NPGRXdwXMT5qAk0O7Y2xXHLNqg=
`protect END_PROTECTED
