`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N78QK5j8zEL4mv6CUKjObBHqS6o2yK6fSP314FQ3p9/F/5hksOgBHnsGxxuiUqa0
WMY4aswCOhU+WfSFKMXGA6hKV4dE91cwhIbFGDcAsEEcXBwFJV242Otah+jCsqZc
LaoJJp8E2yaNtAKdLM4YEC/gIYlZ30++bNMEGQk0VrC+hRIW4wRM4A5OnxuqvY8B
xzvNmJhBEZz27/NlB/UAtLB8mMjmQx+FZ79k5LXUQ6nEW5ofZ+ylsme6qjm7CzqE
kJ1qFK3oku6LE6EV1YMSO867iR3fAg+xvNSaJEvrlgBWRp/Z+R0L78jXZBgR15bM
68clmo+mndjT/lLbKrOpdp/L7pnOKNtbqIzgwTxuRO4DBSGA57QZO472RFv4Cwj4
fK9ZNWPRKxoQX0zDX4/uUHrhIH2vU5DtgE/uXno5M2AY/kVdaizy5F6+50aT3LCS
vPINsXbZIXXtFBJvonQ8mHhd1b7b+OxR0zxr7XY7P6dO+88Afflbku2lH8NqYnQq
qe2wJA1fVlx2YmhewotPZpyNc1ex6KkdUJiBAXX8oT58R6nEoDNgLlEx5+JpfSfo
f+09br34epa0BJU17G76lw==
`protect END_PROTECTED
