`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QBYGlPniXawyjaLvt7FMkhWCn8UTx4FPpIhTnjnouTD5VvpuEo0HjFsCa/bNOsp1
o/3EY6ePvTH4PGcCV5HTY6BF9EVyBZzKIRH+WXDiS+1090HyNxfIKHvW2omXdu0T
o7gIPwYhZkvxlI9a6HUEdPN0Y3+3MLO4hZbr9eHbWkgbSxHiF2K7seAY+e4t3bhG
3bUiHolEPg5h90+A4jdq0nipX8DF3+bm2dIRGFsyK/0CUP+WavSWgJfU9pVDpAF9
pmY3XipZyzLuVOUBQ7l9NL1klyzF0aWQ2rC+QrOaHKa9N1jZmO6/P8ex7kFk5F9Z
39vOvpmneAIborJRmOHg03VL1yRNKIWQ59+JZimMPfcJsZ23ffS1/gFPvsNtuf/A
fQlKfLYgvuCUvtuOqfF4Tkuqg8q/mbdXUJ8KZPNpPo90reuWSbp9ECzsg7b0W4Wr
Epz53t2iIlNUoIRBvKOow+6UiUftY2Pxkj8KTBnRAX76URFiy2IxC80Cg6bOjqSN
Ds0wuCTDqo5GyfTrqi3FVr2/lZfQjTuQ7AgW5l+nViGEHI7QXSTKrPsgxl7owH+0
gk9Rzat+KmX6JYzR8jHgDhVAKuAFfsdQBlx5D4CI0xv5KibGF1pSb7ESkjnzTLMD
DYR3lcAd5amHCgSZdD5Fq1M49yM2ukA9TTXIQBWGGCYHQTeoaq+V/1bZZQf0uru8
o2MH0CNcA4r2R7BbiKR4yTBi4YIoA67zcvQt/5hzUZ+MK9IUrRBmJu9ijGwETVVl
nnnwL56QbA1N14UFTItXBKFEO4alEQTiOQtdyDT7UEcI0rLj/WJyyzal6yOB8YKw
QaX16Fswcvm/5pAcePfNRN5taNAtoC1Z0kfk8Cz6IqpZtiHON9XdjFcOuf/hPiGb
9SwAKMidwHYshLveWqKVfuZiWHTstteAOG2PL+aLoEJMw2R8omSwuDOZNq8AYQ8X
kRap/4MRIPFfpzlVvxV2wO8J1i8/M3RjTtldh58vX31Z/WrRRfcK4dwh4nddtcO5
t8RpBSKivfISK9aSHjP/Ff8PNChyNlrevDFpVyIJLVBye+gb7/qlTPX01yS/yONH
4/qF3isQx1Te5zglvtFUtOvULXFMhky2H0H3psVsEucgWV0nroe8hGl3KuY8Ih/Q
nuawjp5YKjQRhWWbekMdsuIrFkwqNF0/o6w6V4taWDc6r9C/KxCTKnpwCWhke+dZ
8+qyFN0zeTfj5Qymvus+yEnfebzpOvU6UtK+JcwDKBe44zOtiDdy1OMkmTqR5HRv
Ly7YL5E/Xh/sjNX9mMzZBhEI78rDilgZRQy1hBrtzYxbne3W1WpxdDVL80MIcyNm
NkBFQA1abXOuG7ooFGmIemMRqqYz1ZiE+zCNLA/vr/PNBGk5cotMp2ujd3uGN1GC
PP7J8o8QT84X8Bqvfckxl2skb5zcLMzmNzuBnc/FoSImH55EsnlL0NcjyBInNA4W
EKQvrhhn7jMrKufdi9fWpCtsxfvPG+AfKRLdg/I14412PEjogcMdg+9m58tru7w4
6sjIX8SMU5jNfiUPzlQ6+/1pZSbdRA3uOfZ0Vti0J7DmsYo2+XtUggo6wwLYydZa
JGJrG7WnsvvwmwGopWT7KEpNjsxFr/ivx+JxgCqA+uTDeu4laYQyg3uBdgpfahtx
25m73HdPqgMgwEM4uo9O+tokCaMtofpBFHoPo49KBKIoLQs/OG8EOXIW+XWJSilr
zkiFoI/KPTyyUP5nyb0ralWsHFOp4QYpRXHgAfSxxuP9U275TUM8Q6v8K1yMzxV3
gQExLImRb8NnxB7xv47XFkuUAGQ8x2mc3NeitAxziaV7EVWWth+Z6daeVh989Ne5
BVNfvEbV7UMwvN+HYiLqqsdDkWYqT1WPHcZbeOZ7ON6LT0/IltWxNKPZllNpvuzK
aw4JL1cMg5fq/BW5fi5y01CQGNNzB07sDEIQkP9PeSW8ODtraj/VdSt4HT9N15UO
pnEVtzryn9hkgtlbjOzBo7umMfMkaZswEUWTVvXkPuhOWU7x0ioDY3Y+t//xj0GD
z3ZH720BfylgxDASmu6LEx4vPzLGSJ3rOc8M1NQ+Bjynoc7GPRghnt8XHxnTv8Es
5eYQRQgjOG3Zy530Ym4/J6aWCk+KhUOix1jc4m4PA0AsjllDKhZBLFA1FvMwAO7U
jaEFmDrmT8OIiN9zolv20/xSZ4T20zMC6VEipkVFW6uq2MqWEaJdPkZXOwLtB3Xs
K2SGngVUVIbzDXGn93HWXNklVzWMW8nK/kWGfzKPK+dOG0l+HVqWCZZwQWhsP/2U
jiNvx5VGycuHx357pUiHkE3o3C7O+q6Rn+9nV/6cXv0GDTie+VHQ6SKJC73LSGA/
AryIKLnE85aaCCi6smNRHSOa5tOJP5ZE9jyXr1RIS66AQqOCBu6UI7WPJOXr2Jqa
aiAzEINUemWQxZ5xTWT1SQqp+ViYKR3hWjkSly9PtlPCxyttm9ogqy57ZDFTczZc
pH1VVpTdglm3IxxbSmtLtZ1x0eqbMpHmrR8zRnlbO3WdLfZWGmRLdPaD30/fH4Fc
uwuu/9X+Gr9UhIM0pZKEVaNMKnU26a2yP9JPKprhz7fjfaKjS2emQ2d4pXfjt6ws
w9sQXb6RjLGWZofXEPdt8Vl+v2Dv4aZlVzugM+47d/WVAO9Wl5yJjRp7ftZnsWAm
2Mj0bRgjEONzsZayvAW3nRWPNer7dJE0CDlYilaTliEFL3CtenQTbmNTjqttZzIV
12pTePQvtImIBM05ty73uuqgmik/o8x2D4Jyd1kZF+VRRmzFINDdVPqaErXLL42Y
GaunbfyMdf9xy5lgB7jCNwDpWWcdKJ5XfV4S9EmjHlZz60WKIbz0nDcdFa/Y21bc
K8JhrLG49Q0VUVMwSeVZMlyDskPOaT/3Xe2qdCL12D5/mu4YkqSe8quLbyqnYKCe
M14OSqa/xpC8CUWsADW8ML/XWscldr0CxLr5rDwIJK/uNn/SkdmlN0cqRULgxpAh
hGRGsmsYb/ifjcxbHh21GvgG+zPaJOSti/9K4Mbhd6GR77i+to9htfnKtlaJW59n
f3Sl1o61FG2oL/aa/pTZ5MKfiEcLPVawp6FF8Llq93tvAkGRaj5fPAJ84VSrFfDh
AbXx02nJe8YEwh0Tn03m2vrL3lb/txo+2WL16eh6tyXf690SnVYnBIWArOOJzxVK
jfwm2tcVtFAV5blhY8/JYd3NelKit/LVd9ANg/ZunhYfIh5wrRW8pN15BResmKD4
6La/NRxxqcF9LDcIJjpLRO3IvIUJACzxWDP1B07GRkbwKX4bfC6KVsnUEsDhL/2P
OW80w3zeVSlUeJIRH/2SCO35KFL4/3lmzmWlubSJjWL06LSQqUD74D7d2So1aZp2
B12+78YWwC8/BYdjZFhzSMDOzYkqObC52qBboONanwQH/CuxeNeTTScjLba9Giup
0Bbkd/IpXDFox6CEAFRs6cnTWuOYUditNg037OQRokXxBIL9YaNvZPbNlWe/Lo8+
yzMipNwXX2Yen6g24dFV3ryy4RY9AWmVJ3RzxDY+U7dE/UkJ08k2lEFT/Ug7d5C2
TBy0/j+6bDou5iWU+XPjmWscHTeknK20+vb4zB9phGOz0l406NVwg4z1Hu9ZG++g
ECj7lyeKa63IESHc+vMMu3gq5xz3f7DTHeugw5MMgLhUnRBnQgRZwUJ2vXmBnGPa
hJ6xVGIR9QpgI/rjBPoiG6AzAILomW/7FGaW69l18a+aWZ6otGZ2QbPkEfPfO/ev
asa02Vbc3m/BEYAzqpgFHHyD17Nn9LwTn5WpAaVLht5xZf3afmfE7KyD+e3UM5JC
TTOr4MkPTJ1ij1WyJtoErpd5xkCcr53wenzcrfLOYInNt4WZUpZatpUqEFdwNwf7
bzHWZtwvy/XJINAol2c8qap0SAgrbsWDiPg4dlKbZlNSp73af42cwVdfzsnb2vDG
No/2k0tP955zi5BiD/UlEohfGOz3eEApt5u47v0MIMxfPP6YYYIVBB6PgfAcsNr9
5o2f7460aZFvtIiDpX7lYn4oQqiXqUCcxncXOE2JbkKjjKhWJ61Sv8cyBy7Mvvhu
koO52wSwQdK9FYr1KLhGbE8IdNacZ+lY1FnIMjcS9S/t6iuDYJWmR19Cx7zN6bZa
hV/jcQ/K6ejtTb6k4H+sd1Wx1g0gBWHXxUiShFe6f4dr8/gkCS4IDG5E/s5oGMUj
WTyyw/hNZLZ4h1ZNDR75h937+9mOiYFQfUtqAV0JPIqE3H2hErb9RK14+WGLvv+y
PNSz4H4J+xk8YriroPkH8J9rIWHxx2iDrfDHJP7fSCh9n+bsMs3vIuad/2KMtRou
Y1NwsZo70H579PlehzMneTvbvM4uWuViqsfHhfs8nCY=
`protect END_PROTECTED
