`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fldxx65MPmxv8vL/RKIoAF7oW+1BnvVletP63WAiio1JL5NeUrSkfUVCvCUzrZb/
MoYXgHvoPOmRqCAITP/Sr8oTP5CXVUIIvHSwVD4HFjYBobeKcxqqoxWWZjpM945W
zG1neWxHtEBUJhUAPmnlh9sB6fBCTwK5Zp43iLiteV7GzoQySlB7SckhH0Q0mMxL
iNQsk3rUavTE6nF8tVfg20cvhmU6M448depzPHP0jAh+3nHrG05ql/jdSOevMQps
gSmUIzjg9GljhBsJ5Q+fY0Xn/Uc6HhfBgk1WpLROy9yQLWm3S/VkdDebGNuufTqc
8a52t3hncig16QOXQeXjFhCkb66Y8Z48Xpg5bFhtsixBR/1c3snrIYlvy5kDBhjf
HXRumCUHy3Sf7W6/FUfuCggiRn9Jmgeu0Rj4ILZKVW2MEFqZI8CjnwQP8ClGaO26
zzIZ5A48ae9XIvq+D8MOwwAyzw3wPmpPkmEAXkGbtnzfX2CexVh9y4ZD00/4YuCa
CnI6rWF8Tv6oEHpXIXXEFaSvXaG2PxVcD2IRejoF1u7e2ohqEUOUV6h/lvQZ2l9R
DjP8C59skQV7YKPlWHBGYtR2OH0V3ZxPFSthvXVc7Zv+Oc/kclfIntaZuiff8Pah
ucBpjP3dx/FmF+hYdt3h0i87oYcFjTLNaSY7tO8ZJPzb4HjgPnTcOy3Ogp3SOI4y
tP8ptQpIwnxhipS6iPIVx8Ar+pWfoh+6dQWuirxkd6MwpOipM98FNlzXNS4aVAHI
AK4cexmofbri7fLbCnwsQ1Pco68UotPVXtEDYWKfjknr69Yksaj93aKG+qmhvQIs
dyhEhQBw7+HLqDvFUtLh8hxE8ujtcxJzvQ5v3I/+RlbHD4/ciheKmbcs+eTFMYC4
PepzG6ujBSPJp0pVDIKvtqxFjjLle+WSQcf79pfVYGHIF/WxXgBMsA+Xjqj57p6x
HvX3VTsSaivirLNm2c7/MUbjz3bHVTNoxMVuiFKTgP+m4NKtH471eXsWcScYn2IU
zf0gzV7sKf9mHSaL/NWp3IYwD43ZKP4CJ+M2CrFDtdkrs3W4SmDMhmf5zzQ8gnOJ
bo8FpJAket1QVKoy1TSWGob5b1VKs5rKkWBf5JbNzpDD6JLzytQIm64dmYMPyuqz
0f3SuLrci7emO/AByBXbd9odQFVB4xq9jfO22YXDu+rR8qXHwvOxGS8z22TBG71q
eXUOsNO//OQrwg9HxItbog5MBpVrKFDOD/4WDuJS+DJ3IA/zvw642WWjGTws+jVJ
MzkMyHpQf2TwuaH763EY1E8nFTqeFYHW0nVHidDyFKCr3UJ13pOzZZvrDGCpPHrV
hEutcWGF4j7jLEn43d7+k71W/toPF9nAIeAKv8ICXBwJL5jS/c/Pe5/P2hYOBHgz
gI1+DKHCpoBBgiWuqATJ+gOIMcHVmZKV42132TkAxj6v4a9ViDb3AAxqQeahLnbZ
5kBO0A33OnZ18lCI9RSd7Vxi0RYYGhr2pJbBL0zMqZgglozs8UhZU5AGGld2cJMJ
tEQQ/2RtN1ihXLMhwE/gUX+hX9DOsuQgmg4Q1gUfCaSIeF/chNz6Mu5DAIWhb0ln
+90eQoYtuqlp274RXm70Ex97zTPW97E5KeqVE2pI+hPi0vhy+U/oUPrWzXSY8NHk
po8C2ka10objUK3ewVyAo892fKJXfPtvXGmjI1l1a5UVIMR5lR7Gb7C8mSkE9ueY
QcTfgb05EVi7UMFSr6wT6QyGKphgM0g7obTSANR5DI847MO/fNlNhM2i5JP7zkCe
+FrpJg46t3YewiORQWCeQjHGztAGPMTbUWdzl85h6MnXX0E5BdpfbWaBnn7WBsFi
k9Yufj40wQ6ORg098eNTg/Msh21kKkM1zsICqz+BSFpBLtdygp0mUZn5Y7ekp0gK
Rj7fzqqPnuxIMlpE+VSGKt5FL+yCLfkD6E4Aky787FYULwihR8LrSDpYFfNbzixa
nn1MlMQSXHDbkaP8OxKInGYJHNShtggUqHxZaN9SFRe9ko9J9iOv4SZvJM13XtP6
sUHAPBwaX+oTAEQwwbZafQtNK4EchG62lrBMpLj+7TpHHXR4EBsY7fpuTGe386Uk
lkLyWdfIWn43p+5SgY5bPNq6GzxJxmCIgOZbM46pbLA7rpUUtCPfz+R8CDcxSKoL
kykgWx8/VRtMjlSmvBUeJFV5pHYqNBlVhHhufuQ1TacMy6jvWPHQa+ambOB5iN0b
uuUBCoFvAYZmOsAVgdEfwV9DGwQRgX/sDbVhUJBeIWdmlnyKR1JrF7Tkk/qeNRkq
h4dcVerNr8y5ufMMw9eeUoiNLhDIWfvFuW9HO33X/F6y8buB0OijC6/NkilqNuR6
fQA4gFyYGjStPQz+L8+LIROGjnWvrIySpwyp62zsqaS5UVEdEOowpy0VbOfQwsnA
r8eversEoWVmnLBIqx7XjpLkAI8+49jUZTXJHRP4GyFmMA82GAZcLX00cCnIf4M7
YiJoG2DGfCpOSWQCOnFIYC/74V8t09q6WrFvXJCq5SHIMJgzpjkBJ4Vk2yLeqJnH
nMUV0SMO9h87lSYz0QR1NdWtNmcJqaoxldw8VaBRTcGUqp8wlnhWQeHHR5O9834A
BbKpJWgPbxgBMFBNtspknYzA06bpc5Q4DN+qnrLovHqLjmDUf4NtZOkOAkQdE2eX
kZH2fEtl7G2wODpcznx4tDbqj2xmpM0ALwA68HDq8NjbSRFKv1NIoLhOpsl5yt3l
OJnQWwxpJI2Wt4tBY8y3F7SHPeVPlGUZ+67wawxXG9Xlf5/EsBZA/vlY7vyvYAIA
x/wQZMZgUNTr8/8Z4DqbPhnayWJrCUPyCJPIZ5Af7d9YycfCI5mCnsLzSozWs2sA
IQuPh96TLhdqK2lfpId62W29OFQJag1/lu1VAm0ZL53KbPU2VNdm5nFlq8CvAJGI
e8Miry57Dl/NOw3omxXDQMQ+8mQw2RrfWHB0xwmbCIsQeicGCIBpuFjqEDN6hrE/
rNFtQlpRQDd3h2ApThVyyJRNLZTUmjpItCT3sd3JVyvYC2+s/iO8T3LQdYnF2zWQ
MUUSqmL6L6ttbgWL96bOSESKpX7lGaB8SE5o9eU4BG080jrQsedKwzgI5RXH8PL7
veTyn8IrS6+YtnKyjY6mYLmDWLhCXkaIq1ar13FpCO2mfBpksYRpKxbRCdlfguas
UL21ctbSjZsBQO5hNw7mREibopO8e5ct++Ez3GD7zJ/G7QYRQmyWryMjTfCMxySE
TDPmu86xVnAOeZ8iJ9rAhr8mXigyJU7beElrIb2tTp0jCfo9vRBwMO5Zfcbdse9l
56iaE5paXBpvaGGie0bBjX+WoOYsWFJC+fhT3jVWZg5r4LRJegETaPslM5oQ3rJ6
wyHsSPL6EC/g+DCLO/KpZnJBF1hu5lrQjUbBT4CQu8O2sH6UQ96tVnnCu1gpvew5
7uKH2qzK06kico8gYhZ46MFWSe9Jb56ZZzXrCOcocJOR8mVSeuDIzz4S7DygJCuF
cVtraj1vZxeSA24Hr8QMXOIs/KVL6ea/84NOpnhdOyCCAQJQfO72mCF0PlqwVTcj
6j0KwFruANtd58Cn7FE7yD+7hPlaV5Qae+NEAerTaR3zvwNYsR7S2VLx7wc2o4pR
gyQsxtiDICla9chSzZFueo3gP7BhMny2eCtGeMFgCvpvd568T/5lzvYpPjzZoM8B
0Gci66GsdUrVnVuc7/Fzt96MS/OrhzOdmxErHpUqZ0dShCfJ7cMSmq8sUu9kLeYD
h5/dRBfUvRJUW93pEkx6zBFPHRkIbbsPj8BkvstqPfOURgbm/67lN0RkOV8zR/EE
V94Lobtd6oA4ivTO1qfAlgHUD7ZYZ7tn5VUgLbfm5zjEwaDyUw7Prv94Nyu1/S32
nYuwOhpr+qY61D0aGhyDlXF809Y+n4ynppz2Vd4YbtgwOH5X48blVybZzVYOT+lq
FNij67J0GmKAVtpNCkiPckbWaProHBYN8w/hNUjs90KW5Jz4SOOAUSqL9KmuSZ30
+NUGJw3uK70GUB9kw/J2IIxwwHdik/3FkX4aHmFPLiAuSVib8VCDYoLy+wUbNj2f
Xslxe9UKXFp1RzFxqT9raN5iGnzrX8tnI8R2Nf1MvQDdmuGigSuhBnHleQIg2bpc
WkUFcRfbTrwvPseq+s1lFobSxgj77aZRyHQvEHcyBjFLT5vtux4ICMKNpxyzNXaK
/2mbUQn3JWjLtGJaVyJURkBwLw1QZNBOeF8pwSgV/q9s1i5x1DJmmjv1lufksNBj
t3gAcIIFEp44l1rIWUxriWW9dkOm0UZAfsBKrixxBDUXBvaik+kTSfMj3Kkmi5sd
yasJHvcoXOd8TEz6oUCAApT21Y19xhwoUS89WX93h43+vT/vPrbGYaXI28D0XTHN
LlEm2HjCTnV5OkAAzzZre3T4F5JuohpFQ6TiS9jb8mzlExmUgoaJernYpQQln0IW
yKwPK86T0FYtpDjX52EmFIfF/8/aMQNjQU9xmKJ1qcQ=
`protect END_PROTECTED
