`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9iCytVxuuMYfY++cHaFBAgiBt5SCz6YKzlNHshGwe2qHzWBmB6mT5pQ0euS2S7vg
VpGRrUHtM08AmxngyfgLcFIQxEZ70QXdhQtlsKrMNhjaN97bFIu46KXfdrEuzCKW
NKk+fFf8OObLE3U29OHjK2Q/PrH75MMLrDStWYqMMMEXeIkbPFbpjuVZ1bmxknRo
d58C3P9L92e4UVsWn5NBHVG1+qhCwyOVKxC247aD9oA0c6chV1SvtbISFqMzGtlw
GS//OPufhNvILr29pyDCOYFLwtLpzrpQn9ryPmwX3y91BzioR6pJFUECjP0QqTfq
XRtjK/ksN5wM6kF4Drb+FTRpkGwljlNXpw+cfLEb/QR38gM3NR594PCi4F1WCOea
I+kX9nVxQKyjmQb3iFrKoJBPLFkWAWwZm9qDO2Ux4tjjs++SijzgFeOCZMKFTtht
YdNJtNpi6lm+wsP5vkhbk5G/fgGmk+aIscZTwGKaX8KFvHsVohLh9z4cWtAqWOU1
SeWB3l3KCik+yOpL8TJYfUBK1PK7Cf9PVt/mi7r+l86C+074DQOdpC1UHcjiLqzw
e5T2xVD6WQxDmRxNhMhoEdVeQDwRL2RFnqZNa6ZQ9HDESeyRZbc6KNFvMleIahYk
OgV3R5ZjaNOXiWtl15Keia3bIaobu+OzlvhHQri6YFYdawPwwNtYGfu3wBt+ZWXa
dk9quqEpWSeAJyT+GqagOBQdMSSE2nFIgRof+easH9xiBg/bqz3pNwE7V2Bk5jhW
20n5MV3sMHYg6xf66DfvrkLGXfJdLXvj5L88xR01dUAsqHZiFI02fatBao31yGc+
SAhVT20eapzaaU8v+k7WeYJbeo9FoimomLQjcCH5o5dvbZGy0Id/bouSFfy/duZW
d59zMkR9kOi5uoWxkIUfxIoPfqbUWYhcpCUo1ppifqvFKN2apSrT6q1jVZWjvc61
cOqinqi8mkbqBXXI9A/+MMi/jTpVBHKIW9pS5qc7P15M9yIhAjfECJQrL2bQeJAz
WQL22dwiEqnAvzfv/hqFqm9WC80m832PFprguciAO9/gdFGEuWQK/aJhRfOzB3Dn
d1S9nICQecaUTYb1p/6+U33EA/IfE8IIq4TDY1v9UEIzGhHUfyENRRY1ftuuQP5n
dOVdX7xuxkVFWXTQNeD22nHmmPpGbolEv8/XXnvcaEUPnIJdSaEeFzAD0aQBpop8
`protect END_PROTECTED
