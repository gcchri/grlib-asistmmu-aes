`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZtuhWnmkinSW10Fdgwd4oDbWDeKPx0EApsz452rZzFNpCjjEFt8rmlNzRMtwtIa6
u1pc6bFKsd0KpuuFUQmuSpPx6u6Jo87lptMaa/K+xJGK6TDSrDVvmOzn4ybbvuB9
lfCchUpDyrpg1VzM6VZYovSIM8Rl/nzNwMh/vhxqQcT2Vks/1q4d+oKPY4F7p6B4
ka/1u2RwQlJ9izAGNnhgth8N03wODgHMZ5anO+lZjhSWVj4WPVVYOMMv83k7T9ls
lnmVWwMX1EkowXeeW0u8VI9ImHo1gtO7hty/Z9C6EBFSWCqvW6zMRPm8/h/pKiVC
W1qGsAc8GuEYuVp/8aFKYosNJ59hZh/er9OJm0a1cbeHLQ5SVVIAKq505Gvg4cW6
9ZBw/TW4z/B/YlL1NLQjwbkrQpY/NWKnthdLfSAWHGo50DEMJ2oCbJFBJw4DT3VI
I2KuJXFhEsVgB+oLlgveEKm2AGtppVqXej+S4kXDwY0qArvxyHuxb39zOYAObxsu
`protect END_PROTECTED
