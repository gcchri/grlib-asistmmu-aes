`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sv4naK7wmZDqYOwfowtCs7xL0U3akEV4i3w48EI1EGKwwnDi0L0wQy5AmmxJ/nM/
TUGFXSNJRG8ZE8qExhwG9LCoEHqY5WjmhKe/YiD4/pe/p+XCw1P4BKz9kWAXGN8O
XRqJT8XXulGzHsExnDkHa41rQIf+0OWgDoWUueUvoc9NP3XQ7peSnG+g+zLPIbyf
UFQfZpUrLrkU0w7XkE6GfYxtcqIDcRs43NisTr1hdZ4M/Ga8rwr26jfT66ah5GvR
xpbg8jIN+eY49BuF17jcrl0I7KJzFHBWaiA3Ig1e+s9pu7DW4hXZhqYI0Cer9QVA
ldunAFH1vxJsrgQ3z1Ptwastn636e7Te+Ra+7e2SS0MU9UuBPuaXq96K11vRCgDO
WfG8ui81E1O+AC8024fu1Zj2XzBF3a/COeI4Ccp0pMm5E+N/8sH9lck247zXzsMy
WlFjTQhqpFrGM+GJsuwtMz8wXOpoVMgHOf4WKC4cW4jKQR2B1L0TBrhU2OrzJeI4
`protect END_PROTECTED
