`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dKgXzR0GMYVhUid4O8AS5hIPyJAyvIH2IXlMtvX4czZu+QDDFUwLO+aze3XC7kiH
EVXXa+S8JMyDSCaWkSVLT2qgXx7XDHJr/nxkbFOTgZcoHgtWLKu/u/a49M/hOLo2
s7nAKw8QCytNoSHG8qbVI64wZnQmVimE0JzUUsH2Img9YBps5ooCyp8SFLTvRlPX
a5CtKYRCOts+fH8Z09BGMDJUdfMtZnEc/fhvsLSnMFkC5ehL44u/XJz4p9fgncs9
LAzDoFp/iVUHxThumG00emKFw29wWMnQs3QOIx+OJqOaSuWo2+4bdQD5K8v7lqO/
dOlUAokggDvvmRKTT2LBxTM0UOVgsDjswEDOCr6djnpl2v/nThCVQOmMuqo6J03h
XGIJBULrxp8Zjy10MwXvzfSIAZ4oLk6quMFA8cvr7RVOaOJ+PnT2W7NJfefH4RZ5
dM8ZJ033lJhDrRV51jAIPPVwmTQ6tsNyHVngZj46wjLTIGUI6zU/KN9MDfITEsFH
gbqLl7J4ybCwtGeYHyKHtxEzJf5AggKfL3EiLpV7HaY1XfrUHH6i/6TfN7mduodP
O642bH2S4Gy53vruEsuN6k0BF6v4brd6mbo8+KbWnp/OfeLZcCH+ThYiN2SX5+Ry
LD8eh+QMtf/A6g5k6D31NVKJ5bOFcu+s2nr8Zqm8NqqrmRob+C26MwD/+Lq53gKw
6FrRev/Fio4/DQ16PDq99rOjZPSW0K4lT7GgF3rGg5W86ye8J3NEXZX1xZqBhREW
wJVtNvVcT9mUn+6EFn4+ydGGFmpL1ZFy2bn7TM6Cp1jds0NPyj2tYDPeyD0feWDI
NRV8TaNt+Ta/HKu7NHPnimnXr1hNvGx0PbI0E5jXAt9T4VGqEjEW7HNBL9cWlPTx
uCyVv1dD6Qw/IaDqjSbWHesr8WEQUiH1W7Cayh4w6FS+n4RuIyhIbB7Ud6iSY/aI
mNy/C8rYwX8wntMnOFnrr0pzyJzONjkapH/QT+MEhd2SnsEf8AE1Z2CKSsdybO8A
JrGYBq4lYQhHEw8KrGf5a/j2H/2dZ7aXtROSdOrdeZDG3OUGKCGp4xpR+cAhETPI
4rL9byswhJ2ikSp9c2Fbueib8/OD/iqDaXZ3gpHTstadplrlkvt2b/B6hLm93ZWZ
Q9AwZUnhkYMUpH/xndE37zbF0wk8BOyd61MiCSln3ecNpP8wmF9PfN21JDBJZFhi
7rIu5PFZzGJtvp9Yk62WWEk5N3cdGj756es9LX9jA5UjiyCafgpAAm22wBrKSJLa
wO/kHnCItdV10/pVwYCGek90zogxzq87IGt1aqUuLUaxiv3cwJE0pGeJ9mbXfvN5
2k06TGh3XlEDT7COkeXMqTRb2fZh2X3wl9CpXIE2bsCPokUXTOipYbMFR0cZb5Ow
1fHkHpsYDrpO1Vqo2VSQTnsSxW3mDme3vR6/cyFGQRf27QUuxi/tfruX/HkgYBuk
VXgeVBNbgA5iONJIc7Cqh6c9FSOWaZauDYDGYerMfQ/9ML7172imnXYeS0oRHnl1
gFq+tYh2bTauc0q/CtHcN3BB3fiEKDbqabD/+c34xgkbI4Ncl1DAHZFH29UaMNhU
XntawM5vr604Zkac3TsV1enAV2OFIMxI4/dcd4E61r5qOddIrP0qOCqueBwe2Un8
/URs634Am81Kjq23us7xC4EYseaPOutGaFkHEQRjVqAC4TQ1+lU2GdVnyc8cJk3J
KCvMIx7QE1Lu0NWbGB/SoXR+Gi7ctDcNztvcTKCmIQd/IYtVMn0ZpBYBIibH4OE3
q8+Uu5FRg+/6CGkTreaSONAJQP+AqJ22I1jI92fTJ1eIvnXm2+gsTfHwpmGnZIdi
/+xVKK6GqLBoOjS5ldI1aACjXD8wDhfSx2b3gd9anGKJt/f5DmdUiL1pqsUhAY0f
RqVrAXP/MAtOnslTJYDS0w8iLX0yafnVL/WUtfL2vXtpBV3DQf2XfRlAMSOfIWdC
RphpA6O7ie/b2xFg3ck41STZPQd1IFST7SI5TptnPpyj4px5TaMxr/Y07H+VhJw6
itxCgYNTpj2M4Lh0KXKkDjler1tyll38WGrYrN4/xbwyednpc3ZGqb4NE1CKBzLX
lUVPWwZ1kcKMr2FYbxDdxPQRjJc6aofk9iAHuWUaDzh9GpoYKouuzj35DZVElhON
PxGTAVxTaeGm4zeCOSWcgjKfF6dejz0hWoTFBPJh1XIBymMHtRsJ83zkgKysdTvK
IgpDOPMgwR7/52Pr8JFUDSNPVVfhLIgx9ZPn9CUVxjxgOP+M1tXAsuWtJb/vZ/AF
RxFXfR8CMKz8MRzcLPIMd/HJV70+9pau/3pttjJWVb14JnTnTm1B2HmviXn1re29
wtuC0eIznKjIAsSpjPTTL0IWKbFzIdzMSDkjvvRpVQ0bBp9YnqIuBdAyZP+HrXWC
/ws8Cf/+EfTSPCgX/B+AUMoxUMJ8j1UKTGuqxoH7+t//CD6utNWogUNT0mFxFzJm
In9e2UT6m/V2BkbA2P5a6PhQTArYrpg/RragVx0snsVvTCZGPzmrv7dFGfvnLIif
WeSxxb/h4zcaRSDo5pLUqkX4xq1u33U4zjipj0Er+JRlLiUWtcUMOu4AcyWIAOqw
WEwrxPBc3jCigVtry1T7BVJGoptAp/djDotFlzSkTYqIx+LxcfXjvV9JwBABTGvR
EC/gHPVwuG2T0BId3DIfT7SO5lU36pXnPLrZV1IXhv1WiJQUw12dRoSx3X7EpmWY
Ci9ODSYfyEcuuXZW7mIy1LtlFyrdj3ckjwEX/A0BkcbJpFDX2r8cnpEUTIYg+D3V
ctfchzxk6ETqC1zpNndB1nTMEGGFt8vJNXip6QzYbTuGCQRv3Vyupq34WiHaPnq9
oG+juiXwfhw6szH0bQ0fuy5DCLqg08ZarlsDLPKYvTwEWCdU/CVqfGUjUiUpJSeh
iGEtLR1abiLPXSIzC9WWdYv7zoMdwd1w9nuxEmm+ofZcPbKECIIFQdoi6EygofQ8
N40LPJriIsOVkyEbcm5m/uTGOVWWnpI7ks0KmdoqVBKVExdZGPwqTRAG0eshhdIY
hD2jL3LQVRysKb5l6F7hsv1F0Jix6BQ11K4/5KNIF6AD/R/VUDE26j1PngsjHsJF
CM/mxrzKKKqdPwKejn1RVmZcgYiW4wwbYDAGscPe8TG1SlPIVVmU5fBRtPKnidVz
8P7TUMw/n7wEyD0ayqcMRrG9+SoI/a0OMC1T1u7wPb0TM4Jmw4KOqiDONtUFALgo
zChY7KPaNPTbzKwYQufTK0ksiuGFue3/2yn42tLwILxzU+jrwCGhkXRDQVpZplt4
eQLBhIlxeYQ2tczqBBC+ZxiMJi35IkTVkipAfEIFZ+IXojjW57jqWIU3HRIgv9rC
4U/ccvADyXT/EAJbdypKjlqAD7wR0e71omf+Olb6hBtIt772oRnSwT4Uk+xrNoVi
GIydERceIM2uki/d0GSbNsPScBHgV1P0fFdVfIvgtqqthugk6R725QVWH29M176Y
Y3YxOOwaGbX/KoMLO69huQaE5kifDPmVZEL6p1R2Ntrr3CXdu27i1eYSyvMQuWnJ
JerQ9WvRtYpIAoAnkb3qrHCZ1CrvIhnhIaNnCKhqx0l37kPxgYzuKWERbWcRwCdN
2aeFgWfGz5q+wtZXoYCELkmzLbEuXmKXxTgd1SSVuN+d3rm+HgsABuzL6lsgOtS6
Ma6EEesLZGefxXwurZyR13u3PvIsgcIIaVAylSKI2TndbBkq39fu7fvN+6huTbwF
HKz/OmY1T6ki2po8yb0cTnbBXEO7ZlgkaBalzVbs8t6D1l7VVWECvcnpiJDyRDha
H6xltmn2D63dTkwb764h1enxo8yK/lQ4p/H/36Dzy4jgXlti1dEueVKV7CGTQ5xR
d7m3bNTzQv9L1AA/nKv9ZDDuxAKDvi6FlfXQ51gBDW+uLxGz5CohmTcDn6FvK8no
YP6AMNxU7b+5svj0EkxFufvbjDNC0qN2ZiYHKRyJjtPeqlbwYWajYxaYC6eIzHFB
CxFwSeBvYVafUo1Mx7FlIbTVkICgeEE6rkHsZatls9FtqkGm12kqQ53VS4//d6l/
KdUS/kpKXndwLKP0kPZ09Yig7Suyo6iA3e5bWkA+cUTaRyxe3i/WO1tav1oGpcK9
YOeAAQjflVOtRT93l2EanG6dyswnjEcVKbDIszmP5hxsOp3U5JPjxpiFX04fuLS5
BHqKCnRyLtZYflLoWMGjBKV0fzEkpZ5eiQvARVB4dJeCxYIRCcf9anBeFcrOjj2D
IC2ypuqFDuj+sgW3UtwMdex6jUdQ57xT5Ox6WBWclH/bAnTKRxouCNbK80kHy+c6
ZKuVoebvOP0COysUlFYVuxiP/IN8lbb6lSHun3q+LF9mUfN33joQAKZ1X6d6nb1r
p5JhzgPxCZRXAS//TRms80KfzPhjb53g1uym63u21f7t8kgGJpFuWKbEvaVyFE3k
BaEJQBaExkWeDs4w3lxr/G564fDSykTHYLA04eMacsT7f04Dda6GqIFC5SSrLUsJ
bsGlkylt9AmnXu/wgbb46ixQ9sPIjzSobXMEDX1y2P55vHRfp5DSlAgcOyhoxP26
yON+o4IvlIDvcce/yjNaM2u/pG2lffNhTY+av52wfJcLdxj5wOEKYbngDrj00C+l
`protect END_PROTECTED
