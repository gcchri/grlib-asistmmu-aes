`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p+gzpZ20ZetTxNFca93A4BqwSmHCfvYVR9hf/vsXRR5CYUD7Yizb8dpT7vSMFYua
dgJSwBVt9r6C4dE+5mWk+i+zXYF7vhqH4CVG/uFK54MfC3qPHMY7VXAmyVixpsU2
WF3DP5nZrrRxnAg5KO/I7sHQIYla2dpRAikE1nzNiLYS41gGx2iTr/pd/nR+avGs
Kal8NMjV5JU065gHf8HQ7sPOFIm5wnkamHA9Bwm/zcJQ1PLTYhEbRGHec4G+Kt75
`protect END_PROTECTED
