`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZJcsDKMAEzixJ5V/9QL8alitaH1uCPN7wL2m6gTinqBEn3lME9BJSK37t85AZrx4
hKumJLSvegTpychD6ihvfnZ3uZO4+yIFmI49bfr7NNtxivEmZR3PHzblnAdy1ybY
55KH7DVMteYcFJe6IE+SACxT6auk2AZ7ek/oZTSx+h68qdQPP/YWEG+iznU7aYc/
t8BW5yDVOtlxzkjhGrY7gJlGoEMJfYatwZ9zGokdbB300S5iZXyvH3kVB8o8sAz+
MP7ut2FV6EoBVLjL7+uJDGEjuW9c2YTUyyPO+p0hQTop7v09sbxyTSuKsYU7t9zQ
vk92p8kQTJeHFGOuAtRflLavEPft3LOvnL+cELLcDql8DhqDYv3/+xB4poGXnklH
V8ytKnJX8yYINeotisBS6ukcNfWUwOzJFYo51FPB2D+nvMk7tIYosJfaI1dyRLbu
q+H5plLoE4k4sWop5DO/iyewAB7g05oc67gVp3GR7Yq+P5Z46b3hz+Xs8r4wAEGu
M2Rdbrnx1utvIzyIW9oqOX00PzgLso5/AfvRplQaDqDBiYwodAzjFz6QcYWyDKGb
fSfXAk5ks3OTKse6zIri65iLCV3PbEiPAPlaR6yQxHEHpjTJ2XURVbsLaraKnQ5N
ZFX34TNYh1FLP54Q6sFuPTLzLx+v+uRa4qbJaeR0M/ydGkvXuWu4sZASm48xFUps
uZS/k0F4cLD8XobqCqTCUwpT7nsnoh50eFhttRJQq4vzWe8kOofkEHixkNlfeTpY
+HcB0S0Qxvc+S3Gj1/oU4w==
`protect END_PROTECTED
