`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iaSqrZf6Gj3XiBfO0c5gDGq34FaWCEAjW8pMT2h7JoUyJkXwKCCbNEWYMTBERz9G
8bqio8/0RywiKo510biEUjUl7HQJKQYTan4qHPzR3n0JemJG/5gMsAwdddE4VoKU
PateUQSrxd9lw+ftzK+tl4Xbd9FBXTS9hxj9XSJtd2Lbv9FNjit/F3ZxUHWTR0Dy
D9+r+83iOmcpnG/K4YykWLqxeAAQvhSP/FoHxHWydSEbaXLxYa9Tph9E1VyYAGmc
aI3jmSI0uRKsvDGLDSxpNQJmAeJiLJpYSacIxueDw6ju9S2QZRFYDob+cRbq6wGr
lgEWBBLEn9gXrdDlC+XBei/8UrQyVDUTBAx84KH9nOYNX6E8iziKBLLYiNk/F/aX
Z9RrrOLZ7VYBrMoL33zfqA6HAynHC9rnM4g68Z1rLWoEODY6G5dgfN5tUlvW7A7Q
RKNQ2ZX3sUuo8jmKbiKUHCxBP8ri3pQrkQs+8C4dD5Ubj9WJj48Ucz0lDZHAWR6I
`protect END_PROTECTED
