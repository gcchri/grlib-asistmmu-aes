`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gzHjqpwmYe3wr6ez0taW2gpyLMjoZk7NKNzNv4njYAaD+xknQK9rGtioJYjqJK+2
WKjY9qUidWgjKqOMS+CsbR/yWOyrkE2naXH0peKmO3S4a6imJ4Md2kQR8/WHR15y
071NXxdyPdhRb/f3h7V54T2ok7Ep+ocox7m2/fWXm5VfAFQ8Lox4MdWHoLSa3O/u
jM6in/4p6SBJ1oaA5vMFNgKy47X6+XVfhO+XfMRz0ijFhAUnt0S0ZSA27wbuVJRB
vBskadGcna1S4DOe63W8o6qpqQVoxwkdmSlISHGUgEE7/KC2OAvWBEFiJdHy5ZP/
NzunbTJVNbNBGxvogtfeVBr1MAciCkp842Si0VMcxTTQAHaJt0OTkBRXmQW/mvpc
zsLjRp0bYjcZhvrv6Bv1h68HilQmkzeaRqf9XOn9mOKDFeyMhUrTwbughy1/aVy3
xm99Z9KZxfWhVDCSWL8pv7vFdgdeLKcO+oc0CxFhognfq7GPxwN7HXnDpmI4Nndd
Ykj9bXYdXXuejcWFRdsq24kUiWJ+YH8Mo2XN43oeMUxy1EzokGd5vg3WB7RJ8Jcn
nB2wMlxnRwyWpDtTiilv9SQAFZeS3oKo67yJxeO3EmBGLkC+8G8NooklT9ia8osW
vC737HgGlnP29HbzjtGyJU9Wh85rcXLs8dZuamrOBkr/+kpyz6kAizf6NLVTnABa
+EZB8+Br7opjjuEKUubKkApRokzbEXDPDzPj9fx9ply9fytlDtKSlZUptKblMneo
oc1yJtMSiNnGd/KQbI4sG/2yPSKNkNUWNnAcaG6o9AEVqfbMELu4TjNmdxuY5yz3
ZyAAjh4E+n0j15/Dq4nPHOLiEjSj1dSzLLsppnYJhd9KolqDrE50FUdNbwDYd10M
u4g/U2qP+w/DgP4LU3xpDE+ZY3dT5OuJUKL+2SWg5Bmhk5dkYyBAJZ0Y4JufNKKt
ZyA2KW7KhfMgHoQVtprmNBk2KohXmKhH/f9Tvb1Q3o0HeKeOs/dnzgqPmJbmk4uA
eVrJCB5ZBCdroWSMmVnSi6odYzwYeP8i6zJz50RQPJfdQzC5Vnqb26G+3HWo+M9a
pPzuX5D6L8XHc/s3Wd/Fe14+suojyP58njK3qjKrpVyh532rKDAvsQEm7ehgN4Ya
wWW1toj/YiqybINQsiuX4IHG4XYSblvdd6Nda3JQ4EZTTbdUnYfEPlJwQ/Pd60EJ
dbsMBqNv2E3lVXOD0Lm2aDMcWTggR0YaspMZtBdyihYhsag+aFoUdLMh/rhHaoIV
chZa0fIg3T8asE6/uUvQEQQXVAITrn4+wNEy0RC255btVRHhansaMge7yY2Zfw9K
ZYN0UCRZG0jVtU5yi7yJG9i2ZyjwU1qS30iX9ydj5+H5B+uVwH1OSOKvJeCmKmQa
Alt8U9Ft4p7sv2bplwhC7XuP0lCXJn/voUTIEe5gQGg+o8pAMVDW1g8x+dpsUDuT
LgTz+jtvC2KlaLTz6GkOnGhOA6IYQnpOMZOhpQ9STI/t34bnHK7dXG61tWcNy7yn
KS8/SUn6ZrrezVI/M6VSqq9w69HbcqtTunmG7uojZzEycRr7Jc+gjVMDFKjQOiV1
iLnBGjskKD6G7gQSQMLIzJmHsiCp+4aIvDFITZzlP8kDYW0ZXBANZCgGRT6zbySF
WOalhbDhVPiuTmI0tRbCUIgFnI8NARYTgSj8mUjWBS/+x9KnmbS/WIrM1J2Ix8kR
EKFGRFn9n6SDzO1tQcvpsmqFGx+C9PWGS2AOzmBHPdSb2KzaLp3x5P/T27826eLf
mhwFGLo1Q+6DMsNrjrL+BF2O7YYyJnohr3XeT3kOE5GFKornBl9T1U55oKXaEkVB
mmlBaPLTRwlC6uXQY4+NvxDq8cYdeeoxFpPMbp7O4etviqbi8jKtgcXnnOtnhbRC
CD43TGJep8BV9vYHrP1hgh1752USwtHsbIUTNK1eRDF9lDYN4Yifxf0oida29e2/
sU6u+4KC8ZX6rRmTgjSGvCbq76Mipl66emjIz5jl174s+vn35hSMBXIUHqG9cfBO
xDfTQDfii/mgt87pviHB/CB3q7Ac04h5zTgxSWsUpZnYGBn1OrikddSI7Dn+dL/5
OBRMgMQBxkXjq0U3RFE/2CNHTV8lAItcQUfYRaieNUzfKd2KVe64d3/WHrRPGCwt
hxI6EG2r3SJDOzNuPpdI8cUahktXNihapwiwpTr8rFowaPFUg+pQIjX+EbYsulTD
io6EbrMHeaA/213rjj/Rg3pozakBcj+4dlue+LM2S+SzTzWEVSXGjEDfbg9gd8sx
pvz4USsVq8b/9pxQAo6tjhasGwSWuqbCicLNtog0ZDrxbQX4zQTfWBOUUnx6VfWT
4bpzlQCG191Zb+vAufZTG7DnPQfaSE+YcVlb9Az/TxX9zvci3mj5O/a/1zh6UoU3
cvgJCFHjQ1cDSfDWuBITimTpijYZRtcTDLntAXacbGQNzS3jnOEkUgftPWSxb0bB
ALBVmkrg2ldqEROtRaxwIklCVEJeMsbY2WHUpthFOwOxJy0oN+ZIAM759X437ZWh
3JM5sXF4Xe7dxSDUpv1ja7XpYhZ4OjINwggf8tMS0V/wlpPErDM/nD5O6ZsxG8Xp
o/JdQauUAqj0rxurvDXrWNlP+jKDQUIrW7mKdbU3fv6dywg2W9KQqkYkeNOt52q4
+pfWzGcewrNbTH2xIv/sVZpabGoTYE7GRTiBTxm/taD0ovOQyfmG+P6H+I/5JLTQ
2ha4TJuEwYeSjIyl3mt8rZpDH1FncykHukfQ8Yg5U0z8kmG5T86/FJ1hxiTpy/h2
Pfp66LCWJlDMcyhpTWsKYvMrYwygjrs+BeXwY/2vfGYCnv3VPk3r/TNUac9+ljgd
w1eGun0hu8XbSVakVE13IAmDa6XaBLPMIkb2HFnAUYH6aZY/t8pSQqf1iQ0/xzbV
/dtz+TzTj2sD0EFUpJJvaPcY5dB5tWEoR3BQtzlX5GGG2A4U15phG+D0IN1uCVjP
7Dks6epJWhBlpeftsIDhTvaLEVF1NL/G7JgXUr1A9GPc5rDlMCJarI/2ynJSMgu/
/ngqN/wNYp778sJviB1YpYIcfTN5+pswVLb+5cv8/vq8l8zqoB64ggBe2+km4vhy
BKGOF4gtsus9f7rJMYNrqg9DUiK7SOJqarGzGRNydAI0bGgdC78WI0AA1XmsL3x9
005OeHR9LOAYdgD3i7JZU6yVpvtqzqj/QPcPShv9/MfGkbumg02mxeG3RN+FB26I
hnAJD/Q10alLXqP47HDRjInlm3iuw0H8lF8vihCBaCdFAUx8v/Ri+rCXJ8RuC12y
/qZJJl2mg7u0De4I4WEExNKy3ScFKZJJ+IA2pGBse9oXr+iI0Iczifyy4wRXQmLu
9pPcq4Kgw4VQ8pJaaNxFCYOYkqYkj+eMMoOX3G2P2Judkc++NutpzwyLeYHprZAB
Ftmr+VcryF+cRWHRdsuBP2pQBgdw3BrElPvzxfTJY6XIxLCjQMXPt3gtKP1mGx12
3Z8JzcNgbknSyth6QofhdmXYNFcYRezl/R55ms4V035y9jzJsNd0sZrtULZDACTc
eSUMa0tFYJ46Cewip02JyoJF7Zh3ZN/NQV4E9QmclLOYfR6W653Jfq/0heAR/l6Y
v/T6ZGHGO7rLaCVmS9hlrsewTsU3Ccbp7DYikuyFdz5mdf8WJX+BaXvYN/Tjo2iS
PReQo7vuiDuFk8Hl6sHSfOD3KJMVAF5JaVlhAd+j/OI1FqrlkbN2QVkDIAPnzrrr
ADWBL5osGwkIrcLUnfA4oEVAHXtVXGDqfeHJBC83js4PPwEa/DJJbxQum9Hx5Irr
rWcNha3B3HUBBaRF3sr47UknxntFc2dFgPol1fQW7ET+3GyeZe/npUg9YbiTg4ao
PytT0TBvcOqcvXkRihn0+rDe0K0ru3afr88WP3izn6OgC2wqBiG7eXptCUM22yFr
qJseSIh7Ase008+odFVufQ5FmCPhGUsj5wHhGofCYgT6IaltwwkbAnTiTLoQmOpx
N9bxrXtA7z+zWE+CzQXiU5bUUbh7muvn00BiEUXca1IAvcIfM2lY/2fEqZfJkoDj
ijVK/infORmRS717W8AjCb4uc4JiD0QozfmxnxwE6Hz8hlw48vgPgd7KLoJ+a+9S
FNnwCqDeQK6VhwsffIMP79w1sUBv6IcBjAT/DN8sPWoDZGTXmuQDjxvhWp4lCGkU
pE/1XsZcDHs4crIYqw7jIHwqYK211Hx17EMnAKxnpEHT/at8VEFCVPC3FAI1ysIy
eCfwOfXQnkKxA9zUEgUQYRVu44Ack13hzQbIfGFIupATS7Xv3vqJwO9/aISjTq0h
8aaIQgsrVBFrAiKB7RwNFPrtFgj6v2s6JHqgszTZNS4mOPxbBpnGzq3s0v8H3wwl
sY4WQGdS9dC0GV0JmgDvEgPMN6PqbN0X5sJ86w2qJ0Pavz2b/flnv0gNsyQVZnat
caUNuynGlcKSy0W4WkxoqBQRZXc91Iu6Z0sPNR0QP44nuaInDQP921KyilZ56Wav
fIzKU7Wz/kuM9vmT3rue/QkF58vrnok8j4OFNz7mdkmNPW3DHAzF9sTeYLWyZ6R0
jVMKz6/j15taR1jqY/Oe8BxbyhrpZdkT/eZ7TsvCCcH6ZVN8sicXEsW0tkY+NgY+
9UjbeJfpPN/Y6H6DLQktSkKOOsWqgGvlLwGkK09oHSuZkrwb0mSqRBUxYrPhq8Qp
WJFZmhsDqNVOmQTz15y1yWrl/8YIZxbWB7SyyZTf/sYmMqVNgqLbeBFHI3xQdygJ
2bQlL42ciNlS2R++j6uzJQLbI5wBJOUCmxCwZeFcrilZX++cHlNcswrh/rq98t5W
X3KlBCq6p1rf3ETUB5e2xKvGjRD1x2e4vMOuFjljQaKqeQWdtgDXx6wWSIQlU2Fx
h/R4rdnkD0REPFv7rqwuGnaS8fMn4OZax1fhbsf6j/25cDjAdcSpqGD3nylea6oU
0HcGUQL8hZzTt+RDqa90TTYc9LoftM6bVEK9iBCK8pAJ3bQzS1FU0X2X6TJ8sxSR
4UxebmHtjZtv5D0NNTJztZ0r9E6/CBPqFf3jVLZazd4pemCS8cBNB7SpBF8siIQd
TCJi91PHavu7C4I4lhcYn2E7MF8bJZDTkpwuIY75FIXSSRJUl0HSB+ZBkEzLPc/z
lTxadk6MTLWa0b5xtTl2geMLi67tylYiM8nM1zMaLpDBddraHzpwN85LowNB0rVe
BvOKyNpjYwt4avy+tQvjPsAGUc5NUKHXVMl2Ryu9GA39EkrdK50M+nQxX6c3rJRf
QAO2NcHQeKeN0TJHlygF25GKMkJeq6rETLtDOnah/NxDDSBGkR0u5nVGMpzT9OWu
Nnt9fIg9Dp7DC0yJ/sL4cyriLUivPOmsAO+hmks1eYK4qJBYdvEksuHoUKM3nXCb
rmokqACsJub5Zga3EVNThOw0lVDtVaRDHhuak2xIAHiVMctyaLiT2GUdAyw2Ksv1
G81huaeSbeiXtS9/vwdRGNG12b1cyAA+Cz8HEriHmBjunh5NDwAzvFNyp2vhLEQj
CdSL/NF8zM4UyHvw9zazTh0EHVja/gRmm6GPiDvObC29vRv3102GI3wV71BStytY
Dqr3WDGaNhZVRPQFE0qR8bpUSdEep0wbVDniWnxO2kE6E5oBdAlyZQdZ5Fs3/2xT
L/raG/J+XZSIJr80iGWkAZ+4vHnlcbv8A+3CclFquWtH/z6KXTNDJ5WMksICJk0b
WMhBTX+QNdz+kHxU3SrwodLGn3BvbeYWEWwm5WaKmRMQWQRkhsQPrT6rUn3cV36m
kbzHQLUZhM7XMOYECm/QmaOGrxAPkwaNl1IScLSWevxtrpEVlizsKwt7TaaOXmq+
+0SeVM7qCbQAWniU+IqS6vwCBG1qm6Lh4pHCmjSh1szTUQxwYmjhhsRWaBcoim00
CyKiDqpir+n1eiRlyI3dKvimHZcukYjb5rNV97Fbo4EtUsZyGZDC7o0ocfyRtzV0
4YXwtLBSh9yLkERU1rnpSj803XodHQbCvHZUJuhUHZ/ay2I+qhUauSvT/CaWX1f2
JfaCX9DoN4CZ5fG2jAySR+GqyTrrDcgxnDrODkaE7kx3ybMi3vnc5tREDe6c1HCU
Hg6CQIJUpVQ6oTobN3z4qoQgtzy7kGlah3C7JCZyHpsWNCGJ1it4fIfE3OZhpRiM
WilH7st38lAYz0FvVpvFzPLRVwqquLm5PgSQ0jJBXC6Aip5V+mp7DqJsbRtWsi0Q
gzTmNLfij39Ny0OkRtg/gGFsb/TQag6x/an2h/AXXbQqNvund+5yKqJR1+dih4Jr
3GUk237r3bPC7Qgoq/hytAvaKxzNv7yx/HlxcyNAEIW8KlSLkmXE3x6Gb1/27D+T
yQTxHyOh0CmoafVbhDV2IgLARibA5R1TvjtkICzX3WJxlgKflh5lUD8ypZqqAprx
uQkY4nyYN15w7T7WEIqxWN31cbDY+tVaQQrrF+uaW25kBwnFqC6kFYI9/s+xBypw
4M/qWko9+Pn0E6nennAWr8dpW5S2ZlRnD9/s1B/3ADIBqipNsPec8xtG+73u79ho
7B2LsZvieQS+2j+tiCs9nDFaejnexAaQV9S0+sKJZUUMIgsfgKCkP89Dck3lCK2b
Lazdw/6CH/VXe+y45FcLSjEt0+IJoczh8eLkNMlZ2zfyvWDtOKaZUmeh7PZsu6Td
Y1BC/kqk8nURr6I9RMCnXL3vx88f+aeaMBmAe4AxAQSw8yzrQWnv59Z4zSDd1VKQ
6W+5rUC4aiI1JhsUOeTUeHtN9YPZhhWC7QoxWn1+of0+zkRqErBFF9n8PPfUq44T
vhnoSr0s7+4lfm52NjWxhkGgZHjfcXByN9WZDBfRgEby5kUaiZ3+Vd5/y9mibd89
QKLaFhGFwaR/s1D9LU2oHEhLGYHy/IxD5Nc8X0MSVEU3NNCqanDw2jGufJvWdlqi
a08DjHvU7B2lx08gnF2tRTvwqxDoHPiiinq6QEaGDBKz/zc48AkGvLh6kJskFhER
PIkJzksMfa7F/gHJsAx4fawRaszWo7F1Qdp7fVKbE3hyo5GYdcvBGPNLToJH5gbw
4cFy+I1S1KaZqUCNLYDPhvA46luPhadOd+2+3I3UkZXkRxktEgSKVQ5TvfiQZw3y
kZrGKlVc/kJUaQ055HQVAivGgRHT4ZUvAF2HDM4R8WP3UUSQ9xuIK86jwgZa0lKl
Z6dzY/pKdflxlJPOpc/brQzcYF+R2QsDLaRfZ0nJqVwX+myuE+ZKIucwpYCe6riW
NhGBbbKSH0S3foEshIRLasO29FaH16OOPTIgPNsGQCITs0laPARbKA3nn7flGg0d
KTTQvrAB30XzHXMcWZ5wU1xKBsGbNaHLgzqoLmBUl6B6n0NNaW0H3e4MyRE1p/kZ
R+o39V08v7v4omsCEzEP61MGrr3dc61YtDTwEKQDTKrd4TpMh0nt32a4c66CSeG8
ToyQhN0WFC7D5wnSpuPMTrJIGItEx3YVhPFaElldQjAuFVgzNX5tceLBO13KNfyo
ONL3uVBIJuSd2q3WrRBXeOMDTHvR6Xb350qSjVtNrCSOVOHmqpRK7T9DYtrhU4mG
n6OjFwKxuc3F/T6g9Ryam6fg61gYxaBFm4835xnxfisQIUY5gnCoW4TG1SaWJa/P
d1TaJT4oCP+1lnkuRLTWzj4dfkTnKTsVTmU8MXrR7imbKTVgcM5dP+FJ+aMPBWfg
JOP4+fxTVE90X9y/4D6LKw6KoAJy74DB2AaNW1cPaPVBsHlkazTvkrboJFoQIM4g
r4eU/A7kgrnC3Q65s+Ge3ZjATe3raMwpBhhvgMW5Uzv5dPvVG3yWSa3wPioNqhxv
g6eUK1zRy+0EpTnZt4TxMUeOy42aiKeq3MinLIV0TNWsLFk5YMP5fYsMGCzjgkzj
z6uQX4q2Rlb8XNSLXoGGtIQrhBJjqJoAdIT2lVE7bQqTUlsbw67GwixZePWksZSU
IhZRdvRZDx50L4ubmEtI03xjh9qWy+g3wAnk94NIrITSWeJcK1hEAvO7we2wR0GH
KcULl0fn3sZjmp+YOnJGV1ssNlH/zG8qzA2H5L89BufTFGg7sdl8L+FPPhv/QZkU
QUPdWwecsNhIupYoYk1ZVitko1p/wHY0AbbJcUUiyrTRsS73BxVfIzdp1kJx2/lH
X5JzdGDjz0FMoGhxhLGX6TexGN0dWV2Nkxb+0lCcb8piVMUAQIK9Mf2jiRdRTgfm
NfE04wv2TMg+JOCaTdNY3vQ6EXituQBRstNccRavrzIKhW9bxu98h9WRSOm8CH99
ehkCtnJ46qWFHep04EyqVsfsBurG7riJ11H9ta906MC2SEbvlChFO2fH/4GSGmsQ
kAQatT8DKLrSrJWFbtuLn33ZRFa2QPdsH3UQY8i0HRnMvxteL35CncQdMPzAVC/9
mMAkIYP6b2z6rEFkTBu+3OaTvzZkGqyWK0ie5Z8e88HnXNMieWxzpilzQbwHiDop
EweCQK7n7sTGILHIYKvaFkX1xuDL2U2xV3fJm1gIAeX+t0MDwkmH0Wr3uiXhDgs3
bOVvzXkiwJxwjNFj3wYuevPVe7cesM4rB2RIkag719rGUaCnSO+4v8tefBl65FYH
Zx1VjPOibip5lCzZQ2a3vNbIQtA4Se5YQJazbkhmuNQD6GvogaCbzGAyTudkFhlf
cnejtZ/1cc33P5RZZKnbqnTlriM3L+ExmFMCGhlc2G2oUgANZV1QoLc/f9udlqJ5
6aMwSiGi99Ug0ptbr7kkY1xER3ICe3fAW7fHR57FiPco7qgyBCJTuSWhI/lS87lD
tKXxEMfqGAYUAxO1KDuKB0EnlRCq8OWSmqaSjA4azUm+S+7XskNcDtAyDPrst34Y
2Ob4NC+GuLP+fF9sFMQ7cwwSVxkzzQUdKouIGPad6c3UzTx4XG6GzTaIQa9izH3E
KvwwJM66LbwJcZtUlko3CZihY/zckpxh/z6Rx5VwKVnU7bD+l9Av5cbUImQIiVRD
znMvQx1/NZy/1A+rSBit94FBlU4RhznJr2aa4tQ84nGpibvFKom6QcQwVd10emra
kNpUpWOGOPTgFeaNk3PCi1O4lMTa5FlogmdpVUFt5NEtD0hXQE83Polmyceg2TrH
/Tvt64Jd2N8Dhq84N9ojqZsUE1xF+ovSaBk0rp9HAAnRbO02Ep2euxu8aHF/s5P0
w22dmKhSCYi1PEvb0pCY85BboPjtwzlJu9fMoM/J+XiDh+as0QmzAV550gg21JV+
DLw/SS4VRd9j/stcxS9jTpUt6z1brQkHiI461MTJrKh3biFkErzYfKt58TIzj7Yg
rqdz7jCusVpAl37fExHvJeYwBkia2Cy95ihD7UCOudL2ghj3dVlUYweYz9jGYBwB
Yg4Htk2xRpMD+vmxhYTLi7VbukRoiD1t7su7G92hebsu0rfk7WKOnQLlT6dy9VpR
Ahh3i88mMX6OLtv8jeKTXYoLTaCAnJPw8GnVcCW65YclszmLA6uuUsnDMgxUWpIK
mx1DrcSBHgD1mgt4bxnQEPA0REa/X+aPceHKBZArJOwURZSwhM4p8HR2tX0dP5ey
kz5BmIZuSiMKmpPgl9XuwGNJtxycNIwX5RNCRh/AV/TqOSxz/L4//s7cwwea6F8V
2tOc7+f8PmTmZpfNn8BCsxyHVUUEGQIXyvlWH4lOKN8+Nb6jJpyf6WEZhFxNmvt6
HSesovnl+gCZdCLrm1Ts9JpT2uDRjpxYbUtr3qRTg7g6JWKDdW1fCCxRljJ2XmA1
a3nJDqfI0A0lJ4XCWohNw4qoLwg+2N70HqgEg+tSmw0I7JYmKTXas9c4F7xjJGxD
kBG8QNlrJ4AYCe9gUkjkQwFdpwWYvqkCrv0kPS5ZxN1qt+v9D+0z1MvzBV2zMaAn
7wKaYfvZZ9UZAryFsRvp6cv6zMhfJOb9Bgw8Q1uLxiU=
`protect END_PROTECTED
