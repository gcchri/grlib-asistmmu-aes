`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yI/RIO521tVAVu1y0zVI76czgbo4H/AjIG92eFFet7LGXwIVf0YwWQZvSQN13nxs
TjjkqiiMHnMcz/r+RaHCosdYeYERdahRm4IHR8oxxQxszy+eH1NL9YLIFKtOFW6t
QeKsG55KthP/gR8wWjg/oHIWJpYp2txOPExbjpwMny6wGQK34A2JhN05ddYVYtwX
C57Kw5GAGQF1eFVDjScLHu/gkR5ud7SYAFY//oxeo1xOzxsQz4zhVhLEcSlJBbVo
q+dCkvQ26K+d3yRR7WmFUKQEaKeUVhZi6ykOCr4a+DI4usGCpVwqNap2TDczuNwk
Y7FjvSCc1v/gAwX1i60JaiXQKc7L+6YNc9GJ7EvXcSkne5fSFjkVrVi+8Y7NgAcF
US0j7HHQJoOO+pIi/9mb97juwZVCoRToDaq6pjW8vzseGSZjj2p+j7aEvGLBIGu7
D6Wc/Lb+rVAsbYup75SKkxWUNQKZqwfS1GObYfO4LqIf0yPsWcn/rKad5jT+kqFU
yMbYinUVxjVSOgN14vpkPGFrMSaD97J5zwsVUFQHv4JZtMSvfGkaYQvYpprC7ZPr
lCTWUqhT1dwCi18E5YlwlNLHZROY/AAUXLt8i27fgdd8qgfnaeloiCwvhzXzxQr9
Sldydo13xWqaBic6/d67WblWd0mZMSe45upG/zp2Tg68I82OurInYjBaxfFz8Gn/
sbdJw/cYI9w3cflTdh38FA==
`protect END_PROTECTED
