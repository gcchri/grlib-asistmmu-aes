`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
avCMQbhZH5u2P3sYm97g+SN2OC7VR2Yk3m+59Jm57J3usYhhKfWBUfqPXE6E+hSb
JCD9P/aUMZ8oWJTvCR4DPsYJq4mRtAVe3gXy1ydsgPIOgZhePk1z5Bh2IcTARXNN
beCOLqJqoMyHsDme575Az9m6wW/CtlpAzv34BP/E3kDEKBZiw7x8qEPfwnj/KNA1
SH9J/UsXAS3AvGK1VHKl8hC3WQuaSgr+7tmcVhrZ5UV8G+DylzomfVNFV88gx2Bh
ECoKCTzVlKIHLXTGWZ6sCg==
`protect END_PROTECTED
