`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
78sc1HVB2Xe5yKgJNWNj4SrkotF6v0a6FO1KLUg7E+ccZGZRJ/tXaIATiiiRla6m
ihSPCpaMjFEmYd8+N0RCKekGSF9tU+yi1v4+6H4832uzqZLlmxd1376CmBDx066R
NyWxKfXy3FhUbKacFRc7DYsciBsX5DX7VNn+yrbNXkONO1mhn2lSVNiXBq3DyLLA
ga2O0erHbxKy7Ngmj0cYUHtYqGkvm+1I5CZsdBcBrSAsLq2FE5dqs10FFzW170nv
ZyhfFL20na9N/Qqxvg4hZyF1kvkdJovZYc00WmFBnExxx8795yH/cHK1mK8puD5M
30j0dD90VpGOhgi44A/2kGyfGDdRqcy1WsV2OzxRl+23/44yXYiDEMiPXN/XCUXN
wFY0U03kyYGnEzi83ykyQkyx801zt0W1uuxlplInAod4Kx9S92Y4PSON6zQ+IZ4P
m2K7wlZaV84xcPTDCI6vTzSLOOEp0JcX9GOBbBds96Lfe6AO2GU9N4SQ71eSrQu0
rFiKp31poFhbT/Sw0EwEHaY125YcChiII48GgZhUNscVyQpFGOzz60PZxPqcQIzc
Gk1AMQZViNSv8/kbjtrmYM8donLsmIYaRkeX0x7BbymNsR1tpJceNTv9+N+mAZLn
lEmhooi1wiuMrO6D/MjMRkU238ucPeZoYdm/Qim2xjV0x0+VoqJJY1D9tBUR+k8m
vIJUDuQmHYh94Pk5H8msoQbuSZB0KnQTak2ngQ4as/lmUF41nODKONkWpqbjbxgD
LVdTBQqfG+YOpc2IiU6naJu9dcXJDvtxOWGZ/kG3ERfhUORha6oEXKxOHbSQNaEo
gQ1lWCviMfwDAn0wQ8GaEPSY9/StQ2QL1XFYcvFaQatzTsh+Wt4Yc7irjr+zVml3
IDqmBucFeHSfqd/o17WfEoqMgLVfHEMcF7apSKY4EpXTOEZjK17hxEYnAkQxex4h
maj+mQrHcIEE0LiCNk/OpY61jtMRlb0oj7AZ20Oasa5gkSDl4Kv7bCz6+Gba25xq
/n8Y9/t9t6eXSFzlw4R5et540cQjd7uFppHH+02cBom+nxjBTubeAO1LUio9vEEa
lqW0uvRJkIhN5r7GV7Er/TeY4ye0qmauy0g60tlV1T/dOhO+wyF7k4tIhL2gRmI+
VAvg5DdeRSN9UtnxRJzZ/Wg63ap07++X/Eqo0p3JyXDXzH2gahIbe85bVIDk+gbE
SpehW9deGLENBKv2I31CYotp4qflJEn05+vJeugJgwU7AkaxUKV4Ptpm3qd6yec0
+Ob/wakc3OdvJ7oqDnsmJ2/Jvok/Ckl5yhPZfqRQ5wavOp5UxqsG4jltWmtxAqUS
KMiAt1bng0PzCF9qoZ/sKAH4VIuvQsi7c1J23mS6ciAQ+Wg+NloyFlgAHzWuZEd5
u3plXs1QMXKuppw/PQv4DA7m8WVTbf12fiUXS2I0z1gGmc+qmKGSCJeibcvE+vch
k7PU9fBn3fYTbFssbSJv7v/nEejZqIfiKoTbS+RRq8qdkQGfD29tz/EwUmd7gp6i
8X6vLQu2wyS80eIeqc3UkWrjCg1f0z2dbAVqZH0js6w=
`protect END_PROTECTED
