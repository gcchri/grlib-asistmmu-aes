`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jR3BGlG5J0S/yQDU3WQC8Bwq9qvLb3CvY0au3VjXQQgib7zI6GpKDdNgs2USzoqc
d+D7JiYbKnLwxk+6y5265FkTY06ugX2N0S4URfe+/vcUnKKZzefTvAO2YaX00buy
hgw8aw3qNjGOaNp9lSnrsprFD0nRKylM6ggcINkvLQgVB/MPLv4w6i+3gbedXps3
UR0z7JPhwh8bbkO5+zmiwoSgsSdxB2VopnTlG0SM5u29z5YYsZnr4buvQmmrLvv6
SSoW4CwKC4rbSCoPvvZgNWqUOQeFxekPA4B2I9Yk/BGAoVQMHL27tVdEREoEJ/dQ
p5Ae1bDX9VMCAWCWBvjkbmsTQHIy3en5/+gmGCRR6gzTFRWWIvbQiZ5Ya2hbfV2I
`protect END_PROTECTED
