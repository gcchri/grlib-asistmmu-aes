`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a7UNSrkD2VnA38USJSCvMh2cFbenn1UO9MzPf9hhNAkERfMs1Y33mCqCkM0bpoZR
QzQmbyJDTWndEebI3SZ/z8FyRbmclomAnlqL7y3B6Ti8tpDAci5dQKgpKCvBUW32
esbgN7kujYwkPYpHFRnS22la6OdGO4EhCHPv53yxYIP+5NoC6zRBuqfzOREyNNyi
Wj/lLp0hvEtRJd+FnsDMk/yPtuLeqcBz+NvMECf7lGIf9WTSKh92EDDtV2XVMt3m
Ef+c8IjKJLjKorZ8oF+yDCoEuV6vq9ZFOQSDJ3FBtorc5N2N0Hs4ieZJ2RolYN6+
tZi1oEwyqSVxv5UGE0Sm7cDPhVp2mbeDqreVUltSuE9Jak1CQDH1fYR2O7I0TfOZ
`protect END_PROTECTED
