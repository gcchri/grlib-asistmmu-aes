`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UzAp+VLp4ziyY1G4u/NUM7zrq3s3LC7jzZSYbTkaget6LfzkwaANl5hUFZ/8Zm1N
lATOqdxY7cI8SFOEklNMFl5ow+v+WxD7lmEAWiezZld9oLinUxBzpb0s0sEqZIwZ
+TnKcaurx9i+IlCH7GOlAsHSvjcMF+TMUuUkBJELPqLoUU1lXfzaNg6Nrzd/GoB3
iw9OXkJL0dzPcj/AcCxq5lhA38yDsA5NPf1qJnW1cVw57U3hE0fRVKsUIKHYaXBP
cWqRSnWobXPYyq9niiWcy3GdV8gkFCBz0VfY38rIUl7BvXBY2o6tHWZ0Ly8UwWrR
GvEGeUCLMO04GE6u0c8T12UnJkQlhdSQ7p8qKlHPnHwXRIdwLQnRxuEqMhawDdNN
ub5D0MoymBkBd57NMiE6zEWlBL1c3CfebcdJF7MSyr0Xr13QW5lMPz4atkcUmkBp
tSNVSwUJOwnZZc7tWAr4b5xDUtOQWAmXGxSXnnZd9RU=
`protect END_PROTECTED
