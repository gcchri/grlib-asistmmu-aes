`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6UNOL0dnV8xT55poFw0vv4CqH4A6FfVATAWQwZRVZDEwHS1kIxRUFa+ilwg6rIgs
0YR66U5jltjZea+M56ea/eUklBMoVvabspYDwD1qBwTY3fH981vHicOW9gsFKsKO
Ev3vhjnzOHRHuLf0YoJPk2wAP8p7M4lqj/7bcHGabVw0wpg+akYRvUwCPlLMqtcR
UEihFjb7CcA0jlgIgmmvmmoc9G11dCsxBBdRaL3cCRS5jUcxFgkjBPNPT4N1XuYj
Qs38hWDkASq+WBZRwRRRW6wxh1k5Kt46IdDSlH72hru3jmt+qPodG8SNIYbjncTa
wUVfffisArolIewJ47KNqO9s88ih0Re7FCDpoDA7EZFMyosCcrzdpUQUfoNF2rul
s3elkjTvnXPWbQfNjLv+60SLleFHjGyRtqeZjW9uzVU05D8Uti9WHya7HmD/2XaN
`protect END_PROTECTED
