`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BTNVvrsO1AqJXRKApZzTTtPNMUvUtXq77Wp9hGgUvsxo/0G6yZqI4mCkVyODDeif
vMWThRj9onDYo/eEgIgHDKSgVZfJx0uM8WxCQ6pLrldfbZw4GJx8SGRJrGISHuzM
ab4A8gqUhUQkCrA7fPD/2UmBQi0pv3NOpR2uFf6e3cAUKwkU7kB08sxeVQ/chjxX
7ruW91IJpUuYBQjZzT0N3DPscapks4r4XKsDCUMl1fEqTsD8WDn/xaRv74LSDxYl
7xmNWnZ5AUcVOQN+LjXI1xTnejMtKz+e4qmw53CPeOXmo/bwIUAKHH2NaA96AKEt
WnJmxXrkvj4b9u8LqylbQMSVoBEQxgB17Y77/P8vjtwzbCFxC2Wn4MyKtHWjRTPF
3Mri5AGfNob2XUVeRYeSnK8dFqu/Ows475748oi8zKA7pHcDU4+XZAoATxVuTMQA
VGMeUbumBMVRZ4x4eLaE0bIkr7HT6lnTLAF9oez1U4xDX44IjVs2K6EncYU7sbzP
UlD4MRGY3pcv2cME+9pthT/EtjHBLCk8NdJFwRGiPOs=
`protect END_PROTECTED
