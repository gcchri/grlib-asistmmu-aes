`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O1GSNfUv7t2CfxXYD9Av4/4Ge1IxPOi1/E2wWsTYTCxh1q0Xoooy1mLsvOCi9WhQ
/q4KaVf0aoWix2fK5tNcV6E4rwb7AtWP4yquBFxq31OIGa2BlUo2QIFj457sRZRb
/C+X5z07VhAtnBz7ojFtYqInFNj2UTsqnlwJmZOS1gO770xBxDlAnNSAhmJOALmM
v46f82izdyu79hScNJEPz1jNn12GVf1gzpfMLJuHRfrm8ssNu2eIqR7Lr4lGqecs
ML9gtsIx1zvYUZWoa4HBZ8PkyDGSKXkRr7xh9IZHFBhYYitereXw8Od6aMtsXnCo
DTv4jBY5ybLeGzelmskXHM9GGmfAI09ietmSNa2LYGNOp3iFcrF7OoYUXSj/yiIc
3pAehTV/tJryrtgXPexbqFKIIBMxAUoLlc632+TDjPV9yoxkvX+XagS+bLzxuMow
l+m6NlQEWFqwQeijcW87JRe5Z0ajqfbcy9QyfuXDJi9ogggf2Fc9oIe6HfUYQc0W
P4isrx7st2PqT31uPhriTwSrrcy4IfKJLsc2izWgRqW4ABlcYbSBxcnjqozgkiV/
69JF6TTsG6aor6c7B2b3eeAINT/BPOaL8y1K4fiID0QMi5w1/fS7ppYm1Hx40NnA
T00PvhrtTa9BZ8R64WGG8POD3h/xjnrPqnUfASRyBePI9Z1MykBEIJVebV68bEJ4
myOuo1J1U5XvwKyEUpox8kR+eAZagP8/lyIcvwGG+y8+mXWTFA6lcmIivKWFHfE6
UKnRX/P851cri75hiU+xEJbNpjAXr66BibuqD6QlYPnbT3HKZxXOoCL7BTNwSMg1
AydrKgW5YpKBnYXej1zyvqeK/80poIty5hWDjFzqTe2RR7XA/w6HsdnV/gZvjGfk
xs9cnp+rmw+SOkJfl4CHciehgZHizUrWkfRb/ihh/iRDBJMYfT7Zh6MOFpbXGF6B
2vkWCWblrrZLO2d+Ygnalc8PtFrUvHdr4zBi8TrR//gjRKbt7hiJXyo3vMJnlyLp
VT6nazIdEVC6qfFe8tToFtwTXymrzsOituiXLrTZGT7UKRquEd9S7Z2cmIOH7dwJ
2nLLlHrfyYIPbDO10TFOMhaZLxda17LrhEkiKwzTSaKFpN2tJsr3tzIxlt/SqSkv
P0AO3Cq5bN2wvxWWiB/xWH5YFjKB8I6dpyVd5bX0dQ/oyh8NNNilxaBxr6l2vLC5
y5W79LwWY9e1s+GBH4Q6mP5UUKA269njZbQ/PsNr2B1DML0oyuNJBh/Lxi190ToF
OZTY0gfDzFu8aqaTr1HoacVFl5DlUSLWNGzKEdYmOgi5Nv0C645eElJ9aHGJxUQt
wAFC8u6ZG/KBBb1W4RuAO8FGPutbxRAqRGflZxIa8nhCq3TnA7rT3YWrYdOgVxR3
2/X9cakgGoQS2FUE2V4nIz1mA3ofC2j3fd0G78FJgY4k6XtNLP6KKjX8rodIWDee
bLBxSmxjEbj4iq0rF5PyeFfOwTrr3vhaCAHL++5WaRqle/lRuTPKU85xIHHe+5sH
3XAokhiI1JKb8Wn/mwrI51eKMpuCdmvK/LnKcT4NNdioTgbHwYYClK1kQHU98Tr1
X1RPVZVwCe4wtvulvxVJdL/5ONF8n1R424znIioQ6VFiYZAB2FNgaDLwCKlc5GgC
GldGrDUsqC4FHxvLcCL5Ve1Erh7iEC3QawisRcUnJ455hMJ+UugxbuiPnjwVf6hm
cCZbgNtSqifbgoYxvcNq3kxlg3EHKmLei2olWDJ2SgSMbRFgRrvhJH5+fFof0Q5t
vtEh5EBP3GhwVDmlYqn13+YmUwG8tymJ0oy94iW1alXzyFSAHjR6SD0F+Zo+H1l9
XfX5KXAsW8umHbcLN2LMOs7ixIU7SPOKqG39mmSkBxLhjfj9j9NhUvfRpH3nJHAg
8Nlf8py/fe4Sp2KgBKnmwHpR5LxRPCTuw2tBLWNsGZf0EXswYw5UFdr5vOurY6Xz
N6HT8tYgQu/ZhSrcm6gnt5H/tGNffdXeBDGH/dGMJjl6l5t1nX0Nfe4PJnjWafoc
XN9aQ/VoMUodAydSbYNeRjeGvhNynZhlzt4bcLdz4s71QvQePE1nfK6tS4yF8BAV
uoicE6rkksWOS1Yn/FwVtlD/GYy2lvMF4HeHfyfpwl/o7gDFsUN8CvjqhTR2atSM
PBB0oXc0vxLY+XT5X9hK52a18y1TLvVz0MagP/EmUqR8fu2w0fST0Ytg9cDi0nY+
DUrIDglbcV0zZiML0Uv3my8fgeIBUSMqJYROWpoA0zQ+ZcuMWnr+ZdfnzZCXCGpl
VCM3GT1tqtjUtgF0oH6XOOzWn5dJ8NJR/YCUu9AOiTVHYLJ+nGF6Zv1liqPckWoq
ZMthjd+1H7+MbRUsjEuNUTl92fGThZnPM6KnQM1WU4sjehmrt3FbHwYXMx2P3oAI
Glj66juevjNd6821IdJNgZR8KXFiKsbh8as/hfm5ere20IdOQB9VKRtp/jLA6de5
IyeMrCeXt9vDSvwW7SjVfj4IXPJRlYisj8PjeFo0eHeDs2LZa6nI8A2aD17MJUpL
FHNCkeoDqMmuNT3rJBqM67QIltFRdunHmSdBJZ0J8VkfuVNFBziO4FHiaJz0Bn1W
gFbSD29n3x8PRaocfD43sjQbEXixZag+kYVkWrT3rREd9DpDxWbBO7lK7WAoR7KK
X3sb2rCYRz0+SEHIgfqWFHCGaTSt+YJiRlEODEwMKKEkbamXXvo0c7a4Ss4QBxin
jYlBtFeHTyPyNBvKcigSsa5vHshlijjT/3pjG7wmA18gjtptu+Md6biKTTBt3Y2O
C9MxFQijnLVa+bSYPuI4z5aCHk7+xCcwPNAgKtDhtKbKtjwwfdlYNOeVZucQYqAa
Wi0IErjcWYmpbhbDvgqc2b72t9OmgHkD45qD0COJ4yznArTQ66bBcfuuv2qdKn6E
WqQnKkLB6WIdFNiXf2tKmBXFx7k3ztCqv/MUbNIaZZPgc+3wfJnvkcNJHI+tY7S1
bpQJ05YPKMtMcXOInKqbnsP0VPgznvtj9wwUYeRm+63VZMGevjJUZzxnGfcnFxrA
UegQQpZfX/SexxpoxKMTKZmHNqjEnNtENykvhoIRcCiMJmpA8cIEYu5+NGWRAA9r
cwpLDkAZNH3oCqqklq4jsUEQ+tBGLUFizGZonM/8wsPPMkwbgHp/zyhEUthnT9lY
A4734mDMkz8uzTerZf7jvV1lFO7FhdMjArjrezFl8Y+NPwCGy8t08yd6YJHE2YBY
ox8Bpio2MjURRwHjP6nnJny3f5vweKmeX71oz9XndTJ1U3V14IMKDQzTbr4R7RMI
DMBLhP+lpU1BnCUUN2TtcTIO9NkJCrjaPl+VHSiRhL8FbMVDuWZaJHzPsOWeAcZr
a2ASdcVD9VXuoI4IloWskmDoVqyHsAcRDU6p90x5T4Y=
`protect END_PROTECTED
