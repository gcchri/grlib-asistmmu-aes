`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hiZvTgpTKUsa/ZbDZrNQTyBkPVhs1L5PfZAq4uczm/M52eF3PcA9iU/8wHIyBcXm
q5+AW9flIqeZygA/xWwNC8gxRqJWqi1j/WZ65yNQpfdfl0xMgkKN5lHfwVj7gjea
ffL04tZYF8l7ykyGdI0HAzGqSOwlR7VRzrGXU42hTF78XDTPNl6kmfH+uE7F6FGP
2wzH5O8WSxe89ciRxMYvWK/893f6CFodSrg9XKSopflgdwcCYbTUvFKwlx/K4RlL
ULjTppNOEZVCviU+/wTwh7IKvcqC1K1V8m6yjrtBgikB6L8JhxTTSUCA/emcVSDq
BK2sACmBQSV+tovzRWxKLNQV7EJs3t6utDgOtwLldGW9dvKtGmb6/VTsxq8KtO8h
`protect END_PROTECTED
