`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
boBcmVwbMblcRby41KbWnK4eRyT2Jdl5lQgSf+5LNlUhqTpYPVuMgJ3bxdY4x03G
EoHTN2PuH+zPGAUTgebD/oF9cOxxHzFJMR7tiLnjd3VV54rXoA5gHIgddeKh8jPH
LfDMdwR7WZa5c5lP2QyzcHJJKVMrKSr5xGtNc/bKiwYVDBtsqRxdXiR1nt6nhBz9
nJ4oAoRzims/uQa0GLMrwqSIwHZ5yHmr3v1Qg71WcnGvbW/LChXX0gba9CpzFnWZ
B1UqDBvOil52zLlbFvJAzqFq44ETkbnoxyI2KoQiO97aPADUR27AQaep/P/Jh0jT
rQuSPEreqcON5aB3hEX4yg==
`protect END_PROTECTED
