`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/zvAy+oUF5ChF1/K6KQa0CPpM18z9wlXVQDdvgLVfwxMq019JWP3JEIfa3aPK8+S
lSEGyTwikXVdYrYKZYZ8ZafrLGw6RYGQ3ZN+2GawIAXSljdVqRiRopaMIOxiwQuC
ki8xNmQ+nPbYVZZNtOGDw8gpju4l30rPtWtLpqaD2TYeUEKqNb4O7WFRsbwmik+7
GcEufaCt6xAgs2vrO/QqB2bT+/Hn/qnZAIGanc/EK1MGN23tPXFbcycIATJNzHb0
Hluzu544h8S+v9WeZGPOca8BK4o+5zcMHBHFSZxevjtB+QhsnepLm3CgpoIFkc8f
dMoiv+LTeBVkJtC1bWgz/XXa4nnmk7ZTpKXXu3rtjOfDzbldu1JjXF8ieEnxPRjA
MdXcNsA3l4RpHcPs8DPcusMnckQ0TSWcP0mR/XQ7K2915g/AZMmoNcy3bPtrByxw
xA+c0bFnaMC2O4D2HmUt0zxmImYczkSndLpFtUA2/Yf2Ip/QTnhee0itEhZtHdyT
`protect END_PROTECTED
