`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qFWNX/3lGasV+4P3RjJiSv2Z45VqHn3VsbmO4zvLB+g0/7l8h0DoqIo3HdYa2iR+
q0NXdRNZmY/8PWWr7k+d3mE5EzzAgNeulgxwSi+mmNg5WQ6UIMnjNdls1PiDnmJz
i7KtaWY0Kc6vfwQlfzHMgI5nFobYaSDjcayptEvnaTxS2iuq66CoKQcd5+vDyNKq
cQ/N0qTaJyflmd4uWtSsLzj7QNG3+M1Ki6AKzRcwjBaBMgW0VJnDHCv2Zs7JWIQz
QfINngcifAstUcWNme/ojFuZnydUKJzwC7ci0pKR1haa0KWroy2FLwYiJW+wEtzc
H5/cmufnRbZbz1F/RZIPgv3WQveBIvQ8y89CGwhdxsv61GQRIPogE63ZEhOhWd42
7Hxs8Gq2P+CEk1b509LzMQGMYy4YpBaZHZbA6nNqoRJiUTOAt5HzO727enMMmDl6
LUmiZhooS66GMAnwIxvW+/yzDdv77uFY2tcBatqcpWRCkHtk+vUNPidPsBtDmUG4
h6pzOaq0XB0hWjm7kDKqSvxFiKmEvFkJfJz9hOGCf9/qHf6elgIEft2d6dGTCOIU
v1rj1BiCWkch8v3dorHFkwCBkdgrbTMxu8YQom7MoeBCdnO3g7m1RphaOPK5pn9k
Wv8PcqjrCXbQbv5PRZrHNM5t6GMZI1Zhok6KuyJwTREjF53y65jtYRFZjxEMdbZF
A6ukG7W17GSnwyYqqkKww5ao/0bwAXqFw/yTPISLXBwwRxGD76TV3rtJro8hW1Cd
SB7z7oVHqdK24+N2FJtPrGHV8UGbfUzyWGfT30e5SngmD4ZdEhMhtFSZ3wip/D1j
uflUKvZQ87L4+D+6exIok6gyTFczNYl7kL1xIhg0h+BTxVBeTGhtqD13KGZOhSgV
07xomm0ow0vg1hrITnF55rvWzOkFN8bcqHmF5RmsomIj3MlxN0GxELPOqbENJkAz
`protect END_PROTECTED
