`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7D7oBJFuLNDGMGoe3fWpu8f5YCHlKorNm4S5skSNuqrDUaf9DjBzVPBOxNHjYcry
Tjj6MxSXPmm/ee1KhNlQJXCMxo7ALmFgegvHK6c5uXUwPEbq19nj/7Ir9sCa+4Tb
ibvXW3JW7ZKgXVDvYZW150SNhvLykBFEC/ljdj9ReeiYuC+O1rWjLicUbj0GCYnu
q9ltAIpn9vNqJBpZERe0GmcZBpThawfPuBbU1VSIyjRtXdhkJGZR5Eu4uTkz1NiS
ODJtITEPljACY62t874EeIMv7Ogz0fCp2DmHHXNbazeZgfMGq2yvoxXMuWtyX7Mv
jAjwc0vQgtCEYH6nAZhF58dBZOose41sNUXb4PDHpWFvSx3XMz4kt5auzxS4NFd/
1PqQuFO13FSaCFxCgO3r6inwIfYBboo2CG1fxDRXSn6usYaoC6CU/bxcGptueBLU
1yeBL8TeYozoY9bgxSyeh71DFbVIcqb6wn60OJFiD/P5JwAi3WuEy2bFh7ABwBwH
D0pilnE3oGqVdYptEh+nQMwv9ouP4cvcCcdCQhc87X83PoOIeVediNlUbXz2DcjB
zc50PzkCkjQ/gHZfF+Rzoxw7xVSJgSFnbomvTnNlPkIG3QNHIrOwuQez+OPfxevZ
uNDk0MUCZLOti77g4HVnbBb7XbuLEzxZihXgei5AKFCc26djy8AXreICgfadjPCW
tQvOzxQycgkc8QWbBNsmN7RKUimcm1qlBln7ksOA8VrxvggoYw4UuwZlPkAeJ+bY
lizPwM5n+qPcgM2qLjyUty6iSZ+LTKmokXPe8KAB0WzxXw5huGWcJhtu2YyUJL+l
TRGYOrU5daSHZ8qnphVph8kFJN5RqussXCHcEr+M3THXKPMILkMu/bgQ8xt/xC/v
ACP8Rk0la95ezbVfTURIxVd3T9Eh8Ml6QETHY3v3p261y4LDW2bz30+wmuktu2Tr
qdIsbIBF0be5zZTV+sEbjgz8DxWVDwsdrW2b++pTDSTM+3wWX1gs0kkHCA5qz32+
X5CqhBA/OGB1CwkFfqvjNTkuZiKHcOc2CP1TFHegyVKIuD/tWU6IKJwWEEudExTm
Lkth1s0lwbRRn0X/q2nTAtF6TInDDZVo23gdewygU8i5sS0Sw4DT5GIVjjW5yg3Q
sF++yXvs9KVOHn0I1f6cvNP9xwMspVmMhd245PLhREuGGwIvzoGpBil+rO88qT5n
7jkmUVb2T7fwMSd8cjKI8U9fLxtZsEEe12os7zL0g+38haAcKRYgHFpmvkL3gnUT
5OR2NksRta7TDmSjbSjunrG4xSAume0/b6AlD3z/+xK68jJZ3C2jQnbNZzy3uASX
pl2c7n2e4BNjTb+3PR85XK0FhsjXjUums6benG8zd+JEVMLonTtM+0MAyS2NyOh5
8wqPfHPjrUEU2fZgs+fCZ+v5TMoMpBCVORwuGMLLB/HYso9vIWXbmDAe80m1gOPt
mkhNMB0e/6ov5pOKeXvlp+kPLi3OaPhl82NJe2yJ4wl07PssiRrteVyuh9TIPQ4t
V+eKFxW+HV2GNLKCfwjQ9AtwdDz5BNjNcj8e01Y09y19dXSfRD4HCqlH24eUoZ/R
PzxUWRfU4HKheqcPpHOxHU3x33k8tSXvI5n0TkNuAdwffdQqKEo8b/J0nt9cHcaA
eI2sQVcf0no2WHpRWZZKYXKtmtp0thM0RWK+aYv4jxaWHM//TSUdTLYKytBbMtYP
yy+mMybeDB0SiH4mCUFgDw==
`protect END_PROTECTED
