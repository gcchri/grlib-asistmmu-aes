`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ifpGRUcy7Lzxbkr0PZ5Cg/2hS6RozpYm1cXG7ZoyIRYZNP0Zlcje9zws51Q2/En
vJDMLTZ39USZ85qrS6sfKqQuEE66JW2FgIGRE81qcJY2YX/WGCT8fO9q9lbtgZZx
rhf2zsPhyCtYrESyWuBa4Nxzrz6jE6vBfvi1DCMTS0Us7AKV1Y8UlLiYC+jFJozA
OgBSM3aNejQjglEHIlxAoFXoTVfszjD4dyOSVFuA+Veg3UZF5uPCsBUYUy1/i5+b
RQRUtamNYrGtg3Mj5jjF93HZhvpghA/aC3Ck1DtNFCzkDm/pDWwYuYhK/rAaMg/S
E5KIWIVbC9DtjUF26bDN51C0n4OVvl5rVP3rB3JQdL6Ls0yUDXkC5w2z1u3ONBkW
Odepi+SEHUaTKl2kBvLTm/zkpQXg6MFLs/DKI19UCNfSBCbK7JHYtOtqVzjaj5jS
DZ7yuQFPVkse2FIheFBCRA==
`protect END_PROTECTED
