`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E+W9WN5zaPqvvZUFSSVle/9dCr6wunrnShWNxAzAMVAkOIRMbwd5U4EkFnX7BUKU
4bu7y6f/9k2HWKtrSl7EdEHsGy5ViuvX4KHRXahrqiAUeqWl5s7a49pS4dY792jU
t2wnH+x4RryvbkBxwlkzFvDcLppIfV16zNbyeSsEI1AOaJiTS+kZRHw3Onue+QUk
BuMNnsou/hP89RqWi+XLAA7Xp2jySWEwT6LwGE6Z8XUoOiJAEdUesQGun3Dcfvu4
pDWq1F+sOWE3OS2RHMue+OSZOK4cAuuJZpNsYY6g7ibvoxW7/XxArY5Q2Q0HwNHx
hUEauy632nU8h5nZZKbtp+zxomxSW6h4ds/k4+Np2r6m4DHjzZkIz3sH0FZCpQaa
5f/XWK0sXDV2/tWseb6YvU2tRbLk14Hye3Y8JOzwV00ZzvZ20/mqFfPEC2V2OblZ
dUzBBTPqau4Sla+y7a5LmqgdHZuZwXAxae0DfgxHPfO9QfgNv0OKoye7VpUXnmWZ
wfMk9HbIzvOA+biLYmXCitq7suuTcurvcdYPGzEKyJcmRkO940Zq97E9685psbd9
cBrOUoK2Rya03v2CflGisihQAkZoEC3YJ4a2Sd5B7qScY4urZJCPKzse2jXHTQ9V
mNxS5W58KGl5yalnZmoL5XY5FLBB1+/quJPIYB0aasBISVoiRBSmw0O7uQEO4XAJ
6DhcHLJZmTiZFviEdGF650ua+Y82ZuMvB78My7EMTz4kLp/tjN0uC2Q8TvWC8t+m
yM0f4MJPYw+oED7ae35WKTx6IxAgHCNVAsr0a9jWn+GGrBA4rWr6iUpN5AIDDM6W
Qadre8X7urooQIblJHwUZ2OYpeMC8jjXaGV7ZzzDbmTbnYAssLiA8bRlfdbwy185
R4xymhECpWBwHpq75Nw9NAhU7yFDUtSqLcyLKKxLDk8QCWWibTeWiaHY5uhvw0Un
eyaJnqr9ZzFxxl0IY8DOZVky+4KV6WXYyMNunBmTtOQC8Ox6kuPLLtx3bZRhNAmR
jcuvHsbMfHF7PgblqcR8m9eawvRH6W5t5R39mNWU7rdCf11U1/VnMJF3ozTUqD9A
/8BalpwFRRIkhVDAfzoiaTOGW4FHED9noWDBW2BBZMax3JO2T99+QEsYqH7kTnXf
uNFcTQbS2FQN6mWragD/2ZIrIJ1qYLC0NJGc8DHDgyIHTOF3JVk0U5ckDnB5TecJ
n5A0nAo2MmNPwI5wBV0oUyEb4/VO34mPo1u4GbQ6eADaiwqA+gjyeU07X7+mmgkY
iWx1kuut3gU/OtnJpnnEQllRJwQFa1Voq2e5komJ5VyWQ4wvRmXinuELwvTPmo9W
OmmGxuecffPJ98LF0wji6Bj0/l2OfZRJA2bHZentbUArENOLt3UQVNdK8GntDrJA
u+nAHnrv1z5DJN+IRegenA/fj4IdSzbdCjmfzbPdjA+MdMWxG9lCC7RpoQVh2bEV
CXaHQsmIRfyZefLQpTHz3eU9pnTH+GfcwvLsNLxAZXBfdABshiEJrFOpWoe8Wufe
+OKw4LFf34x10tdL/ibCh753teuLS5D+D18GtKyYbz+cXUIBbrQ6n5D0YkNUSPsG
8AGc1Ngjxh8gDBC8clOtrZ+o2r+bHXMIXPYiY48fLbFsByiO9DZKAsLPbFNApUOc
ECRlycaKkxXpbs82lUhsVsandtR+DtQIUWmFhOTB/dAjQ+Q90wEnLvDPFwaB6+BG
+ss9aESYqhZIEUwiBFRcFRQ9RLWJzby/1MsZ3IMsbFkmE0UIgDGyYyFAAPETXMew
O1AbUNsuZj22/dmi3IQt65ZtIipnYvCjyKQktGjB689IUCAcDDZ3nCcmHgtM9mhj
fZyr+fKwAz1GNVR4qmgTh4dmNndG4Yi2ln+DlkcgMSZrhi5JW0cohTyFWEVhps83
z2eCQsmTcyXqhM7+jrXkqtIhJtrokbJd07SCIFzQ+CyJXqc8YlBZ9SjB0q2LHfSF
SbTalL37Vr/See3mq1EVu5eGJNWcW5JFNlP9ZClaHa5u5/Vx5wYRTiBgqp2dKr1m
ZfZzcjikMltJ+w172wPef24vnLcgJ5HjVBm/cwLS3YzeQA3xCSUQH9uVEMsOEt58
kEcv/8UiyPy76lCryS96XyIumFeQOWc0jva4bPDkwu9sR3I9pp40WBqIjRMOfvdh
14/sva7X54HuVN4uwuFCQE+sYJ/lgMsHmyfS6O3qIhvTc49qUjrvZTJtXD7/krXD
9OSaeeAsBPe7G/KhPdL5NPEPsK0/ZcO/R7WfE/3mGVYZt/Kn+GUJFfB87Dv8ZYmT
TYCGIfWGVAZCl6Xil7LjGkQVMHNFkj2cqpLFkvkhIxU=
`protect END_PROTECTED
