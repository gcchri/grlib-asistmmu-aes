`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V5jeLv6hW8Dgpt7jCWWi4ux/UD3NJdv6KAnNzXhiMWkiij00F0vJaAxDIoQwn2hb
pkHg1p5eZHGtshdrso0QRG0+avgMtvFNiqDfxwxQWpgw9uDGigj5+eaW3GKluDzr
ZVUmakWaWG7/2sAH8FGfaREer6YzWXvofpPKUEzwHAMzqM5xhjMn/0c+qwFcsNJI
JlTX2hZIlMJyzaPCPMxOIxqParKuAAwQh6hXiutAavCWEdkauZd9YBOuigmHCxx4
5tzxL2ffWoBB82oIwcCjK3wx271JuZw8BM4kZr7OCpQwgIdavCgOsj0/ZpyWRxuZ
iAY8LHV0pzvGp5YaJ3Ha12HMT+EkiFhQZw+H8D0huSe4GCeFzWC10cuiVePyDxhH
USJmagz+uOrPRTuVMVgnMQOUhLTs3aHakRHfO7wPu9g=
`protect END_PROTECTED
