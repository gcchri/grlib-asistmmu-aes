`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PkvtHfpIKUhFtQP5zwQNwi75mYjjLzTCY0kcCxKXp2Lw8irGFuC1TsnueHm6rUgY
4RGaQGROQJcbE1E7RpwaIzle5jrHlXexedrxD4eAl+EpyyJi67KyNaQ/d7s9IuPA
6kX6Col7UmZGSjOFEkPJYlb6EmkHXX3XfejXbxrGvWcPfrn3leWUGBHSxM68XAHy
jVGCsVfr9tQivEY6okz4qEk+TOxo3udVIEb97JAR3zAGynLzD2Yl6BHtdt5mWMnx
KNgFACF9RcMjKSrWpLbfKfjZX2zWAoppSphq2JkbC0uOQID3YGZrD6UUVXqr7KAt
8ji41RYMXYiejY3JWdfWDboCo74gZ3dtK/TIRE/UFvAAAMplYuE0+Jqsbmh3vCQH
C/dURmzcIg/q7Amawv/O0pU7l8swuzfHJT27omQRP0QcagITDTern8hwtjHP/mvY
SS2i6IQuCHI4DVkp6Humjg==
`protect END_PROTECTED
