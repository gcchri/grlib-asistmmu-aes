`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8iUQq1a8ClqGd5RhCtpTn5l3d4Zo0YTYHJ8JkBbJEl+LoCxeK42tLT6rV6ZUGVcB
V0/Agk1gNmtuXZEERhnvzKgI42ypag4/FCW7p8+tOrs2QpjTpSivSj/YQHiS7Hm+
0KVNv8VA7o554qJll4SfUfCiAWlUpSrFgksZVmzFizJHZCuu+EyjIz53grKtNO8e
Wd0R+oJSHKE2galmsXntnIvS5dZWvVIoGkqio94/fxo119N9OxZMAGpqUPJmhhxP
TnYuOCBh6sjB+iMfuIGFkRh33l1RCg2ejvynjjlQTqa5IuCyxa/Q2tEjEmL+VeuJ
Tp//mtXHOs+jM+gZiYmueqZGlVi3wOuq5T6qLu9gYaslDbOREA/XeZi0gcpeAMKZ
2zA0UOaXp1duLEO1YEjShuFezFD0wchfoWcQD+7ReliOmX/5gkvz/FAXZkeSqKKi
cGAyhefCTZS73e+Dm3tJ2Iu7L8XJNRHP+XK5JhESh0AKbGvDraqicOjflzQd04D1
CapVRxXZqCW5SvS0sscVMWTl4YFvSTndFula2OKNUQmUl9zSO+5PqHdPqlP3bCXS
eWGlvjw8YZGdzHnxu0C8BMvUeLpNDR+S3Y8j1HXrfI9ZLTisowCZ4QFVCnm9JPRE
8unKNY6FVc3sstinOCYoM81d4WX8VtVambupy0ztJ6ZXZAvVbY2JmiZPwA8UfwHp
qU/N1V+sQZGEtJb37gv4D+aiCzlRESNXOE4cLOM14/4Ex1CNfVBIjy86krXRj+Lm
0as5pp4wD+DEF8xk163KOakRLQ9xYYM94s11ntXuOEbGHlknbBUnrQH1UdWysiGA
6U4laJp4QVOwJ/SDHXJ9h/A8g4AqsBjwJBDvZolcPyrO/t+SIlzYTakzVy98n67y
swBW4hW8Y0vNWUcZVwB9Js9x7P2uRCc4+3shTxR42Cwli+PcsToYzyDXZmn0pStX
08dJmeiDR+zRs6WLYgA+zL1SzQVYMmhz1FOfJ7XSdubAzDG/QAtcDDk0lwVhu67d
NnlJlVx2xTWIth/oZZhVofnnlKoqeN115nKSnjBK1sBA41wRhXIuzUxtNXJjnuUX
Fm0ebMy/0yIDAr9L6J7oFqKGNnIxXHz4j+QF18gpWQA=
`protect END_PROTECTED
