`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/0XVRVo4kGXfQNRFdPG1AFDw0czmtuSejK200Yu5igpHLRVwIIZ+g2tdyuOQxC57
oP70yaklkRimopedIqURS8DADmZUMbyMePX0LJX1iWwNN9T3Hx3lvR3R0wROBHko
AkWf1bqbtE7Eh1tSDtVXbwUKNpTGK2uiLxzTPO32A/zOoQ6+G7tOj2HTE7T8KN9j
Fq/KY08U4XXSndqsKkYBveR0/nd6gtx1fanjVv5K2Ro2gkIWf35zR8CeR4JHUNLd
yXYgcEZCHWSdAqxdtqZH6m3IocU6vHge6w4UsPFsisS9VgvGPvhH8RJlY7NAjrUX
HMVBL4pVbVSC+llHItfd8P8AaCgn4xSOTh+tAk5v6qE93oo8frGntQEI0tzK/1E3
uCIKJWoSad3/gRt7UiC5/r0r+I9YMBLVPdYfehfvcw2ejng0pJJS2i5QDCC+ZOHV
CwdY4AbLeU59lwOR2EX1veJZK21tpGpVnPC3ADzlCMZnwv1E5ZdegN7o/iAt4qwj
RNbAYLltKPiQ7K3zrJsPjNZbhT0eBqRAQSOx9YoOjYmZhltxyQ0FrDsd4INg0CZS
iyEX+9UM+4L+R8MERBmK5/ciptRjXF7qq2uEtpie5X3LeS07VJyFCj/IDT04fvCH
ZA5PUsUQhEda7RXsGo1dwJGRMKFrUN6DFweZ8nCDdQUbWgyHtPQudH5hDhZXjG/h
3v0EHVoAePvRX3BvLAmS0uyhYCpOVONV4cY06yns1PkhSASDidk7wkx0NzXscakC
yml5nj1TGJP0BSKe2RJPMMmnMi84RsGPrqkbe8ddwR8qyfk5l8PAhz0WSlaWmcz+
Nq+MGjBQPj4FE9iLcmQMhJLljWYw1aDNhoT8KY9gmHydEv3OqGPVkAsmakLxZAVM
FkquO5IjN6DROZcwnO2uGxwloQITvRSOA+k5Sqzj0Z2X9N1IyqST1xH5Z+6BDAuw
o9/5CZ+ns2Fo/eBqRbsHHw==
`protect END_PROTECTED
