`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0QKHcvqH6iHAQQxfLgsP+htvEpw7jPvYGc3Ul4nnsg14A8hseaeR0BcIZ/7zwA2R
e4zxRoreiijdSGwyuXYR/DRYys1/9uvw8y7j5kHO656A+5G9b4ARNYrPw+Fpx8ty
3xVSc2lXA7wzr9LkmLZ5lmdua0uX17fAJM0337SE8xQBNiMnX+HEtxBXGrudRIU+
GWOVbJ8bEKy7gKw1qus9HitPkC253l223+k+95XPy/GYhzUEDuRjU1IT3m7EMLDR
wKQXQBAO2DkmtO71tQy2jmlnH3uzGbgaVkJMtpGE+d6nsPIPpZtxm5K9/642gXik
rfQyZTucuQsyJmxtd2TnyyXVoH/q3VcxA+XuS5iP2QSXsweNYPlUYYVT2270EKNt
5+TCzt8ZK2kJxP4jqRKBDZqQuefb710W7IcksTvFESI42+BNvkQOSgzBAU7e/HR6
c56ZNUC4RV1kO0qFU1a7xsDTfeLgvmXrHxTle6rMQMmPFEa7Av/Yafdie5ERAzUv
3ad00N+QBc9qsMg9DFlt3bPvUd0O4mfcYXMKgYgniiXHN7sqnF2zekLUx7pPFy1F
cde7Gh3gWjxJTXENevzjCCxz9ASheqznOt7STUK1j8lmZlnJNgAM0jbeLWJinLgD
yewsEsu+BMIL7zl2jk7MqA==
`protect END_PROTECTED
