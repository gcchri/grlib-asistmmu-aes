`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JI9ETen6g+0bKS5uaCsSJEwWTttp36qf/fRyROtBA7XHRYJSMqfNXptxZ8EbLrtF
xmGSyBDjiXsajLKKfKO1+sgonEMPYGScaJvRTovhimc6rw+sQAmGIqSF6yMckDLI
sSkBsoJdjEU+e5djYNDHRyHlQaypme9vVJlYggmZ10elIaZ7FJgbSD4lq4NG3dj1
8qn/AW4d7ZcXZczBPzc9+J1t6MYbK9BSpoESSaScyfiHEAizmB7iPVlrnCsXxe+5
2fxY9WgejyHYyN0DrYodAg==
`protect END_PROTECTED
