`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bk7dmrP8WWMRzRyf2zfnbyssrFpdTbAj1h8IKNr1zLV4b2D6eZ9P1kU3H3rkp2h2
ZhTgC3fjuHFllJg25Q27HxzUWPFaRt7USH89yyEL5gSRdNS8zzUmsIk1ZGkuAZ6x
pAd9SSx/SJgv0nniFhEPxxSJI5OykjV+pN4TVdLnFvdaUEK0AoW/NNuPGsTeZZJg
EH8GXu9IuwUQZM0zKNMlF9msxV8P7AaeTuqKzt8QMFI7qB01JBAXxMskMe2nzL5p
WvyUxYpOJHEVWpjRS5ztJLNGA/W7kjiuVTTmJ8YvFZ+ymqZQRSrLZK9qCgUdho/P
BfuKIgGWYe1WMO1ArP0spOuF/0/3Upev42MMojO7KMUMIpuW9643caysMkzW85O2
DcXBzvs+/rye9TJ/X6V8LzX8YmUYbI1J9Cowzzn/ZKLs0ZgZ1YLzf/HoRsgWhqAP
mAm/ur1rZt8Hwk8eZVbuu75nR3Ryao8/CUQy/DivvGQ+EkIn3Jj3yHeLNx3m4ny6
0Mkkb19HdMFFKw5xRwSoHcmAu6Sss62h1O+NUFGkLiPsxuoy7Y0Fr7g7+0NJ/40K
iGrOFSbrWPXJ0Bvm1y0XbKv3LzUV3u4P0hesQDii2/gwFtjY74q5GuxxStF6W4JA
geVKt0/N/4RADIlCG43Vqffnwd4pfAU9FGqvHq4/H2hIsEtzEqbpBsx8hkWxDWwG
13dbB5gnFb8M2NaowGfvpMcT4ZWB2BntJfyZOEboqqsxen0yhwZGNCzxyeQjQXpo
NRd3zhteSoMyp5Cz0DW6M18TzU8pXaNebXcXwBKKbkIzvihX72HdQ62XU1DIeEn5
n5mDOEmAyheWyD304r6VKAJzsgwTEkFyeKHJerjuou5OB+IOV836A+fTaqmF7G4C
/w1kavw3z4gel+nujkaKiHQxO8h2GDddxFZ3xNf+0GCdYlmUu900IN+Vu3Filz4M
cVhbwwTelGuWdN4KAh5MVyTMk5shOZN+ouxdbR8IdoBZ7v+TbzUciC+pJwakd2tz
wbB08LBszrdWfKc3ZvWJ9qprFd9OatMBfcK2IkYhgpb5j4eDW4MBQR4jo/51Yj1E
4Y9zjTVZa/LtGBlg4v0hLJsfK59puJ+3pOCCvaSttIM=
`protect END_PROTECTED
