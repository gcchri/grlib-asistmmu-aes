`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AdyETIObRFVdlMJzXKDPfWd8TFmL8RHMB+nKcX6fTfMOm8Cy3SqQ0vnwO5kEI5+e
9tq2D71nw+jWJxM1CQ43iJC/orCqStn3h5IjEQQWdcuAYbOz3Z78GElZEDOsFQgf
l5RvJW2ReX4Mb2r6kJ/dzLS3V7lkUnWrWDMAzedVQB8/ImDOG0RxTVVrIyUw4iCQ
gj2xH0gKgxrEhAZSm2oRKGbfw5qV4cWrk3wgY2Jc4dm6U95u8K8Aul1jJOiAiLYQ
F25pmMNvNgA2YO496IhCMP1UtWCwVawT2GwyE37a9BWov3iIK/7UryNFL3qTbesX
Vui6ibEsaAMm0705OayZW9rOokmX/ifv99PtkfbmdrPCM8YssXHUjuO0dKmLFyZ1
TpiNVDugsiD3VMiB/8T2E9ZLqdlmvMymzhAKiGHfkQ94od886+4efsXO2b8j5UBq
4EQIBp8kpsl/3r/dVeB+NI1EPRlAopiRqOQkcQJdvXAxKykMLuB29q9WyIBd7GSa
4zcijk8lx1O/wpHN7FNRJiUIM9VtLD/+h6U+SRpnwq/psDsz8fUrdT25Aiu9s1yj
13KN1VBEloGe0RtXPonaYv7vGSD2UMiNT7gSTzd2hTT0dZJdnCSRyRP1iLCR6CvL
C0XUe8F1OAfhknfD3ao9Bpo1yJj4h/tYoFGKSdLx3IzpxEAKM6e9GpKMBskMYGel
oicV5jReHnbG6XhXdGM+ED2H9e5KXTR3KB6l+eCRZxNVxjalSYOKxbIa8udTEjTF
is6nv7QDJcSR/2CVQg34o+6yd/g/XTC9oTguor+BZPBzbHYRKWE1WJKLjRUuL1cz
eSRPbC1lZlepYghwZAU4oKIxMm5Zf5M1lYxgWgpuPS2qK7LMlTMlPj92jtNDlYDp
Hqorz3rdK0GkF6ZjmMAmbi78LUf9p0dt6nJrrrVqTMFEtWwzTiNkIPMKiSXBQ1+Y
WIEr8rdnobjGqiG0/EBHhWEMuRf/w7COmhcBzty5Sjkda8hp7E/fGH7MtRNiS73T
Ob1gnyZHv41uaT6pW12HF+aEFQs0ir8C+Sz6qwKPg/STH8glsjo8waCcR+yzm83m
bMjThfa3CjFtSdOD1Ci2kczdwAdYSbGfTMdOO4mQPeHFhT3p4JdP6X56JXT2h46E
p2Y4hFUgCB3E5fAO3FEI+SHiKYMN4rAC5iBgmECKWlcwISaqTfjOrUK2+3DpBkqq
7+FlBKLlSKxf75W/d0koo0DEYRnpLLIrFUigGB8GpNtnHxK44SFGR4aU7yym8oAr
`protect END_PROTECTED
