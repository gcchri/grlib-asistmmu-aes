`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TsHHmy2bx6By8U9oOLmbS952plx0aTvRFAIzfbYOPQJfAzlQdu77TVn1UUwdEHlJ
kzV+T6qQ7uCi0ZgHaiM6yxIXpnMjQ+Un/+pKnDioASMEe8COgIWgRV2EjyfZAVnj
DGsP15tmD0l9/MAxAFwwnvXH1JhkxJY5JTRUBtgiGmQFgu94zS1ifmrpxfHVEKSj
Kg4oRccPUDgSERlY5DDsBiXSIRgtCAlnx7MeP7Ee9n42ZEZHAO7DLtpwdN32Edqy
4+39UQBkKljRVlaUAFqaXiGKCYTjsV8LvNF0xTHn9WsirzM2gJid69Ay4LRkZN9l
OkVOtiu6/3MZ640So7iopQjKa79FWok2va13Ji1GPwMcF7Y7bhwE9xD7e5BijxFf
RIwTnWureJpk3i5G61PUGSYYKKkkGq3OXV9atk4E6+iOFjnT2zORa7W5Hr40E2oY
mmWY1XcP8+hGQBHQkdV4AiPc0Ek9ylhR8pKCByQNHOWc0ZkNu8oPDZ4uV/vGC1QN
1ztVWZr/tkZWwqpobSu4a4u12p1LgZCMTlklKJUJlBei2JqlVRNos7SLhIlK4pq4
v74hObagnHLqfcMx50o0QsevHIacaTPWugdZCr2om4K94LuUJG9RCyv7uSOFRvHL
wKOYTGqpT5xdrigWuuMthSYQtWjuHUtkr8MwwqeUJ/TtWtsidEbT2jJkBF787xfh
rd/LHkdcNmdKMnfNmRr3UbZET7MlZTxuCqzzFlgFB8SscllsxgkIXCN0eqRv9hhs
oUzIwDFSO1HWxdJO7w3gf2MHxU9kPjfPAQv6bscfYTwvicWG3et+4HVHrIixBW25
t8H0TABmS6vyhbVP3UayWlBrGaj9KRxbtqojEDgfDHvy4Jp6y7srLHQDgZVsLdLn
TNwdapW9wf0mts2YWJrV5MlVel53Ioj/hkxaTzQQbda793hbXIdSZIiJ+ifh+eXA
Br9MgTQvBIdrc2JrnKqTjEAfg7FsI/90+ZfA8zV/UVXe5PYaEis4tBAD1stVrsi0
nr6gXPeRo2lnDSjX7N8nRIWUMdTaoQbJs/DcQDnFUXKPwqryO6XLoUFOJ2q4NGGQ
Z2gmQ6cKYcL3iaE8BmGXW7q8dGAAql9olgWVdNYLXnGpEQffqhsveQhZVJZtMUbE
hk2GTOCr69YpL2BfBOnqwaTs0PW3EQWNnPc2jCOfM7RedPm9xb+UHYyHMAIGLVDD
Ve673ghjcdIt4dGhuLcRxJoT3+tNDOyhz5X1mBh6VbnITLcWJiJNwkwang7tCW9V
Is90trcyhX4c9Hpi9KmNqr9TUzEgZceVeY5rC+Tz7HAOu01B5I71I5VkcTi74+BH
hX4wmFmJ187HBmh8v0Cg48keGrroWiH0qLJU2XzoW3/NNPjBweCGtRfemnI1T+fm
eqSjJVAs811Ro3OhocRUhm3PPuhwGP8iG3VmaAzWa93JagCg7gsKdE9giFxUd5Xj
UuSJ52llvzMBSVPthDCme1TSeO0hwdYi6BORL2U+0N5BoTahOxNIVcqB81lQpBhC
NUumSA2gMmeKEZTDsAMcg7tiYoTDg7ufUfZ0/j7Sfrr0NiqFchrccrm39TZczatZ
4LBxJ0cN0EzlVSpLwN9PBppSsF4F334pyQuoIMD21MbTqqKDOjU7ZM7H7fLXVzta
MHhvYuziYr+0OV4SEq3B4W9WJqjlsNzts0rZDIFDaQpe3islo/itPgaHohoR4ShG
gIwLa6egcrCninoPD0rxQZZSrZvG25M7RY67RGQgcioyxoVjzAKkEBOYgyrv0Ydu
eigPxV7ioCtzN/9UyF44tkJZutD/lzKHuUnSLVxVCIwLRb4MYIlB5R5umoy2hX4g
f+YFyh7W2C4nNlrOb2sSt54YQjjRxlCYT2sPhpnuoznXz+fTr162yoz7AJAIqYzu
4afyVsRHNzonLiov8sw8HzolrI7R1auGxum5NOGBDQRfMwB5ZdH6nT73ZIMWLipf
VWVfdtw4I9p0kkVbZSnlaoBX8w91aPhBa/npWovElfSxKP7DziJF917CiDpAcq9o
7AugLMehA8GgT1hl1eMK6wJNR4Gz1ClyQPGqEcb/vUUycfIYZtjL8zgRNODpUEG/
z4fZ4FUzomTuL5RM9eXyyWVdm5vRQzfGHQBID+eRUJr16eDPXRtgfJBaK6ti6uXl
WXogl5yC8rRY7Y0NfS+Wm+RYMeCuq5O07/hK19XSS0YqUP6SW7/tKotMuYNTOIWF
iRiY6cA65gLY/FWKEW5UnrXt37RrMsDM/qa8lGE7BifB1dcPonJgWQJq3GJ40SMQ
D/ufVET8tH4+dG0firRHEG4OolpgJCU5KO+atHLfonY+qICWCF8lLWl2PtBQz/0m
VF7Z7cNX+7VoWWKBXXmwLfjzjCWd/1MXxgOVogibDNmoKdNYVeONn6/l8cgIcWGt
YM40epU1od0OyBmaRTi/ffisz84Ix0ZHt4w4Z7R5nG3jYq5znmOwEkwexv9spubZ
zn7xMyhh+LfJR7AGPKUwXQ4TVzJkQNLCzZOi4o6tLmnJwmEOY94w961a9B/8vADR
3zLRg5Kg/XEC0VZyjrkL6EZRp1Nfp5UwgBf4uDaxOGbcOnV29jIbsCshPtZAWvec
FBJ59Qw26Oc2HvvFIj51Du5XAdV6m2vSrZ0iySsf2MWEyNaFTWMAcP1k0ozyWcG+
/PpwOgoILI0YmojbN+plH4qTIR5+VKih+w2IRAcbVtNbDlhTRoKbD/MET0NJhyzE
dl+zMW9TpuDkYtN69W908x38EGXBSb+PJcNJ3Nz6e6qm/yyahI7osPONWbKt2lej
7FVqNcLrDdenp4IWrMd91qxz6WyxlUZQ4FlOcAlMDufoQu0d6GegW+byI4iZAxXX
DqQF5NHRY60l4uQMWktu5zWk5nz00CqhkIJTm/aSoqlAZnohUHRHvdIZ1ExpjvnW
T7yzzUB8RCrCQ+E9GT5Wrn3D9t+MLvA6BbdTmkF3h9AvrZCiw2YnuPaVnkh+850k
cT4po2YzmrYfosTPSO2gyDIo/qCU3c/XJyO8DsySdRbqlm9GEjBYZYnl+oPTKPH8
0sSa2vBS7V0nhCJhJiTe4DiAbTsS8mAsac2LUnvBeNHincd3WEWjJCSLiKPeWp3k
tH2oBAFFJclOUIuP2r8DrZbzIEqrHs+Y8rNVXEheIHWDbMcVnXPPqtMx0LpUKzt1
lqp7i2KB1XN6uBAfc3ROmVNtHEF4odk0KMArPpfTxH4+Kfkm5kbUcEUPD9jLQToe
RH2FJ9MS+/SsjT4zDYETQxO0UReLts5Me8VHwamVad9iNYlzF26FkIqeMO1HgrO+
TbHkhPRMf+Ugc3oEkUtjhohQIHMQKgp2L887STiRSA9F1wAO8nfp79CXX4rAPQf3
/uJo4BPs8t4i4H/6huoC2ib2grC6UUkiYV/JWEoMVi8iVGej1TjqXQYHrxt6hc/I
m1LapjPbqEhkVlVog+sCXxydAZHHOvNhlj1mp29vDd1UPj1/M0gppfZM/c2yD6QQ
TRGfwa9P58ukwzQhgFq7S2LmIcN3ZSrdpa5/mRKhvMHP2JG1ajRz3SS0tj6CZVrx
rr+Ps1uAsf4fm9uDztS/PSu8Q7OOLq5xNO5r194/cW1EL0laMQWTre6IPw+N2UxR
+jvnfdirbNu/fsX0Nz2s7yMQlnvJKmPazis7L56EIjzg6EY3+ziqi7wF6XlT47T7
RM1UnpXbi1bV3UoypLMXtt9KCkmcPNqqfEOszNdfJm6R5SulYIf2sST/ds77X6Ku
IW/v5xUTNONAIxAfn5ec0fXRnsUg5a13MDwiDrW/76XBRk5sa4xWqTuS8eJ3XTrB
7aEjOLwEyLg3bj8zYlLlbfErB/RiYYhaD78bVZVuyEtTYu3IarnoTbnUwQQ4Ae9p
Tx+A1zJCrOlxvY3QIoZBrxj0tqLsrDfgcygRMua/6aYx/omyea5vzIEcVJvC9vBP
1og3R6pUMGL666kvv8RmaQnh0DG4byOsDyU+VdAE9FnfFNvwOBQd+OC0FHO6lHLS
ERVKxJpU2DKl1nF5IGx+ND/oa+4q6u/RiLzy3ZEo4DZhSw4w66XAtMOsy88E4ASB
1kwOUC1fG0EhsI8MnMUxrzbEfuP0QH191BT7lKV/nQQI/k7KKv/KM33FJLq0RVZT
wlfoDMTqWRhk9fIomBpo79rOpEZa3dPXz64jlDnqSZUKAAupZndpUNcANa2/m36I
o0WMKw2SQuAFNdSqeCdVMokUuzyNWhB9BGJi7UhR3kyiWR2++NPpd/XRSuNluPW3
FDXV37h32Vgp3+0SSXG9fGiF2oL6dU0zgnbJdAstVGiUw824EYzapUIyk8dSEEn2
ZQIOwxTRXFtz9Ze8OcRqXsMVlv/MzXOlv64ey3LdWE+aavvXmrXykQCskKO7YP2S
m1y6pDevc535P5xdExkshH7ek9cGQmSODiEhO3wp7lLnC+fW+CBf57KOhoLw7S73
yW1tbMedB3iVkm3TTZP+YDgw6av7kO/tNLUiIiCHTT1SBO+ZNJvf85MEnvJFqGKD
uBbWrs1J9fvZJFfxphzUjQX0hSZTTTfRRw5rjqAnW4WS2zO26kENlVJX5fqxO85e
e0EY0Ca2sKVuAH9kMKOX2Dz6HE5owrXG89qeYrxL5RnYK6zpEsdyoNKJTK7azbwt
eNZQHN6pwymq3Q7IEwp7GbEu4ZpiNog1/Uj1wgFYdCsoBZzP6t3OtQIep3EAGstB
VOkkpkKby7ydT042RNpVCpojh9xw+JIa7twQvYuJcPuDXHd+Gh6fgjIJTVu0pkbD
Y1ha+bTcUFEv8IlnV3MuAbKyxvw2EV/3jIAeaJ82swP6pYEM+taCba+De1agTflQ
YWEtKsZVcYbo/E4K7uILlYgrfQl1c/WalZMsOrUGGjHoWzqUZDEbmKhFWb1v1cxi
fbAMDRl+8NG5Ov9nNukPkUf37NJkTcuPAv+EYgLznZ5SY6Us68W7MFV5qRHerSLF
GAs4zQso8qZ5Cto8z+0bsTe+IXIexecmpz+/Qw7UndoerfWapSicCFzGKaFbI9Ra
PmHDNC6C2nDqDWTNLwvmnTFj5aQpjTfIRvmI0uufOkyPDQLcNDhwwwdNwdsBRQK9
zTqg/iSI5PHkpB+XuXk2lIo3FMrN68Z0NdF/1eAY2R94LoQYspPFtyofyO+ai6Ov
j+SxuZllNG8v71s3vWmAur5VWA5zm9pdpjHlZ/RfUjRPZcAFms+6Smy7EXWmim8L
4G7pmiQqMuC2kLTSyMK2vXcF6C7VAeqYKdqeE/bL3E2qnIA0gqmTpq0YluppoHLl
34Z5SYB0Ly3v6j8ys0N7IDdhXL+PdpwAvwjpkQwBlWH7S2X+GHjQ37eyMeUWmMr5
SCjznqtyxv2yzwAUc9qBFDSKrGnfj7nKU4Y/T14t+987jxv5FqJtEdqIZ4YOTp3k
IRIyaAMG2C647A/tUWOxSojuTjvDg3czpvZPXnlkemT4LzEHTv5RuaAwBxIvqLIj
zpsP0nwdlIsz/uMyhTDm5QIKLggseQXsNAeRlmPGVc9d/C2lHxv9En5tDvDT3K0r
42kU4iQ+7FatOiPMPRrugB57VP2Tx49ztvoxypr3O/4fekexPiFZBvIP82n6LWrG
RadAIXrBp20o2mZNIDMIakKMr16BqZmgvLC27H+R56NxdZs85ra7qhevYr2o7mmj
zzuE0Gj4JWWl70i4DFPvepSmwm3/l+dHWD7A5qtHvKIUr33vMlaUDcixxLDrTc3V
g0wb0glzqC7ROffsadLAt6vQQ1QhO0XvlrUZFLK0SfFkHdRdmNl+Vrr8p29Epc/G
kqpqk7O1nB4PjMUSUmfmcFIBnrn7MiqlaF3sKMGrHLY79BFgY+eMRFeddLiaztEU
q3rVPfquOhWeHe5w8XZjGhjH9V48AQWl+KlTWwPPB3voZs+12QfKMEUTbfn+LDkY
+MJPbOXWaLx3NVqoRRlkS0eOD7XsMWFnw6e97R3lJE9PsnmsnL0YxDP6sxYDBK6j
v2oCaFtIUL9UXLjo5XDjucRb7KhNmXaq8lkWIhxDG+7kVPvcD2qg1g0eXyJRIaQi
d/5rsbQfixY0+rxRdEEX9MHHYlYACyH03I6jnuqPvndNXBY7K5qYf+KRKgQAcKlO
oIt2F/YaMR92KPJMQkgqbjaqABwy1GZpVuP3iC1zjqEzfp7wbabDsqCImcBjAGiP
FiaeW5C064XwPMGdAHOg/ZVgGUTZ0f8QjOqJ0gw0UAAKiC8wfK2zet+MgLD8aXek
jNGzu1FUvbKid+nfWczGayQv8f5xBxInvkotrRL83ghs+JV/HdnVZ5wdxp4QUUbl
mUwGJry0ikntqYWYN9A3AFA3Gtkng13EpCKKYVPLJ3pwQAM4+HOmtczbgSSm2/0z
2aSTHMVVWh/WKw3zLFUVZP78N+OPxvLoRf4RmTMW9CeB0hlIgnk+69GSX+esrw0E
/C2qZNZHc7XDV+68sm1q+MxeWsqnTt0+pidGyOmnBLgwmCCO9cVOjOBqA+UniR+a
N5YSf4Pw1zIzqlqzZfyUvDNA3OtVVie94r4AEtGTFEoG16Mo3wnblOK7Z+l1Tvzt
4Xjvn1d/oRsc8pW+GOO4XDDfdThGCwgIdCPK8862MasYr/MSzc+HxWGFjUN95gF9
xm80u8B3S3LjX43InPnPrHaczrilITBDtnQrF2+tVGuswOCqbTtj3w/i5zGuWMER
R2lB5uLDn8GyVUb6SY1IjRVwnsW/jozlCD9lkKAnHJ1rHs/H9Lg23t3vh5EPFeKE
WOgn167e44MuOOJOmCUiuVWU06Y9QHKyi6f7PA9sAkr7vwSnX0bQARNQ4MJ408ic
M0QLkr4DG3nIvJel9eIuw+qo540xAD1Xuj/N/H1Z1vRFDSQXV3km0l29bxTVz2Tr
h+lZbRwXUtwt3hniO5fNaxOe+83j3MBJ56gDgjLrU10YKeC5KxhgyPaZo2OLlNiK
Kx/l5B/JX+xNfh2A/cqFefVrZ2VGP/xt3gDMQag1WK6Vwt0xFJxCi78Cq03aWYgp
oVVsLA530Y1JwX6kVfKMd9Xp1th7bunAZ4oMJsrCFTWujIws1ceJ/LCsCOnkjdTx
CuY1dE4ws+Qo2OIcPufoZjkS7sbq9rlry37yQ80J1t3MrS8e2fabt9fuVAyRwlFM
wdyY3XCdadFYwsmJwJ9wXf4Njv5Lf8JCaEk6P+VQF0A+yR584ZUVI6648dDKNWha
xiDK2q9mYL84g6oKBG0eI6EFiOIaJDB3EowpYe7eVYLTS21298wGJNk6wKn+ynAb
cEv/lH64ULy3nG+Jp4OCay+51CHAd6UZoNFfblwAFZDEv9pOqgRi8i78+GBguGuO
tvix/1dOepxRwDEHXNjLjCEAvSUiHPKKwS+w2tI7Ao2CJQW5LC9PP0rvkTgMubxt
tLL3nZyvufcS11PKqTZAPIShmbUwiVTKwcjmjwicdB4uWVpC+UL6a508vZgknGSe
Lw+IvQfGB5d8I2XTphZAsQx5vQZqZe/WCdaEaIATiUsXAksde40k5JRVP23XzrUI
eyg8mHF56EB72fOqh0/X6eWqg9YJRJnsGmtgmiPSvQoR2Er8nG8DGC4Xio9o76DQ
mMIEjifBED1s3cgxL6G0SbgM+xAVcn3nzXzsiv2mmuAs5ExOHLIkVrCGncjJj98H
m+dgjefi8SaUUtayFOuVegQSMEMQfylZnJ+3hP6F9+g5a98PRXCIgJNnDzTmugEE
Dz4WvYdLrWKGCVEkJRs9P0TEFiihH5QheBG7pE3yUTCTk1Cg1zjk8R4yW+cls6Sr
MWeuSG0zGVcPPiwFWtyRSDYQziJRsmCpQG6LiAXitgJ4kb4aghb9ShjfRKihWAe6
zd7G+WRkihhweHwmlW+UUNw+jccy5OsNJYZQxo2IRhp/Afwc8pLvEJWhzN+Ghdpe
S1AuFdu5+TCOsMGS2z0mX1mxOzSwNJJjllZOnucX2U3vJj/YpN44UG8oWIG6iXhW
LI/KY8PVju/Ta0pj7FD2LmnoxN/1Rj2MYa4nELEeOiIU7elNjh1ChuUnrIFghC0i
ZcGv3MSVZYhV2rH+/C3xDh0L2UhRHg+MXoEovRYGNTKPVH6E4R6jkeH1oIZpeGvp
VudlgeGtbeH5F2v4z9ocvDq7bIzNQOdy1JiErApVNhQlJE3tkgH6gBR2dMIN/v5Z
8CWq8qyc+TAvwD+9sgtRZAIUpPgJi37fYPjmCz5HSKHYa4SZHJ4hxN+7ai5hH+wZ
ll1ciWyh7nlqCK7xNZ+pBuVSiHLKCn4tihW6dXILTd8/rWM2pVx6rESVlJdvLA+2
X+nkwp28RAu2GZbU8ZV0tqg62RuFrZHsaXU59B6qbdHaZlLqUfWkJklnNk5LpCKR
11Kkv6iHkm8TlaWKaeRunsX0jDiVUXwOWRBPDhC075A4XHQpozj2K9mZKtWtj8kL
JKpPcfeYrTMEj16OqGnnwiojDIUQ8/8yCa9PzW3WA71lk5tmDcre69LhyyNUv0sC
X/47nxw37h+xKW9OTXODcRA/pvW/y0u/vRQzzil/tUNDGc9S5pKApzuraJSnmtS5
7JZ7aWQgDvUKgBjAjzvnTcugVvNQZNTzrQHgqXPCk+DAQKEJFrnLdLpLq5ALQe0H
61AAk0cXh3KM9etQI/d8rz8JTMHzfWcBFGy+qkhE1bXKRFFDHUttDSE9FN1Z4CVP
27QR4SxBxkA7y26keQ/321VzpeUmmhh13oE/F1nGxCZaG5upubn+DwkIocDfbwU5
rBjC91DMzGydPNrHla/xNS77KGR6K+I/zJG/5zzfsQqmlQiMdXTDPa8sFqT31XiF
rJF+ZKZpq5beBLG32miOcHUZG/AO8NR0ptc4ioZBZFX+VIGllElpiGYRuL5Iaqan
9UD5FVvDViXkKk1vGN39YW0Vcb2xBpCq4ojo796PqYBiwZ4Jbm84vdYYixnsvyzy
5Mah4behSModm7xwJjZoGlxfW4ZHRRaa7so+SNPaDn9iMMZEYgX18smqaf6dPkDC
Zpqzm4B0j/Ia7MxJznuZto6NZ0b7L+bW3EsoZWgta/+yBQazGmp4Pqe+CY8dXpgh
IIw+CSj+fBg0736fcu+MgdEE3BWRs74NzICcFSecWPTJ+RKratpHCbA+OcuHJuvK
fuFXGV4ag36UUNqxLG/JSVPN/sjiv9zZpegUjYzlFUwQF2JNpx1Hv6UTQOOddIdZ
YKQzc5jfTNIVh5lEXEvMjkjShP+dqD4ebxGuhnlX2ciEOXa/w2zeAF/fmHw0oThQ
AbERT/zSA3yFcORPzeKn7Tfk3T1Y8hO3K5ueGHNCWvHDyPdKE+M4L+U+TK3FSEm2
Jd411cS77NvJUXlXsMRBbuN9Yyn7RxYvsRl7GQqAr1xQI/dgAuaQzRXgTIp8Nw9K
/Pk5bC2kxFWumhCxRFT2CrYCQK+feogpFqaHFcWDPEtpoopDYnNc2DXdpLAARLTh
lN2PEPTo9f074q44QTgIkVcaMzj4gV8G8toRuDR0rJ9uS7rk96tHGS/B3cpzJRL/
2a36eiSMYsTwy7Uodp1gwnVIlhw/2WB/dkkD5q4v22T3eFWAxDpta8hRYybDTfy5
Af1K1diCqvnqgRC4C+TyvUuU6GzXa7sJCd1k0dkbrat9e2fSqyG0Sf+5PaGWrMWw
9Bai2NJrR54tAE9w9/sRaxcXeInlmJfDdYukC9WfckSwKky113AtzJtiiqmz0+aY
Vo/pOzbRGhWQ1PSibqzVVX28dt3aDcHToZzMHHQpEszZqvMahfpmLRswvl6juF3u
V0Rfz9LS3+9TU4fdFgIXxdagrU/RGQeL+DA4OYrWFd8ZPNFJTOHk34szDmX4IuQ7
T1y92LRwWN8rvTpu6VrSF8y4WRpBJ+eAv7zKSmHrmCAbIs+NJyw4Rit3nxlZIhup
6qQgR15Pyko4XFfq7+K5SH/pLbtDyfZNzoImjzW7cDAunyu2MxImltobWCdk6k+V
jRqgtJ5rGHGZsHMvBv1vt9uPG/z2Fr8SaX0HqwWPBzABKilDMGbW+Q8uXGWktqTM
N/D2MaMssI7qJS4MXsXAsK/5gNfrohPJH4NCD1iHs3x0v1X3JWf8w98TG082DucF
AJBrNWh8PG/sEh58cPJGR6P4BhHo0woD8KgoPESKbjAWcj9tzSukcgpKqIltgRDv
OtQi54g3vT9XR5KQCeoZcqlQhYo0SSt3tafslqPmH+qExkhiTdL8Ben4Lcxwo79x
RNtLGtooSdRDu6ZfbMtD9MRzHi7mhacWpYMNyJPry7Szle+2EXoOJI5G+2+f5fIV
fSKGhYMVJuGyST9gI9l0GC8L4rOI/T3WEeYwOYYHPkJKbtzpdJGEE/TMwHwej2yQ
4GSLgwo7AtBlotstsNjyTzH1XmdFoZZM2jDrO0CejDbPeEHWXP3fSPFb5XXAb2Wd
3Sm0COOY3O+k2Ze4SUOrHcwbTIdfKKJiihyHzmiXVvQhcYyaLcLmZC7TSn7DJ927
IHy+8OfF6KM4WWfXxRYLkW3TQzl5UJ3/LhOk3ogxjec3zqdgUwKn4P83e2uy1bNg
u1L7zoXFRf0SD/QSv82txSZg96viaww7g862uJRL4CWULbNj6HYS6qVg8DDTZWXi
uMbLefUAXuCZAlnbNUlj3aKSCZ+GApKNTN5xd+/8BQ0yaQQREOuXgvVy2eWHvor9
xnZMIzViPVYv/P2kEkpLWh12svaxCMZS7AErTM9Zjz7N+TLrCrsoVhzsx1tl1GDE
6Bn/8FEg8cEFScKgcNrnqkwm4s4WgH1o9jBftkn7zbp0hoTIWzgcNlUSz/gm2rKB
24j/svyAs9A7NdFKvjSYoJcJDVjIKw6Nz2sLoxepnbmzc9KxXOJeiPfy3XnOxq0B
qG6ZyNRSSfXA+RWRivnZmztf5bJ7m0hk4h7WCrsRVCOQs7tLymCG65Jx5IdprcB8
QTb9VjKhXEe6rNQlqbHXCV69GyI224teH9iBYysARqaqJL4n+7KmvBIsBYe12BwK
bmY2VEci6rtEVCs00ywKQfepUBqepVNYVAz+3X9hygwF8l/Gx/BxTzwm/VJfBqlQ
J/E7OVBNnPkfIh7m6CcRfL0uWFnfcdFu15psRSX4B7H6U+m6RDCSxyCqHCTM8xkL
RTyXlYIQQO+mMZN4NUAWROGKj3JFM51zSaGgk3trI3THIPQFnZqGnDb5sJxHec1N
4cSia32IflTPlyQhfumogIB20YirGQsyfiDxU19xOZUIezwMX6vjalC4nhrKLCpf
e8I/OjHBADz2bjfJ0Y8eqFDijC+RpqfMtHZudqdCbbvRcM3jM1C1nMhs2WmAe36F
XRmUtvC1HeREzQz6z7Kdnses2ltsjj+KjUEogUoS1g+N1dC8lTlB7g+UtZBjh7W6
ymgA/+lRP5TQxRYBmhhwV6fFXqqG1GZEu+LU9ZpR7dOnCwtEw0tPtqmPMbKo8kzU
YjgYBijpnj3bUGGSbdpVvUA1PoF0j0za6Csngb2ijUD5H2FUhjUZ8xJ4DBPK1Lw6
wLIc3QNjB0q4fd3Ug6iTBc9xhPq/ejLbZnKmZDIuLqapqIIk0Hza44NDhPZEVtTN
W2m5/OSY7tznd5S6VP2nzGo95UwLJ+ugIAXVXj5/Fc6wOqkrXhgEy1OiqNBHNlkT
ASUJq+4+3EnCSObBKdDNq/XPsEsQGLs5+6O1toXQ2+9NBNATNFBqtUcfAZvd8ORw
gpciSth1urzvx0XVa6urX2EUjtnCskC/yClUMpu7Ycvxp7jq6cEAhc1O6pkB/xdL
/pghzNjxxBZZhMJS7jxtQVjIlcYhLyK4xS7nnKJMHNG/kQrI6nSmBg/kOx92pN8R
chvO1I/6pgcku4XS0HEWvjNI52yK9JoPq3+nDAGn8/LcjiXeVL7aJq+OCKm1d30p
uLtB4oohr9NmmmkA8YBCL3RUknvEuEecBaU3jKNg+WUdW8b4pv0K9c0HoogWtMHn
3/82d9e9VCUfZTMvWaVtyZgyTZuGcI2i/oqBzPnsFeuHhgvUt9Dramz5Xhhv3Frc
tiIhpIQaOcW3Zyi8rq2cyfhuT6Comq4LdqQcVvpEzHyuAWxWBbR6na7wotkNYFtK
NJ9qV33qalkeupqqRvFuUU0jWYFns3ZiEPISC8rnzwPHEm2HCAJ5U8yPJWMXZtSS
hNta6ARNpUQG1s/jKPHjDknsypO26isBTMdYFvuyKEEC/LgMXmardr6iXCFSOU6t
QnwANngTRpl8H9a7i0YSGTck7dMs+pFzcCjovkz2JRvYbbZ4LFOjxM+dB8lJVEJG
jr4asCXL+F9j+8ZGdWS3wiauUFrHr4/yQ6beqV3zhIRPssH/qseJcGJ1LNrQ6Qw7
ZTc4MYuwchGg6Gha4O4zO77p93esQ6pyJETjGLdQz6bFKPmOt0AQ0a3FKDur5Wfj
vshLfWAffl4n/1lq9QGV7WqkRx2hiOSoE+90lclNujX0VRGM+wWnup9PsxlwRvl+
j7YobYHXoL5gN3fKxi8Hr7g7gXUDOPn2WUlWdkclLH9YWlfEUpL/X7hrw1draZe1
PhYjB5+Yvzori7bBZIf2DXvdTXuk0/hObIugK9orFBXkMTC71R4lKV4zWb4TYxL9
rif2NbuQtpcnXvg3Coc5qRYmi1PjkOLyeLkxaOCv1Utet4MO2M7TmXqRTeJrAWdB
anQeWJTZtN/brz7wdFoe+vowoaPeE7h9CxuSuL0TQNy1a3Qp64JsPnzNwYlyHiEG
DlcAP7DH7qF7Uzhrc7+CBx1Vz8ayatMiQrv8NleGamBNqurNaz1RHDPJUqAIzd3R
B0Mk6EUoDHEZLhYAcqZsJLVaTdj3IngOVkba/p4p7+nJDG0oA4tVvYACMGeG2eIh
z5P1jw5VXbHLLobTkSC/aY5ydhF4Nw5TMRfvsRHFwJo+V4zMspXxRBR90i44VZkX
fwLUZAru2LE+pQdoiUQpY7JDzd3Pmdhc0dUBOnit0E9DdmGzCp/P+mLe8cKk0KZF
16jZqrI9um1eO9WV/8S6PSlurGNwIfGQg9frGzQkS+meAdht/aNKh0ilWKO4tnNS
eWCXDn6YOGoAH4nkjsHfAmpDyFCLS8DtiOaBu1q4cR0rDID9GPlF6nRW5YRZG8pX
HLNoxlLAXJ5NTCkVfQaZp8gipWxZp9CJ70lr0doLBSa5biccIfS8j63LLo5O78ll
H1JY7Uboq1cvNzGOJHLVDGjS88CyMQtyjaOMfsoc38sfwtB64Z1FLU3mIF05HuCQ
PyM57DMqc/pKG1+5tEz6Yyef/PZwCl+KvUFYCWL0x+2c17RoaTJ2kE3fzB8M7JbW
pX8IBovcYTV5MxDmugI9ZBEleAD1kkijGNb5ZiLqIf4Ad6Gf2tFuL4ktJmtlJ7/0
YEB5JCUFkUM0JL5a9MqfuTinJCi0j50FrsN3zcSQ4tc6yaeMmyEbntKBkPsYesDN
/qWf6zmyXETsGPzraGVd8gURZX2K02ocx1b0uKR2pvZONgt1YgvhHIS+pnP4JoHs
GqWpJBPYB/qKcFkrkUN5H7rgw772NAuDubT3ETKXVgXxNv4/PFucc/fM0JQwPmTr
r2nYSpTX9hA1k/n13uQgb+1a7vUJMIl3BvPh00Rby3lsxQ0NCNjo/R3YXNhFNv0u
kqj8ibAZqm3thIs54KX9i4C1OQndwWpzxijaeq5ZA1roWq0cXjT3H/7kI7ZEjsUK
i3YTQ7pHMCp7NvuB5xoScEqdiB6YMm4SNLD6gxUjl1wKvZ33R0DxrEXZNKtKwR/X
F+/Md03vIhURX5ybg4nJU6L5Ipj9geZWp22+/mVu1fgzqEjw3jqR1GI05pY5MlLz
dbaluDuRGXVNnYGSLLXMSLI6mNwwdFqZbWg8EhWsRQSz21dsSDjQ+69H3vyJ5En+
odOaq8u3wtebmI4DILAfAxlK+VDBLXEjhNjULc+qSewmFshExNrP9k6NO46iysSj
emvTLytR4ApDUPqLbcD+YY5xpm4uIlAHNWvaRHLK3fscfSfDanmFFl74ZI4Tf/qu
4+rOW3Qufx3511VdhaKWAlV1dqBda+LbDyZm2PClC3eCzdi8kSdsqdNwyrhV9228
Kteo0OT/iZfxRtkGJAGDDW2invXycEPp5tNu2o7hiAppOm3Fwl6EjpWwSABLkCgH
IlT9TGAYGTrehvd1z0R753/ADfgYA5TlBc54dY4tLmFwGWGtyqv4Dun8S55w2rKY
vNFH6+8ThRZi4DcyTswx5ORydnGiTQ+BeKKd8YUS4IjHGcgaATCpJ7J3969aHB2R
/2eB6bbVHfBecww26iWgyZIcn7+NaljIRaAezSXxdDrOMLuFIBdlejE9YNYtJWRQ
3CaW2gmnDhwU366zRX2xspbCvcHKL20iX7g6mllOwzoU4nZCyGzdmMoj3ZBPLEsk
AiOuHGB2s/LPRKVHT/flU5OhFvdQdKrbsBLO+/xU1+r60NXaS6+937YTxWUROLap
L1SaqOEt6QSOuDOKESx5Bi7B5wnyiFPL9XwvwT+dC90OcElvtjahyRpwQDSIhgHe
eGqCOiRRwyPwwwnBg33U+pY03XxlEDfWsOO2SxXuQWdJydbYFdJhr8JmGJ6f+r1Y
CzowmDECuHpj+kDqXyt4DGBdxXxJCI5jJ3bkhfVVFMEjoioSuaoqs4/0uf8vLjIl
J/KiwfSzujaV1BbqAtAw6qkD5tNChCKShtinfC865OqTfNr0BmjHTj0b2XbmJ1tH
1qszm7OJALY+pWoq1ICqYUU9c67/aFUMols7sqmddkGhJP1lQM88Iu9gOB4k679C
pYJrCFztP2D0IJfSHDYjIbWmI4GhxruVvNGjjaqjTcuiBQjFWBYfspBMeAKhYCE6
y6wuAAf2THmkjAGmk7DY6I5DCjLDlgfrBaDG5pconpu2CI2Fvqcv0bLMJY961nfA
9pgadHGoB3fUYV9dJqrMrwucuNfYvosUgM5t4tZv7a6X5f5FqCZ2AAwhNGJ98W4S
B7f7wll1Kat/NOGepTdmV7296aKpx2THwT8mHaEeQi+/AMFEZhuHygh4AVDJPKIW
fTs4C0bVYnoZ5H7fatfkvI0J3tbdHi76PhP+iRfcu7WHCUu2sR1pyFShqyEGAylr
1CtLrrz0BdRSbCXZXiPHLCk9z6t7Sw4J00H+rxg48BPe+zv0Ldt2L4pnfCHxcPrM
Xe9WlrPeRmwfqZ9QR58Etkka6vYjP399KghjNoGGRmJ0tJVDlWZzMEb4C4wbwN4F
LERL+QdyG6DvG6XKmIR29/K+nDtrwfu/9BPbYrHsUrsGHoRebC+Nrh9eFsgq/2df
nSJfXeOIoj+I4ZZ5/kr16FsFC7uE7YiPFaA7FdwCIV2Hx6fp38OsSbpt4tNTFVP0
VYhRTaRBqruwRPKEKKVa5t/KCAx+x8vlf2RNlO/4E5xAtQ573tIgzT5f0/Laz/rS
ITMbl/g0P0ZWFA8KvsJiouy0bzfni+iJRJz/gas/oJsSldI44TV/i/t7nh/KaBrb
PVsN1dboZY2+A7KVeO6TbH38jpmxOOQkEd96iz+/QOoWYNRU/ygMbt7Ohs/3boH4
bsRwsIuUxNPobH85EK4LaAn/y441e/GEr585T4IMMC4wMB8SUsKTsiMAvN7nK7KC
jEPdNa8eNILf+D0RaAmlm6c5offFeNJNl2dpLaJelD5q4hYD+vFVN+LfKV9LYPPp
+U0dTOp8T0evFlobN67Tb0nCXdvlpyKR4dEzwVde9SOQg8UibnejMdCzffnIGzHA
hZtqdb5v+uGw+XRjvpltluLh/cH0KQ3eYa0IRBDSSbLcUMMyKHMmD19Vl4iyp0rX
Z9zK2rOuNoJaA1jwd7o7tejA0phPdATQHQpe7iILcBDbjWSG5WXp++W0RGj4GXgG
+m3BAVDpJvhIQn5vJO5iLp4PviVlbsQDFUegYU+lvQ8BYOF1+2XHaHFeOVBYJEtB
KVNia8HJKzi+tWmXyxmcCEB8yTZu54j2W8G1l+VBpCZzcqjL5cU/JiDpPGz7Wlwt
HkRDU84WLPnlxDmGsjr1W/FJUnRlzmpxUv9otKbZ39HoSJV8MA9I65lkd4TscIoW
B+XjpM3kmjdMY0CIx3aPxodYpNiAG6Q0HZfj/n5PXN5MR8CbU+5vM4q+TLseRHSu
GUz3ycATtS9CwII0yBmeZu2R4SNO9Z0Ktq6Qtj9o60aSwrE01YIanHsbhNehgmXo
HYAG5/LLaut67N7VAv9nnPC5iIEImVUxnh79f9mOwVi0vMlkU9xrtX7aHit8hB8c
iag/XYO6pbFCKqKlGoappqzVzJR2y88PXgRyzv4rHxyybgjHydfYuOd/uyvatkOq
wF3WDCX/Mjejqs1XlD0UIF7S6leD77vv/QOqTA+qyTsZm9b039fSQ/FB09IKatuy
TtmI3CDhQiLyl2ocZv1+9RJk2vw6LtBKf+xH0ZjRqK8WVdGTujVamqNpT6w4qESZ
pcGKFdYzi6aDgeCOkuHDwJ/gWI/6E9i2UhyFliDeH3mMwiFDICUszTr/M//+uRTr
56o/HlEXWeQsw1BDTBmkihYNiG8o2ccMMO8jNguu0nyHCcAcOSu6y2qbl17qYznQ
cutHugWmtjP0Nzo26s4tc7sYlhcT0zvgy5ckLv9lmXr7EZNUQofdPKv5DFyI56fP
vEmqkETQV7/QMJIb9JrolicptMkN9f7Szb1fZyKuXzMKxQzCfJUS1O5dM9Teah8x
qkJ+h1i/msgoaY2YZR3JHOWWB2KKNHowFmkILe4Jit7pPl1JtXVZzNTn2BECrudp
Y6asIA/4aOETspLdVBP3u4okTymcABWuoZIsrFJaswPmhqJMUtRRDCLeNwoxgtmy
G1t6goTdNcbI3QU6cmqOacdbtZf02nTnxa7RcAdwUMFMF9zBBFeoRlZZKTCsLzM8
wYOD+8w1OVL+mwDJdj2QEt/tH44vOvbWHQyouASYbz3zLNSGtWUOwtDqkN+EhGZa
rZscwosIPOnZTnxLlewVpr9L46mx8HZUSrsvp3iexWzThIkACYTPc0f4p4xSyePV
G/K95s7+MQLJgR2mOT6QZTEahataHX981SZaZGiepieXi+JrlXX1Iag4ccdHNpIS
46F6e4kaA6SbteP8FpzJWqzaqfz9UgOBVPRUModwZixzDFqJY/1hZByPTA/9Cgqs
3ZYJtyXd+rdWncJtY870KUzuYnQnmHx+LIQknH3NMB5XhMTohvFjyAwYdiUalYjs
RrqsL72fC+H0ZUkZ/lAixC0ddHWIp6FAKYRCt1b8qy+Zgikv3y74bDcUp6kSHNg9
B0jlDckzaTxMChlsQcuTOMbT5ZqA9xyratGeoaU6DRUfo91GafgXYFPPTSvwqp9f
gJrcOzGIWsVqkK90comtdvKSLYJrBHh/zighXp3ew659gUVUj4Yra/B+bFQUmvpo
mfhfbDj7CJHN55ycmxhy+k5s0Erjorzr/iw88oFy+w1kTaFZLC2nF764fPcF3y1I
HatVwYaFNxF+CaTbvm+LNMUObyntobPCdJ4p8KHJz/N9NQ9VGaUapb2DCYk/OkfJ
R4slwvQgFsLcuhTHSI0uRYwfPmVQqawC4Z+Ip6Y6S/93CVfwtpbiKs8uSLQyuAJe
q+9jnNDMgloB4dDElGMVAZfm33v2SERhipIOh1Y4LitzS0PQ1tOsPRoNMkCz8g2z
/F7hZy+cTfxSmHxfM3nAExueyA5RBL0d9vwnunv36Xz2rVbJPFIFnLirWLeJN6ke
sjjQw/LO1G2Y7t7B4I+L9gInXsaXVR9ZbLTtp62p9LA9zQ96VvmIAhfRtA+NTChe
s6nBdNAcldUCmRBDgQ0Afd4/j3nvOnWntLp4oqGQVl5OJYNkkC9tn7OOE9SvxW3c
TD2H79XwvAQ9v2dIaI1Sb+n9Sq38Iqt7cre2YQGVQwfguk7OENoUdPkq+mm8uibl
2a7SuGLPUgut/HS9VbMBOCeosa2M7QWu/qyNC0pf5cC8sjj+O48sSe3AjiG6Wiea
71bDdPidY4bwPWhMQxkGSV2W+fKiW4vYzgjPL+HIgEJBJBMEQ8oHjw2+fcw/JlBS
z3NFfmKbtW1odpnp52VHYgiGldm3J8gow8Tck6J/YIo4ILfIq5OvOBoTboKw+i+Y
KOATQ4yF69+0fTK99vUyCD0yltXi5GVxoxZWa86xTiVAcFIGizaaYw/+9GQ7Lsj7
DBluXqaZkuAI2kBULYIbc+xuGKr9nkodoB6ieU45w0sgOfgmHuAkpCf/8a0ogwTF
Cun9p6mh0gvScyYM8MzLLbadxQRFy2SgfCtmUb290OSw5uwn9/8KY+NSGtU86Rua
z6cFZaHiZ+OGe9Gu8NwJqghDPZIweVlA1YUdvJgU8946Q9dYz6ZgVBFXiUQzgq72
94BEBJNmMLOb4VMcdR9Ls8i5Q4QaxRLrNmFUfxL/ZJi3vi3VNzpekmKBK258bjbk
DueYlLrxpYQtakVY9SbH2xtdkWjCP9VuRC90oETpbqXi10sHok6pqtDE7HTcyHUP
5p0rzVY5DLAVlWGL3uvum/+aCW9J6UXBDCiAipo5K9AWo4aWV5Z3F3hgq79RQx4i
ecuTwWwQ6690DtEO+FNTreex1N8JpPOjzuvYJwC2wyxYnbp3Z9G5b/wSXXpXUfGy
vI7MwyVIGGvqB5EmcIvOxWw74ER6pOGQgQVOrVtDF0+lruQ1MgyYpvlM1v+lEz9J
lhCehYBd/blRlFzTgBrkTLFTzv5ZvRAVNGFlhQ3g2SxksDd08r4XJDW5xSpTiceS
oCqZ1diTfaVt4Exg+GI4PXN/AAhMOBZ+uxiAErTt1yymnGtxgJqEaoqHoNv0nRxK
bnhSlrtqEyqwgA7BMskG+ysKuPlYEwWSRaoXGJhX/4Si7xN7Fpkg6rlGwg7kz3/D
t3ir2NqTEBOYs7PbZcJhiwC8tAIK0tzcKnExCL3UKLbWAUpo7h6/Dlti45o1sDOV
zsJGxS3f0DK/3TmsFGMwfXE/1TKkIp3wAHwAqmHMCJBa7FcTxkR+w9PXCZ2fnwn6
XIRcasF6bG+z5T2QT/8HElOz3bD9DJ0OYNTCjWT1H15JpeNE1aMb0NO9tIV+qeq+
vooUX35GalNTiedgmbUXDjEN/kmWYAlH85OpAWzboLtknjiB39PJ8V54F4OOSAQj
soYX47Ks3cf3PcDoDnFIa1RzLybRsSn2lLMCPCBYWV6H4MCN4TScpbKbhwJHmH/w
5f11OhgX4Df4kie1e434TamV1cTQj2CF8yjXM7qQpT6Kdq7K1iPZ30IkQUFU6TQ8
oJ/AcIeUHLrbFWZcEl4ew7KaMWleyy5wqor/Oy0CBRLkEFv1OPMssfSEn4+bxBcF
cJs8OvlN9zkgo5xyhGlzFqowuKjZfm4kzL1XHV16g7ioWxG1isY3edC1lv95/GuZ
1V/y48KHEtRG+OzqexJJUQss+kQSAezKDkau0fqfYO0TPGP+Kzez2brVSTDX78LX
CW9NdHOidyw7QeCWhew82VcUdSfiQVZD/ajrPwVdq7r1psrdGUhWTN9wjUqSKQLj
mMiQrZaboKhnsd8xRoHjjcvnzT3ar21ONuphnlxrtzFQ4QVM5SICxy1QG4UYSmsj
qAXPv+cldVuMAZFpr4bygoivEQXJw+8C0uKZbT1CW+HsItBRzRequIksodamdmif
PLC1Qq2yqgau6/85k1yr3dD2Wdvb7gLbU9vv6kopGlqJQvRPgfj14gjQYuIITuPK
S0/Qa61OpnOdie7lpaddhXBwiMx26+PnTSCoDSXO8lWeGLXaGltr3D84V85VDs55
6STXt1lyou1SdVykY0XDE4zbGF1VxCk4ooal+iqGQy/APmSvo4CJ7lk/gSDZDrap
RGSX8KTnjeiE5Tq+CN6lGJj5uXDm3lsJlvRriGpyRjsB11512omFrvK0aoGftFJC
TMsEHq7wyNdn96ZIwCFtKjjwl+NzApbrL2qP60czpswYzqBK0uH0pSgNhAgUjiYr
WyIu5pGIYkauabrfoqc/s9QR9xYfYVoFxBy1d0sAk+n4qU+EFYew27Ct9WZ8rbv4
9BhrvOnBLP0sOW/3eGYHpQmfRdEdqx58r19NNixBF9Ull/tEdOR6vLcYkMHq6fOo
lUgPITv5NzM/jIdRvOB1EqNR+P8443LMpQ0stNhRkMc1gG2PxRlKSbNWetmFMqyx
TtAs/WglxNuF5h+PaDH6GbNQH4aOFyDIS2uckIUUmpO9pMHl5iVCELvz9o6qVsS6
6sQIAgYzvelP7J7piQl2eePUYYLi5Y2NgXn1MiMnavIUkOgI21D6vwcSaBGzazK8
xV+kF3IuZ9fh3NUzPz4R8qNRx6nRISRdXDeVquijLU0J4VtNy1rz7bYQ7fDuydE/
Jyu/v7wFOZRTmFBAFVZDc/9KWCEKLKW0UY3Kx86ZycRRYVAog8U8mnTWcXObX0HL
wwnPYaSXcrBqbKEIGYUBqemZb29zov18IW1hy4D2p1wT+dL2OAaHW/3zMJ30hOTG
cBdss6sILLqQK+Q915POYtRu0bKj6fWtx25GALZvMGDI4N3vHmwEaa/W02LM8LGk
A0Txm93Pjw6rkBE+d6POD5DKCUvL7qrVfHxEh/gAsa5iTWOG0b13+U23mahc5TTM
4j7394xMBXBC/083rmyakdaEPSvaa6B1yhbuYmKVU7S0hB7sKJSUAVJ0XKc3vU7G
ytiY8ryVQhv+REyV4jfPR8ZzKZrj9wyxGzEVHgsmKs4fn0KDEqjzyllyuNzgYl2v
sq8C0I6SB5WDxNX6rcJHhpPvR+9OQQOu8EF2phBhCAkf2BZ7dAKzRFhSEjjf9w3/
UAMd8k5M+SJl/zpq+ffGEL/LBIz+gixAyJyKLAgc6xwpjcwKoki7LKf/PpZNyebj
6HJ3/0awyro8ndQQ1Gb6Owknm4NqLhO+FUsvGe4zhruTVIar/mKWrYwjzPAfGxLU
2+LGSFXoEwiBBvJs9J4YkNyqGhX8YrtH3LMoVWQV+ceT4czo1RXq87LforqAXgHu
PqDoeQLn/+uG8Qa3vTib0DrWDH1tOvYQTxHs9RwbXj5iJymDmXsTOeSTnV2mIU5q
CuoH1FOcTFzl8eb5XlF1ncu6iep9NhuHYvGPYmy72EZooUu7Y3k9XosQxbRoRQNG
oYBSmfRhKMbazucW6Da31pd2oI0MD33VN/TJSsJGNzzMYEFEt9n7bsVja6TEqqUO
gvrdt30ElxMKxKuquNUzuZ8mdBnfRYYt/d0J+hBhO3GJmzLOjr5LNdfJIRKAkya9
4yBFHX1xz7nnrVWRj6l7Ag/+Qktk6lUeCzBUgA3cDjB44/CTHm/I+s1yZaTuhf+2
N/gi3dakKi6As4i622k2UPYE32fRo21dS0MaxMFnTkTlBY6DT8ufQ6GjQrQr0/4z
hILMLCDhRb9Ovc2gw38gd84NsZUhqjbBwoiBq6bTsbYgjbkpn9Bb4Ml7+pCxVg15
4AoWGZXkczhrr2/RHaMiw1g6uyEBThcJETfMpMcXzXL2Xmw9NkE1BAg8SKcl4Fv+
qQLSNO+NyCUdGnzALprJ02fJRA+Cb74t8+/Eu1uf5WJZ9o964XWXrADFyRzh4UUl
MYoi3ruWQ9C7cryMy/CJVKWNXYFPjuFuMSxsEZ+IXstqJX1zk4dcRqvavN9T9WFr
UWJ/hxp2dSqpQ9nXmtuXs8mX7Bke/5+JwUWlI6wqYhq7N0pbWoNqxUl05apjAA4s
SfAHtbv+4rwDc9NcPEQHe0e0MjOvcRp+EmBpJEHYLJ6zi9sNef/J5wTgxtvZow3V
FFi7wLsqeqHqdX87b8UnWBgNLpybX+PIY+3vbW/yIaEaCHQU3Cl1O6Q1/LuN3mde
74JhtL3LMG6KIIiLXYPNvl0IEqvXkNNAjEW+zhcZpUqCJir0NLxvHceHN2t3Wa89
zbIOord1P3M7buJyoXaMJwVvyt+7d+1wra3k9aZroM0wqwTEomVgTMtFFgtgcPw4
joquwKHB9aUgYR1LkCArgg8uzMHFIVIew6IShkOa/QahgzpapyQx9bMmZZf0S+Dx
hkVo1XZ921tUo/gXbsx6JWcl2mRu8PNvcgFOUlKEdNHqhbKOdjRRkdigCVYoMZAo
jFX84mbh27vQPiqc3pMK2xoLcKssHnGUb7knCkeu4sjJ2eDTxZShS864PSVoLNEf
xx0A/Yj9VU1xDGll+BB8lcnf/ABPuG3jFGkmGVLvTB/XCaAPCpqFXu0zis6Q1bn1
q0L3uFSdC0YiTen+RQphjpUGvyWY8V7mlQmeUu0lf+gB6o0LAudzU3Ij9EymvUxC
okp3evyqKm3roxqnWij/v6/hhRQ8yhnwrpswG45T8ybki/ghJPmkkSPhJS890P6B
xQR1oxgE8HRLjNzzWtBhYNz2KBdIHFEba0lthampLzXRUOfAZ3ftQYaRHbso0ngb
451l2gpAQImcHxuDkINkW4u9Y2+QcZy0RvZ7lICeBMdgGyEhC8avxz29FL4hZLxW
dhMgxFJLzl5A7I1lL0wVIfFKNKL16n8/vl4AHuNtvSRXI0pEoN3J4T6jqjXzDlcz
GYR1cFpF56OoS1Gc9h0wTeAk0eki1pQ7VGs5gTQOS6lC8a0f296h01cUtq39vYh6
JUoKzMTKnR8V7nfi6x4CtypCfZGR98nv1SsKG9sQeRTHz/aG2pFFDbiyfxtnmEZr
gy3WUgn/TSXj/yrOz3bi1nJ/X49zHSykKwAxWYcGQZA2K3L1yTYgN6vcnepz3tzZ
xCBCr1QwyAPVwX0PP6HOXeMAq5aFTQQr9itNvSlUQHGUuPHRAp48HZGMawF5QWNu
egxZebiCdIyjk9udGsbQ6+veHO6pxYIfnfrU5h3+WGcd805Gf4UnJVxxBphd+e9O
T/WzXHRTqUrizgFK4Txkh55EGk/uCQ9lkWiQ/4PAw2VwPUNZcMID5Be5nfhzSim4
+54Qb2xrmT3S4mgvf3MWkqU1DPyLpFkykl3T4DynTTmGPsmWnQK3fA3z+74jUL6D
9+7yDclc6Ls8QcAI556dFCpEZiSpk1RUYGuhlXiVnKtPydjo4VF2w1/+EJ3yDzKU
v3F+R5VQj0xci31kJth/gmcspYFAp2U/oreLbqgHQdlRiWcIy1gqEr1EkIeuFLQ1
I8WxszkX3HB/h4GBjy38qwsoLj/wfPKBoqYxzC+gGzkkAT4YK0HGjkcAxV5Upaag
e5b1OjFfDDIv522JUOJNa6zxWFGxBoyWLziy2R0n8jNS72lXUWZl2Lp75GluUn4x
HaG4ckonIokVFEE5sB8uHB6EPN5tzjgf4ypm54VIMhY0Cq+CXDrmAMmmqDsnBBqO
/LKWeHADKmt6i/UK5MRigyAs0/dLggZbVDizJhe2Tc4ZVOKz1w4LCxsIpx+kzOA1
eNLttMQg1rE2KJvm1uRHvwJ6woWxhvAcv6nxNdMi/J1kjavf7zNmZ1W6d3ZpxfIU
euBXecklOGbxLjBGMJQ0By4EC/LOEGiq4FbCd1bYptZ1wIuUCL006Y2bljcLRYWJ
oATMI10HWai04B/7+5kqxqZg7GQFHFh4Nk4JmpJwWi742qkjIaPkPmS7H234sZfj
7CZG94fB9aCzD6hSC5aNVLBgQI/gqJO6v8dCCx1O2oLQpykzNinQ7RWZXZUFd/1Z
4ILhnlLzdr260ufO4GCI5jHKJd7L3WaFSVXGP/Ubd8yoVdjZYUzZp+Xn/f7b/Z6l
EoUfoPYdy++qXEc1Hqt3Q2x0DGZoK1fI1BOodbMkFtX1wx1CE76n4jRYa91utZmd
W4i/COpdYskbOKnsqMA4y0WLoFC2tPQ5kKEw+MdMTnekaohg8zxJbZQmGCT6cdhn
u2OWn1VDRKFOFf92faQHLbC6SCV/hE/CvPSDz6034E/E0ZHRGO3iAXUsi+9muEAY
DIKuioZLkX8svG6plpLIhB+PQn0FNWl8hvJc/L2h23hPVEBCmg9hpmidCgpJLIrd
ATMv8YdR8lHZOU6aIA3byVmjmFpfKhUxUBdKofDFhEcSxzQBRPS3QhDkz2XGyGl9
VaFQZzywYx+01aTnvjbtTakl8jIQDtpU2v6ePG7Eo5kXmLkWHBMgpv7YgjcYwE2r
b9ebmNFc2eI4GGFHyFAa00JTX5IhRU2qr7NvB3+rkzL6cAGcrh906QaKg2vybyY2
HM4Z8bkpwfNEnZfnS0zi7lFK9a1ccuvRlZTu2QkpVEdbsgSihGWxp7s9E3rYrHvz
AusV84EgvehVj/0ARVmv8LolEaoJmIAToHIwhYMG3rpfOeDbftlzX3n+V5ZRb1P4
rptPp2sDTPiruekFZBmbLPQEuahbdAKmy05KPKqRGGLDQgpLRsVxIf6RQM0BF1Fj
yw+dG2YVTk8woBVDihDFS07d1AzvIZG5wl3clwL76Po1PWWsMFaTYMOevG0hox6Q
zadKpF02r7PRIiBx2hHyF9e3Y8CMp+dSdlJ4gJIJNu/KUiMht2oOmxyQA7dv3wio
ZDXlwFnp+/hkCl8eWQsfY7VlCxENE4ZpMfSRfYjra7KxU4OWB+vOZHxC/VTGpb6b
cy2s/L9Sq8WzpZWrGwJgn/PzJCE/NhzN6LxWnKjhhp6l9LN5qQTPaan5lty/VR1y
fL6x9n7ULcHtWzQ2jV7K/2lplBDrMQiSqxQUEGgyyJnhGsXc/35+7QXwxeFZssH2
gNKnM6KEGXye23rgDjnHAYQp8Am7TNq6B8VBPlBKJ6JdiAnFlhvNLFAw/gt9vedP
gBvyKSWy6DVRatX8FbQJNA1DcSqYW3qlIoK1QcifjIIBiAwwU+fk8TKxwwf/cK0e
IF141Kg5y3ovfzlrdHAlpO4PWwNtoO/La8vS/r4RwPDTd3S99hGDq/osPalkm7oa
8pgMrX/hg3zf+dDGITByzTZUDYuHSWF1WYEih4iV/JB7zHcRzpm5XsFsJt/mqmIS
LOka92Jz1ez/t9EtfRGVlxOh305AUtBZQebrsv+vacvs8YBkerRA9JOzuBXwvjvq
MOXFRTHrw2SqF6jkdyuP76xFdNg+OToiuuRmFAlWsUZ4gSaW/Mx3CExLyACL6v6T
5GXGN87//Ea1RvMZhgvY+KkTzo1eBt4mTbt8m6d7XpiSqT74i6hia2Tt7VWMUmfW
ult/Unw8N4CCJBvhEHnaCkp/3dk+M+TT0tEQDNafESdqTJLuMm8BmsyU1DFVous7
dCfPM5hctZjlQSP7JGa4wGMczNds4QBq2HrVPul0I/TVCK5UczJme+QxaQnUSakn
gMXmMcK/cb7pgKni6NDa9qhKqEsWa+WJLCijjN7qSmwJV/vv7MPG2UlXdph3RoLA
9hrA7fZ2C1tDhEq5BoNa0KpZ289mNc1qTxkP5ZLzObf84npJyzZKS2/nGnv1mYNp
cNJV+yk6OtIppxKuUdVVyy7ifWSBqe5QEdwUsvxSfIb7PUVAvtteY7/tOTUzOWjE
elW+y3FjyQRKZc+GdgZwjWt79oC+u+rYxw/lvjaY/xMMW6K2C+/EGUzLB+BZLSL0
l6S6uhQRVeZ3/7uszcRCEY0wXJoTUGN6mllfJQqlO3VHn7qmjcsCux/ImNs40F53
kzs/1SjT3//gSYcDjn0fGB0wem7qLncEIuQGy2AlbKRYkEEUsufMY7HEG3sLSTE/
g3tL0f28xOY0h421x8nv1AR2JMys5j2W9NYGbEZLRQKgpON/0nlMNnN1Lp+XZu7K
h5NfusAPVYq2PMZ7Yj/20pgvf3RLKdnLF05iHuCQLUtkkPOyl1nytVRk6plzZ0yV
u0ytBkHrLS46aMW0Gq6/afVeWtkFoEdDkGvKFnqRD36tZfdl3kkfpAyBJp6JVfx2
QYc2PAYl/DAxkRAjFM6Dm3S5NVwW5OU7vJu7TlX/uDcmcVfq8GHgYWWSKfdWk0ae
chQvF8sujkVS4if77HNRtnl+Gxpvf10BJRgqjssQ+n5JMlhzP2TE3dcFGb/3s3me
55y4QecNjZ6So7+0ugyFCaIc1Ih6N/kuZ8lCnfZYyiv39QXqGtpxzARmLJjJG+ES
php8WmDOkn4D9+pajXEzBU9rPUMfD2ONcSznneyIilyo5DY1McdbYm/WQUAaPaal
dKGoauZA4h/806lklsl+keV7l9GsrU/l2oIq7xbO3V4M+mueVpQkU7F403b6QSI8
YLrXZ9133wOAhDEXEaidTcwi8yriJ1fXmq+S4YC6c70VrNi+wGhz/F1hpTDha/hN
5VHUCjDFwqVIlpztFEWe2gbAfT7xMY9CnaVeGUDCB3DN70g1FX90j2GV+6uaKhrK
68FkrT6fiDQsjZcsh6XfNnqjkVAbfYaaq/KFHAbX47QGfWY0N0o6Um7jp7sW7Bq5
e55GaXEuNVX1X3Jr7/0IGNCLC80sAN6Ixq762ysUPIjNjjuoJrvhyE73Fa/UaEFa
omaUyynA2HUt/ND2bBPDxknyQ3bNRM/mVrbbglrQO7PTPrSXd/LCfmQ27td+JFYG
r+Jc72HR+JjfBPII6C1h/jM0QB3dTT9k2ud8mtwUx0xxKSpIg3LWQzMDQCTCrhOK
AC/FQEiLAI0rqpV5Te/ZetDfb/wwRqYa/hDcX0qyKTL3ZaBwvM4AqU8VrBxn1fkL
nKuBpKBEuJFSw3XSuRspQMjKrKq7w7v9UM9dEUzVYJqHgRiNLh2i0zUFiD32CVWz
ScP+42OrV75VelvOadapoNnEDJqqNF3zw/NzblNnRz6JftxF1jEBtn/ffgydvOMZ
m5BeQvC1C9202xqVlWCkJkAqCDZ2BtvO4QmJ55e/9oiP4YYgXW3x3dVnkpDikvj9
`protect END_PROTECTED
