`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k3tKkkOJOLtOAZRfpFTT7WfTp63/Ug2gVFndEI1+Hn0VLDl3J8BKhSv8ZUomU3Yo
0DXDWkdH+hNV+jt5GyNQaJCwtgaw0n8PrK/RUZ307UEhqW+lg/uVzqnw/1p9zFYr
TLrDFi/yO6/Q3PoK2tTNR9/kuIYNciK9OPh7NiDxomUPpO8pwymwtYeFkWggUitz
BawBIAtMLvEdJgXUvWojm5xa58CQLuXz4KhccozkH0FwNTmZG3eChIdvVs+o9kqs
m4ApVexnXvqdE5DyHrfn7Z8BHqjAHR0hB+RIuDLICFVAVmaqN0hHE8HfW8N78Lv1
UOldFGDnpbC5kp/LjOoLePF81hvltquDpWKtDfF+SKerbqIfanD3Ke0Y8wK1uzVu
M/JNLz8RBsQY4IJMFx7FiBuEFnRrLBFDkttk5JUOeCe/9tF2W4ecHsIm8KL6exub
3odEvOGP8lUV72LZ6CsBdCNH1g5AVtvEhXMdtkqRuqUj8mJlxjVxAyMjh1+iqQxb
IadZiUtiP2b1COyiXCso4J/FuWrXtH6gldnwgy1UtXcmpZYH/tLdo51N4da8zgkW
uSk4/VaXQmuDGmANjbjW8ujOn3oHbT+hCmZEGvMciYnFc0pj841vmvJu4v0Pojvo
kiQcefW4mZE+47ERElIWHqbShaD5MgPAwb3NtC3lp2IxNhX9SwgrMmurNm0N7fHl
GreZ7GHHK88CsPf/yaDAJ9Lb0FjfWuBk5lPBSDsvNJ9apu/lwT7F8HMOX69CQLNv
tsQMeSqTusHgv1i9nlJGmeMHbSq2SCGeTbp6EmG4A777kAAHhpO+qSFHB43MtxBz
wytT7OTHI6Pie5DMahfXNBFv5KYkyaxb0FPLnYvGEBn/dF1r1z//ywS9M+8+nb10
HsN8kdRWfCRMIHGK0zuaWOA3FNtwxEltEj6abuzyFp4vWMbHyCQo5d6IC30tMdvt
4JnoP0opW3jVNMKWBoBOZC+CLoSddXCm/92ua4HIawOa/OmIUNx84wag2kjXpVlc
/v6UXYBMrjLbb/1u99OKSPX7kTfyZjMfNgslENHWHdMjJYpHmF2EyA4GL5o79N0c
7fpzmZSIFtcZPVh2mkBdvwwtRV85Qq9EK5kVGnFzvt+eew4hh0CtMd84EwEEdaxg
FkeFCycaY/wCo/BpAzIdZdJseyxCofEF/wpa4tFJj28yjFokbJzQDQFTIo04jRMI
KgH9eJvNvqeURGfQ9MLWels5KlsDkqhI2WACUIdXfJQdrZboL3pkpJAaVpyG8C3S
WuQQ4BGc5Dw1xempTdOYYOp5pYmeqoS3Fa3ARvzx9DUFm86WP69Ci84CBmgIaRXs
Lmvxdec7CoX/KXgNNDBgxJ6Dy4jmXh/TFx0eKORcyGAA2jK9MOyjOXgoU7oysceq
bYEmqMsUWnMwJQy6baQTf/nHfAarz7TWWRgk6yKG/+yd5wTRMioHZbrq/GUrQ1U1
GIpDZqImWTLrRFK6SXhPEygsJk7RN3j2MLgUIGhJiX3dsRcxgny3lQ0GCZKUQN5N
bpTvigYINJAv8Fc/ZmXqn5Og5eCUKJ5ADZskuLaQg2e+d7SmUBFMYXnXLamDX6lp
PjzzKJhnRKLaaylRm74WDkUjaeVL83tV1we+R3naUB39Zi5cUtvQhJrc0K4Pj9Bd
A3PbUdSg5HMVHH0qa2SVDKFn+R84qlSIlcR+ZOW7ac4NPs0JjdDDxTNTDE006qR7
wmZIB03FJcpOdV3EvkFSHbsCtB9SM477BJ6Op3bO3h2VHxFEzF5iTTsCj82sYWKD
W5/xy+/LX3Glnv2Vud9g11L5HfBcgvR79oxBHM506bUsEppg6FSb9jAzsmJhOkNi
VsAnkCmN2MSfXnIkTa2Rk+DSRJzh37AZVeLyxzLnrjNM3NcoRG5r2fi2HYXEiP3i
g3PajLTbsmi8Wxjuo65uqqlzNv+hW9MC7XsXYbXWu3IMmrS3C5AwM9dBqd6JmA9y
hA3JTmN3BjZUKcLo4m6ySEGDn1VHY2+VsmuxzUvDN6GpD22X668/vNrD2HlhaTqv
nLV0Il0oaltJFNsdZ4ej0kc5rkOZ60UVSa5Qxtep/aSu+l4bgK0C1DVmyPF/yGxI
AQjmSHtiuDQy0YKueUrKeSh9knpAzboAeNl1AfQ+9E4iZn21X+9mW2NroFPL1lzA
cSmBtClVMNHx+uHBmF1Rpm63SwcLNDLXtXxRkNOy3LZGSBHk2ITa6xPESmQKws/H
0GzYRuUMptbVaQ6f85tFg7OPsmBnpHS/cYY0KNebDpcYUt6j+u+FNa9+U1km/IXx
T5SMWUdlmvxKgmbYYz+O9tZdCN3L+g9KUxv27sE2EZua8Zj/0vOyiqsxP7umU0vX
aJWbHEVKZ3L5cvmPeuUrjmFdBYWKvQ/e/PPw26QB5QImS26pY9T3VHDpOmZtcC7l
EIseKgfZTPM39qTEZUk3gkm0378cdrLBsShupJC9SPTDCT4kxQU1cnpgmyLpT3sD
ovaPPV6sHPRUx8cbaqT/25n3KumsKNZDhTyEE4bLFpmgTFA/Rnm+VFb5wAOh0Kyr
cMlZN/J1PXCPIa0bxvEoKYi8PrPo3eC+wK6/atHmvQhaybJ9btBLhUwNFwyRMaR3
LvnccysnQQ5GrSpnGNnUdpMpeGxS/OeACdXXPqSSN99F5RsnfKNlKF+SKP33E1ZE
cClJzl3R/viYJnmhNa1rIVx7ENq9rbz7cDAlyWtP9ZHHEBp0nW7LAHZ2QSyh28SV
jk1Tiy2CrQrLuppqUrtbhVjDnZfIPntvJpcAyysnxXMcGjOXJL3OmigIHnMQLQ2Q
8GNV9krUvJNx2ugeY4bH/PMziDvT9JLRtAX5G69/m/qhNKQgiilWb+QY/RW8sADu
V2MygT2dZqPfWDOJOCFe8bGTAxFOrYajKcbcGhwo6uhxp8qt65Bjgv40dLA8nLH0
WPfaQami55YWq0EmLVnGbMO1UhLyzxVqD9bMw6zZ7uLZxlJsPQGv6D1PI/RMRin/
KzdXgcp6rFN2dALxcCiHs2a9iV0n8TYK4jJOheLQcCOvV32rBvY+b+iUZKk4NgMc
zs9Qwu2UsRiHu8Ehyibz5+R6Euk8d4U4KTTDigWNB9JBZPDFY6lsNuq1ZgPjx41E
i/+HcmFaWnShq3Av1JTgb8MvcQfNVltUNWDsSI6ooYPXJzJRtcTQzLa4sJorWITm
htt9XjRMcQH4VZ89b3Mm7W/kFMHMOzvPRy387eOCGGk2kwcXVbCLS/49h1IJAhXD
wne57QtzZN1btetVPPt4T1XCW1rb+cYm/OSPzIKeUvD0WHsdZCwdXkauHE23bqqk
YCbwz4MBwfLEjNjZbKp/1dcxYE81SfxcV63PfqbUbG5EN5eUPJAurZ1PRux6uggu
vU1Op/XLpZ3AxneOFHaKPV1PUL+BLREPMGfnAFo9Vcz5FyscbWesN5BcaNdXeRvt
kxL05kGK8UcLIsWxIAJdcg==
`protect END_PROTECTED
