`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q53UtsFBc4LS3/nLBB4XUEABCDAEkpru/lV1PU2FoXShk1sJpZIAMBvE6+kbXcwg
SpdcHQol0c9B0aSVNxFI8pXo8gSGKoVeyezpb3rgQ+O0b0LMZYTYyvlIoEViMq+P
Ji8ebu6Hf54cNyMmgI78nuvHGg7/YNNiMy65PbuBHeBVEZ2aRXgGUSV0Wlg2TXyz
LZt7DCuKVPZt8f8Ivav7hpQptdMX4EgIgALtIOqtb4iOwzyimW2ke0Q/Adb7Dx3F
6OeIGoS2103CBBLXtFY04zyR5hAk+C/mbY1/axXywuI7FZmOkOtmpT1jZmNYX3xt
7l4gXOTpbIZVc+gbZM+fr0//wg0H5bkEq4QuN0qsUhxXvH96VE8m25ZYlunqP7CA
MJIdD9qBsc/leDYhkYLeR5LtP+ZbGPAn7nWvB7JR0PKS25jdbcxotiEmmy7n1Dwl
kDkL2s8Oun5JSOx7Kcyo1g3XWF0dUr7XCSQ5ELGr8DYC+aRJ+r8ebaifEh1bNJh0
yyYczadvVP+1ZBSO2KvF0US3/y7UnV82kUbKBoLKeIjM9jFtGeRgFiPMRsBIydjH
6pFnA6ijqWVc3UsLf7ChuuXWqsya6FJ9Y3YTMFCZKUHsPsZhW+r5Jyr8VxQvgGfU
cvlwrX0KzXR35a9QajOPkWV9AiZOZomp2Ol3X4phEFk=
`protect END_PROTECTED
