`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LtIlUmeUZL4QqwQ352sCEOBB3ImVI73gBNPQOAwrilPUO+oR0pxpCVjmJeYqq1Gx
bfcpAa0jmsV14tkjGqawMoN0IiI71FpKCXx3Psh+n5pm5+LIkvfOGJIk3buVixYB
VGVA1Kst1f2YKuGqIu1n7PnFEb744zNmUjzPzJuSaElulILekWbmZMRba/06FI0X
H28qKx9/MPHrOItRNnVbwC2jVC+6i6zWNV054xJQfzCpfiqAh933k9dxFISHMbz9
EcEn5bf+bfWG+9z1xLn1o2yswb3zhim3bhztIOan/c0fouOiALj9+dtUpfK15Xrz
vJyp6VzpguCmemhufvF9MsbjFW0aN8HiXoAIaKSA8jof2qATwlnrWRUWJKcVHEo5
FPuKVNkPvoA3wQZPnW9DVYFsM/lLIA+wC3c2M89amwtzke8gmabOPO+koybq9+hZ
LvZZC5HWMnVGJJiHKLEbwbL0utLjT0b1Dk4XTjqC1bXjYirDbF0YSvXNf0wAUeQF
`protect END_PROTECTED
