`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P/moAYg2n3B85iIGZNmQLJSrDUShvHylW3VZh4t/A+r7NJk12feYlP2iA6LgkD4s
1fDypRnOOCVLjW12coGEoe0K0XrGmrb+AYyWwuQXpE0EMQLFMZnGCgbO58XiifuN
6yV+Bsfc3FWSvXLJajAnZn0/FpQ7wo3ha06DXVcI2SyooW0J8jaMyuCCZw+ZgFgK
aIuJdReUFwjHF0GQACycMPXss8gi7WxkinUgQ0nZI9bDFYi0K5Lc/nLeZmL5NI8w
4Cm8mq+65VRwHOxr1wZeYrqvrn5pfL1FUbmA4QpzPVEBJlVqOATT6sAXixOuCs/m
OOoYAZQRoRhPMZMGhQXwzF+QmbcvTykiIYw0nH+0S5kQyezkQcP0Hk4Wk6cYo4J7
Wkx8acke6REp05ERGdk/ClXT+tVMDK1tVQWuZJmglk+yzYxOXhMmO88KBecKdGcK
f8wMFp5u3/MX143b4UlYpO6gicwDcBOgZ7rYE/3k+i+F1doIScUa+4n5WRFFihhq
/U6K4BgEIXcIBA5f4zJlUG2OqP7rcEtmKRgmIVYjcS/L962LrbyQ0JkQ+RWnlK/c
v2iYIXWBTv/cz+o6OZvU3xmOeSIeoWWsEarHj6pA+7bEEJ2PoHFbEliqyiyVKRLg
BnJNuuQMM13j+C+jcgIQ0PT02mziueU6zp4PssmaHhdz84KLNHfq5hteOtJe4KHa
lY3m/+u8I9GeDkJPi04KMA7h5GSdoQ2qBG+aRbM7OMdd5WRQqxPOzROk9wpEXvuO
UmjnSIoohzU59Clbm/FjCg==
`protect END_PROTECTED
