`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CJAea6USZfnhOtADHPOxBkA52hfhjRmsSbW0xWu6bqsyV+aKtGH9negO4kj7UkPM
XKaBgZ5/5f9HLt0MxN5NY2cLmGm79/jsOe1GTSiBQ+NY/wy/eOY6/srlRRL+WOPp
KqhIUdzZggVi2j3tDEPGMR3PlRxvrnW2G3LsR+0AwN+jvc+5lN8a9yHsu6Pig7TT
NSSpVyIhXXfpWiefds28/r3lcnow9MqACaUTrSkkpsPdJ5S0GhAlt+apCSmMJgUy
NcDM5Dy5Z/gmRxJaPaw6pQ==
`protect END_PROTECTED
