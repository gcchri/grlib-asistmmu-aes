`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RuFhfjqGY5TBx+OLP0yWR3P6nR4+j/Cybz4aFo3/mHbMRg3PylsPLXGVs29MtogP
Z+6S8MYe/YiWZITJSsULqa1X4XG845iYbCUInMa5esRgHtOIC3/Q4hv4BWv8aih5
QrgX76nMPRMZuHmS20llEgRByQd7KpY2zw1/MdTvZV7uWhojfYHwamkmQd0Y6v2X
3K+gK/1nht278XIRVLqczq/JM/Myd61JWRrHABR49M8+3GhU+2L60ZK4bymG6efK
`protect END_PROTECTED
