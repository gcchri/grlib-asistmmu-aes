`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gUqLSb31g96VVPpqDuGRS6Vdlm9rw1OS4xPZr5eKt9A47QdfKaep6I0ShW6q7wEO
bzedyIZ5J+HJBqvAgkY5mMJuIb3aUo2EU4svEbofKAMRuBd+GrCI27SMzc+pFVRg
V8IjMq03B6jLbol++mdO2C8c2UtM3WM3cD5WEctFuzaAXbiJ2cOY9s9XoUiQhGef
fiQEjgho0dWVLRBGLxgkf6+RkIC0eb0kZ+gOOfGm+b+SYsT8Odr4qTWaP1D2eAHF
fAOBEcyyx2fE3j044doMRNA4MJy6k3jFb67Mc04Q8o1AhYKL2WbcE59jeuoIXKm9
5e6m83A6rKvGy9osHNW3IeI81h9JP6+2D5ECAcBqej+uFDW0DCOObaFZYHYuhbVy
3HSjpQnpi3pTz7l5ChWXiQ==
`protect END_PROTECTED
