`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mZmsni4hB2fqkU1hj5PTXDGmlwv9q+XO/n+SOLfa7SYe4J9UXqIsFPhJCduK9pDH
8QFvCfFZVFW9Zwp5awGMCM2KlkZ2e7jD76Fsb/qJ1nARgQhGbT93hDm0Opbh0w22
CZ0u2H7AWxNCMB2I5T108e3aj/A56qviIhnVmBQ5ooFNPHy7oNwpIVCKC7NEjgQC
JYaO2JCyQa+qy71epdRRuTmoyVGhjnJNa6DzOZyJ6kmDrm4iyr/zFSjusskhNz8f
GNqZ70fGjIQkGxxGRlz91qYjmR2i000ZgfdAqEb3Tfk=
`protect END_PROTECTED
