`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mCPFhvwZY8Y/GRJN9Xo6YMzT6EQW6EhJ3qpobE1TBzX3/gbrzAtpHBquENTK5IJ5
mhxF2fQjGO+I9qJisgshj8Sb3B1W8TW4hxCM7iza58u6OdZ+vbPh3xvuVHkEklVv
WX6BoyHcnnTrtQp0U0B6nw7EmkvtcpvUH8XwzuS/sY2hXpfltU5f0mukvaMUvNvP
ECsW01q1F3/yibzjUUPspkQ3bDEWI+oiaughfZLZOgdNliau2E1ojIk9EmOEGNq8
66/HwH0lWlhxUDY2FEcQdPaylI3v9PGw01GjB3eOvlWXhcARCckMEPswvErPa8cX
XlOJw2vpRLLS6dUzU0I7ytt9AWmHOBdXdf0C66DSfVu7el2oVgTLsrYtiFHtP+RH
Q8Vw78MPTq0ifx9cO6pJ2oI+1WmRhgWr2Zbzf7La5kyt9CI73YvCVZJEq4N82gZW
KQN0lAjpXJESsDBHYbKWZwqhSBv9oFJnB6NVaGTdAs3ARmjQZPSpAxZ6vqFV+tZS
F1iEBDtHTyw02b3R095ws2PNLJ2v9e/Sx34ykrnv9iUMdKRAMmHnnh0zDZd8jN07
371qXF+qW6ove+6K/XwqRcUOPzPhS+/Tiv11EeTsb81VPVoswgYgnex8Ak3+oLAF
Urn+ICa1shpXW/OTOf3ByIoFF5bJkzNPEtCE+nN1Bf7bSRVUyiPrrZE8DhpFkJGF
Fm9/hka9gWSg/7YE6RRILR6b/rVft6GXr5v8GKJ/Iwu1WopPsgryQ7xDcsEAbrk9
tbspDM0rWRdSgXosO5Hpw9572oVItc75NbxDmVtV2FTsFXbQBwkcRCcToMoeVBVF
Ow3HRKVFtuE1J5cb5O2Pg1rLFh2bp+bJUTE/wRxgpQ4hL/O55Id1Wy5arRfPoJeq
Zn0ancAVP5kcw/2F2r3ZeLG7USbmiMNSIbbuR2aZaQ1IOQLgIGw0W6VNIfya70rK
hKKuHeDXxCxq6PlgN/db8bmoCrKkTe0nxvU3g1Z2ATZWxA7HOLO9dMkrSSQ07ta2
V0PeiknIXv9cjCZH2vtYPOVrY9CHFkKNvNtYK+ChF+SK4MHL6cwpUrzqGb703hZs
NMf1VyW/0Nb9oX0yLeV02TgrW074ztHOxVChBCzdINZVliv0sazuFl1dsGYB/RZO
abwjaZO+ctxHGAjVIL7LlT6oWlgADkPXB8CcZgF11GQkaxglyYdvHkyDKMOSLfoV
ovKvFqPMAv2xNRPTl1qUfqTtrV3QA+ffdkV6EsstZyikSafPXz1xJ1Q54YF6YHcL
KrkyZcp81HzNhD2IQAdfIove+k4bNRNzFcCtbcS0jFnIEcZLs/rzkhQcwLqPZvQl
plpxKOwM6K6dVJ/p/YNmoXsmPV0DdvlMfaTVvL7VjX0ed2PhrCKWsK/EdHNK2g+B
yc2SS/SMYMixc9ETHKX+3EIXIH9lEpk/8B7mqP3mzpfZse+qfZr/wd7IvTVhBHNk
eYhqzwChVqGuXg3ayATEjwI4qVD1SDpNoqFyECMnDSeRk6N59TMcH+U0IDGsjaT2
tHX+TvmYDBFohLWOVa3vUAEmB1kq0PgyDrjVx/HidZwCkQI3e/92Bb7alrZoUR6f
UCI3dmvFK4aT4w/G1yGvKdPhjLRKgg9CN2ZE/skSVt5GpS2Gp/dX94VskYjKOe+7
am085saj+s4NTP+AjwGTVz5oIoDu47jk2SPygKfCgC240ZABgmStyKKQbbWd5NKz
3Wc0s11yyoEGwk1zrlgY5cXX4FZdbn6N8gxozNAhcrnohFziZVsP3nzmT0JH9kSH
JewpGa9geTP0ZtJcmhLAeaJtA7H/ljfvsd9vYqdCMEwuAp4USw1X6LRGlJdjz9x/
842FH2+pOAOBsbVPhaEjdoIGC4v/3TdDrbMzS/vku8Vw1zPpzmpMRZtEWe1Qp7wv
lvbhZZ7K8EhHub7NPLPJQ+hmwuZ8V29dtjdN9ACFqFKUM0LNt43dvuztxvZ5D3KJ
a2ltbXsdMCy+oAC9YvHgxclz/F4aNkht0FZMjsqM8dA9wZm4iIcDCUzjrwY6DDsf
gC+FfsDo4924SNuks3gu0jhQbIhZEZHWi2N94S8ThN43LYoxTmPqS8RP88PZ3InZ
DzBG8M4LewUfPKcty3MvnQi4+Ih2GPyMJnLRN+05WCgwum0ma12qJXWZLPAnC73n
0/nodgn64L6o0vqDuk//FzVFXf6Bk4Crf9ligoGpmNmRazZTGnn2a/40zdW6Au14
DHUuOpVB83yNf72KSVNPYQ3yLiFazowCLr2QWxD8R41orTne9wNov8567lh5iQCs
AyjheIRrBNvTVdhobSl/JTh62sze9wze2hDgsylwxhcIWT+TdApYZGaLnHC1YDuW
HsOsIA6nvqE58FLtjlMcUE9ZMhaYAsN9Px6XGOspUNNmH47FEyjra82gFiJAKrth
O9lUipgbxOheB3JIFDjSOMfySLLpgjBT15fURrDuZlFjoAPd5aIUq0AzLtDBxOss
id8xDoGwmQsE6tKlPjBP8WmrNdlt66q43GKR7nCaNwqp5uZl1pf+AGuZ/7uLQd3x
96WOLcmirElbLRTkAGPhvKJ1o5IDNa8aVz8RTy2M77u1rWky3kexAgK+WIHY+k6I
MUE+gDJP+a9kCKhPpUgakjS1Y+Ryrbu0VFrvZbq+zrVBvb/90yfg3MMcBSauN2NZ
Jp79BSL++C0VQuL2zoaavzcikh6aIdILKyrr30oZ2L1BvSbyE6ONV+8GawoNcnjs
dWWz9ue5b0eIUPU/gYKLfKFdR70aFC31QkTLHmzGqpzBI1b3izYBYMA4/Lzzhnd/
vhk7MYi68ajAruZGtMKh3T4+54h4cI8idJLQ+wZpViZ0GkkAdvL2l02BSXRWLrw3
nZmEBaP3RV2qOuIGnBrSIlgFYb1f7HsS1eFFNC1/apMzUtHTDeX/ukqWUX2iNw5z
gaTmaGItqX0B6cG96NhuwNNUuWnjbDD4502J6QO1z3G2dlO58qYaXakg1BeNfN4G
E2YOAiPfe3NveGih0U0bzB75E9hxX838TgawQAfQLsqtskfMdZxBpDWWmnS6fUcF
m2Cet2QFoQE1fs5W7WE4yFUabwEnFkie3timNBcfO6XGqpQwd925/f2UFKvAkZKl
dwBF0xdebvTIyKQiSkaXDaaPXzzt2u+9n12F1ZhVQEy6XoXLJ070lqfB/lipoHwe
lYyqfAnUG5t2OrYls+OqKvRIPgyX28q4hA62l6hGETP44GctUJ7ZLBwPQysYKqtf
djRYEH0cnuel+J7IWufyAxLg7MGLdP5HTfQQPxZD5tc3NiNhAAICgFBSx6dFJ4HA
to+zivlP25aSGwsr0qHXxDvhTFYSXYmi8wz9Ud5WZWlhD4+uDp2JxT7BNwdYLbAO
HsL/cW7TUyWVZFJAnpbwU/F70wO5doN6eRREYbdPqAwGMg95VP7l5xlZA787OpV/
cSi4p2Eo4OohHsysEZvf99RNMV7JnoYjPK7t18Idm3Nd3flcA+OfaI8TvduaLHkE
rD5ZFmBVmk8kfQBDtu9Tpd7gEDGfmRlk96/owN0P7QujVJLbYukrZaCR23dSWQqd
j5dEvUeLIP5B7qQpfYEl+YdXlQvOcbEZupUAsG626NubL+KyM22aSTqJA/9gtK97
uT8vrfp6u7od5aAjOg+pp8ug5ReO2du/KqUj3wBqE3nlQePynQp2trrKLFJKHEQh
4XTl4E5hPa1NtlXA3IWpyGreUgXGi/IQA5Yw7OTMmX+HY8GaRxVUlttUKWCb9smj
cJISvX9xdfUicv1h7CcnMvBO6hcZ1IbVVecZerLhsanhKwmRuYF1wRFPyPlwpddT
LWlZCkYituelkpYoIgDM5JFvmfk5CYPaDZmDMyGeYiS7/cyy3+CR68iu54FTtV59
27Dr6V5juPh8XZp+JNwAxvB5cafA9M2s2vztWHC/OwaSY+OACTkekN6yXadWYxez
8Cw7u4dYfdk+7b6DNZ0zQk1lVNPALsdNYiQ29DxvzAuLRrRtD/SR75YdpTGwQt+I
FDthkDU6ojsfNMnryfq1HKX+5rIYQJiEQMcxuyQftZU84SvqWOCSN9B2MUfBFygZ
SLuNOg+mb/meaQ5uXG/TIoSIp6cduvLVNEG8KE770vz0v33apySoWwAppAoBkDdP
+0d+gMh/R0rQEJpGx/MULN9coVMxbpvKipEWDogz8Rtf6dBc9wdDw7y4kuM+c5S2
o9hPianodHh8n3w1KxYDSK9H8F2FRsNvj5N/gKPPy7mb2DAGP3DcthPpLinTePvQ
PFhn92pfnfe9znqyHsjtEqauy8YsUXezbSg5uzgZmMMjcLDmKrFbGfFAJHc6qxol
NLUboFBZcm71lBIK5nFbD7ymWElgKUgJHRHJXtd+XjVUapfRTxsKnCes2T45RBbQ
+h4UTQuN0wlU3lYM992cymmzKDPGIOPFnJAAqwsLIZ35VQ7LMENJypiz+bLgCql4
KT1VmLEkUdsioIeNz0y6zfdmZ3NbUHWTG1RlWw9/ITCw5MbNTDgtvOhw3g40MuLc
3FvzMOSmMIAMFcq8dMosw4sBWpRHMO4A2WixLC/ozWb86l3vAYoMUvatx/YmdEX7
Iz88ZbFokp9bqdkhFeSbI7OFjwByxpQkfgNOoWfdj8s9F3UyPscm1znIoOlZi/Fl
h34sGZMLZ/DgaI8fLkRCBuuGcgb7KPYdKcf8o+tnST8wbyOnjGEveuokKeUaNLzu
6VIok6kSKCDI8eUkcbhBvwrFdTQbAiBOuNgDzcrZ2Duv3vFFjd9nhIaBJyxvtbru
mMDmr1mUVnpeZIzClXMID65y0pmW8vVVzegZPsyZbhSjgQj895/YZdsgIohkAHyP
j366BKdX5XfHc2iVg0YyeUf61Sp6lG96JRQLY8Xndk76+zpFx5g8NbMxV+BSKvBy
Nd01/ohXMYxHD3YD/GHp034pk0g1RnKLyXRs9lnEbkeALoshp4mMT7twVE/6YHV0
1hKVhotu6dhn3yZFjnw6Nx9f5tsFkCC2u6vvD9cHYNlxAP7HASsqSPBGQK71JKfD
h3rLdVUomTU8qM9Ft+ydV4HHJIaaSmSxOtzZDeMxSU7zdX/I3aC2luzv8+mFwz/G
TQb3bxZkA18IKsuw9UA6jsaK7EY87PGRgA4WxYv0WyldCRk1UGlVkJOLzi5aY/vp
Zt60uHczIaXVd0DtZcBcju3SwUUeYvgOlHAnkj7N5+mZvsjTfVwbalVmb9gVw75V
AN7hanIr0Z8tNf/R+ACyrfKVdVVDVSYhhKjF2HRfAZUZ9fSeCImi2+2beuks3WV9
vwgnDcN63/3EwuunpktUG3bF2Szz4Jr2PWiDiAQ/CEYiSKfD3Jo1kRP+GeyyXnci
dQowgs0CKXcl/EM13JaM29pMSWLtw25AOze5LzuHh7SG9FCGJ9dfRL48s4N/H4De
aQLe2uaqmA6iw8YG80IMFNGZF5NuClaumzDMBctqEN09TFN9KEZxW6mtlOgq22X0
5zoa3UXEaK/zuAN260B0490yjYniNYmy5WzYmq4XzjdQdK4BvJ3gcta5+483f6+s
MdgYEVaeCVadsRep44Qu5hTJpS0PzDW5OKWEZcKDDzaGIkrZgUL/bNw52D7jwkuM
7G4eFIdlAqOLQEjibyAv5+vhmKsb+mszlxpBRNX6JXWUQWa+EzNQwkRiuev7VL7i
MizGdwec8dSDxRs0zdeGDo8qoGjU8+albM/cOL8RAyhht+yJE8+LraNjxPnXFX2g
D1ycSuhXXWr1Zt5sm3WYAZA7h8HaXwsse5Vv807DjGGs87UhzYRquqmkoxiaZwva
Pac1F3q7yXO/pOPI5qnU9Xf3KUfcf21EH5yh5ODsxRI=
`protect END_PROTECTED
