`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lBvAItCKECLKBEvt3FbmSj8X0txNI79Xqz+c+lqMMe2AMg5OARqPCnBWFGpfbR4Z
3QmZs0CV26rGlJSdAMNT86hu1Ec/Iw/kRxn9ei6clnYvQozK6GxMofF7F3EDkif6
VDBUxH+zYd4RopTRCRk2CUTQLvPTHKsbxnV2roLi60g1m9ibNysA726sULDjtuX6
bu3VTsWzfgeF7EQvsSkL70mkETqKq9ibU8azhM3ouWTLf44iDBNGoyi7pX/IMXN5
fy5NtT/flX516G+weKRUFPURyeyBXye6LjjglOh2WfBWwdApXZ4F5O7SEEtwspkI
8M8rh85H0bVM8YqU/yEc3RrlmfSryEqQmU/O5AAiSCh80n55w7eOXZmkZ2TdwDE3
uiodcE+5ZVfVsre+I9JiuG+AuZMF+rBo8fPxwRtqVvTuDpEM1Q5NGQ4VaqYWFjB8
azmz6KTTmFhFKgkY4qg9Zq4TjWAxpKu0Qi9o68zCGQ/EG5SKZ/vYM5AhjDGnFaa1
`protect END_PROTECTED
