`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2nS6TmouhI55Skcufy8QTIjexeDwQhQ4aOWJRnq5GA2gbM1UnVerFoMNoXvhEMB7
Bode2F8uM7bw1bfqTeaGDom6pTIlHL+VXgZo2wsNe3M4Mp9pMl0Y1pgyYeVezW8I
93Ariq4/IIF3dFb5i3Cd2+45LKw+qnS+7D6HIhDSnYD8Mhi5QIc7eSYWU4sqypkz
jdt1MbmDqHJp6AhUkUQTHClOTS+Rpdw2V4Rc0rxxRF/D6JiRfnLho4p/Ph3mfYRE
tYOpPKY8oR7nUlX7w066fSrSHaQNwc/4MmefR/ZuhqonTEEeilbaKCBTeFTRrP63
X0eBbi8DwFYIQ/peDMaZlmIGfbGhmJ51g/Aovc8bYBAFjinnXPUjEL1ZgFhGDDxh
w94bD4OwvxPJWu0X9rEGRU15uRxanVXu/Pot3QOHYlS0Mzg8EQB68vlOdYQdIlgh
`protect END_PROTECTED
