`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AR8cvtxsmMkfYlPJndapOjOYj85ygr/pP4M8XvdYDGRGIJO2lTVuQh1TYru+f4hc
mNNO0oD6P2HZOnr66n5Zb9ukMEtAbtdrd5sQ0Zkhnc08n5puXBjpS4gAuLyfXkwE
m4BMdsCzk8tZJF3wkkXjuPRv99rkqCWgRSNzmqB4kCv5QRrRrmXFQfAyyYz8WrDS
C6LEZwK/wT6mrF5jjCCUrV1GPIJsxkmn4wIioZaceBDaqvyUuRoAlo3Q28bQPKQV
Dc2sG6cpJaskDn++KiVEt0Kgn5HxXod5Xw/KHSwImGFy0sA1vhN6w7CSrNAQCVy3
JqqLAhUKQP4tCuyjeBawegKxTFmYCiUKvgSvuu1VWBtdXtq9M9FO7LuNt7s4piQ3
TPNcEqFr9cHylpQgWzOvJltpgRq9LvVY58sjdNuXJ3DCjv0A+fPSnB+bUDvIXfx2
kQHqY0usbxVdYapz6BbYfh3Dhnbum8U0ymFsaqSJv7ZoXPS994ZdPpjHHCXYafJ6
ud9+vlCnWfPYwfFQfe7waqqjLNDsCy7pXU+BSRX/tuwu4HaIJiq540YXoX3dtzhC
gmJ5b0nH1SNXAAcPuQNt8Jq3sYWrAlffcnzvxmnpewan17n+M13PN0bWMWg1iQlv
GhooQk+q5oDp9Fw/3CuGEQUN6QF3EOZ1pe7/xgVA+0NWZoLvVXVAeW6/t6toGln4
2ze37uyG9SKfeAdzzgsjbNw1DnS7cier8b40Le8aZxaLg7ByFXN6bzZGitelc5rG
aTQuR4dU6aTCTcsUTevl4g==
`protect END_PROTECTED
