`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Abr+ZxmexB0nCzBAiWiJ0EhMcKbJK7KTylELKn3lPSKt6PKASPxQVtq1cYLavRJ0
aPOxkI2Wn33+CIbFPQbdJOXyNbp+Z76f8lOLO5i1kJK59EQl6ZdXpr99uZ6OCUaY
kXWE5T6eJ9+WU66HxIDpBGYMVNuTYqiz9cuGrk4fE+01HCHrlQFRP9o8csKB9Y/5
Uvw18q70WH9bcqu2syse0UqTs2s3lfs2Br6TED3SIsMlSgoxbOEjMOJJzNhcuVhA
3WBWSg7PGU8qf7uyxp6qXUSGssuunbEAfDq61mt3kJwpz3rigA+0u5IARZhfoqAb
W4D4eZKOFBvPqDCTbeC8EvKKt5XSrMSnyYU7qLDwl3ayDS66jhDJt3RQ0wNI4dj4
XkDb6fFpMdoVOvArlwAKztZ18WXgIEpXtF1xM1werZ9KGu0SY34/V51uVBbIhBWe
dZQfl5pyTcwyYt+oAGGZP9oeXXnzvB/81Qr1j7AyUyZpVN68QBi0hdeSB0iWPTAZ
`protect END_PROTECTED
