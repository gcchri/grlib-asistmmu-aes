`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eLK4H4x0h53aWwN5jmN+ACzKyeLIZ4y0LuxQ3041BihFy1wOzC0cbSg5DSCataf0
81IhHmNCmT+jHEMpbqHrVSYjs4OVdkXe+hBKdEJB32pHa0TnQcJDTW7BUdInsy4B
klHfDpX40ddTDwrWRlqVMdfxWfZJjd0HFnB2qHSzZjYDAWf/d0CDf17LFWE72HKW
6MKNlAP0iTrAGCfHroSv9M6X6zW+9Wu1gPpM3ZsmpymhRf/T77a5tqBIMS78Zg3t
DsmRRXfugelM20PAHk4m5U2vgiTfYM0l8cd9qB+SjR55QgYGm9GTeys0V5A58J1h
Yb7agYbj7v7Sq9XKWUWDB9fMRWAKFn4QymZNmG5MY4D8M927VU9mV5WBwx7GxiRj
k7VUxd6irHiDMEs8g4ZpKHmxSBBQ6M6aV+q2CR634BAQoIkKBkOvyz1uO53a/0U3
+fU6YwQT3YrDggQZyGYv9DAWZX/JDBcLm8yqWhOhkuiYdAaJKj4KtoC24zx9bxju
E6l8sbMiZ1U214fWTuvU4mYRfw6IoOub/8S2o84zvE8RbIA39Pjsi4KERNB5xCMc
/5cNik25xNq4MEpbaryqvWVxh/BD2w/P78yZNeEYAIO/JLNGpZEiEMi8xEz5FRJc
8yK2ZTgIgiUQv37e5KR8f3i3S18fLtnn5qxX8PvfiFGjQzdgdul6I6DkEFvP8u6o
yf+9RapRm9NWC+oN1LXLSXtHKwdMRrit9s0Ge53Yk9t7TBtjLvBduP5vCkEa1RHj
+NvHAApPEHfR81v+CXxujsQE/ttOlsfAeanErqBlnVzpOB1gVhFSc2k+dWMBKrpJ
zfw7WEPlnfbPErv8qxL53BtS2Sh2QZVkVpVs9BYJwf4qXUrbOEDNWEwXB6iyUDrc
p3EZM/jFN0sy/y80crkArDWX+ejOC+yHsWtHPKhkaXWF05RbJ2T0D9xyiO1w6+P8
aGFMtU84JBSxccXEhcQtv/XxvNPk/byZCsyOGTQcP8GXPa4VTLnKIjCx00a5yON+
Dvay0byOD8EXJimKMwWbVYjdIo9VGMirEhsxaGMiPPcY1hAFdnaUHFunT16rxoI1
aW6j2HSi07Eqv0or7aRKHsNxPF4Kd/Xiv1PFoL45ce37D/oB1VKGrZUY0Q5dLhD/
pAn7g2De48GOKRm1U9OMQaSdBR1VTinkUASuvUn1ZEf3kKlIQDxLskBqeaPZ27lm
L4MCeJpzg994wPpkt+rd1U5hm8xyUojDv8H0nGuxZ3Uyc4jDmr2vptsuwaCh6DUW
NsfR7TGgxcPgKIEVmpXfeuYnx2z/ALp5BHab3S97k8kvf3lAEccBAh48PagYieJ2
eqqbUYLk3iGHOS3cHiOfFumgjlqwylccndx8bDDy1V73vJcotCSQprqqYOc1GpUP
jpmpXmvJpWW9ZneWk/wACQI5QGxx9pVYcQlJ2IrUMqrVShOAkw7URlhK7fJgHiyN
NKLVB0yZLtDQGjB6vzN3JbwMc06PTbZ9U0CD2l24bmvfxmnzo3o3qSVeb12H4xsa
82SiZLh0eN0gWNBz1Hqx0a+AUx+b6plCuGHUgRwQnKM84m+mX+MrJt5W59bbcB+V
KKJ33AFPP3MyWbHOxHOGmDDuhpiy2LUPZoHqAWBQpEAMZRbliXyu6HHGxl3NMcnN
THhfNqUkwuPzK/SOaK0Rsmf4aV9isAID8XtD1eXWReB53wBlH+C63OqSS8/6oxfk
Lqpx8KFmgFui4N4TTb4XqtafTYq3KPhuZZaDG1cwT3ktugOzorua7pdfUEcmYPyD
8c9BdYhL/N6C8Oqyt+s3eq1At1za6/r4lHb0ANsfZMNfHEF891kgC0F5xMTN14g/
qB/CtsmC5HnQc4yiR8RLVEjVG5gE16qK5Buc82oqqdroCfNzy/Pn5+iwNNNHfXEB
sJRUEkYeqwoL74yS9sbpRVc+inbhqxRc1vYIjI79WZWXQ66M8De4BbXx+oAGrB4s
AUtfbluvRrAObFX+Fwgbtsyi36oOpYWUtKWuSSoByQ9ZXMawqjyT04gsbHvYjKFb
817iyc/TTudN9E3LaWef7fXb2GyEauQ+swIJ9Ie5KMNJgFvExkhiW0XExdgQQ3Zs
KUhkW+n9b1sCnPgPj4Vx1lsu0UtFk5jtCNyd2xFAdGe9KP24yHiJvjyZtbLoNz8D
zmugDcx9ZsFN4c2TGq6M/3WLi5xpmgeyxT8GEFkR/hDfMW2wl53IZq0JPQCQTDw9
t9CJur4JA5QrUdjDk2v3ImoLGpyuokkFRp6zCRZgnUEhfCcfiRQJfHuhd72tY7MP
oKclvQZSCGiVdiUPtQm/dMKo4+w62QTpUaLFjscg8srYXRrH//EN9XC7QwZqGNtg
pS12Je7FfSz6BE7K4FOzqlDn7aQ+scw4sxJxoM1Xv6Th5HCneS7HgcmKCyCzCbxu
w2PBrDiJSVbH1zSyIhHiQ723uBB+7obxlLYsYrlHLhJdOeQtHTKcqyZrb+nE1A9G
HPS2/g3ExzF6W/ln0dojR6ZF7sWgu/fxzEGSnoUeDRzQ/Qo12AuhytAi/NSuBt7O
0HdKr2hIy/fP1MCuWDXL3LlTjW3EK6W89MUAw0dnoPrFkxVbsFVpCbl0qAAYzRVK
kUBU51GvEkynMsGN27ZxYf3RpazhL3TNQmsTu5ANFDdrBT4t3TdJ0xf5rK1eMqZI
PHYqzFzWSmjVUH8i1UCOyp+pebpp3qmVfnVcihrSUVMIvRD9pudLGgsHIg81vYUv
VPuITZZm6TozvjNTAYlxi0JABotFCMsYFI0PbRHj5RW6mQ7kLH9ygmZeq/qbKIEo
gCihSHU1wxms1Rud1Nsr2SCd2NhxCXWQ3ZABvYbLCiuAW9iA7zUwDJEHXrOP+/05
2QXLDYxgGbKci0imcLeyY+FuHPrWPXaaiUcFmSswHTptSo6N6TCsMoV7YGKAKVH4
obnS2XRDP012PQw77Ht6iAEkU7HADsPamtjf7Y1IsslrzbUTltEeTnqTcZmDucJS
oWHu6Oi4kxnnwIXpKDJOydV2td3OEbO2S3kAg2H/Jtyj04A8IJaacLlHrKWoF7tk
OiPAHNK28U/3KUDiyyN4QDKk4+msUrs3r12mkAXXPp8sYnCH3PWbydnrvCnoo+fY
5yOLMWsq4EDKJC5wGe5yXlPCpW48D4x/bXpT+fThkPoy4vP0ArrynOsonkYH1vgv
dVdw2ege1Z3II6yEDVTdjk67PXuu80SSuVEr6M+OErtTrUW6kvgC/Gwk/H9uUWAI
N0Z3sZ7TsfZV2GbJnAO0oRXg7igDq9Y1yZ4eJnK6RiDs8t9KjZGfEFr/25KwMuGD
0uoWrQ0BPl0cylIPoaS4ts2hjpEFPJt6GARlLJoNXEAJ52dovrWc/+YThNo2lncf
1Vu/FUPrfdvWqoUS9ikWtJ9cUhEnva0tLfoO8/Bm6ZdN4c9+u3QKOMEgiNADM+D+
JdkmAYYKKG/1hgGPoobXWE3heZ5eWD/IX9AjKKYldO5It7c63nmYn9RK0kBNPdR6
Nbhvaneqb8YHaNkAGA3zrjWtKvEigtmQEFHQJV/V5h9Zj4DmFzCkideVAtL4RKeo
SHe46ubJnThPlMokea0yAlueoXbvhgVssC7T+H5F+puY8usKW8iG37pO5CN0Ma1c
qL6J5vFOtqnMOoxBusT//Dl4hvyhz46COtQyYgPCtoYBPFaDgHAipGA/EiHlQ4+m
SGVIaavp79sk8RQVDi/aRqd8P8ggll8cdGBFfza10BOP6EIo0bwcc+rDwYO/aQrC
bED05cnZqN0rYkoxrOjkcs1xsxaOAk6f/SPjILZShJU=
`protect END_PROTECTED
