`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tPqIR+llY603CtbR5W+yIZRr6Xq/pUQrROrK6MFgglKyopaQDj1zpJjcVF4La5Gb
KKrJ69Gj6hdU1Uo9T40FMnymUTsmETP7DVXI4lfWQ+MSeRDxfOn6/+ewKKmxgGPQ
/ZQOXa6bPf3Uans8Z8yvwME1r9eKlIzjyw0bb5Muz+cGoWY+WPWdfQ9/QWOGoL6f
whC12IA5zBWL5cZVw8hkHlCkAs7fjKoK1F7dWEoeip2EF26WDiP9EaTMWqyoWzLP
+7c82aGCHE6V9Snj5fJR5Q==
`protect END_PROTECTED
