`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bGYAzTEOx661xvzGnSDR1WneBr45BpD+vu6BqjD2/1sHYS8pOkpg9hyUzwYirQD8
2WQ/QWbFzuby1u5slP9xtUIdlDxS5WLF7815+izv/lwc/3MBqoISA/hx2as9XgiF
uVtC7AnLMTy+2fLnDKyly81hPq9nkWbM8neiBN3gu6M7Hfwfqhq6o8SpZvNZNmKE
NEpjyR/x2Djsyz+NMHNwY6AAbDQ9weEa3lqDP0ByMYsePOdn0FI2wISJaM4Y9Fax
FxpMF5evO2F7zmGI4YqUJJl1RTn9kOlDEp/3JvhlF3tL4Xun2lC25/PKQ3hQWdPZ
uUNQaUj6MFQnvbDl0PrBNNaD6jv1gXKcrMuHZK/HJiD1zx+w2vI2Nz1O0kjwHL5w
lMAwFHp7v5wCqjLhnwrs+ghoI60EsSt4dX9APdkF4rjmdy/3kNk7GU4oVyYC3gdd
NF5Y3KXHUE1X4tx1SpKsBq7UUfwXXNu6N4WOPj0UlpvsgSekfhuH/RjzAewRNz1j
`protect END_PROTECTED
