`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
72s89O2QE+opqNJXdjyrw+Go+ePC1l0VoJ3iEpRF6tHS/xh04x5Eh8o/6dRuYU9E
9dU7KUMlp33PryiJg+YHys6upRm06uGWeiNGmhy1ecjffrvjTeMf6gK7RTKHdBgS
Xbgb9jH0LCdr28w0O+2HCx7RH2XP6jq04T3UKhICv7+tKa3wgmFNiDzQ8mOS1VrL
VMCQqEW2P3L2iuSfvB/Vq/6u2FLq2MoFKnCQCtnjgCCCoEQ6XRnUxlLZWi7Ty0YA
V0rMMbL3U2huwBTBhl/df/vq4n9VHIc7SDqEFiC28EV/MvZO9Scq50eqwX05Xvxb
KM9UYySUFA1da+uU2e+4xg==
`protect END_PROTECTED
