`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eVIHtVx0HvhE/DCP36iK7cNgMsNXJHeNjwF2epqERwCYahRU2NTUMRHKLPTcqRvS
KwVmXSGbPBCHYExxt/G3HNvsqcIspSZHXQaoroiog2euj9SoHvqu8tIZ6vrOE2RT
nLp4fgadhIyfuJW0sc/OwZpHjTUx7U3Hl+IHx63LF1It1sc527sKkBCx05yFWcQ2
RbuBPRjdG+vIsbpRYDgWWhVpNSrUC/UbwIvCOGZbqvBjuB0uT//m8njUY/VNx1zM
/k0LXHkGwhLQEJvahF000kw+eaD8jhHNDXsJEZglMnlc1jxcjReQGQpGXNOMNTpz
BQ+sQ9gPVj0/ZacOSB4qrdLcof5/mdrgOn1fy/fqcPU=
`protect END_PROTECTED
