`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d7yBLHgXIzb6dVttO+3xwdsDmY2gUcCy6jvAnDCX9JKfD4Z03FHc+hmJCC3vdliB
h/zx64dD9ts66KKm1P2vcMmodmXwKmwz6r9MI/TCEJXO5OLfy2VHId3pwoYm3c5V
6BdzPHUXu4AfZ1hhokyd7oE/jG78zH5mwLImLlOoCEVUBvhxKpdqgbbZOrRO525D
Kyr2IqspMBa3Iz2boj4gAwzZsSdPQsa/wG3k66gd4r7pjDTIIpu7xproEPs5QH3F
5YJapaSjrFAQGxy/DY6mmNirO8oe4iwvOvTPQb59bkCXzjK3TPC5ol5viPXZx/Df
DFNZrCdxWG/1jXmNn92z5k4pN7FUKm5fuhZS5r+MK6n9+k8gMAs63xRXjQ6cdbJc
urZTaVakMp48O310XJ8CJ3uc+WHTQDxRCA4Nx5GMxsfW2ZE7tB70OBs6YtaFhC2m
5jkS/dGSsEbF6noDTrVNBjRoVVWceg8QLAIHhE+IyNDKoMHT5gl7rU4e11DdTDF1
BzNpM2diIaiMUr7bCiZTNAFjgC7hbOEhgoX23TOm6p6fBj9GAsp3xgc2oyYhW27P
2aaftmeW3Qnt8V5okdnrhHBcIn9kLYafHj+ZrEM+lpKXojy4Yg4S1ZCR6bq6u5s+
bspqPFoFaSGRCA8tpfdLVmflcvkikKngDjXvM3iHzzPK0zLTF70RTiRVXaqLE5jz
VvQ4t2Ne+ug1oMf1JxQVDw0sH+RisQgU3o7VTb+1RfeqkEdgzV3QDeAUk/v5qkj5
TLhFcNyf16FPIRZdhGp1REeFSK4AAlkrK1xJR6M0lXFyYywinG5U93Yj/xpW2Fx6
KBbg448q92lsYS36m4SuU7N+BHdsiwCR/5W1v8K2TD3smmNAGibgCC/KLZMrzr5b
h89nu52ndfCy2CUYYfan9T/4QsrIXsU3Ehn06pGIa6nksJwLDKtTLBplUeCWYzjr
1eA8UQdM9NfSQP+YuifffW1b5ZEdHiSNFI8PV2anvZoiyOnZNdqeLc+RacHnCouO
copQmu/IAkCSeUIS1E33CuQdZAfoNHCb0zMG9rm+b/mNdhNcLWPu3R/iXoYkBBNA
2F2e/cuemFQbTodCB8Rlxy17SO/ihz2hgQ4z7tME4KFHRScoZHwJ/mMcVwCqTG09
IO7t4qAKkCTw9DMLNUmSkUiH7QrB2da5dlRjK8xDskkYB7yLJKA5HrE36CYQX85Z
0Ql+8bNbrrYYqnJZI4NN79xXjl3fhat/nlq/X/LuwQQoqSy+6VMpVWM+YLdacj7Y
oGNQSaAMrLkOqaejr3h53vYT7QfnEmMJ06aI/0YZ18JG3PMDSjym5+MwUKEji+By
GRx4ugk2rJQOH52OWVo4c7wdpf/LBsPmH/kzHWfCOyWiT31O/pXBTHEHvnXR+v33
RhNtE+2DWVlzRlMGKmn7TBjjV5QZM5nRgK5gRy8ulOIqFuY3HlJmUlXzwR8uM8Th
DPVeqQ6Xzj9XlHwZNG8gqlzp+iQ2cw3g8yC5PcxC/o6DTFDAgAwSF0esrN8YXO+6
ABUbUDnWjBflKRCHKueF7eRRXTnY+4XaxP0jIyLnYRtrHTERG7bQDM5sSbQa4Muy
vZdidJvaUGo5KD82lh0rNtyDyLl/RhsWlf7iO0YZialGevwEvtOK5mdC+gv8m5/z
y3DzaaVyLcaciFFcTuVvYBHp2qS2Vb+RPAfFEkfBC3Qr8hCSOQf/144rHI+hiy9P
JaQb2zDSy6PNBSOpgwZUIGQmre9CKOaPFMsF6MdESMQ7SIuZT0rOKqg7lo3sEiAh
xk/NzFgBtfMDoRbCZBmxrMAyZXWY3Hq0bo1DdUbnSCa5dsk6cjnPo3LUJyzHnElW
ewWf9cD+cD7ELkS8icrPpmT/SKm7jDkUUYZyIZ3QGB4fZ4xST/c3fns5pdZEN0lK
cqN36aeqXpGZIJ+cFoxew9Jl53dX4EWjENsjUHvSLbQenoQC4V2fp7MzUoIivPWM
tQI2v2UmC9pDxnW58Zi0MhUGvgJ4sDwbC9h3Bmlusr4ipvqew1FyFfhIvMKpLqKJ
LEQvaiURqi/bRDtOXonCdKgXjst9GmV4GpIsa8bO3Ek4J8WbXNhe2FrR/Tt6it+w
tNjBCPzfb8ZRJFMXxvo25sRMh5j/lE4LHckrAOkgJVCXg5i8dLSbDE64Cxvr4bWs
VsFB2k+xMTub4iqXhnQ6bKVRUNoBujwOh9Z0QZA0zSt+5tGd4b8qe9TCjrVeV8/v
/8HNp2gc5D6iM6E8pRTjMPUmd/Mh4EJf4GT8KfG6L6Ytwz0+t42hi0faJYnw4y8O
Whbg45FbEfWL+lxK2gnNqSwdManh5lSPlKVCtbTljwbnbMNKPrx6/mK2UKDg1mkb
JHi/uJ3f/VQZJQd1FQn0m3YvtliyYdXofKPRG+BRYcTcgBtTOZtMc/Y9t1vdSDJB
OKiEQGZJV4pwX/7+JrfXjMlIl7J/ZApGVqi0mnpwPnJh8SN3xwDWFFKFEKTzC6bb
u4l4GMGogpCK2tSiO+xFuZpoMyC9D3tJ5C+kxhCqbjqUBVFCbhXecjGcN/RwQvkH
fn5NP6NaEUupPMXcyAneOVxUDI5AM+pd0AT2R1rauJ74xkDrpmpfRU6wQ4VhNayb
oxS8R600gsKC5IRWg0xAyMTrQFOAOsjM3p4jW3WP1//Ej449i+fkT35Pi11UcdSH
QOBAbXGs2YL4X+Dkm9CmeY3l84kvlUMNI9X6hphslklWxEdKTIOWng3CEmZYz88w
mYDMhAbJruyNRKbFNSgRF+/Z16MJycmbyKsxJyifm7Vog1Yf+xTesutSNJbFQF4x
PgZqS83TFbFpaDRq/nurlGVwo69hqtrFLVbK6IALu2qK1P4v/rgFOdzkaUnrKnqy
KfKl7x3d9CJtawiiqWqbTAeFmTs6KfJ72yMm+cHoSRlePd27pM1T8CLIuV8cqcSI
M/vEcVinS1H2HdRBpgR7oSp3cOq5BN+ZQecNBEtnw4WtpVeHOLWAdt22dUaDDCHj
0kTxqudb3V9LPbtpl0vpZtJ7Jjk+AqXnxnR5my5gC0ffBMOpULrejN6iNBzcQ7v+
i6+qYyr+OwvYEW4D0ynp5WqWASWIOPma8NC9mHmzTvgeph/JKmeBFoT0I8Zfcto1
eqWnH7QtcsFtyae7m1SZuBiR0yYfgNYCyN6AmbZPDCcATa1Qf+Y9+EjMiS3xaRoS
W/pgxQTbiMUikKZMjOYtRQPVbU0WK/4pkfwMoASH+v4HQ0TuTB8csPghFzt6Xvaa
I9qu15gaVZnK7G2H+ua5Qwf5Co06sLQ8+v83nScoarvjXxHq4uCyQ5FBkPqTKd3a
PWwogcnG+GHabK2Y00GBZLUSsOGk4NwxG9Kjvri2umolbqOAFYKVNp9nVsWYAqFP
L7a7hXrQxtQOPXTqX/4xddri7C4Lo7u5oOiElGnmj78jx2he+ByJYN+oaMz+3zrY
DpedZRDsvSXvqYkeXRgXk15yHH5nxSWxAwyHHORF7AD5S6+H7gEU0tQ6piTtMCpU
5gUGQBt+bqgLfnJ1fl5cZ0WLICDa6KKuhZ5i2qghJuum/eN2+3LrOI+8raIA50s7
4P5lU4c+Q0IT2NQ7yyvYm7Hy+AStBGILKSiyl1Tbj7nEIMJ0OBVxg+yLtZi0bbfi
epKZ/MvDRKIRNWr2QuZ3Yr0ZAmxYBpD/Qi1JV5dbqQUeO0lUr/JYRW+s2PDW/ofY
Xg+tr0mkJ9IdeLZGFRQ/gVZt5RejGw0ton7jilSSWrm4XpYHzdLom7PTFzLcWFtX
U7vnrg5yULmBhV8a3cyH1fA7bgUfhAAgU7mMXNDvAHG3jZBuzpgKQbLStn7n6has
E+8kSOoiCK34aOrYAhrLU9KpoaMFfpBoSQnDxgBREedG2+no79vZttJSjekZvuFR
RjE8j8mp8uOuKZ5gFz/3TRlyQLvZShtY8pahujvx0WTgyHZ/gmzLXdbMrmzjU0Ki
BfdnZGW8mp/WRNJslnSAvjpF4LAZldbvD0s5+jap3wMB3yKDYS2Iq/VrvaGpWsz9
5PlnPh/yfy4ONiWLdxJshXqK3yx2Bd1zRrXUdbA+Vv8L2hpeved8qBp6taAGjqaj
Z2iiXUqxQsD/0DdY7xci1MzB6b7qtFLcTNLdzlWj5GX9IH96nF/bpn5w+cZ+E9tr
2hY4WktcwNcnksrteCY+O2Xe6o+goSQKjVGPgPuQna+veIER8NrS5eWmXw1o4/D7
thWPDnH2uONxgoIxr2GWqdWmjnS1KACIGr5Z8JceHLxoET9lq/MBVLVei8dZ/itI
z7xFWzxGq91cOrCY0Qzh3gUXWSmRjoW4d6FBYDNsPhDFNw96eDbXG/TLv3ABhlLf
rzE+JrVx2oOZKo2gMBPzrCdwQlJ9aQPk2Esg7lQBqh2mA21ezaVM1+e0IV/c37nL
PCRPXa1JlHIjPHQtT3JgZQIZRYlbbnAlhwaKBfotm18YUuhtxkA/CD38Nnh++SEh
2q3CUDfOeMoq1mo5Rd7mHsL6osv1w5Hoy1QwDS3Hx3BGY6eR6qlBFNGBfKqHJ6Nt
34TAoFJfGoHyEST/RCXpQhGA6cSBmRoXpR8MDn2Z2+JtJUVdUyMqAR74gvpIBX2G
d+KW3M44kw9OAdl3ur/wjywJl3quCy7IFlHXqfFMDeM4K2vTx2+SBR5sInwl4tte
9FqWGX364CsuJnoN1SaUibO+6fxT7DGaMwnACvMOPudbnJTIYec83KxIyBg6rZvf
4W6hnflgpvv0wMJ0Bk4qTXBvprmUl31udM//OvfLtHWzWvQsgqre2IGoWpBkjPwS
BIrWVggwiJfcyPtnn28mudnrVIczBHI8nyPwipo8Vo3RnKqDSdDk7yqZ/Cw5GlyK
07Nf1HbpWTvUFZ1VxHT/UixA2lnEoGHkpzU4qPQ33uoa5vL1fF/DZ4xNQHhse2Ul
cQtNQ3gKOZ2PugGUR4036g6yXxZ78PJH5ZTf/S2eB/qlHQhHEx2zaamFoQRm5wL4
JsqkNHKYaPGZSM/RGV/L4e72iHwxI0E1AOXZTcExG1mX2X6TYT320WPN4aadBgjt
31mNYINJB8to0OKIDuw+jRkBsmtT4Rfnq8ZYVGjBCIxSFu9AgGlI8DXpUa7QaF0m
YcsxyNlYAGLmFe4FJxk7iedCu6Eqqip/b0KfV/X1b8qLqEI+aG6n6vAAw4CpUF2O
ei9BcOtjKBYjTBkQJfSbkkqc08UciOYGvxVWsqk36ZYqcul1lOlj8/Ln4sB+Wu+M
hzac9THbLsRL98WfLqZaOc9Cj0v5Fswd6Y5fuXUJtSDJQrrOeSHGTuCeATfQRZ12
Ovm/+jJnkxAof62OXvYOYtBCGSBuu2AQ3Pn2kV/4ZxsOk584wZoWbowNyMBUXuDk
TI6f9T6WsZM+V+Nt5g3N+ixLjpdVh/7RGoTJ2VjBr8ZALU9xFvuse++VHRezIC5j
SUPCZI9IawgB0/tAOHSX21Oqikp92bzPqG6zZDOrym1IkLibAHfUlSuGSkQKPOn+
uDrS1Qm7aa/YeHtJKJ0FSQ==
`protect END_PROTECTED
