`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TLz7gXtTnlUuSBYMIyk3yjpA89MC55725wH1co9jCu+K0GvBqHoageiW/4XGawNF
WCuiR3ZMKLtVup4z1PyynMtviqZ7bmtjxei62CjrUdGdk5LfmTPEbg5UQa8Thr+f
OdiOqSrPwsK5ckOW2y0GXoyGSbedKXRHEvo0NLX4onuRpzaOc2JXwVSkBIM3K16a
9LerkJR7o6vyObf1X+ZuCjnFFZDQc2NRq+QrXvKXEjrw/rbUFjbsPMhNBAmz0lJs
ULgLK00kOKKVg1Bf1yo+z2cmxgxr//WpheJD1faw9uB9rHVjvvhtDcWN+f+bXH8k
85AfT5ka4R2h6oxAe/s6zCYIPlr4mK+DG4aFl+SBbF2rcZER24WUdMy6woVu3+vc
5V6nYZjSX9NwIB972GPtAyrTG8707Ve0bN7tZTbR+lNdgpdpLtFU/E76OOt3T91a
0J0QOlyoRf89t+4LevupgL8VkHmIR01mMe3hSrdosnwGOL6bjUszGzYPu5kfiAC9
YF/1Ya1ItB/0VCRdz26Hwt9Lgq6+rDDLfgAHMCxeovkIEA5ykdWg4vNxmJ9Oy2XJ
KhM8d3Z7Rfeg7LZGtuE89FZqFK6EcEWCXSjL8RaQCHXPlXKAtZWGkNOhF7RWQVOp
teB90XQo+C4ocEZMohGEf2NvW8e4e3FTJvFslSoteFU=
`protect END_PROTECTED
