`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n+azJNjsqx0q/46+NALrRBzrEp8aaNPC6CW3e1aF5OMlL+3rYDdA6FMxgZ0vw+wH
Di4AmoqVljXPI7kdZ7S9Ebgnefy8xp8QSWrfDRsCJR42KhWnVB+vqvDWpbnAexAx
Qj+aKWRCO9/aD8+jqDNWgd/VOJ7Kv6wVN6gbY9n/Em0NkuxhHbcyDy92PzE+Obdj
8E+bIdpKzFXtTTjDRomsEcP78ZclALrYnU23olAIZDnTrtTtwh+4K7Imi46xzSRv
UWPSmX5mA+Ru+3rSt6VCWpr0dM3b+8Dg07od2QuIAFUwOD9kzxt/iJ/TY20p5LMq
xVoMuu/HtDbi1ZKu1P2MFxlM5i3PohISco8NNzahrJcfmsULrPcHtl8lm4SGMGhZ
Fjra0KQ4m4M3cWI8cs7pEgB97zc3k7OJGlU6BvfBy9v/f5sPELxS/230w/GFVyfX
Ic2er0bFXt00kZoUwUxu4l0shBbCYLAkzEGmYBj1it8X2KjsjQPqQgdsHGAxb/Qq
/ZZhvX0IAKlLeosVT7QogtTs7Ns7yewHLZlerMK1KDmyYYHqZmMFaYhr1RxFlqrb
9llICO946RDCpuKbtntJbWrIgO2y9LB3OIh+JbWCNsPEL1aWVbaDnnfMCakD1OiE
ONPJD3RZshf+ffqWVBO86klEudq7QOvoJ/W2MUfdKtX+bVLjdzQok84B3I20hSC+
pBR3jvOaw+sqL5efDThzt6Bt8UUAXhxIuPxTWy1XDf1+JoCVRhTjlXHWImjEhNgQ
J2LKq7vgxUzRy6zPqlJLQPyF7tVPv81jSXCa2e1ZfVLorDb860MY0PRXc8Cz7tp2
XhmQO9kgSsYIscXq9HT85+AXl8ozFt6NwKbxyIn5pEQ0G31qbDYLB+T7yigKM6Kr
MR5GAKXFHlzooqLYxoPqHU5WDi4Q8tw2ARSqW0vHgnsz1nDZeAWv98v8h2CbqR6Z
C03wjL2ghrp+13oUJwsSuUdWZCX/eQHlLhLnMIzgKY042Kr0EDMHXr+cd3ERuSRD
P/xb9MbHTA1bc7Rbs9h0SplKBYfWFIo9M0ST4w2S4JnbGn0EdASE9oedgIGzGtym
xlcT+r/hwj9saPDP6jmteQMcWnSa6VQmwU3HezW/ZUgNGj88NYfzLdp8cr5BbQ+l
F1XHytoKksMMXL7UN5bDReX7dyK9WaShwxudsfcTRUoFADZ4Z5x2cJh4Cr9fFDm9
b5rUe1EBTTQz/6TMrdSy7SreCg5krKXstKcFomShS/0vjJKwcG0uztdAhPsqaoSQ
9E/4eu87zPb+3YBTTwTSeAOCAp5MTwa+DOLYDtt9SgiPIb04E9xlGSKvXsEQFR7I
8ztF4z1Awh87/2eLQ0TGG9TQ6q2WXxXvBtfSKOEwG21nzdicwpksPM4EWcYbvUCS
TXT/9l43CkfWhdqKptTfWbXjucNUG4kp0f3wkH6RswrDkX4AlQjF6hFtBUubTHim
AnMOP63dPNoi9gOWiaWkRfBm7e5KSPt2QtiQnPdVxBljW4V3uuPmjZyhp+1XLNmu
XCBDo40CuLOWt22NL1RGF3Q0JGs8jEa3giI3oiRHEF43w/kKzVZe/ict6FkViWgp
LHWELRQ3L7nX3jm8oixb7QqaRbqc20pi4zKvhU8oL9MwD3BX67dpBqaQlkXkxxiA
mZ14Ph/nUG0fC4pGqtJuqBqx6B9yeJRC+Q/YpwtF4H1EWacEC6ppXIApR+JhIuRt
UdKUS1WZYhnxDeb0SXaKtf3iAs9j9/uU302CgLe2syqrpbt+OJyTMQxMLr6UP8QC
Gm6W3klwNkUE4dY97xJpc7V7rL47EMvqcItpJaOyQii5wE6/F6aeWwEKu/2mkHIO
rd4TeyRR1VJZoUb3/yBG1FO93cBC72PvLfhv14Jr8fMt48pTYqEwqzAcFbdLNMR+
frVffEP5Fz1cUZQ7PxuHYpg3knNaoFOnt7D7c5k3l00VGx8YMvYAcEwL+MFvdB9V
D9LtBm/R3nHjTx627YBjzsaIFMatrs4mysSsaEHj14y8esWyqKwFKjm+jKQR1INM
BVXe49WMGs+DEcW1HKvkvr8EZlqznz+xgRwbKMy9W2ejybFeZyX7dLtl+Iuo3fXp
EcE2WDMWEdjdi9RUPK+DfaMTxZ0SCCMNVmY3JU4S/qxFxkO2vrtKaJQ+k4AoiHw6
T8FyqMFv7hCBm7KqW4hHf3CCbmBjdYdyTlSvPtnsDz5OIbyF/xpCOU+8D1+6gm9J
F9oIrZKl560KKc0hl2dm2VmgbK3QmurNLRTVximEPrVUtMRN0cJuRQJMFNm7VChF
727tsT2DwJ/JxLnMfWtBMAGZ1OH9vAyxtJRBJoMGv+BHm7Iz5HlNbwjPwHs68CJ6
iS9s775KQKeo9WBJDdMvqFgeooUrbtL09XJlBJSIZCks4CBua+gjCityxVu6FHT6
Qqn+/7sBF5Fny+xbS+qAFLC1LdU+yfk8L4IqlWZH3y4AWH5Krr8i9Q9bb0h82S5q
HxV4n3ZvD5zLsg6DFZ2heHiddqbtubX3fPXhPlRMoz6v4LGRkQd1QzJMpBa5Jzzi
kbp+lyR9STWhaQxVwKJut1iq/pHIpnpafp8goHZ0Z3aktna05Vis+anIBMTI8fOO
kxWy/54jY1nhbmvPsRYaSHxISTGym4T6Twpr+BqvNVAKzoGkZreiOArIl8M626V9
EP8CbqtPdYUcBUqIDibo3uA5Gq8n9XFcYpHW5ufZ9Mt9TXkNnvIPRKu/GD1q7OEX
E6Z3wVOkjdex/6d4x7vXCsfsMNwUlnLyQ59h8rRduzsYh0+xr8IwRDdzkyfHhZMu
D/GHMP/dxjzk4blOv//w6CkUaFwYWYMGM5D1wkzSKr7CLeQBLfxth46D0vHsb9Zj
BEbCHjmRQ3kUr6RjDPrIxQgYGcW8FHAB0AComGyrJyeeFEIJhfMOdQvISyisGAeA
vO5sSha309jjuN47SYtvoeVvZsPJwJ8pSnS9MH2NHhRI7KvXImlvWIg1MFTDzRxV
LkbND/PHYVdq/WqkCKp0h8A/Cx8iqwhG+8gf6prsT5HzFfadaf6nZexAj+q1XiPB
EJPC+pTQJPqYDMQx1IRVV6N/G6kBBNUB2WWvTNgS6Ozs5ol2Sp+SRUZdsKVQo8ZB
6LDCD8sNnruXYyu74E5Mg0xBvOVHCgdDiiapkfpcR+QG1IcvIc/bzHKl6nA8FVaN
KyItR9gCQwsrPmCtJnvTjGcIhfQ1M+IYkZeJ2DQ2mKJAsk25li1tK/be8GsSDVfq
XAWv1vS4P9ND/f57e3r4G0BmCICHJa6tu9KYBAwmaSQkphlKmRj1LOFbNbNqL3dp
ACTM11YYHqt5UoesglhAhV8aJYKVwFpva2Sf+SkY4fGQ792AkkJNdvrFh15EwOCp
YrcMueaJPQbmGNAT5tdyJZJbdZZPet5HIIF3+SaIp1JQfLpWBbfeMvlP7KR7WukB
4OKBGuFstWIU0CkGAcOB8av6+Ri9d6TNyPzxPhOG4dnpVpZxgIkkrz13PY8eZ3tJ
Anpjfje84f5v4DwAeXPsldsv5cuCh8oalYRmKvGo4puhJ7UHFzNDjNeT5PMH4qTA
Ehq6+njhWAnohzwwqjnjup5skIXG4/Sg2pzPJ5ZwUllgo720dEvn6mTVTUiBlWtk
VH0HbavszX28RSOkBBt4Gb3VDUXSOndkRjnmLtE1FCZDwSGpq4kMjliQ5R+2mNrp
kaylI7djD7Bmfx48H8l9i4hyXRVChGAEGiO5XTX0GuSdSdbn8R5n8/BfFJ2/ndoY
5zXXEQhOkUdmgwrJEgJOCHJS7ZGT6z/C2ZZPXLRv8YI7xsls+94Re3JuJE4Gc8p+
Pjl+7okLU+G0Hmt7bUf0+YJNhXacsFgzcwUuf5GwI+Sdnyf48wxnP+4lFauaXPjg
zAJNVlJQo1qKiUHvJ96K+24sRc1xNnBEVa0LEL18O43HDHkNfxElBJ1hqE6lCfWF
wu4DpI7S5rNqQe7B8eoDWrQkJOYtvg3f0+aTfdgXC2yLpN1uNJIXZZYFwa+TKkoH
FNEGrBeB+JYxS3xvSAXOVL5ULQz2N6+RQM4EEmRUdb2G4y88s4GCharhgx4GOEQm
H3YVNIj1Ix7QO+rSVwKbiPFKB5TV4QwjQW2Nvp/vdju3nxXjcpRiuQcwIPIGS0p4
U4oVx+q0QaHHIgtjZJFjF7osq9m4SeV2dNQHKvTBnteuROfmm3f1pizp3S1cpHmH
OPZ0uTCPi3OQvDK29iOU0RTFvmT47Qqc3gu1xB6YPAE1lQTbNPXPA4fQNSL8zRsY
vDeQdjsqUZhlQqMRQmvcfyDPGwGoB/gjusJJpSIpic+EmvU2f+hEEwIpuMGaqvPd
IKTE61vHYmYvdlad5XaIPAnq8V0flQcV/ZaICEhh1lC/6edjBV+5+tdGGxrIa6lx
kiPHioKV6797I9nwUDDBbK6lYnRebsOgFB/4asm+C/z4EIrBdE4VTCgy/SQJspp2
S/fGVRSDp1ssqoFWhnQmTzlUykyZcERr/QkC++2YgcGX5ZBAiTyyzvtdYzTBZxQY
ApXeXdgrY2gWEmc1cZlmZPSIVCdplIP/N8aDOZVTiZ6oOebiORbQOSrWCxcta2Td
VBbsmDFwOnYWLd8BQ5AjRCpsDHpMT01SAa3x3cLvnlkvr4+mWUmPMAifLkAopbnc
MpCjCaVN29ZMjjRm7+8NI897fQGN7U/7SMfbSYfwlYXkkgd17UPD/dVBjnipZ32e
IuGn5+LDS3NC6rIlBxM2ufyyXrVLmGTIa+B2p7VkMznEQAYsHoTJSSXICta6uAif
FXSLCYw/koK0KH/r+gMymzjgk7BflVDighfSM4imzkfol/f3c19+Kw+3T83HGGkg
eE5wwtGhhK7dj6W7ash3wkgxb611/ByEBWisn/qLIX/a295jeE1qbtSfp5DzRScb
HJdl4vR1Plj4rCT4lBmz0vwMiSbdxJW6WU9up31wuURYn/Nk5XyZnrAwNHABkCXQ
FLk6xQ0l5ENHNSCMJ/t/1+9ES8SvPZuLlnQK03pOKsDzUIXDfmjit6se+G8qpei3
FTfezTIYCyS3zModihcvYnwU6Y5a9eq+UbHCKso7z+hEMGhcIOG50jgyJ+kyyFfp
ofhDFvcVu7YXUGXko8ztmWoWaDVAr35ANR62A86nFPzYiXajj0jhG3c6/N6s6PrK
x6R/zzrm7dtVWeNwt2xl+YWCrxuJnG3hjVw6nlL1vfUl8aJ6VrvPuRxfnS8vcovo
Mti2N2DWh1if9/3WimpisVgQcmIvpOXmLSfXRW+ajlMOiffhODfK/4CO68O5nKeg
Gs0KLlm7w4JMeC6J5FdbH9wpIhIyPQR0lmGTrVc7vqrsmKKMEWCQUFJxVexFZ2tu
el1r3XMbD0HxY+lvHvwZHPl9GrpMJm83bankbY0eVApllI91aFLqPsk8T5EQSDt2
aQMA5HAZb6rX+CBUUK4dZVSw7DehDwSmArCjy+JUNEvpTGQMTxzA1p/WevAUQV0Z
IUT1sbp2krPIWMPbQpwnl83YKGByJpXoOeLkTZLDa1iuWM8aBwrbPdZXLL278amK
hMmpf3swYPdiqINPhuXhtdKx1TY/teoD1UX2eqBC1amVG+tu5mDGr9Dr9g0b5fj+
J/jGmrgJGEuc/Otjiw1x3OO0NEityhcxy4z/Cj7Sc4uJpSN76TuKKfe73U4iu17x
AaUldWeHAR8l2EstW6e+o90kFVGyK3YyMfv5Vz7gkIdGuESsjw5cIepaFnPlZ2M/
63+gyfDg5lQexWyer0ewLnyweQuXoWYz3XEJdxghAXM6q3jOEEJ4K+dHT0vptU84
pnDePfb+wj16Xqv5XUH9Nr9XtllcWvh+pvJkiwHIiBJ4ZPf/zcjqEngtteNCmswa
UiLs43ahnBStnjGmsLXHZGG5izTDTlG+zEuh2rwIC2FNi3ArO18Ucmnu9jk2Nxwj
JazllPUD75bfzgP28kziIxIoGmQSICDhsNmiGwctn6gqXS2QrZjHj65r1Jx7nnIr
qW0LU4aRqeJJXTJPXpemIlS3hUG67p7AhFlZ0ONk5zXori/8+mKFHWta7GZjbw8n
i2uVTMFCiLPcqn3pRUM5ccTi7ZFyqyrTQoNsiOSnIglzM9+e+f3aXTa2S/gaXB8E
3xRIdAN09Cm+Q0HGp62mjJd5Ug0L7/NRsXqaqNwGGqxgnRH+2aTYkEFtp9RNc+kT
fgPVV9tb3o11dv64GTz/JNOCs8tYKdqb7yN6YVenbOAC9Jw/+hDHWEl5TTjskQEd
Yi6MV7zR0qHHEqF4McZrE943mUxWnWcrBZ4eS8DxoZ+rsY6QTZwIVyTHX5N8Z4bp
CAZ3FUjjf6J1WOBFd8PpusZv6QJw+3C39Xe4M2LOXD81+znqo+yHgNp2yoQBWiIA
k/thVXdLCntb+dlrAgTxNS9v+HB93aOjoso+i3yQWMX00s9/N63xs9cfSC6u6MkY
zznyxP9eOGmNqA1zhguoxOT6wFgTAa79xkvbTrjmF6h1xBJf8suPsG+dnN0NSw3g
Vp6VmUnBgDNyLFW4UK3b2y6ujP6PM7msawY5mnjuYP/wPVyr1TGn3Uh861i/Cqgj
GE3izYWvV0GR+P0AEjYVKDoalj8hQ3Setuybs+Td0XaNy0G2JqNoacid45WVUSNQ
LipfwdeHS6ofH4C8GMmsKE0rRaI4ZyvG7ZWprykZPlU4mF26S+z2vU1LqmFfO8xE
EZpdBDcifvAlMkqukQ5ixXhGPh74sfTOzZVsIZ9etbDI928TnUOlWKdGi8slDWX6
OVDad5WNb/aX8x2WQ301kNJl2FaT0viuQ+7YU6/SmxRKTSTi1sie/3tJ95dlSYU3
vYqCUQx+ERssIQlT4J1xXEeK53Nn1vRJU+bpukAt/N4/ZTzXr22w4g04zB9pdFdL
pIADKjgPbuAblVxRYgFo4gbw+DwWuh5RLPswK+OrTU/iBJy08G62a7gOjuZjn7Sq
aL+T3SB2RDW6wFOH+IkWfzskH69qd8L6o9DPb/vxVBC5O74dtJ6t5WfkZER7VN+y
72+6qjl7EWtoYG+ajUnTvMeKiGkeAPUbj9geaOhDFJFpTPU0QMx9kpLpsu6UlMhc
P2y3zcYkQhlDFym9uSyO9/aGmhtTYUTdSA6E3hMDo+nOgkbHpCDxrTefmfuShIjh
vXz9+J8G7bUgOAT9mhYO11zm008eEha/K3MqR6d32SEjOaki/CE7QGFAMLO9j4Jn
IFBielrKaQbDpmh1LFNiAAhvcNFWVjvppmZgpqXJaJ2f/5GtE430VHe8l7hEMU60
8AEGhH9xVwvtghftLzeoqBnuIOrCK220R0Zzjp+HtQwN58j7iy4MS+qkLXW7lmJg
vmoydiGXg5PiLubgicXaWp3LxwaHy5w9tGc/Wkw3JskD+CEV5fcEszsbIQEfWuJu
IrtgMH+FTQLXu3opD3aPtwSX8o22da/02Y+mmtxQksaw1FznxYelPBDEnxhRbRZ3
dn/gsmN0d6Nod9F09Mz1OWBfmF/3giSi4OJAWE+Dg4RpGBC2LfF18dO3xJFMpQJU
+O6P77YwHDQuKf4WDUWeH2H8GfN844h44lIkMAHZH+EoBB2oFN0kYkv0AoAWjhey
Rxa0fAtbukrDm3k+87su+Nbkn0VLdDdrsGkB0CQxhxD9M9OJ/ZNRtdqRAFylZcE8
FJ/qZt4YmccKPVU+jzjOka2j7MW34IyGW+RECZmhnk55GYox4G6rQBsvoozuZjex
dJszhrGIhSCNHSieq2pNplKqVZcGhE25lAu88NPjZADEEPW5ESKVC0m8A9+oVLqd
XnITN4DR19vu7ef87AsLNshRg8fWzCpqlgOH240SKjhinSy8Oipmvg7zsjgx0zTF
7fOqP5vDIMbvmzkHSNTz35HIAKfmluyFNYeUkKPOS1zZeT3c5aL99ptmSbQfk/AW
F6WKxlgawI18JtSA9IzoKdGPtJvQVRo1HaKLZkqbzdrb52leBflLwruRBJjaIyv5
YxwvCu9t1KlaMGTe1dC0jU4MOjQLxxZTGv5e4Eqs+8g+VlniVktK2LutTZdc9/4e
FiAsyTjgiScO5+XruQXHu1ha1gcF0zWqTctVU5p+tU1XmzGrBdfb2n/M88z+nham
pTfDU9Rz4RN6EOrx/NPJxb/xDgH2UVVt/VPeKKWzU0OgJylJHLkg4ned14X8y58P
HbdNQ7eY3LJzePjUpu7fypYEiAl4BmaFcv7dh2hXVT+PhyKupAxRJDVQocklCyTq
1Q7OqVCRgRWroiYaPbGBU4TMUr+BavcZmKaceMbdLYcMtBFd9GhoXl3P4hbUXKy2
uto6VQuanMmM/kipcqQ7wXm1Sax9MvTHrJgESh9Zw1eRDCDzYH48Y77y3Z9gqMKj
/bpuuDl8AfIcUUm+a70t8cG9o3TmLlL8QBDlnDC3iKDApaxd9cbAO/fNGSPZe4qO
6aEQtrTebhdiqZrQIIPxSJtmdNC9dbyZZzPsGcYTZ5/X2M7E5u6vgxkGYTTA89lw
LnsduTomQVRcffKqmXzWZZVBuxJ1IWTdqwCfY7Cvu+GAb6IUo1OL9c/mfMVCFugx
P/lxQ7d5LxtEyMpoM2F/Gt5EI0q8ScCEG8kfXqOlRkHrBVm0SYULVnEsP86yZreu
LE6fB7f8By7WTi0OFQzA/+jlkjjLPq85o6ABs+s0/msyhX2Lr+bo9GxlKelit2uF
zTE33RfTmDRr8qtRe5m+bGl5vZrK8ifwixefWTEOIuW7Qj+z68Hu6MPAiK+sfiCG
pIHgch71WUUZ6zZ6gU3bFp2dCe6WSYAoAm80UlAv4P/JfFR8spctb5QeqSu9l2BZ
rQ1y28jDS1l857X1Rn7hlw8FiY+TV+kpefel40QGsq371nIrn3jYst1OOOqpaStE
eSVQTiEUuZThXTy2siTbX72lw9Ry21iVFNtR4mGgPXlM7bVmDmtnbNLwP/lKwP+G
sV87MtYGtQiwLeRAQoU4FYuGZkHmI3P2Bc5y+u0sWHBJj0Nh/2xZLrc7JwIXMixM
cD2CBiGsmGMS+eBUSn4aMAvEgqTQ6luI/iCjd7VoMdyUrMgV8j+TX9braS3VxhP0
uq16WeaEc+ZKpRQ6Tbcn01chggpWhpHhpddNAjC14d3L/kvoV+cE/z+zvHOQ34Hr
dqDjtfvZOfaF+t6T/mz69ZAXpnOftij2rB71DAaaE5TU5ReraAbb+2/tHoUoPKEn
zRE901rAqElPyHR6+x4aBWxKTSrpu1N/LcoWXu3aljONbxpcUJjo10JvfQub0OZR
CdbNuchR4t9MwP/3kVcYl1xqCNaJdqG410k/Dini0ErAhB0Oo+3SKxtiGJ/0xGer
SnxX53zYAil3TE4SlE3MUbMwPeL0D2ZfKQ0f442JEQW+UFuKRNFxwIJgHCqURudQ
WvaWOVoCpsQm0JmgSEnSuKINT1rhMbU1gJOsu+iJyT8J1iPBr+uJ/lpksAMOp7qN
edJ+k/T+Xrh+EiLZOCL7j7sUjkQvp54sppuk+gTBrhIr3UNOa1jVd0INRvQAuEhU
6Rx1Yrjz5sR0RSrRd4rnjhSZZMuuRMb0ZE6Js4XgO3LVZEUUAqmo/YrdlUhu1RJ0
zJgBrOu962v+mwBDengHCa7PD145DyvfFDf44wcjb5UklvqbFLRHHeWSoywfw7u0
Mzr9gmu3ghhhQdH/6/N2pi8IJRJftpyLNp2ZC+iNXGKxm6F4OfJdN2Rd+GCip3I4
bOyfb5YPSchllfMEO8s4YoCHC+IuC5XH83IwK1dhoMF8PjXnXOGIxU/wkxAyWUIo
Rzoyw18eOGO3G7yFMP7bl1ULvvlCAXUroPt2hodJ/NLJuc/yZmLXimUixRcFsVOO
NCPEEtJ3WXFMwc0Ob762E4Ze6x8qNEDhTWDozGl74hbqy4EylphqyxzMdPvoBwdB
5AiXS/cXWtfPYtUyacD3pUHiOH9d+4AMtsOIhrEa7KRs/Y7IFNzwJWlAXETLnGXc
MUArSrJt7aUezTOU7psJtWG15FKV4u73dLtF2/EESVN3ds5Y9htENRJP/qnEzuXt
a1t2Ixe1jf3NPVLA7krSd/sdlxXyOsiIIm/HZXXTKRrgCKGcAkKIj+xi31vGdbNd
8rykXvttNeZjuG3hN1zSaoyNkvhMT8Vu5BQ7yLtbg4pmiw16II4DVduIaD5QU98z
fiMXd/GZF+0LGXm1UwAGTajeZnYYeQoVI5PxqkDG8HQB04CMCaCjI3HkpmqblLbC
Se0wdrERZPXlr0KuhSA5rT84V0wWW+MiEbY3eatVqJ1T/HoD31x9vaPOVz68lc4w
ajUOtRlOw35Q+bRd5PWkA12e1GnnjI8Wa34fARZH6x1f5B+oyVR1OQUlmJ7E+iSK
KzUvj4gpwJjDAErP0p/zr1mbjOzEHUVyymL9qgVmnf/YpKexyztVxxewcpYiLTOW
snOA+n17LgYZoSWOGeKGMD41IwAbbVo47w6PYW/albCAmJLIEWaBOWkZUpdvffNP
vVoM7VeWh7trI1V0RAru7C+l6arZ2QiWXZN+aIST3KT1ue8YDR95PYiP1TIQgH79
1staX1rx84B9i96umiMUzSkiSfrAaGgt7ny0eOLigHnsONVShGkaLdA5okNUV/cH
/PqJaE/73AG9MbomZtijUUk1ANkC6kEbHgW/l/9P7WeV6WUgkycx3EEMeMqoA7in
Dp+ohMUffH69VszFitjALXmYLBkJueZS1nCvwoU4lf6K0ZvSWZsejxDmtTlST//s
eH1d10h12pVxOQF/9G9YV2O72imjasZjE29Z9b3qoNa6dNDwhOgs7bveL7vHY2lW
czGaH5JSkkIwP6OayqIuvSVEDlhJ1eXiQc7txi22dVJkepJ72Xkdz5i1jvpDVW3K
Klg7tQLrgC7TOhpzsz7/bz6LCV50V5e+dGsOptZJ31P/DE98z8oPdBTW8plOVZZW
wYNmlxJtgxHxVBCXT09pDtLVb7IRRaADAZh4lXPG+GbOZO9qOSpytoLTwafYhtZe
uLd2Ubu8ZCOm8oM3wGuaAKdHpV96oO+6sWbQG0h/xfpboPiR+EDoUQFm77mHEZ2/
qf2df27wIguFP/0BCHfTfhMTLOvKrPojZtTzuayFUtD5aboh1F1/90k3taqTz7ZE
HhReVuCPGGRpQYzxrJXN8KQoU0XhplzqssE2IjNuCdSDaEIyRj9UGOmiBgth2Ur2
0JEDsTtQC2ZtyKPDoaUpRaKt1P5gp4oD2trW8aYTHy3gqKVD3ia6QDX8Rs9ckPV9
dDj/jNIa1SDTRBFxwgCN+l/T0DrTS2CUL806+eT3Bgx2jx4gTcwtfacbbuy8HZrM
z65iM5LseIj9vmKGIXlR+iAA4aNe4Yt7DzSPe+9RUQtX2rovpdAl3jZ6FEavgPoU
Cm588s6ltiIMdlLR/Bu6jkDB5uqw5Bkgw3unBN6r397RIu70hqW8UYOE0lKFNzZM
XR3wQRfTYcOgDot1RaE7C6G85DwJB4jpXzLKmz/iawr/9h/nTRzSqXNPLf5dr4GN
MYIGQBA6PGNlKk7wV51kp1zqw7dJ380X5teu+tJMcvxj7n4+WG01w5MRoXcmgazJ
hQiUKHCVaLItFrxlid3nDcvBwNFVe74hJSMhxnM3U32dyw/5ZoTTd/VzWxADcWCT
0LQsu1x1HOK5pMYTlrZ8SlbR22bZnTMUNqP9KS32yWA2f3LqrT64Fc1a74mXsKt9
PoHu+vyzP01JxRTSxgPSlvPPfXVn05ap1ilbOjDuyWLCC3xgkoaV10xYvHNcxbVT
GhvWSVBGsYbpN07vyl1OzFSYHW1f4cQhj/yBqLghocsdYE6dveUfVYux1QA/LN5F
eNPn5IBWS0KOdW0jCAfhVYEIuBFq5KMatSUlk/Wq2djUFggRv57HP7Xkikj7axHd
Xvf8PJ4CITSYCPwgyUWTU3JhctpX9ZVhgcCcbNhEeJMFmnq/JjJ8182xNCf20KkU
SHiFJFl8AGAbbY+3i9QzdNZSJ32OMI19XhZVVLd2XVRM/yeVQsbA1R6BU88xmcQb
yQ80scwz3Qrj9mkmn32J4MbnzHrqXjox/LcQYRjp8SaKDmE5sn8mIv1qA5/x6IeX
aSNYVJmSXv1/A0KbXe7ULlvvtMDl2uu9JQwNFHJkoFf3cagpUHHPmHLmeLNaaXGn
OgdOfs6dxHRxfbWAARx8VXX2zP/86Wx8DRlcHbFtj6HnYP4nudYsxXkxShgsKfx3
J8xYbSPGbsboNPsSAtWVjBbM9hNzF2DC3a8xcUDljG4vdEUcHFnkKKqqq351JrO9
WlXPjny5j749ow/ni6EOIrZw7v7hsMVR5B32Fq40i5lJYUDC8GkVgk0Q9Ls+d3sr
ZFoAiOiwbFoJ9teNLTntnx+LbR2moWFVMZtyySZ+9UtKSvRgZGEysJrCKCK4Lycm
biR6jJAvHqIGZqwPqO9Xo8AxVPUtTlYuyzwuvpdR2uv1i37llEIOlDGQeMTKx784
UOWrXGl5+JyRDVf10zwqk7S2gHUu0SrsEDIlw0Znkt9TGxF6Z0oYHTic6l1lBsmD
CUbbuhMp9I4oBTyYn9vU59y6gy+xX0VYupvAspXFgRtTBTnd9PckSmMwUP2SiWVz
bhbtQnaz3whUZdCVehc7DO2pTHJl4SyI4bs/W3DY7RPKsUocT01noHKwvq/EP9aA
6frwqVqeUrGmDeGJB9x2m69/id/gPqMyNDN1oz43QjTMG/Pgw2qFYQvHaxJoE/Wy
8V1lrifQ0+qYfJQ7YQqi4ZgDXanqCuKZbvTb7u70GmzL5grmzBLbTn8FOlC0qkdh
y+uFnabLYaX5blz6S1UQCWL+AJdOkLuGQhXvOLn+td+nEbMPTBU58IN21l70Pczh
Y/wmNB5WipZzsKHy4BLdduGohSlc3JHasameTd20Cu925iY0+hGlqTuVVf4L4K1g
vJ3rj3vmBFtAGmdrHE4EyWBkH2g2yjapb1MFy77IU2oK6q6A9xfPkIPGWhPHero+
e3/9kO4jma4HRQJpkwbpJPVQTWPdGz1g3lyPMDA2VnkL2nfYTZHG123qUI2qaj4I
rjAPTooeMH/RxqG9Z4hLxYiwnhpIcCCjqVObnOCc0T/vKUGdAIX/TDCMOMe+okEO
D/5WrJmYaqae1KfA0BAJpHCtU+IJbiS1REsCLOSmkvq2J+zuU5+uuaz/qtRmVPSc
O2Z33oq7TPtRwU9LivPRIfAkCGHIWlDOMfTvP23ZxwiuFR/cscGlu1H+EzM2Fskp
Fqyz8JyZmRxvE3PhMJuL/aXA7LGzpddVb/CNCE3FLhMKTw07G1RixJxJIP2smf/l
wL0ElTP5BgGRwDKrOLiirKAttZkVtw/y+70nRHQXYw3/CB2ZJ5Rr5AdJpqQQSj1d
p1DKlyAwgD+k4Nl2cAO7V0mwYX0X1RcrZ/YUo9mVicYM39kQucM0wKjNBFtIMQ/u
qSCljW+9jToDK4/ML7jY0dexEEZe8tFivU109rNKtf44cHusLoPof0KTRKMbsN1/
b+Xrai9H6wrDBaUff9J5w8S4K+VgXNse7ugYdH3vwb9xdtjiERAzfcMWPhOMRCmT
mG6hure0EHFEDdWBq/d2CU2BEmj7+iJ86Vqa/LAyv6its8ruuM8sGFOBzgw0w/cu
j1+BHyKLglg384x22RgrbMmIi/DUozeBTG9AJeOzeA9wLrq5eaR9MgLTkKpSnpbt
vDkqd/bUhyKUZ48x4LXoe49TmLMtTR4ViRpvoZMgvbysNJo21Zfrha/XwDejamZy
mBmpD7dR/PvQ/oT7QEEJ6Pd/CRglDLJTOKbQ3XFheJYjH2mJ7Vqk2FbD8xHBND7Y
xI+UlydSuNwJaleF1mbvi4xyWgDL2awIWA2kUeIsgw4pfwNXlJnTyc/hrOe80+mS
fNg3E3dJhszo0Qqb5INo9o7HvZ7M+pJzSuJ2zvWk7XSmmZLo8phvPBisV2l2aR+E
XzqzsPURrd78h9l61uKP5hEtLo+AdWr2dgTfcmVB6A0sqw9lRW0R9zp6H+fSqAsT
iiTzrSHemD34MjUjmb3zqZB9W5eS/tgyMgSPBKDaiFLCFuY931jfuEFIgrEDv+Kd
QUhOjfhnqgCyHp5XyESzuNvPhMoV2QQfmTxDtoY7DaoU4SDeSP4jd/rkt8bQRBEG
shcp+pVWvw8o5TwBD6KzFVID6UWJmDMJbbepicrKtYwU/4LGy0zOcw83UkRC2uAF
F0A2CTrBhMy14IGx12CRDWVF4mctMkztRmjQu/KDeX4HlyWun9bPywTwTroIRbNq
fexRNgbdiems9eg2IshQi+AgobggbKPGmmIhzDnY0myAtsgJ4UW32xL9GTieGqLu
2rv3dffoAlhfBLWcc+LALVzHEyHdkOWdfnepsRnjLGnnXjUtRxg8O6K9hjnyyDx6
qVZbTAk16oGRjXVXpVXJoifnAh6HTk7CQyLT8SSkZ6j3R9R3ZgGAKXM7njC3KJOm
ciTnROyPx+JT3FZ7BjBYfBK0XXXlENXcJzkMeEIHxxrY/raaw+uL6uAprTtPzkPQ
DaPdTqE/ahj+VX9poc24tczdZ34ExUzs3iUwCKyfbzhZrp1/syV2B8a3HCIiOwB1
G6Bdj7lr6oVZRUkRw5qQpgkMd8PB8Jmf8br5/3JcLM5WFuu2CzuablIJEG5JVQdb
+4pZmzvWRChtAJyTa6/YlK/3ZvSbgdKKrbRTv0a+POUGTYB1g6mpKisJEITn1WGm
Hjue8OC4sn54h9RPz7r8cdz/pNW2E16wN2pscZzo40tvkfUIhRRQUscjDj4uz9h0
7xeKkxczorkcblk66ciB7v0UXaPUvdV2RJbI6/ThP3J80F777vXdZhVptPpY+++p
PT0lgyARNnh8obIlATziHJP50jEs0FRQSh3MJH26v4se+8D8pMvozGk2VpZG5Qmb
mbdz76ovWPa8W/aloMNgBpakc6uYGwTdvvVauTT4KPHVwLXOodZjWksQno64jwqy
G4Bhv6GuRIaSQ1+FbE/EHFOuAicRHL4Q1/X8e3YhP7lyUTVgWJ3WxxHVwGgomqZI
2c68/ESzK1qjQ0YKLV2+PymJ53xgWrM73W3X51UuZozcdAYqmGWFfQ9g37ohSGlB
datRZj6VUI4lD6VSGPHxKoxKlY8p4qVL7O02XsvAoLzRwsQuVooKWxC9Tp8+gkuT
5cnJFnD5h9qjF4L4pcm/UGTgC7av+9LGfUYPh8Ql+9DL9l8I9pJp71ljYkIw3pYQ
3DS4t8iDtK99hGFTfdjlQz9/hnSMSX6l78huumpVeQV5a8/IpQOtAuUMQ6jjI2uX
JgiBEoLiaoNTIFY56pMcnQl+K3Grnq6sV4vjC9uqHpJYDd8Vf9TA864Wo19vMnJQ
kJrib1eAPFjvSIG9VLsJWnpazdD6TWdBYH+wDRaMo1v8FK/oHoAVNmAEW34NZAJH
uKZ2z/LyaRqGc43SVO/c3jbiIGBCHm+gQEg/UxLKzqkMmdehyheaBZWnVT0QmfQq
HyPvfVEVUROJzaBYHqXY307jE6cyLZa8Hpx9L57C7FRoNdCSMVElbC1pwzguOvVG
Kf5QBPcQ/LbnNHMFOGJmtvUpJZY6zKZt5Koep+IV+Agcm+pkgT1/k/uyUnqXozZK
SlQk5R2t3h465KHoG+80IqpC1S3exZg81qPOIqf4kJ5rrIRm4gBUh7lGS9yPZiQM
85+EL+sSPQt2cpZw/olKuHvZqgodEtVrFGo4XH3tmyaJEzDB3JsLbos9NkRH+bcb
yJ8cfz+VS6V2+NwhWG1QKX8eO5liPEHERkCoycLpYN0MQuLWS5fLUwskK99kgjOb
bUJDBrcjgNlHRMoB9WeYZ5KhGpKLjTiuOsaqGGCxfPb4Ps3EoMRBt3Pmu2U3zz9Z
XHzYh5IvTHCMTOnrgY3j0GUlbr2VTodo9JJBLgmDa0WZGTr5uFeOXaXLpQAwFq0A
2FSb5d+sSl0OeO0xNu0Q2sJHL5qDKInn7JWSj7Zt/hqHP59OAez2PVQjRmowxKRK
YrltMP28QORYtgWPNGB/KdYpud5vuLvWKzluGd/yEokVD3GzuJxNmp5uL4VyN/z2
cRPIIevLcR1FibDhzVV90AsxuBDC06nuM+1V95weKWJoyWlPyv73Si6vG701yCGJ
trmGvrWom7apKCw2bBYWhSENb68YN4u1CL/IB2NWSc85DtytyWfCLKc2RKgWTdxG
cL2WkEP7PvH9BBACcq5pVCqQnJPtIXYgBfikvyWSZMantPoEJPg709g/FL6FubKc
5o4U98nJmqkzostb9Njbk0hBbi0J/AeDACPbcBPQFJFvyr7Kq5Qmz+m+82TnKttZ
aSgwWEDhLpZ7OY3hJPwPe+Zfh9LJt6+ohxxjbof05MQZc+2z8mMjHeWenE//r+Vl
g4m3gb84UHHXVYWR01Yc9QFYfgeH6FrPnjJvykg4gLMQvNn66kkieJclq9Q0LSKM
wif0SuOyml6f0aqDOO+ADNar3c3rd1itSGDboy8nBhMvkQ10NckJnCGALb+eP2dz
UzCZRb+i+Xa2jt7n+q5c0Dyiec4rQms6+i16jVgCwdayRYGy+Dyd9MyZmtt5yaWc
BxPdhOaqF2HCLvc7m7S1ENHA+Mh4ZNOx87sMXOFndKVjErSYg2a3uSMigYyHcbEi
5AQp1NgymI1yOgEZyupaMgxEwD5M8J6FIXIhYIPHPCSv/b/TsEgBWeRjOcOVqNH8
TtsRHvTbe9NglV1fVfot2ERvSIMBkf/HfBZWT4WJoQRPPz4jl7Ivs4/fRSU0bgNB
3eOdz1jlmfzKltzYS8PkafxMla2fPs+yQs2Wt3+KxfMXggh+umoQz4kzICdEsjkm
u7bzttVW1B+gQLUZkwrwKhgVkeSuMuzq7vsYrvqFgEU54+Zx/PoHljfL/RER4ui0
afhrc/9BI60HT2CxF7Zz5rldGAIzk39xqUGXNdVsJ9BSVyuxWqGzVlyEvVOJPt+z
8cVtmvwsgTU71DzVKXS51CCw13jzPhR2FbElU0PV5708s2vXnVT5nY4xfzIYstXd
F8A2PMemGElCVLXHssw4kkysEqEoCglq2tnn+ajH9jDU3DTZU98DGUtgD54DQpjO
7bMl58+D7TfB47gOCvKMt8pVzC1Nv/zXUJ3Og4JS8K4IoCSQRnQcNmsXBzdZBhB+
tq4ejQTmmem40e/SmjqCg92Sw9AosgyoWGlUGm2SqDct0DMuncFLyjje7uXFTRPM
zMb5Xb0R/pWpEHAg0CA8s31MmFQrg+hR/qQCpBJ5P6bH+3iCmEn//sfqH3d90xPN
eJW1aqxiX+TkgPGD4UqlrwH9P3qMtp5a3T69Dz8zdRMLn7ojbdXbyjmXT+WvN/Wv
r693xol/zqUvEb0eDtBDwMTK8P5T1C26pWVQlwohS+DdjzQ1sTrHuz9r5E44q1By
Bt9N6lgPf5zBMWXj1OVMtwUaAzKOLxlz80r4bIKzst1EkRahr4WKOD8NArDwOVYt
W9wWTeZzlh2haz8vpU3BIVy6WJzaD6sm1ctwbSQrGbYvW6xLsZe7hiqakXU/zIos
5hohDdkjD0YeXAnmdf6wPR4kay6+ZXdeeNHMrB2FuHGlrmINP2T0pDJ45nF75ENo
bkRkhn6jl+JiiUw/Ctv8yR9NMyaKAU4Uti1wLFoQPHGqbnrAxqw1Rrl8FLgzyVny
sI3fSro7909CJL2Fd77FiKHwaFk3Jk040BMeavzmzueh30xPsbS7OHDQ3DxAcD+8
vs/A8Kn/F+IPlATeJZDnMFwtJTaP/c0jbrDhKgv4suTkGyTOivsYz1VeDF/YgK5q
rlrBan01ef4E1z5ozNmu1CTojZ8esIfD4YS7wqVEouccYpRn7q0+VytSEZJncNhM
zg7o1hv8RCejTxmyvl8jAOwLq7BewmTF85wuCI+nIGqHQygP47rWfqXyKhujul87
E2aJqaKMTu9WfxpgAJiKBkE9YBfjUkm+DB7NGcgbuO4K0KKZmzFMFuP5H0OciokH
hr0lNBaeShhL14OpNIC3T/JU3qbValxttdHmMCUSEuiHBsLf/5Gu7KbOQq4o2AzF
WT1usj+/o0+h9Kl2wdTfzDx76bRQsDa0ykrmZ78hHkjl4gcxGhJCqXoRDqvsGKih
j/h2ikcaOcuN0JizJKc3Ur3Yuy7ElIKEhk1GbE+Q45t+L/V55I/gx70WGcIdQgLT
z/+B9ewHY/5YCDZ4J8VIK35X4dbjhxrSfYrdNbhIncYrKpS8YOoYAC2GIsPq6xl3
tpz92dT0RWwGvYP0KHiI/NH/AeByWXELdOGZ+8S71gwx64wzN4TnWzc/2fDBkI19
rCPntzXuZTeAWdj6D3vLMN7Y9LJQ+zu38uAkwqCGrE933oLwmG2Q462T0cUbOHPd
5lVp+7M3v+zNLIjVOR/iHFtbyBUuwJfVALBkY9qnDdR+uSbUoYrRVzgVCPAUdyVS
oh5ObrS+5bhoHKXWdPGlGy4LZB8kZoAP4hQaZxjb0ekTzIMpAom5cLxoSU4titgK
mbmLrs6Ydo2ozRI7bRw2+/AyY1VBiGMu+vBK9v3nyRXoa6YGE3eHSn23ae/nEoia
0jmHB108LLr4Yn+DbFR0QLGb304m/cMYJQUfehhwq81mWqeKLkOf2YWC88a61VMy
ykcAwmM9uOZn1iCh/STHRgG4kyognMDIHYiwhvTld1+dgL+9R3MhwDOZJKaa6EuV
VA9U0uTr968H8nOEwuVvAzt9qHXf+5WQkESa/t7SzmV9zTBWWKiipq78Yte0GCNx
G7ygEbbUwkkQpyS7Y1cmJvKJYV4m1sl/RRk0EkFkVzpJZ+W0DliClR+WVgi6RY60
suDrXd2eiGEZZuZBBEttfNu774r40iX7C6Wh71FoIi5G3/LMXaYX9x4CfEtAYAlb
M7ggn0jyRi1jVJzt79RLRzYWg2a0eGG9vzPXPSSHa9GD3M6V4pAxEwHbxphIUvch
aD6msdZ4UqccyMYmfXq9hKOLlYDEkOidYtvyurxogD7s9PmQa14Q+3K5AiTqOVW7
6X8ruf/TB4UPMRSpm5EwSsWC9S2tfljU3yxNJdl/OYa2VY5XdbqfoOwOwveF5NBZ
c2viNndxsmDXbWJ++fSQmBf2fJH6Lh6SHWphi+wWFrObouz2kWyjGTN+V2n3mHLg
aUO6K5KCOtIq0+mXzHU6kxpxbSyPowCABVoPH6g1A6dZW5sFXRR7+ks+fqugTL41
TtYFVDNg3fgjF+kH5mBSU0PKhwF10j1h014ugZv8f+gM2XHAZq/Eb3Yx6xQkmX4i
o2KiCptQ4C9WsKxGAfDPApsZrMKkJOWdwBuikHKzLlam1bHQOR/iBLS3bEPvNogZ
+taKeJDQFDImHHC6U7HlJbJGIF++IuC5A6xniwZrnUvJotfxBQWc44n+qUVqJTox
ZVGlrbGKqr8/n73vGL6IjaTyPoj3DIRO1Uz0buAKWgFgl8CZXToVKMd2wr6pTvn7
lINIygeCF2H226/hJRUCnTIjEqX/TkyDP9TeWefG0ui7S8EBhvQ6IItdovX/KmeL
lhYogCvWTGfChiGdc/D6cL9C5cax10165YquYkxVnoeMCgEIH6XMDYIPZQSuQiTU
yr1m3taO/pfFsblcvGaOcr5nzz1NiRe2VtgBdmkunhHWT32L6Y3Upm7B/FkheLsG
w51s2/MEDick6bO+Baao1ALA8/b8ey56cW3lj/ihIcUNxsDUr66mfEiH2i4CMD8J
npTIuQdCsJA6+YHUfD1fmV6Ek1KwodlwKK/6mzDNlRDcnaDavFOrobRZsV7BK4p+
ilxljVHYur4X7qo3B8ZWk7YhD9L/JB3ZpTG8TRxt4M50Erv2M7XxJXFWQyN15wPv
V8jLRbDC5Ox/RN0crgp9ZMWWoVYV1OMJG/9QYTIYkj4h0yD/zBSuIk+2+ouZlbqa
SDJgXRP61f364tALtTuPYPBaOwVM1CPzbDb2Z9gP+JFsCX7jVt0g0bU3ZaZtQEZ8
Fv2athjM9h/Ewa+28aAUVyLpG+NsX7U5BxLR4i+aJiWR0RgmYcCuVJCVIQyTK5pV
5JZ0zgiT27Y5UcnckKZxhvLn/pn3mQ4jbUw2nUoxuksSl7BL78xBRxGTBJMxAd7b
nY1fgPJae6DUz+3bP+kv+kDKA+dz6yde0vH3z2lIKQJYXTKRDIPOObABY3YFpFUf
UP2BQIjg4YUc3QHhgSYVbowRVKrjiC0ujwNsjjmK2yXtR9stGPSnG3KZ9JL/oS6u
nk4YLvqQ/7nDnI1iMXRsqMbUSMwMKTGmHv+ZjqX82My79bsRFkpBhYPEGkrf3ag+
9Sfx3LSVCPoig7QJwdzGaelw9H3zjrgptV1ZLO7QKFEbJeoKykUwI3lBnY2NL/PR
M03krEnr5/vRnGxsBvPscIkBW/powAUkMns7mqRGmohCc83oOQat/rwkG/p6hTGe
uoO2kEiCgU9YWrPgT9Y4CIFQ2I12RXraJtsf8GcLG3tEJi1qPNF94cp7aDo7lIkm
6I2ORBHEUSrm1l46RGdNaN/OvVJ6oWFh4aKPxSlGn3HR4g4caIwUyC/dQ7PEcD6s
zuaS8bpJ0UP7qYEM5bZNQjEU1DXxzchtVEDsH4eqdmr6eh286wp+sYQ7i9QQ7HNA
ZZeHrrfyUrI4+0vmxwAT6bnBUQLlijlj0MHbcKBG9t8ZwzkFN+iu2sx6v8Rkq+oX
80i91GsrPdgg7UZAxYgVtMi/oY6DC55AmBOd8QvscibaTw63Jn2OXhisw4F5yJPp
WYUoIHgg2ld6pv6gLe/GuGWAH5g16amZYk68j2vErSEvBAZ37tr1qTAfDQLo/38s
zITZTtfLmXLyB/Cgw0GNKPxkpYQLU/5ReB0bDvbyRG/q6kwxV/AWZsndJmxef/Jf
oETeakeM1bumQaDryQA02wK5iGCp8+eYlWemU0lOXF5AhBuam3A5raaDoErrs4vt
Qj0qXSo2fY+acJX1j5dAqU6JW6/qRJ+cDlkVsfU3hjI1Be7UKqwxg959CMXNnFOK
vnrOqqYomWOfKhw4RCJDrb90bmBH9F/fOYa0JH+Y2woyesEm3QlQsoGAxMdZlUcP
SFSCutMm6alaTI5L0NNMYEEDYRrqkkaH/8o/fkxsTWGwgUZT211RuM/FJsdZQDNQ
7SrA9O9MGrLMrCz4Y38F/lIQVs9eSkMgsLjyils9CA6efLOXnzxLIPdLKbyHHxCR
y5R5aZ7sU8LtJtglmVrTtojxzwV6ZpOGGv7PzV7N9+q1h2ho1DH2yNrtPXWw0Iso
8B9TubY1piwIPX07PycyqJUMwXEQlrxO+dp3DtY27jSCh9D03kPsv1esMIYJqa6P
Ex8CufyYZwqCQ/DIWBydFoEI9auL6Oax+CwXq2FzonW6DFpPvXmdb3d81k4VQROE
Lkl/2ZPPCBgLqmq23MntHLviKq8WYgjRHycqG0pN5meiCDGfiN6rLYPtFyilAic9
N1N1RW2He7kCZ7BWXwTczxAxdh1BzDlzyUywy/vAoYVQeRFW6nuT/yTIbDx8SLKl
Ewg6kOz3fXSvito0vBzKOeflVOKLZLkB9c8krLE9iG9JDrwBbjAwqIZwpZO/HOYl
AF09D91rTK6fVXlf8YBCmImLH5ndwaO2x/acew53MPWH0X4SMMpGkMy2l9aOjDh6
HpZxPve5DgkfITAY3yUUjxB5JlRys5PB+2CFzOvBxCupoLhc7Hr6MhWuvpq+lywx
Pk1LfKpB4/egMmvZ0f7gBNquroSc+LNTyOO2oOavzi4EBSTmkrFbPdtPqCVRRKiu
PUQIq0cimsvSDTh1QNyfnbByJzOP3vah9Cz0y4w9DxkJAlPEnY3T/+ngo70OoiLd
AOLiguzcYbZOirJ9fr1UKdELTQXrFxUdurashuRNYTpU5EtX278vcEKQ3QbxZbiE
gPeC0LvHw1gUfO4f+Mq1V6lStDizRa4maS7rcXAtnsOMDqyh4BHx9CHkfnL3mhkE
BYAA9NdIsnU3+VMG1EC9Ic/dJgZg06e59iOIqTtiNAhh2pWia5HTVnSr1SzaSWxk
L2PPL4PVozN6u9iODxGe104ABnRLmlcLB6CkHOKOY2VFp1fWgBDrKnOEB7M/D+M/
RyIFcHvtwzBQSEPSy+sU/5GRsTTUUzSZBcgROqMGZIWbr2XZauVLGnbvsncdPzV6
wX//uLryFE4ATN1+tJ08QfHV+7oJB+I/5u0dYZxqyqoZDkhrS+T8gFaPfPs2MMPA
ZcCeKhkov3ow9ZoSBo46DfiCSWsdG/X3dCqIDZ+yha/9T37EH1ThfWQ21zof1+pG
A2SO/RVMA6J5K4R0VgqVJhZ2+OhF3QLMj9/3N78fq57fsffWlqoiPKu8bukYIKUe
vkuGRWGXYMoDPdmRdDBXynNg8HF3lpRwt+ugYOQS0dZBQ7c4ApQdToHgqnh/UJmG
+jw37vvUO255p8L6mPASRxKZc4+ED4YjsQVa4Y/s2Edi9Beh55Os/AhCvDghYjud
cgc+2X8YuhHMt4BOGvRrSyoa/GoHxe8VupB9kFQDFX+A3BsncbGQ1uC9JJ/utbnL
zPuNsEMdW8ECDCQVRrbgPiHbh3Mw3E0NmO2HTCmHcIeeYiUP0UM0zEgo6d/Xj0of
mS814oyYZreZrR3wg1isbp7gCyRQWxJpXklje8IdRxdPsRYzmVUVl3BqY7l6oJEP
aP7K1QniyvzpdeiMrm+o0eqjW+F7lkXcCAK1lenQbuAdtzvF5ViBuuK7U5iCsNtZ
wf1k6cntvgeYC4+Qhz6XxEXlY4TasO6EILHNBySms9l9QMaZYLtKoGWKKxDB1Js8
t3asy8NLuaFlLrWcuFXJIqarfwOLX5cWbdX0MAbU+fvUJk3RwEIZqZz/1ghzXEQG
krZxYaPXddYptNu1Z3mq6S6wSgfojF1ttXb3gQtSOrcxeODounelHj1K8vTteKvu
8lkAHDRx43lmM+gs0dkIHiFyasY9qUMkDzKU+SNj3sZPIYTd6uD/ZfXLRfxiHRyH
3biNXwMbA93pVVH8c49kjBJzkEXBekGlCyoPUmbu0B+SKv0RM1XbbmH7LzJcVN7K
AVKoTdnt/LepMye9QFOiCQwhuPlkenH/gceoWnrf92fjv0zI3G/OHZcPANCLnQ8I
YgJd9e18kQqIWo+vU+IVZk5m1o8okF4E5lPTGhtF8jFh7C71bhKJO2ausQ4KDbSe
1j7Q12nGwyVhFNOAQwpjykxN4dsS4I2ONon0ZOHiejtiGhwVyjtC7FNYA9IKiDfs
WSnHHMIIE1FyU7LIBjPZCY5A1v+7Za7E0ZgnBr+eePdWlz8gndmpR+V8lui1dpkA
gDzbMNmFgNDlWXQVa6KJ4bV2XzS+ScMW1sc+ziee6Qi5seH8F+Q3Y8ZgiryYk935
rqPmpZMpzj1RdlAoNHANe+t+65lqFqZhJ05h3QK1joefj4ec1nNRUsa6ggm8iqLL
CkbsZA/22YJvlS8i8liHnUuMCCaaUlDbJJYQBWiStLucxQTZezrgenyTjek/6Rcj
R1F8cjDeazZe1GjkOzFb0MKE2chwW2G2dFiju0X3cCB9GUJ0wTMXXPB5rQdJKElS
Vp3Pb403XsI8YN7wxv7FCGzgKx4WdlMqQ6d8jXzV/lZg+PbuO4cKRJS+befCMGlW
sUBCPQkTH7PMw7WRgs5APDY0owUq8SfmTTg6jc7IyqA04FKEOyOp/O+oGZ3C2OHS
J1DTWixh/27CuhSmDW5jTCrQqsCPmNuMyoIh9bL6Ohz1bkgB8IJXAISoghH0DdDA
Ed1OBFX2fgdE2r/2vuMDFpbs3WBRypy69A3VJW7dQjYvRgiIgRC9RG8Zv1ablEAS
0hA7oClRH/rxu0ag4xd4+a8+KgTRS2hRO6Al+BuUOCFDmDAV5MmjxbpsLx2hBEJa
7USNoK5BIfbUZKpSh4L6u88KbyRMKMf6niPAuAIxXtMqAwDwqaN6ab1RSUYjZc8g
IJfbG2cccUb4TdwWEsoBikY0ae08Ljg3q/e4YeklDLLLs1whlmyVAD5wR/1Gmgc7
fFAd04FRD/nzyQVdTwTgr49dSborATGqySuLRJ1diIp2B4k6zmpslvYkMra0XeeR
439EnUWNuJMH9BPFEcfut4bZYeg4W3DwXnUvbZe+NPED2nfAvWH58G4bb1346DXG
bDOjKmEJ0gQ4WNdJcoSxwdP3VUiJ8V+5MKqvFVebgqRHiT6vI37FIqyFwb1mJcUm
FXuHiUyNvnwSj58iO6eTzU2lwTUwwYbUyo7UsFNfAcvtRGT3da1pQI2Te87Qbk1t
C4+rX2v+kMAhIjXP/lSBeXDEsMdxEGhJaolJfAguo0WrqGYxfFCa+SYfGu8GPz1N
vKexWeSYUE0viQ68tjKWA3Rya0NoDBWEYuvjzUJPTpQ7dE5juFyZ7y9QcKk3jrpK
/Oew6pQKgetsYuemdnqkiKYCHmbgtZlfFy3mdNBYGk4h2vfgLvKht9BNm6kXvV7T
Ws9Idpayh86Q+6X6aZ1rJyllK7kYHOmxv/sB/E1F4gKyFUYzQglAT75G4fmGOyJc
1PkPcBX+ZdhF5y7l7sMEbewmYBhyvEkGXZuHallOc0DLYob8IOgJH/+1ltk9Falm
9M50kGYhGhhMO5Sl3ZYryYyzkOoUNXJh1utsYCjt1Dj38tAndIvax8YwmmX5BeqZ
bujnWmudklgttyphz2jjyio1QjxtINcrKIsB/HdmUH/dIC80gK54FTXSgZ5luqjy
qWbqIcCi3QDyHuJimdE5s4/2mAmH71u1vsYK7lGMk/tkeeXz+o45UWLP692jQFde
0sc9CyolqM0tebnVtQC8MdFcr3uuAtejaou8VbXbGQxX9mF5tuiZV52VMB9IRwuT
JhDLE9XVxDL6VHNNCNGdw674ladEsli63LeK4a8I1Lvw5gSzHcwvsspz5ZA5zp9O
4bB+1rCEiCQC8dGHwAMkDa2Q0DgJYebkPqBEqSyettr+a/r3OSpNHwTrYbEidNZD
9I6bAgjaIykJJUxfQVvUKjQYlLq87WgR3ej2BoLRyYhfozW3MZ8oQkkQZHPvau2S
wl3kKPghKkFHJfwv58coXbQEjq98z0Nap/58vcE+WCnmABItJz9kUfhWHG4bsiwK
kkDxKtzB/KWBxcRKF1D3y80/Go79ax7HYq6SHhptYZvOvaMu+HBvnU1EcLQbM4o7
PbONygybDuIMWmGmzD0J43uS8NJz2bULdUmLPLLUTvyzMeLspZQC8JWtAGRNz1/T
HPAzTsM8jQ0Yufm05gvHbQXWiMWOE4D+GiBrBMoxNqwd3YSFjZDrmE1kxAmCN1XR
5z1kN5N5MPnjDYxPSAx3pPIFkWltuaY7NYyw59IYrhzdSWQsHm0qi43qATMQ6vLr
ERAjnMBszSi3VUIX1fK8EyvsQEYsHqo+0ADcOrscmjZmuv3sK926qk9eKkw2NxHX
sxYsmIo9GuQ7xr+xRxXfruBGQB2uuX685Wx+QYDAHwy8CL03a9TL0OXWbIWG1QMk
rotEfeY3h/F6u3Fd6dg4cZ8VJeX4i75HR6WXZ21P4oDsFVkQ4yk29ZGfFi3rgmMj
qFLlQozQGTrVw11OW/JzWn2mXs4J4+d4Aa+zmICjOk9kiJuXJljDkqtZvzLT9tsL
3KXGvMJ4NfHqyfa/niIHhuZqeltan9zOtGyF/VnnEqtGnx4P5+tWzJ92Tjoz/55r
mKQLAtHA/Jd40exg9bYUnAPmMECxH5dxpGneBhEM5QSz9XZ5WZQj7ZRMcfVlG0Di
pQSu5xTcgXzc6Y9FwZYYZ1R3j85Nj+DZiNvlPvPGyJ4t0D5YafXp2Wge2NRbPyQb
ZTksnUzROTaMIS07hx2GVAhb6BAa+UfDBoX7myQvZP3SgiYHifLXSDXdjbG8jwjg
LQ0CvsPbhdURdzwnJgAhjGWuNypEEYKDyWUX8PPisUM1wu7DTSDnQmy6Qt9QH/9R
7U3p91SB88S8RyywKCyp2e4Vn2xRRO4r1WQPjoRfw71Mq+OprOGr1tOKaszJXF1L
VoY1jtgtBMrrl7FToqp5Ja/YAlx7F69d1eaFEv/ZH4FNovUuUBLMGCyr17Ugo3Bx
Xt3UsHVIJfOp14f2c2xTCpdEpf9PwseCoMxDTlJIqNIhDTyUgop/ljxhjrpAJC1t
6UeMd0Et4FSWDgoKBeRgNlIFj2vRzPxNWXs+vS8drZijX4WYTUDZcYStD8u35G1R
Ti3w+Hy1E9PMOra6hCINnGxqHxODscqUJctzgUKhYUPXEgFB6/H/+amaCMCdiMru
TxnrpF0faQ/44yXRGRmhRaM25fPGm+MmmEfqKhZXaypPTidekUenCMLQBqCzntSl
3SOjc6rDM0vguH6F1KO/5WhKDpwJUI2dlKHUDkY/ax/jQvYq5+S2opyxk8urDTn0
ycJU38YQ9puUFeqME+wqDHTI2eVx/KBZQPRSVY8EjcyPsTElkt7Q74PhM2fTmtH5
n0YR+bkdLCsecx+cV1SGqWpL9cjRkKQxYWqA5qjcpIoHZwnYsGyIyY9CPZ3mtZe+
WAjwjgMzXhvT8C8jdOgZ6Mr0mB0tstj7XIClXYmguUtb3EOcbQ+ZuOSVbwAMk+V1
ri7x4Ys8EmsA3YNvrGctQtsCP1p8111Ehae6sVtZXS6Epm+ok3Y0KcgGrlVTNaK0
9L9Z96gxwZuM/uzS/jFytwjQIILKxLik37TmoOysvmpjLViEd8FJ1mR4FZEVHptg
130/+FLz+/vjzYygxbjEyZoV5zcNX5TZGzzmaCRLF1sx2AUXlggsm7e7xOJpMlSr
BQ8TO3IIdp9bzmr+w8hIfX9GeUhrLvencRAEAeIWN8PpAWM7HwD2FCv3Sp1WsZty
BpBIbQaBpD0Bm3RGdYBSKUW1PHffBNp9/cIVL/+ytliBkmfMYCJ9qrBbK7IlEx0u
JS9iIbJDTpglMkAfDKgyvfHOmdWIZm3SSY+fyZN4vKDe1YYaSRA9EACICSB4nvZM
HSYhhfuHJicVuueeVL2efGtO+GMMKFX4BzHjC+wZ76m5K0a46N8PFyPQmnqKBUl6
b1wDpc3vEE3zo1nb06a9nahPvnjMDyBKshA7BFBWGf5mWNcEO6mcbwEJ/pigIPDU
4JHHgeq2QGQXNkNQpesh+K1lFCV1GprmYU0gFKgwtPGB97qmeywc4MD+v6O1x8kx
SjFlxbTzF1FxER2KLTSMXUfhjezCFWC3nM6L2x1j5f/K8wTa9MLxxRR8R595D1YS
ShGdCtyU6bQrn8iaoLpJaIToYkbWKSt/VJKJ5yqsS16nekTUonpTwjqJVWK9XOWV
inWxwMu2kR/1Ufd5OL4ewmNSa8lF+pNid5spEfaGmOg4HR9OrAMvRMIK25RxeJAO
BoZZXOEjhzhS256AlI3g1Curnu+agg4rKZEIrMCTL4u6DTX/a49KfU2p2CeiJ3tB
ChTtr4jdKoOAudJs/O9iwkECXfBLcPmRA1ToxrCy/G+WTc/A02hDjWOr0azBx2Ov
n57NdlhGtLWWTShy/dJdSq7S4mvTCgda1KU+51h2dffjHFoti7Nb7u4j1KIume3c
wATPeOtibTDZb/RJs39YmXGlPelmVwBaqG7+7dYL3a+s9aYgbVGmyKVCC0QnF2/H
XS8WuXYg1qhd/dGCfcfHVMGzyLP1r0rkNIc925soTZurMIrGV4D9lY8xElZF+M0R
gtBVR4Ul9KU8fbRlppwYHhlLDFuviONCtLcnDejCRnAKSfKHzK9XaQoAv8EjzChJ
JPK5jqcXxHr8pv6tw3nOXhvWKmgYqkct2hU+7H1emkRM2V8x2h0KhQA+kIzuL9e9
TEjM6AML4gHp1RkoLVV+osqb8SATCsmnFxwuEK5jDTbEMiwnlrxTI+cE2W03dvV9
/yN/XHpJoCvXJqqxoJ/DWUVrz8EU3OIL/GifQqYIIATgVquDZ2y/f8XXI06+k8G+
7meh+4/CiGU/j7Cd1GEtilJOLW8EDxs6fMuG/fht7RQxWnOYxnZGmMuhW6nwio8p
wEM37zOk3YqaWHKqnpxbMdq4s1A9F+PP9vx+lHRJi5iXhnz6RfQkMdb+PAOQoC5R
JTgDePFa0C7WLiNUH23W6Ue5K87Hd88NCTXuF2Dzf4NRoq302SPTVe3WkmcpNhvY
HSGb7/twPn3+W4Xq1Y7jtQjepJpySebB2jWaHUr5JahkWx8r9x3DdLePkRpQznfG
mASusfllgmT2n7rdp5qI51KRgnFby75nu7uEbiymNC2qjfu0n7wRHECTx26LeT3z
0ef3gEkZ0iwt+7+Iu6QPJIf4VjDhqcQEhkdR1JiZLR1whOw7t60CKD+Wiq4NL9iJ
QLITwfGQB169htSHCsEZwyY0JbsOWwQlZsZ2Wf03iBHiuiihXEtuLJw+9r9kKo9D
nKnJH8gMv/GLp4y5EKZs73xFFFBQ60Z/lIjlbxl4xbA/3u8nFbi5YefsZQ+JKY0M
IjJpIjjUElZcPZdik37/lei0LNbygth38CEan/z9dZs3TGtHJJxI1SnbG+Fpt1Ug
Lv/0RtxzZR9L6vKl5KLK+kb/w2ZEL0EYQTxJK+Gm986ictP8xx4jq+SFL87kpnit
QbLlKw4O+HH/Dk1tfL2EvCNpEy5XkV4LOesbepS6Fl0CZlA+Sp4Rn0kQNGyDd66j
rAvPV5KUs6lciGovnPYc2FnrtKbxvpTfKRsKdOQ4naSafXgPMQywqDIpZB3+z9wW
FXaCW2WUTzY7PkqIlTu8J0WGua9MzJ5y65ez7kgSRxRXVpS4WUnkqi2Ww0915DU6
dzOTK5gTOuZrggzEDhvMmUc0hT1kn8fEoJshKPAPsU7hwxTrdohStdww4ChM/iM2
qxSCOvLajkZZp3zIqWDhxUm/B2xuelEonxDOCAK9Y6ZxLb3Sa23VH+l2DfG85RwA
tafskHq6LX29P+/fs52IKgAzi2MsF0wIsDMDSrNFXaEi/6nISaPvj08j7kTHR4X3
UMyuyjodNm56VMKd5KWj7S4sXCCk5gRT4GG9sj8lmYQe2FQjoCy57kUxx7jUmS3/
T1ypWRv9qqZGTyflWNqtNgBJBAl3yBw3Y0oGZZMeQElIgqqHpHmIDCDWOjFW0K1h
XcE1v6D9enrSlgAbdQWh7V2ymYlqBWZVJ5F18iaXk1wMYKqnLz1LA1LGNbDRClAv
NsQAsdYawlPqlbKkkosBxHJhdJ43HKgrEfxBPvS93vb5lzHorvfyBeAZ8Qfmif0j
Rv3mi90riuu07E1uCHDVq4KAGbsxEv0kPBnLOS4ygyCTFet8hzamE/PZKwb7xSlv
mp87xHGvdrK+BGa2G0JuMLjy1fvzJcmLmEfL4QKOPFYPGO4R+wTRY8vCYzaBvCLs
qVRg+9W/79Cb2LFq9w+ONFrWtytfbtpgerjDyB3yhoyYNM0gtYySj4UIHs8Oev15
zZ6zab+AgnCfycBQPUEWg9tUDSHzLvgAWQ+XzZglT8cBHZXjzX8+pnN3gLlxhpV2
hrjAlSSYglKWkSB0ySBwoWSZ3fpx+wiOWf3v0qHDNanihFDTOinlGU2GPASNerne
g8vvvc6H+93A4X+9T7CnkQJNzBvCvJyE+9cj/VZhBeme3XwMn3im/QWJAtym0xqY
DeOc+mc6UkOODj/s4kpVxFkP2VKTvsXL3iPfqYrOl7IzTLkeRwbGHY8ad5awI1F8
nLYQ3mcMqLGyEFDfvD7zE5HNOonDbutHsGvAhYQTXgYTC5XuvnLnSXwjAsJR4LsS
xZkALDG2Qkhe3bskOmLlSJJ6Fvs9dpgAzfbqjlXwi8YEa7UGSugNpbVPHOjuOgG3
4yg7LYE0jyp/y1sBs+Vu/wgBBySTDVpkIaRU9q26CfzUIhGSO7KxugXD4c7vhs5+
MM3uBP4bvFuH+TNtCWA8fT/ju+rDhnS35saaI4YQ1gzMtsfrKTxe/sBpPFbOibQL
KaZYbzAZY9WTk2aLKk7ArdiY4UcZrOY6Gcf5nLFdw5q23QNRFCIBYnK/xfk88qsq
dl8N7QgsJ42a29t2t3wrQj1Z7Z2p5OuX2mQ+GRWMLDJ/XqXYBKjl1KmXdgUZZGNC
h9ruEGP0XmqURUeG90MQwOuFaqja/9dJBfDXq/g91+lkdDLwQhvvs4z674zs0m3Z
wIvaXxQ3lf6EPbajRb4BUrslyqHwGR+RmslODcYQy2VOyPx9QjiCqj8l7myf2Mjd
ffDbtaMjzMF4mJfYnHyt1tBSeaj6KJyhtkWk7Qlf/llW0WxroNBPkdXPOhGqoYQD
U5tUyKRpwiahpLeeUfGRJctv9byd/Ns06yAZj/Q/sbCnHBWN339fcFle+eSonsJ6
vGI3XOSCm89Qemrb3ivijopTVtq4B22Fou2kIil/yXObiQwHnoxkC6NXxDXf3cgx
lOrHvQxG6DAvjRcevP3InYLdTiJPnyWsnYB5Q9dv1txDrwVm3DOXYNZFcWOxYnzp
V2zksc8zBHw1KknBktutLKwH0eb6jGyqdZAWY1X8bqZ1kqd9BthwYlJ5wch1cp9G
SWdAbYTgkOz6g6z6sdTwLNNz3plJLcVSFi8rC1qwCyro40BZ6eGnsziInnq4DhxG
cN8ibsw0Vt4bHMdkQQEX4GM5PRgVPBcTAtGLYAuRzBNOas2OAXiPnEhY+Cvn4/wW
9za6Kl479sAYDfLm9amaaLt3K3EYgdM/IFYMx9QIjjAZM1W5K8ugKuevEzb5al0H
4YIMQdTKPDm+HnJgK1aNrVHbWjZlmzHiVvHhzOaEMGAmpf4qOlC3SySN1l1sCwRM
VDe6bEEA0BVucOB6tn8YkHvcccQGYgnt1VsSmtl9hDt/n/TgdOaGA6kLrVH8Wcnu
oj/lJ7i1ql/UHoqHwsYjWunJ9tBw3JG32joIe15OLxlQUXSvNVMDTdVvRZvhL0wp
kbmM70MRLkl0+/qfCYaj+S+cTm2/1LU4ODVJelQMOqe8JycNAiqzoc6V2qE8IYx4
H+Nwlq82Kv6KWZQFMT20SJadlLf7eDwZcT0be5SsodOOtksS4hpIhX0lvrP317GB
P7ACqTaDhZAbXkbxPe/5ao3MG7uxHrN4EBeYIG04BAm/tmLKTNsA8sc0A1OwRmDt
m3mJYgk0CAtn2JBShNCeXT9uSWh4OPzwzXODslHYjWPpWZAyD3TYczjWrzh2Ykgl
mcT3clk6IHOS51vv4xIY1kthaYEEiACg0GhKhfYT8vYN8JslbQQdIEFzUza28Rjb
L/AeUsotwA1xKvEHtmaXX6OzAeSHamqJLiA/GdHfRLr4y6rU8/IbyVq/MMwBSYUx
NGqqJFEYqoAzQBLkRx+Sqg5DKcx6SUmwWzUaeU8tLyqRUPGb+j4nUyNFujjQx5Hi
vBAdDpG4By6OfkKjXSI69zydZ8UyEE1XUVsulizeZIfwihtW3lanoMlh/pCDwiCp
oKquu8ZTl1+LZkRUGCeCzWutsza1QbbA1velq8sXlDbK6fgz5mW/l/Wmk9eHYf0i
dsN6Jf0I4wTJrg7F5j9YV6Li3oAzY+YQXPlZ7tYb+KnoOsNbaCZE26ZdUurb5h8Q
T1n92NVKKj9ID8PwRiXIUWg9CLGeXj2vxoWBeyP6NsWEEoynaviQDyIGVUSSaxl6
a0SjaoVK8e6LLKLuIWUWsZLXNZf8oh/NCxeWGf1lnuF5RxiqdHZZN/4fu6cqQ5Qj
PT5bypLE+KXddMhsksLcvAxYulne/kv45NxvqKor8W8rzL/a8eYILNoX4R88PiO8
kp4Syo8gHHkLlWlzwjPPaQCfhS6y/4ICr1ysH5/ABJhArgRR5aC8Lc3JaHiPO1Uf
3on8AjN6Cev2MkPTRx96Jb1s8oVY/28zUtQvvxwfxBZGCTQ4GMLOAifOnqzFVU6D
xti1HIegdNc5AKXI24MpS17LTI+nM3cNP/2x98/jyEwEyZ36nH/fV+2F+WIyUFIn
cezkgb62vxNBuDyLzoJNoKQOhJg555ENz47tggBHkVweFLRcNIDWNcR3MoWNtRLe
dzJRedjQYkymPp6wp1sbIleUd+0ZPgTfhvhYaU1dnt+SGpAFDRgyrbRCr+1Ki6HO
fczxAAjvbzWiYK0eyCZzQPYGmdhheekiEJ/kcxjdgMJPHNqT/S8rJmS8qqU44UPR
RhIUCpVgpEOxOs8Rsr9JXtTT0QfgjdrLQWSeEPPOgloaXE75iR+CdY+acP/+AMJS
3e2REPNFM6Y9Lngrkgzcrl5nbnXB6//coycjYkQniL/zEEFwFkf8SwjLxLPYbX1i
yiyECLIxn74rPCiSh4bT7SAFY8yojNWAyq6IcIaUdpvsHuLHJmZ0huEheuChusPP
kw0e3g3RCT7MvE5Alp/vWrcXEps5ax7GwMRxA88RW96qD3GSxn8XD6adp2j2IB2t
vIngBWY8ash/PY9bx6mwnL9JwVJ/M/qRTo+gOVOW8RtcfbZHLwPDTr3dJWit57Yn
JKkdIXIwUYXwa+vNd8OXpsSAuzV4cKOU1VZl0i+/5j8QCVqiQrwcrtdcDisS8l33
ickx7+bhkB71SroYh9ju/z9T991KKOX6gd4Zr91sLiBeA6HuE7S0b+6sBhJ3+Bdi
himojAcb63pNryhfMviKxf81xmNj//xpguHnYQnozp6XqO7q0Djbd3TtslgBPFU6
/hELHp2yxhK4zcKneZzjzP80JDQKwlD1nxP/z8Jw6BQhUueswFxQqKL2TkNaHi3z
cjYy/1bNLf+VSfVoL7Q3tDr3pvwhKbrSLjEX+zEKPyCD1buQqvtsrsry5+lYw24+
fhyFNKX3x/bCoWflReazk3wL7pNlywhd7HT/pJsH8I/s6ajPFoWj4YN+2AEXmDKd
BtpvCW8Fvs72GXlCpeZ3imyGU+ZZ5qUfaehba9UyL1Ye1cq5WmW+UrvTLG8RgtXs
AKxeeBJ6sSRoizntxv1KoXuR4z7dDWg12XTp3k0c+q9tBQlbhK2B8xylLPjxFtKE
8APxUkWpdKaDpYRPXdv89hlxJghicqJ9FIKvDsjY2t1Y/cyk5n7sBb6jAUJ8Aw7C
Gdbh0UCcgRQdyUEqm2zkG1nTQy0nxMZpt0bhwp9maFCbUOqZT+yHndChIwMBwRgK
fl3SLay89WD5XAr13tbZb9qQnColay1WPUkniD7a7BhOSrYce5EtrHzp3RBX0dQl
6uBaucQds2cE2e4I2bDr80VcAE4cAKlTeIRgoEJVdHkMwtI9jb5mIe5O84XrDVf4
aseV/vvdCJJKXqZZZvrmVAGn0yfb5ijOvPqqxZUxkkz+2b+2RmRxv50hKG5a2jhi
zJd7qjxOZ46bHotioalplRDweVReM03moRXnIlXdVR73ANcOevKRoJ4KnkikUpsE
++savPBdIiCJOkX0TENvxqz9qemb3vkqdBqKbsGmksiETU1dFQtS1pilE7EeThlq
g55jpF23xAhIG3ddebgS2kaw9fMPMlzqImVurlKPeDPi4Yy/MLtHiGQcQDw50eTK
B07baX7hgMIpH9pmhOHGHzmg3B78p8LplCriVBdid8sgT7DKCSsF7ncovRqOei18
RBcsU/3DCGBtEigcU/Yh4DG+zIyOVGacm8Qe6DIWGWHvGXkWviMwiTLFax697HcM
ZMdfq/rMa1TZFrhNc6SiXIYlTi71iOXnU+9RNHk36o9Bp6UJdPlqNz0OsfGEcy9E
YE20yYeynrZfyqxDM9FAUSXDp6giKqiW7Lh2CZixyPwQZIzChFDf+HIEF0et70Z9
iZMoVW93QbtwrGb3z+WKp6VYxP6O8Oz70vKWXac0SxwpX90tnDJYjw3wimAiY/Fr
mhtYrvghAi6IPPmeRsiFr5crWk1/CnvT1VHjzInPeMtumexksKt/Ue0WgPvS9QZV
IxlM5bk6zKyODTrlk6c37Q+dVmZ34PNjIB8rtY7a+5k8119+3PLSJoc+vFRb3zmY
FzZTEnWfA6V0tlomnc3re/5TApYi/ayinTGyj0tjwcHGBK6YJiqfbDM6DUN+WjSn
vx1E1l00f9onFCyeHXNvA3dH8aykZ9ZyndLFaN4W6gQuGz/6mdaUAI0OYepEMU5j
HoJ8ZLMAGBXBDQqJ9qaEuYJUWXI+Z87REBl7Un0FutKCusr0cJ5g+mnXJHiFL/0t
ex45YlvsWCsY9P7rydZUQUXvWJmg5yULEAepcOMZ0CyBqRJxBm0mJo2JDMRXlvtZ
yYQ2MS3WXJI1jbowwpQo5uVptMxrOnx7flTgTr4lB/nf2nYdTypooHm4UYcCZhMy
Cl1OElYI/JDHIHMlWd9Jqk17kETZHHXxJRjcZUlATq0M+WJU9dJdUUOU0Sw2ToN5
+Q4ASejusmEXEIe/0ShCv0J6qqhxcHtvL1N0HxvJVdBtOoA8kyD0YRwFq8cGF34L
ekvcv34eqVARfl4F7EWQWJOF026hKvSK06H6YpHbwbjjDXqGwIuVYdSIoj0IBB5J
cMVZQaSN9zfv7SsOFupldAC6r2xu/Z8+lXewLnJuOFKcmFy5NfhLZvc1whjdw+pP
xrQR7z1W+QdVO5nTHtla7xjfmBJOBvA3mzxy3JxRu74bDKYK+lRpaWmkrRqgm6EQ
DBOkTe513AgLttShvuwm74pRNSRo3OeVbkdoIdLj4rZsePGjyMVK7JQ85TS2j1mx
/nrZn9wmlgjMe0KeV2edfcSSNXcicwgjHC/QqXPw4Y/wTD4M6jTTwdoAz8IGQUxy
tk9Ee6yps8i5PyUo0PoyA8Bxe2j50KUpAkChpX5VSr36Z7ADjkOry0Q7yWZUbRui
LoZg5bfk/pYXoqAjKrF8TazWNuiv/HdGMV7LMNiujRogEKcGx2Rb4dXWvCted2TB
R5zndm7YL5jsBxti3weWLSbO90AFT5tYYi9Os5ZxceL6ga1fSrgjRWs4qaUC2hLq
zIV4Y2npS0DZBCsc65fHryCLShDK23ErXnbtalqeOWpzH9eaSBheXhqXl3D8JZP8
spudCv8CdXK4WsH/+5Eq3EF0c60Pbs8r2jewmiS2XYvEj3YxE2Y5IiuUSqOU964t
EVJcViEi5vYhUoR30OqOw3i6DqGvlltf/b6hquW3vuK8HNz65rtNMnHkjCKfzZdr
ZNvg6uQLtB/16BDQxFDMxMxk8qTQDkWJe4OFZ/asI9VBwGX47DeD5Yx4m9mQfuMa
90nA5IzClE+v/upR5KfLMfbSQYQ6DBf745eASa3FIuN9PEDq6cgBGmAGRI0/gW1G
WDJe98Q39tbyy5Vs9N4NBWY341d9G/S7/8Jg1Yx/Eb+0suQSWMzulQNrSVyCPADi
ameElFKxRCBKQOxUVUfxsWwgClK2jq/GFkXYh2jS2BTRIqBQx6PUx7i63Bw3+6XC
ACiB9z52oVt5tRS7DAAjPMSdPYIwSYAEB0ZxVJK2NpTLsI+RSKVfe56kB6CMNyld
REPFY7fEVJdT0ktLsS9u4pMJUTxeiKbuQUXR7dy1cd7f2lahQysWqqd0ueOxm/R0
INvLV8jJlqbtENKBHJx1f92WXi62Yy2DwFThwiOT6f0rpCixuK/3vemmYGVfeO/i
ceL+BQn5AFWKeTFgKLJYpUHbdCM1eG2SEUDCNhE0rhn8RGr2DCj/9zT2JB7KZ98K
im3CXqM6D2tIsgGLGFAKMOwnOwvsGEx+yjqLvk1/DGaDwWXcU8T1ltdIjgPM9l2L
xXbHvVZepaMvmnUchADMwrRGkc/DRu117hgew/QuMTrIimUE9UHVBgpfn3LaA4iD
IqZCqAYYXBiDadLMBKdc54eLvbDNNIRRbLB5zJ+tB/Coqly+uDsLSZLplpGH1Xbq
PNEuLrNZtXDMCDqwbi+9HcMUIwKGNAQureMJCEH4n4ktNd+t7Cxcf+DSmkYVGAce
IMb5zGrGRuK64CjDpFXTrX0SzGsc/s5qEooyT59vl/tjKyPG2yQv/++Bv7l6cvok
tMsxyoGfzFkMJPcX4myaJu0n7UNoK5TLndi1G8mdKu3GmthyX+GjnvEBr8qkRivG
LP9MoMgM2azuKkzSxTRaDMn28wezorB6JIolIcD/Y7VjDGD20PTmnr6D1lTbGHNc
aZ2/PJl2ONbnTb/H7yBlm+GUSMhohjHrD5i8fTS5TTwmymBcBuHZnUzHKMZe5XOF
2Yta2Bm0E023eb1QhpYRuKVojNWXXEqMAzvC/cTYLukVPe+d3Er6KkYjjxq45Ey5
YGJteh8u93aMYiWyjPsWBTnpzx7SS2LGiOQN9I/EQeFcRgx5YRo1JadVZsRDBZ4t
FRcg596ERrJ2WnRFUC8pkFlP40RgEosNkDq6AodstorNsrNpBSQVtXeTUXfecudA
GGaGp587LyAR7N8Lanv4QAFIIJWZqlPLuG4dn5QE5Z4FQzD5jj/Y2bACNDmynXzx
iQ6ZHchK6wmJG8EAy9vqVIVrZU73JQzxHu7iQug34fX0cYcrnNRcZ7phKzDtM8S+
vOXfD93j2qaV3y9ro4T5673opLYPZDWsoSEl7zutntRbEMhE7IoCXRv5/iICfYWW
ZObLnHOPZqouObXE4vC+JOWsKXU0JVk+A8NWJfbyOFnFMvGBzxRZ8rabRKJYLO6F
vUC6x/BFiZsHjJRlQEXNaS7F4mXLsQ+yJr3fvPnaNIJqW+j0YNP4tzhEQQDefb83
BIPbciasQpxzeZAZ770Ygw220RsTiAopmZ0aybBWd0mE65kAXiMLBbYc3RQNfDLn
RYyNM5AWSHac56cLywjyLHADCZWu2w2sUHwZdwld47iMroDIsN7OhBAOWBU1f2Nu
+7d5P0cOwaRzvbNlwnvi8zUA52NJpGG7w9rGFjCKzfifueGkO4tm7+k/+wOCP1VK
AFrmbYeMfaJYtA+sX3uiQQAVYuH93PGV6jL+MCp1uSoGB2gqZegaBt4m0+MZhN4I
UTnu3F4v+qkcFdbwH9UFgbGmsfSyPs5/yetuBHBj9CyIddey3lwkB+8OTc8vcXG3
+ngwRDY+mCAXtRJQmTEeMdHn6oxkZ5UFz6w1gSc6zumbEPL3eZw+n4X5wVe8E/TV
NyA/o8mqGlCnStEYpIKVuJDshkeioZUOmk0ZacD7gJdH0UiBGQ/pQHRpbWUObuFR
olggdqpaHdPDeIEyv8Sr9FTElV5g1TXFFBggRmtoJ0SSPcnq29pyIWozZR1H8Ft6
73hG3p220BpWSv7cuUNoJgF8EbAdwUL+LB3CjEPFy7mq3Z8nJnu4a0+ytaZ+EpqT
2R/GsgLlK3KFxfSxELXM8gVzUu0WkLjxeRNiNVFvOjq98KFTeHiaIhR1DDWKOZ0S
Iq07nfzAuInsTRIZ82L9H7cM0LZCxXLNGrK4+QMUyRN9DSOY+QQc6CMGYJrjikLf
AsRewowsMckdxTHHihcwpOp2Ud9jxAjJS0oFR7YXb9LXrrnEJ/HkaANlXOc5eZ+e
bfyzRSkOFUUH9iTUElcM1G/p8hfn+CftLNo7pUwE99aCmY7cvoFZAOBiyVYunH2K
m61ua+QCxncb31LsmnuLIod6UglSbts+WI1VJAlUSJayrvvGk9dpfuYynMWEppat
GNmoSCxgJoUQ6x/cNhW8y+yG80FBMZFMLf1Y35jEehADaUqeEU9tIr5uPQNqL24g
442wKPbNGayve2eMcvmTeHpnvCP0MmEQelTqwA/uoNoJLEkLcIeqE3DdHrZOccJ1
4ZJYEGin7Ony6AZC3l5hm4i99MFXWu7+ZjqBzXP0ekjHb7pODhgXTHMkg64fxGkc
9xRs9iKN98lpx19oxw058E3cHH9ORU1+bF5Sv0n3rfUUHQtYCQmZUyyQXC7zOfOB
6OxiAppymbpWJlVc7UpIR/FLKoV/5h56Vk4AysO94n8nPKRuhPP9MeT0SesrcGOR
Jb6/db/upu4+l0yBrCKZVfALBffjrZZJoDucthtg9lLT0W2fa4BtPwWe1KgUopZV
pH4GT6QIiJzi2xBxFnIeTg8U4+pKm1l4/x3528bii6w754EGpKRfjeznmDZ8Brlm
erE6YciOq8A6udFKC5juykdDhlDbzhdEbjg8WcOJr+MaKXEmDlQ6/RrdFi2dME8H
V10atMRVNFjyXOcRWQYXP+O4ChOAj01Lu3jLobUpuKVl1c/6nh+FN37KeLpYd+z7
sB5cVqFlaa/HfnVNEgdTRg6+cmj/aGqMATRfIhE1uqpCwZw+Go995txfAHWxFrbe
RWfkHfvQ7gkZp1kDNSefFURX1HxvFK01h+ZlCNVB1L78WTNRGQViem6gQ/cZeinS
aldquKh6K/rh1CMhVdo+jQTXoyz43gVehY7TCX5CxfWXRUNvGSLE/Oo5UPU6mvM8
gK5pa3UCHKZ2o2qpfiOIxsgh00nxzxOFq5lPzfY3ARyJWcV296V41ZYNNLFHSRw2
spnD2G7z5Ds97HXiQUIhBtDu5ls9gGVVNljfvITA3vTJs6Wp/6J9oxGUGZ++tV+3
5+EhWyIPxbfWm198oc41Q8OwzjAXwO65uo+IBRBAjF8+4oavO91YRQ/0gvm6xU8t
T1p+DhKKFHiPA1ovgvzLNg12nrRU+YpjSy93Iv+Eh1MVDZRx/KJy012vj5FarL6Q
T3DRLFH1D6IXWS+ACplVAT3NFw8Rd7DCcZD16hp4EcY9Eq2PKHw8qHGBm05blvu+
DcmsU6N8YzakA7NGC2nj+osBsVGvwQMFoyq6kTPvKVhwhYIFgC+MAuRAZyI5ty9s
21lnLjOR2bq4ij+oLcBYj8r8oktmQS5v79xkbmj9oVqvKgFjyw/X3vLXGGNbTk9h
K+dyTELlFQyY2/eAVPB8S3a+Lb5NkHvCsVlIBmRUGXYmWyqtgAjcgtVhL/gjXiiX
rfv+bNHgx8mIigykH2uok729nr+oyuEfHKva/WS5GKQJgtVwRHDFP1mF47XfdgVH
BP1ONrRXLxBnl2WibIt4zQty1EaoysFLFkp2BMGvlwuhkthgD4ViU3H7tSKcuFsh
/dG1ZxJHjrkEVeorQXIcQdhTu9ZpVZ4ZpA9rWINoWTvSRv2gutpV64aSxiGks2zY
F77c0Ho5kiZxTx7ZlFrXjC+zpk29oR4lbRNvHAZc5AQrOcDakDmo5C8IvSKB1fgU
KQ/kIZ+KkBD6NoKDmFaFRq+xQr1lTAcKRLoQMhFn5QJv8hnOl0SsvTZLYe7KuFbu
3NyCPGeUAvUANClDTwlYb2seBVuKN6jYJkR9ASegT6QrfxwX5NM27nIxOGquCB31
lvZydZzGh2cEmvxl1VI1pkkRZwKEeHxz0jPmhhWBej2XSE+ghn52LW/2U+1jJCuP
tRb8etHy3M8v6hUgIqAvt+ctbj76g3gjBdRQ7Ml9TsjyedU75dXbnrI8yp55Jk0y
0hf8tKDEG4lMTMiuiYdQhRBys5xxDTo+2Ju58NimolSydmIptbAb2MW4tqjaJIkf
to8PMQeadYGKfucgL2HC/ZSQVwSeOgbwhTqeXY11++lU4ms4UbkG3h2FvuGDgggg
GlYAjpJek4eDSISHMWxvriUQlgW4CIqujdP9hjAHF7pUCptzJKR3mwmbiXvREn9g
dqGL5GPs7SsCCWSUvDSpEFWfy0Ne0Snc/x5EmYfezHpFyeyF6iAOAbvlkrgzTD6G
yfpmbHkIGzZojN1vPClgHt908Lv5SMGjkxQWOCrhRCrXEGQKSjp44oI7WkuUDlVp
76okFZzR0fgP4aa9/wGHo/GPPVTmepeHQTyrxo3c1bkF3KrrWDX79wwydzGljkoq
a68iHEYjl8TvHgW78m6E/leq/xssQIqgGUCAslTk38rXsahZyUgbpio0fcAThYu7
M6PkSkh8N9Q1rJkZmu9e3BDhVJJItaVwyoozbzdsYQtfHMbXw8yiUOzr28B+HZy9
7SoxcZhBMzuejq3t7qvK1GL2XVUanpxKb7HOS3ZhY31FWqT83uaWVSHIzwuGWlO1
QeFyALS8iIn/O+DEw4PQ4BbtYWR25UrvE9ArlmRmer43cf6gwswJ3sWP4C4tJN9q
triKMphOSBqZ4tPSCvapLAUYJFJ/ctPPQPy6tD0SZ+WbUCM4hjWsLH0RYF2ZPfg+
LulfAkER16Q7OwCUehicuPQqn2MX9aDBVrrBHd/2L2t1MtvoCqvVH0vb8Groai35
dBUUX+5RGou4KX2uSp3c/MKUmtf+WB6zQdFkjkpYUMcMXw2WE0x3/LGN2M1qeJ0u
PSvqmgaQvXAADOOJtyuvT40jo/eEkw7AU5uV/pyYu1J9nHUyb/vsdyUoaxbCqRPQ
zaq88irjRetqecfs59S/agXlF+6+JTzfB01bJQ0Q0S4YVEEFov3xRQUeopPJdQ/K
WAWA13MZrpCiCNOivY1bDsFKCdrKIleZIJo+DfDiz1o6cRSfuevn1Y0Y7WWiG+ac
bIP+WaMW9WaNBZK6dILE47jiPVCg13u1H5H8CzwFyfltRxd74eiJGiC4YAuuJ9Zq
DudQbVyv082hoG7TqddFuI76b4dy4Ea5FpPBc5cmfwBXpiFNYJG3ZqGIJbaZPM5C
h1Xcs3ITqdHCywpuq5FneXxDWvhE8aavuFZ2ATuBNq9R0DXxcJD0C7SFtFKE6FkD
zWtS3HIslqiBooX8px+3VSoH41t1n5CK03KTefeJ42ja57uLuasZ4h1wyyrRuMm0
DNPfDQY8SK4gN76Zl3Huoa0Im/o7LuWIjjeZkkYgy2PrGPEqQ2TkOiEMi2nNpC6U
CNh6mzoZTyHs4pIdTZ2d5mXSqWhiSd7IAJV0+7WLg2QI0a4XWj1hmSNazxojOyRF
5/TocNoB36hrGOGDnyRx4mpbNCYk4+AN1bgwgR26f8mNwzM0wrhUBzyhE02mAvTm
/CGLmGBsnGa+A1Rllz7+k6HqyiYa24OJYlvzoBixet8AF8byL6KaH5iUcCkqLJuV
uwI/t+Rd1kBLqdTkKg/+cJGSzJhJahvrewDPy/+xmpLzo+7m6sOjpotCl5e8WDtN
yTuA79DF/aYHkO2S8gVJ5TAelxMY8oPkL8yPnI4U0GTQzmCeV+FgZSqdfPmxNBFe
A/17S9XsUDhd4t3PQ6OEdCr0VNKZnwqFueQj5DeJBS2lWBMT/n/qQhW8S5He7Ma4
kh7gcjrNZ1n0jmCqABivKYUDkdJt7FygBqV1zDTIPeJwSGMwQas60GCovQhKs40A
aKOeA5r6agUt6eeKBdkAJuWjVUXLkT7Iz0bORKbQuqXipZQsl2eJkQIt9LDUHRqO
ydQRJ1dSkS+SGsGcZLaaOLprRtLkZZ759fdoiWCwAzuv6M3eZv47TobZAsUu44Ad
SZTU2EC9t9IYQ8Sr675G3Afq5DKzbTJAunmWvRETapdjZIIA1+Wlja6uuyhVNDhg
HMadnZ6ezJ3Ou617szYN9y7eVvur4MNT6spSYcAfCmN6xNbUkHwBkifzI96tm0hb
Tru77sdcXXyNyeiW2drwYlazAvSwILmLKDIE4yMrgqEzgZ1fpM12Qik8PG50iieg
hmUvX0Pv4llou6PIxlpHKqhtnOwcHxyPAxGyCcP6EOsAALTsrU4qagRq6KbKD79r
BGaTyzo2b4kgYaO2vy9kH31WONL8aIA/5T1z+j08Hvz71/p87QHElDXRfSyAHIbD
SWS8wQELteO/ZgsQFCz/YqzEP3aRPGFQL6BZq+VfNzEyPTnw7jwlbquvhajFYKvW
DHG6E4tlDQWL5kPfvv/H7aaWJBdGro3+Bvk4+nLhZStA+T364/bwNlpTayQA0tnF
ygQR3Awrf538GY6sRmBy0wSXfNndxD35ggylJiRJ32oO3ZhnHnky1+P3zFYa1sQu
4vGeL7UdyhEuSms1myudlmtI6p+9E7Qnws1vqLVXQtSKxt5/EJTP8NritMMwUN6x
BODXr6DqvrW7OIGkpp6OjuhYMSDusya8BOLyRXY1Ur9YdPJVe1ctZsMWB9hEengS
ItQXxwSej/UIvnwkJg9X4XcQJlz/EvV+32HU7jGFry8HoOl30RGGHwlB/RDUVa8X
rHdcUQjj8AD0dNmHW4wFz7t7UpWvJ0GLobeOu0r+3qaMLOgs3DR6917mRneRRMQj
bBWsNR6p81b84OlD7xKSJwT1G3QjBUpLwtauRXJxN28amyYJb+2p51TYD0xqwt4p
csjqgFZ51F3/0lQagtr7lhpayRr22wUm1ry4KuFQ4Hxm+njRN0Su89hRfM0XoA05
jPG7BkwInQMiCZ2OUswNw1Oz8s3IO7XYFok1jh7rw4xq+Ry2XZj+z1nSFfdTYTfj
NDVLoNbO5rk+ojhJYme+dUpqKOi2RMsXAhJN6P+2W1ExtCdIGYIbsP70Zb8Z0/Mw
bYAKcHmy/tH3jYZRhexXuR7TekYJjI/3Yw1P5bklkz2gSdm8+ATwJ+0X3R9pEsWf
gb+d2NsyjsBk7ph/Y4FJLSCptbauEN5hlQXuihBtcZjZ4zKuEMUyD//FL3s5xQS9
+uc+aC11zc/S5e6xjxoyxc2t0JPIHu70pXnB07zaXvjrthNxJ2SoWLGiieVxmZ/o
twymmfMOjvQoWu9iTa5m9KkFMqAphZ3CqUztaHoq+oLR0LJgZK8hI8AL0LU2Iqoa
H7+o3e874MViyuxo/7zKwsnBhfJY1E/ef2BJiRQZj4u+5bmCxnFRazm7VpaiuyTF
Fk1869NowP6cZtJh8rgUpOWZVDr6H5L55bocg9H3R1fURzF8eebPpk0xSuZvv1Sl
EotaVkEWDax+l/qVRCz7We/UqkNZEDStIB2y/3xP0gGZ7wbn8pXd0z+kXuz+Rtd+
ZYQU8DuBX+xPrGE5YHheSidG/njrgtHqPhCMgVdycjBwzDlzofbdJbhaejhqMU7d
9+OvC711Jz6y2+dpPY//UO6wemEHUrAtS8zRCUOh2pKw42qlppgQj/irtVgdvJj9
APW809razqO3rWbLiqkZidHG+6sJRoYNzDADJ9yNFbk5H3x4OS/ZZ78kheMCV0+z
4tMukg1fss2j2+BCVEEwAkQu5ZNsguTY+f6kWpcJUz7M5MYEUY8GE7nnR2nywcz4
IBQWSP7igYdRPL2+C8WZFewDlRns724esvBFXAl7jaKNJTBVTgF6RqLTYeM0a1wy
+OcvFlAMqGLSgJy6wpVitEoK7B3I3G7JCn0kytmABb0bsRa3Bw7uOhRs3U4Nxjkq
p+2/1EK24U8K6zkUKKDZMjQRu2obK2SLM42WTHGdSgq/B1esbGeq5e7nuk/a9/0W
Gg5wrPiNMumq7ovDLoY+JMkZqtMOZEH+7/RuC6Rr/cDFv00TNN3At7vt/OnyQuXS
GhD4GjC5dOnLp/igERf/igyXW2bY/3tSLgCb/LAJ0RFWNWtuSzR68y3t3r1h4fRp
LtHfpkoVeDdlFfUnyOMTf37MUP328BI4+Ke503xlSHb0/21iVEnKasBmWODIpf2T
tO3fCOuJMMVcZj+MBIvzrdWEpuJ69ZMxJ+rkxKAjBVh0kpN144DTaekTtlx5oWmo
CHpcr+ye6PgdKshaXlSuC3U9VDq5nqPOpjCCmGiTtUxOaVjKxUSZlgCQso06TSDK
/X0AB/7S/AsNaygS8UIYuy9le1cae+XuKHPpw6enR3Py6CEX33l8bjv4XMyIgSJS
h9yQ1QD++45SLoWqDzaz0MzwJiEQ7Rn550DeOSfLN5qDvomwmRfE6bRA4aeF2Egc
zhttodrIVRHxOPM0homAewSoxO4FsK1fOBQYQ3Mj6FKYhfkPzYjh8D0nq4NTqIP0
tdp8AYhpmiQHctnsUfd+U64bsG2ZiSC1qxnwLU+I/jHjNvaqQ0lGnN3lDAUrti5Y
aVMR9fdhKjbXwRKJQ9sCPFFrH5IzkecmLirZ4JJKxaSBAvOiIBqnTso6cGrREmik
I9A2fznokKm3eKxw55NCBMGSRgAQqsSNN6m++o8nZumIpp1UN51tKivcW2B0xW7S
s8jEJQbsxz0biEzZjVlztfFhKGojL7UzJrpCEXz8zvuTB1H+OSxo+Beh0szSzamE
3N/kyVyVsVPhiR/rL4Gf1dqAeVS9nhMkH2b3ISnAyC/Ep0Nqq717IiOmUSEIvsgQ
FlyrghYsiQYIZbARiS0LoYM1QZiC/BFwRzpo8G2GgN2Qisul7dkL9UDkQkd40Wfk
y9ND9PnJ4979+OEEcmSC96UTC/MUktIDEGohZ3g+26zs/7b/IgVV5fE2zlLMryZc
GeQeMEpF271vCRuLnnK0s7jlFQdry/w0UmtAGdkf+vr1gwm8+fjHdtqZ8OG51JfO
LzKFebWrLf9R9pwWfMu4+OMgvOPmlbda8ulUNioelozXeNmCXAxvSmLk1XK2vBbs
vIUfvotUtdS4Pc1QkjpgM+t9sdJktjyBPyYyVccuuIEuXkkuw8oubx2eh7ea80Jk
6wg/WZlNkh/xPdGvReRgNImcA4jRhEMuk+eIl8TcbOggo1DdWRWcxZPxgNQTTJxD
aabjHjLyxDlZcKDOEfKa/HWejA2i3Zc5ZCXQHxaeVCtzWxNUy/n8NFcm4HICC1GW
bI6ud/sVnrUhnMvPMb3Sag3UM7X37/J5JVZdbleiz7li1DiDpcdIdK4x32XKUsWh
FIfxoUm9dj1WMPPGzfbZZxFPihCRr0ZbUEd9hJx0gLvm1nYcxG43p76tV3I26T3l
Ghl8V3NslnwdH0TuCxFZlwP7Qc2WuTBuMSBCUTKg8yOkuU3z3bIY2j2AI3nlWFX4
jS/H3U7lY3D+GU76AvtujSi9KYsmNGwMi6ivsMMFTHBqV5+zsK2ycn06E4F3MPRj
FTIIajuKI4JMx2jo9G4J6WR/516+1j+95AyT/HqEC8HT72IfmYjmSkIF5X/0iCXg
jEOw/il4t4SmSiJqcgwEFX1xMXe+gg41ju0PuhvFnFXtUUTpq5EQAOcmUmBlZYHC
2v/VFajUYxUR68pmC0LMg8YImIOufwLEw5l/nGP4kg7eNe9gFq19jIYphrkdu7dB
MiHYa5KRs4N4+NBlSPxBYgb4HQ5bfWqA+0BlsnJtpIiTN6kO7ZDd84jW4/orQs66
9Ql4P+rVaeHsyApD6By4Tf4wd+HD4hX5q6w30BdnqJTv7YzeV7/99L+oTLv3vH2Q
DH0omK3k0nmRyYJch5tzFxWh2JxGraZyV9ZCKc9A4YCNMZFDMJwCE/4t1JKRhArm
OhWczd/9U+6KEK30WxqpGSD3XOuJcAjpScjvMDE8dJUkry/2DaCfJ0myR+oC6HW5
zkrcK34d6p7vzH5VvVF7UbWkmG4laZUxhKWsZsT4q9VwHbnXolry1r4NwvL3zBv5
iwGkUzpJZEDOjO0T1pJAwODI3yUYb2X0w2ZESALnBVBbvTv9oa676T0LCWu+Jp5U
AMg4OA334gq0LcQctOjRzEHlcDwqTjeuQPw5F7EiCmBJfyjB1vbeI3RgBbFEbXWE
SGriDSlhvkaoHI3reh0fz8r1sJuVCgVRMY82Z9+dX4caIctAPbFNqZsqtyiU6yqe
KAs6mmrkueYpNTkG2aBruiraBheG+EJasp7pMF7xwgH9tj264LEmvjVuiun2IMoH
ppSqVx64X4rP96wqwA0smLS7XWscdT1VsKYqZsIziwnvDznlqhHBbdavPDDHiqKn
0gJj+9yL5M8oc9vQXr62sk4oFoeupdcJjdp9L7J8jMkHxgZxl+giukb6SXAVnLUK
6qgaEn5npv9XRhboAFyoy9fDV1tMsBIeXftnynGug5KeT5gKoFXI+5smX678shiq
nyrVa5Pd0Im4OUljqCVyeVw5X/T1DkwDT9pz+gBd6sPLnH+jZWwGqLlKuvyJB8Tc
aycGy2R3M3S0ZOey9Fhq8LsZXS12rkuFZqAS/KQ6Jvy2trQWrhBGVHuW+j6wWqSP
8PKJs6k+f25QzQ0O+kqed+wnwefwYdc/XWmchDgD2YKVD7MpLbe3Y/Y99CDuoK/6
kkvB45yVI3pk8KDXMxXTIlp4vbUf3zM0b3U2ukNCdH4Roc3sOfcQfiqTyoAyNv/9
BSFoJn7CnBDZNW3rXbM0tOxrSB7+VQv3NePWjxF59AYvNWXDjUBxh5ILhHN2U0sr
iQoApb/UCNzVRjuEn7ERcSj4YQEl2k/iTLsjprI2dtX2CZOej+kh4qcaKg/2bflL
iYS4tPfl6s+ilvlnKr2LmkweXEMAd7y9O05nCZUxedClBjjmUE8RFU9oA/tR4DC8
rWT559cpODWm6i+XOnpPufJxV+JsbdTsitw66kCqET9/23RKiAyPAUz1LUDZ0VoF
mO0Iz3L5vMUAUMvicgr342jDEMWoHSHvRAkQQj2egl29IfVCwC9FlrtsLsWl8vna
8L1CievdeYv4wXUxQjZ0SgGTBy5RtUdYqMWK9T+dfcxp7STUMyI7KplYQbsK4tb0
6xM9eY1VidDGA0qjr3u/9nmL3H/BYOrdC/vFjSVhWRRjoV8s4ImRQrxg2M6RLMeg
1GV9Mrt2W5F55iWmZIUI3mf2Go9L7AWiFQoyRqIreq/gefmKtLvqtCwKB4EzbfHC
WTXW2J+D+n4hu4w+UxQntet1koYOd+npOvbI5xRotfmbhkIOCZIeaAy/WEtTaXWd
epCQHQleyMMr6nSVYvm77Kn61yWikvJ4UxlLjpg0vGjmrO/xMvsXBf3isdWPcIId
Xd6qxMc5UhZ7swQ2I7JVHhib5vOdIl6o6B44DH+6K7wJx8fY37yKjf7M/sTllNql
kopJuABluLGoXuLtBqNiDcAc+dVZnPOeATOOecA9chUrwMLdFJCmpvjGtmh823XE
Hxrm94UU2SKEbLjDIYSx5s1/9YmmCD2hShdoar+evL958uI/98wKQv2pOBGZ/PGB
8khTIX2IZlqeKo8Qi7gfeqF4RyV1IDsMOjwxd3/U7+HksqLcGIzZsBaebU6Uim5c
LGKiUplXQw/5DVpJxaECuhsP/rk4pjzc/hbewqld1wsFgj7QuuFdF36cx+MWipVp
/UGn3PHhJqVKz3ZpivS6MaJOdIWPk/fq4L1RE2OUnm5rM+wd2RPO7FK2AKX6GYZ2
JS7c0X053+4KDXEysbqYNuXj8IbPc92/LJiRkDTzhVcYiZuTkbm/WimydeU9Vrib
+PVN4Nu+IKODUgU+XrRi/KKe6bNX4V1MtRf6/MwwpWz8IWA9PZHZCxVUHFOwx3Nd
5RBw6AE8McNKpHFCHWhsU79JAZWKpEN2X+DnOzp0pEv6Shw9MF0nlAX+iCbigHPL
tZL03nhRXYaU9d1XXVXx80tEcXqUeX3oreYbEVDScG2NgjBt1cg2h+SSY2Y70niy
EysbtJlzvD3EQmYhGseugXdjVjuUawamKF/pNPczSV8XUHl5lBmkPaFSZSntegeD
MDMsRmjyk1NglmjJrDlo/ZEmRcmNhyBwU9kHPCCY/EcK+GyvktEtMcSI6TPfy48H
xgGZpi4Mexi351LA7FKZoqBFR++Z2axdNXNNqLzjoAVbdAwK2ZAnfu5PC66KlSwm
zb1M+48vY+tnlonqVkz38uxxjnopWWJHjtMAEC9lbkoXS3haMr4s8lWEUISLuNUM
qR/WZ936eEthRoveYjhq4JW7s0JQwqCSqMbGTjtmuaIa4t2c+GxEeMgnEaeEW4DO
Ng7WECsiOcQTDjzoGx+++h00kRLQ0fbJNt4Hs6ZblmtgRX314c3uxkvUjGbEpOcc
BI2WEEc9ua7sjcICUzD8dfpxz1MsZkUD/SZZnGshfr2esdoHL5XTsu44NQbQ/pFy
SM4CYWZvCmggSNfIbRdXOsRjYCl+99fSZwUm128+FjP5ti6gWzRmFaEbGhbslak8
8t8GsfP49CURDfr3kD0h10jhNYFA7yO6JhqZJh4+xsrjD7RP/NLsxmM5EzvOlNhe
YTZssc4lJ+RhfB/r9pfio0neizK8VdNWK8URgrdONhqtIkuy1eUytjc4m0MFOIT+
TBaK+kCluZXzKwSJhrk6hz8jCf7N/eSJcXe2XR+HySR4qRrLiQVjioBasUqdGt/v
pR9acgnIRbHvrBEyK2XSLlrEua2LcXrIcY8jtYgjrIhVk2IB7CfNXRiD7zuVzTWO
i+Uu4LHBlcAVCKTjcpdcOjFW4H8vdtqpFVopb/P1DOmGVP6OgwczrJ4PF557CVw7
4aI7v4iog7LFOA9Hrzb+FsMu7e2C8Ee9PdzBqkzL30YBIyFp88GMrcTU0I8sRFtH
GnPW8PkRKt8k42ybCCcoCOg9Iz6S/d09ghh1dzKFUIwBCRHHcQ3Vhm1TsiINWFD6
+Fj80z2tdU9FANxTw4DHZXqvyNjc/MDMD4VUwke8LEMdswsdtNZu1GZ5uHDwXAw0
Q9xnh/o2wmuz+jzpLB2uUHMphtVySOq1KUusZ2ghaupPu4z7sR7+v8NZGbECswYt
2MwKd4WjnjFe74SvQvb/qUQ1to4BP0KhVRt0Nf5qPlAumOETfQYyWJrSN5hcIVl+
gkTbEc88EUEPW0c0d9RN+RxIAMgkE2rwQ98s48Sy9M3IfAi/OOSSLKgXHnQOCvca
keVfmwnmLeKPpnr6Zfab9dI2Sy8y3OEFRW+Vu0WhoVEqo0YLeYjgVEab7Vpwc36H
lPqeGDFrudT1dXFUI3h8WR8zkyJJ4n2THTQm4ZrD1hXrmh8cxnQn72iYrY1ly+tM
SyESg+x/Ydm7a/L9RrZ5oNoSDxfDtREr3Mk3ix3NZIeUHU8JHAjoL8Zw5ovzIb3c
n33kRu1HTmJvovrPesYpg2lh3E5Ii5Jm/8WBRbB2roOXcAg0QE5ozcG7sO5szPzA
qAj2hNV2Ud/03r1EFKnagemjvhhkxhJDNQg7A3NvuRqLykem33WvcZCxqAmq+R0r
RY2K9vJKI7IQGddyo5fcHwWj3MfXvnutV1XgcivHOrBYNzBW8SB7R/c/mD9lUI8N
7Hqy9XMcbfXaYT7qVyUcGgw0aMZkBaOiWByAga5yaERiviBn/Pjkrlm+2SC0dt4c
7vsRY4jdb9jyvTQ5SEkeRAvhuzbfLpOYkitczyyxjRJ3rnN+YvQnvYVUfX3qLKz5
eth/ls9CWpc0X2eLe5OfoZC7/VwxrMwgNHGHMO/2WJij7PbF4+oD1+8vXa5eiSvL
e50WGr1VSsp8mYHSIX39FotmcC8KOgUKf5+IqRe/iBWL9bab302Z5p6LmtDB0foK
HRSHR00aJqm4G0Ou3ACxqy+d0LUh+JuBxt4x9KEXR2YxycQy7KGSXFCYT6/GgrgQ
uwfwRYOzRuKOSANNC2/JODeOax4LBsW0HXfjkKxBEoitbIhtJlRAxhGDqjC4ohLW
lx0UyDkxaQsb8x4Jb0aIS+BL0kTKrQOZLqCrudRV2xarp9VbwUWVEFfLgz7r7PTf
J2X7v/dOGokLcH0wlN5Y2tXXfsYD4UD9duzaKQ/0e/zJbpjCF6btH3wNDYs8jblD
URh0dquWoMwQfNb/hDcddVwtXhnRCeaVx+qgBri/dkauwJwEE00yLTnmJR2JWIFk
QM0nkl2WsWfGyJYlrF+iUYeCMCjFcIpdY4l9VJJD7GwBYnNY+AAfPX1wLk+jHUqA
cGPBqSAfENgdEnlZZeLa+ZbwoTK+nRbVnSuatoW6UHgka5S6LYUbUT9FfTjS/I4W
rx85epowmCdQusNpN4n5XwQrEF6KHrjPEOBs6kGEqEDU9UBK9juMI9Pvi6wrK20d
7kwtWinZanqaOcVs3ejMTj/Yfip7O1OWKdv6TsLQJolOoEaV4yB4QsDsWEVMN8vg
Q1DIJSt3hrrn/TwkUCFU3Iz5RwC1WAjC83yPkd3wHMf9RRe7fX/nRVxV9x/l+gO0
YBQQmmPud8+NL6nW0f8KwMpfcVmPzwbBrRqAwrd4Zhz7CeUNvs5EcGlyUsr2Ogu5
6KEW4PDjl+fhzs1l1eF6knJYZwiR0pECSUCJ0GNsa1JxGYd5pUR1g6w9lQoPH62H
I+R96S9lhpM6Vmr0pVXmTfQdL/Faa05+cPN8FYs2PsKl2lnCe7n144khAvYpBqrI
LF+uiAK0UJOodmyVICIf2Zcspk/q8GHQjYJtvoM45fCYop8CEMWipk0Tbj/Pphcl
hDL0d1TgJeayl3UcyhSmHlkIQx3DC6TBB1zecqm2fw6aJUaOtbLkI5gQMYI8QId0
1ulS4JJjrgU0hgFvm7mC6wroQM2aUr8219WD2EvzQTlUddGWrQh8eAxkb8Hb9ee/
ZjeSG8MIu9YiTa57KLP5HJOgDC4sjWPM/6KsQT7pB0PeNT3C3t8/s+ndxP+u7KtZ
79h4aep+HLY7Q8Jk+4K/lcK92h7qWdgxo7A0jzt6x8GSyNlb9j2Cv7RMBR8cx6UP
X23JVLB7ITF8vqe/WpSGKwxYjBfUH4N38LxRPhnwjn7jl4gr2MtvpU4zdL2q+A0p
8K6ENSfVGqDr/3TtBHyKHjpIKHzFPPb7uyATKFebe5nVqvPzV5U4KPBAJg+hYeWa
Gd44X4UPp9QDKQX4qu+0gVScBMg7ZSfi60L5S02uxVpvWQmYTDJlZiBR9L2327AX
DFb6yGGLa/EzPuVCB9nmQHpEy8nJNju+YKCr6aqIkB64K4cmfDw9EYh7JZcdb4ot
ir+Aqy2xGRimvPEm8B1IO86/1VM9igqvKQMJiXpLxPrcBocLsEYj6Ehu8SqBSFWk
mQflxywMtOzsZ6+mtQaF2nxtQDcouThzKK20DGx+IZ4ZXed9NiUDFcPfg6qAl9Vv
pT7Y5Zc45DyS6pQ+qhThf7kdHMi8JFt2DP97xipUr47lwQrgaC1D2MKc+9CG07FX
Acuje6w3Bg0xs4GTpdAmOhUzRs6ZqIXDyFbbRB+uE2/lMBRnrqijeS7ke8/7znqG
CJApMFyZSf/4uL738JMkdJAvWWNIgTpq8JpzYQm9sEM+trnZgfElG8Mw5h0KDJrG
Scxj5w8SSeO6YGqcBnxIfhgFj9QrfuLVdeVvxb0E/NvSGzjYAxSXZGUWUo+FsA8D
TLMXgLRUBh/C5rrpSPssri038s/YO9AK9w1vBwfg6TdJutUmtrgB7KI6c1Q6Ri2M
mxRGQ1J6SIuJAuVjck+R5h7LF+ql019Tr8XjRxtQQy09zcPJT4TvnbPrHcl68I9z
9FubsOWvBHR9NMUhxEXB+R3Tcb4oaM0IoiJSajp1noJxGKVjtSVoN5cmLbCHEWxg
t7SQVda5m8hCBzIbbuEfr87wkS1arWk2XCk+CSF5Qc9EgJNNQo6MdvSboYGJB1QF
e7x3NCkvGD6wZbS9vFM+8h6h/vg4vxitySJoEibUeAN5zgt3FHH72p/Do55OGT9v
knyQBN13pbdwVZvzY5j6ClpFxGPowBZ4YwAfKswgOVBU94zIrKxNlWsz0vidWkuj
PA5p15euO67igf3MHU9LDr/C9svngCkU3j8blN8h+NnZpjkBZbn+Yue8F5hXAjF/
opW+LIMYrs0AQd8pJKM4DbkEs3s4wCm1/nxlXZSlaCjyRwQH+HDTwd3Th57pV6P1
30Q4cUZ2U9gRzt/8iwAF+V9+X+naGLCGS2y32dcFSa5UbTzK3v0YUdpopCbtDi47
F5dwzvOWdDWcZTR4fNF/ACIX/pMDL2YzkYsQL9rhK3VDtjIcugGFQQobPDGs98Zo
+MAYoByk2dcw6rYCbsPXp4LYzwPwlvd2PjOSXWMMolRagq8Wr583w4YcPTra+wOZ
5JYFyUXK4RwStOZJ8eI+68s3YIifTRfCgVeiY/oC6wZaRq0WIe4gVmmRtwrhT2qr
p6vGtYOn7/J49n3/gh/qG9lnI/GELGf6chbo7yWGQclswOPJzswh2QMqx8vx07ZZ
9psPypQiA+GbrpHUxLlB5pk1xUhJMsRd2sWxx317wS64dNKvpMw9fb21X++m7K60
WyaBVQ/+5Q+f+tVbfSkgMhRKlyFcxzWxwJX4NSggd6X7qICPe/Wa8J3ouXUGeQv9
X+i1BnOd+WBGrV47A3UjnhfI56vLoooJ1lDnVdJpVtXD/pjF+YlW2U4azinae0FY
YqqoW3IJMVwOV1QM138tLR6oKSN4OP2SzaLzh0Bxzimdn5n9CWFzJq5ADIAMpDfb
B2d3ygyjWuTwUdmrQ+aXty1WsDD+/GwsigIpZNYnNb7AsrmyYdcoxIImW3UowxW8
gMqsIIXehdPyPj5o4i9F4lsC1qKcUT3+gta1FvfRszj5RdoNk4L59tikA+GE0J4n
mX1TPMNu7Qsi6OWeQBJff0VAwxCZ8/ty54OYTJmB8TszvptgXxnvSQfQH32V8CPn
w+T+fZBcwbuSF7u6CH3ze400KGEfD4E59juudp73huu+SMijXbl9vKbmAVrewV/s
T8cL6bLZWckcGe2Syo0mG2vfoGwMvFnbsiE1RiS2/LGBcmFkFGfyp4gZ1DZDk5Oj
kBhkyxKrQ2uiAIZtOq7o6nNfaYZ4w869g2mYWs3BHgkOUWDqvUZy8O0W4vfJY1kO
KA0omnSLcQK44hh9AnOS4e1KmTjl34WKKTEcDORf0qfe0lHtcIckP+Y+Q4byyghZ
iRjj98pCjqolnD1iCafrUXjox6DOBVPHaJ6S3WtNYiqnmJ2s/+2RhG5YuYIPcLOV
Yu7Po5coA0Sck1zmKDI18miBNt2l0KxJ9LKF6FQnD6/zvrugqhUazN6Vn65iZs9f
jGbJvCG4rfzR+GZBUtIARUhQ6zDlGNrT+qcD43MysvRxNGOQOLJVPcrnVgs2rc+V
GCcNjJHyHR3WlIR5E5udUvc0ziFB8sIeZYi7ng3cBLOMcnRH4GP0XPUoelVn+03+
mUoP/RAR7BMMte9xA2kLE204Jg/kqL6IahsKoA6VSVwblMFNWptdahK5Z3AYtmDm
DisHQ0zoLhV3YGuZ9/ZN+YslVcXLTtYa73In+zdQHNPPbWiYxl3fw2lUnoOqosB0
xpTZ8Qb4puu4l6ZmbOl377zBcoftC7zMkEFAJ6ZmUU04iwmBQ+e2HhepYt5zFs/R
JOkow196GCFf1COEyp0wb3URY7gcw2KwfKubWsZaLfWI5LFyD32HrF5gl3zRDd8H
qfe7M7BA5TqeFduab+7tJW1J01JQvUGE6JG7m7gtSt2BgMMnQ1V7o9L4HNvGymTb
fU93PX/He52fJLiqsyDxtqBcJRImeV5GHfsKEj8py1mmAH7Bfy6Nj42ay16wrO/3
C+krgrIzZ95vp888OAAjR7jsthLbRuaRzrKcA6j8j1q8pE2SenTR4si/s6H4YPO+
ILWSqneYJttCvQWBdwNPu4pqdyIRrVMyKOMTDZNJYbQY9X6PUp3wRclv+u5E8F7+
2Lrj4p88iFXcumo+rgKds5gxGgMsP/QawFKWO8mGoftXYFa133Z9g2A4la1baDpG
3MXGjR4IogYbtvK1WbdR9sigGv+IMQYLIrVJg+VMYqH/cAQsW+Rh9Mkz60mpMDtQ
C+WiGSeqDX8MNH9/xplxhfzr5RM4ia2X31ZrJYHa1ajTz0ZozwT2zeYW8HGT61zR
6bxyzfBsiNJFCV+D7DW+wdyVec4JHZPXaQsP6wqYw7KuJRZsG52tbXEzTrxyWecF
8RsWBcgbzu5FvuXk9HeFw4ipMHoQL0vahQ9RGYKoW/3XLUb0mgyeF2BQd2ATc2SI
F4OrY817t0RBGD6TucqfKgeinZ3nUttVSKMwfk0DNGEqItfjBq/xtcCWZvO99WQy
mKwwiHmqcQv8xjZHuZ/Acs+xR6FwY6AiMPYX2KiXVCIHR1NqvE/3Lr0NmHK1nInk
aImaKXoBnbJsWuAJCv1Pl26kMPT3J1rR2dHm7G/tMYGGEsfqGlQAQtj6MJD7RXWC
eumN9U6tCByKMszWTrT68gg1MkOiMGxKTrbezmJTRhPM0oszA5U7usQkMUCJA+8s
9RZvaiFp5Zdu/TTSUhnZY5iP/cjYvYhpi6S4Qa8L//eJsnbw9TtScOA2X+gugTNE
2tEoH9C3yRDFqzg2XKRGBvY5dkI5tWmcnxCRfXn8gRqLFJ+QKnNUM7pi3BvNfg2y
kRRoBznDAiTdsuVAHlN7F1NEdlDzESnQ155A0vosmFf5HWxPHKi7sF2QG4uP1IMp
U8HEjyak18L9q4zklJ0lk3WrrYOjQkm5cUt32M1aLJuUox4FM6VZt+2Glentyt6Z
3vysmAxFwEdi9k/QXIIwzb+8sEnRPKEJJ2J4JNqtNtr6MPqehhitu9Fqy4engI1d
13mV306lawn61eAWcC6jv8zmYcFEMjsoiyYasazpwnsYIqVNj5RXcAKZS62RXFFT
DYp0bCsiNiWMavnpHnK4P30PiXePH2D4ro8rbIPvyeSE6kMwYIJQUMTVedHr5c4o
4i91pn7i+DvSp+MmOsRQWCCXM9r/jlvibPClkiOZW6ME8odjdUj28zNjyYCvgRSr
xRBbC798wIplc/1H4XyYNoILWIp0v3xf4878m8NsR0Lp9KH3u2mztXYGQ9Ao/mnt
m6wxxMxQclyMKqu+76gpXS6m55UC/GrWriOHc5fwoooFo6wK6TmPouWV6jm4bAp3
u5RCe21daqNpFtbfvc7I2HOZTxVhR+QnoS7qC6p3hUtyasueQo5HohA6a/vb1Jaf
5hrXFj+YOA9HZszfdPuAo0DHgWTZtGPRIUpWvIHRT7ikAGSUCY53+/eFE5F+3EGl
dPOMAJTpmZiU0xf7XbEgHVef3YuWn4Erp58eETGq/vuqEJSrQAf6fJj1oxX425ZX
CynBWA5p+uo3gq5LzBxjy4NgFGCp6X4Vp8yUihoW31V2z3puuu5tOvmTe7b2QFE2
rivPE1Sxe+Vaes4SrEm9g0C1MZFV/XGEyoZ5Jsry7spj873otJNhflLMqYmG7rQ8
657t48Gw5uASsGK6OWORS5uPnfdeVrLk9l7VDepS8Z4fnRw1EoHgWff7+zuqe3sl
Ii22g/KxO3Z/WCsbhoKZFYiY1aWBpxSUBMOrjL2tng29kj2Z/ED5Y6YDrpwQyapn
RSW3i4DZ2ihT49tCaTPHO9DiW6rxTxbh19Tvd/qlGXETK/vDH4VAfT8J6/xvDZPY
LqeTqFMkRARh1NZtxGY9ScXKhhBkVrxOZkg2MHSuQsEUuaI7LimXkBPJoSoW41e7
gTPJmY+4uIUGr1P8tK5FmgD2HFAw2/B9+E6qr/vG61BvrIyMXqeUp8tN5yHNhJuk
I6xFmC/ewNXz2jfeWfwvb+MR+yOJyNtF15F7CpPBQWGH19oS1zP7rJqvOfuEaHEb
bfI8tPy4BMSnQyvOCTr8Y7kqVwuqgT3OM2O3ihUbzn50H/cZOFQid2CAOu9rrpIt
AB8U+Acth6E63Ec1jTx4Wj3JKQ93wb2RPxIpnHNlhtKnhe/0HwErR7RiQi9SaC2w
lv7l7BBKCvhjPQWkoM7oZRpnQoDpbe9RX4JozJE5BBzGYR8avxYB6M0MPlnJ0m6u
9EfusNkZGjPQd7ofIxxcNIUYkjyNF7d4vpnjsZLdP26A8tT8jJf9pd6NcrU5TZyp
ezx0As+LHLLlA01b7kixvI1rHMfmdL7dh1GSDBJTcyddxuMs3wRxP/Zm5mfeYK4q
f6nUBLwbIqhujW5qHqJdwDNZnVIOLdKZ4ycO83f8moovIvVXZ57bYzcVae1Cm0cX
t18CX/Rklq2a/43BwdsO6UXCmfOwxwqHjByxPFGJ7URCE0UKfxWCtidpO8wVkOF/
bbjKdbc5g+lZSKoAW8sZ2By/K1k1ngOlsB6K2H9usssvaAisLlcNSuokRl5XeufE
CjOXVeeqbU8ZFN/hj62EYpZMP5cHCcSw0Y8bhDpoKRy70IBhuyKSQga+gka3STZ+
tf7hTZc3++OSyYEF06gxIFiaceoZNUIwepM67YbFJuMNc5EVByJlvkgXm9O1Q36q
0vTmVMzOp1DsyqqBL26Fykl6JyHA+izdfP48U0P8Uzv6JbYsI2c4IWOao/cVF7rv
QbF6y23jpu96rTvK20uEqr4MetCzhdPdIdn+8pINTeCuZ7BPJJSflHdFkEv4oub9
piYDlF7TqX947sP5gWbRwuqdQuUm1PMYYQOfdLrehCpJxTjDY2bxYJC1v/nbpjgn
h2avWmkpBqSs0SFuikI4vUq99EZnOpkutnJEu/E2QYke+JUpzF5/vNm49tdQjDUZ
Jpjm+1lNrRULERj0xxJVABH0PFWfXTd0qYf4l+T2VsyG8iZNqtDuHHgk1brLBEHk
ecFMvoa5Klx8Rn/iy+4k4nIsTlPASCWghJGVoRpTusFWPuHMlPEEq72L8/WnfXYa
78MEbG+vA/xPm6YQ2pgHqrl6EgqSpnHurciWzQuH7w6H+qa44HH5IzwvageN5TMG
LVaWBM47MAuevuUbczPYC6qBxKFtqAAJ6KjKqWtHB1LF9eynOB1hR+tERSYw20vs
uYivtI2C7eZ2eSZRwp1s8SvrP1tzwUm3tV8eaDGrKIONdr9PgabyTkttdEWtNBTB
jx++AeFXdoruo1lQn2h916sPvu0hOT69OyKJw5zsBQoGvjlMdKsHeEVNRCm7U06g
Ncpo+xcyt9l9IX/xOjbwE4SKNdo4SBzin/x0pk8bXtZVRy+2Q/8sPHjXDajM96HV
QYj/5TW10b7PwG4VRHIpKQTVebuSnItZn+KVSEMJz7EqNPUp2UZ4vgfH8vcDyF98
N4PfemgsdrcG7zcjSJhs1p9c4+fjetvkfjLq5dVp94IC1wFHcPT1SXmZ7AwnyZ7L
IzfU5Vrpt19d9b4iMU//Ev1DCKZ1R/SuSCnXTx2/S6hmn80fzQOek0DftLqkytwe
SW8KPd3E0X15gSw29pFvua7awJV3ooz32JXGnSHvnJnGGHXqmMHnhZDqc+xVTO52
e8Z+Sz6a+WZqN6dj2Ec6MHeXDYFNuaHx/oVWD4qCESnJk0vbFJZftv9oYD/FS9tq
r7MBfuf61XQ98QWSYVkMFUdZv+RGrqhjGAvtsuQ5mEPpNplqtRSCZC7LNZpCOoVx
cyGa3xT1/vm0eC4VIs4SQPfEpxVeoPKTtW9xtDun+BQE0FUug6D5b6+Xc+/Ey/oy
6NFWni9PdAAzKdIj7TSunzf/O4vz0vooikqClYudHotGbYa333Tx86MwO8QhvuJJ
MKxerZYgDWsiq6KG29nsKl7h0vfSJErqHmz8IjkFlOGBBX7JNRfJJZ2iy2l9/fB+
tWbCMA/ne8DOrL+StYxYe4vgSpKqzJgqeyxDCzoSEsnOofortM6JGHXVEk32cF8M
uAwrF1Y5bVwTakUO/UuRJdS20+pihoLDjdTH55wD6w+QyR5Ia7efbEjoCGu9IYDc
eJedJZGCD9BpBghziEG03qdScjfhg8CE64A1VZVnAvvYHOxHFU17h0v1XkhvPU9T
gw2BD05MW2tHNgxY04XeuQwQCCr2Do2JOmm0S5RJeh/0H97sh/O3mpHFAsKuYxKt
bFS552tBbDZQU4uJKDv0rLUu4jKq1uXJF+woRfo5KVY4eGFKheiJJGnP2FVl02NT
zQj/W0UwRw9/iibaaB7At120JHRWL7j1EcJxPBu0DZloi/4BGvENl1zgFHchAgVL
ndlXRNGj5/AUWVnAXq03buyZ48VzEUHTh51Gwn6eWma8uxETwkr2CNIyv86GQ+DU
BBidM8snjl0pXLYdmk9rxkeVzgt6qc8KAe95X3Y/jMj2B077WJH3smxtmnMRBStM
sMl1RLw2R5VWIu7B71x3m4JRUKq9HjNEx+TRqLVNHVUCOoD6U4W8gD1WBDaB0m8d
4HuulrhK7gtEXJ1+yPlh/oHuzzPOQEfscxx8MXxkXmoAskcRWexigaKCPuysfIfM
bhBVA6+kQSXQP+VkYeqoanItqd1ah7b3I9WVs6Aaeu8PcG9wDhG9/tZX1imswleS
8TO7t+QKKb/DL9qAhptTdXc7EMljATmXMjvMDrx2qu1ur4w9SGpXR8HrsBNYPzcJ
t2ubH88tyTG0+L1vFoYDvP+Gi2adP7e2+Hyd/UyZ4X1VtcVszYMXZUl7go3aYGZ3
+x+ROlr+tT/jRDQBTmsmy9+/2BtSncrA4C8LTd8LIkq0F3bcFe2aBoqf8yBvzbp1
iVaXPCVbXxSISACir1vdsB2Sq/1dSChHcA/0zBjaYVScBSC0hTSVqpxvqFh0YSVU
E1VLGczziISk5BSxcvcLyaK97DjpX061XysSM9YpN5KjCbenyKVVjwFm1L+rzdss
4qM/t2HxuRIRilIJb4qzfqSUtDXFrHuqYoOqSMaIWLmaq/4+tLEjHqdQXd5gTjSt
ih3TOS0tGtAGWzxZ7LuHql6CMl8PQzIxMYdFEjhN8b8C55TEQrVmcqo6GfJdI8NS
dIJoEfvtJmyFCWbmxikTCaMMYpB2onrvYxSaxIMExHrK2VH28x68p7thudgdm+4l
ETNJlTTVy7674J7gEfVrOhGfLPZPAxWxDqXSv3+J1if5RvqyLx3IjlfrQ8ThCZbc
nd+aLuWNzoIslhPq0xttdalm2MIqcsTLNz1uF7JhXKyU0fRXc6YR8WlkrIco0neW
bHmG9uvpT9E3m/RGlfFIVIrpWQtKff5zftcuxKpZnv+BdAe65nmlea8g9xwiMX0c
RwaoJssloIuYIth0SiZgBezwC4Acqrmqu+09B/WGLCjr9BXKXUsc0irVXF7aUJda
2WBKa81tL9bxkuPZcml79pXtHx+AOXxTnXt0HO4+czdbfckDdnetEUqb/m60GAbU
Ju65GlSGEk71cpf0jgHT8QDSRAul4Ffiio0eRFxpwYr+c9MpXsuhFXUBtC2fs8zM
Urgt/hg15sGTTTGdcUTO+kmrSxh7kRK7x2ENoifns/kClmyNtN/cuuhg/RiI3qjD
fhvrCOAkJgIU77Aqi/iE6Jc36silOgC1UJ5O93tQmN+j7okXco9xTUmsW3wIdH6E
SOxkaE8ZZukVEr5RBR7Yui41YkCFiGpCoLdBRaLwPAfnMSZwW5uN252Ar/LTeHKH
oWs42IVkvpxw18hxi6OPaWwIz7b0Wh7I2ASxT4Vtd8YYwXDFVu2SGi5H9J7N6w4V
g3o8ynioKClmKirUKXWAS2JVj+PRB28YEJF2Ya+HiFyyBDKtWFADSIU/opomnzQU
x5aGsRFNIGrmPLa22+VTE0tA4YBe8dp6rHoDKHV2aJP9Kttj+boIoE/Ym/Ok20QR
BVzmYhD7Y4WShY94OfhaGQPEMiYua/dNbEKAngZxe8LNCm3iCZYZkPjWqWb8bM2N
7tcH8M8KCuSpMZ5RRrdsA29Kdc0D3kgGF8tqFFw3YK/FmWuFQDmCpfzgQ9Vlmy0U
I+P2XEtDI0oOoP0EXRh/+87d/eriz0I+HHUqfqhtM/XqD/5nUCp9gMQ0osrvCdy/
6BAjhHL+fM1VQ7NLN7C+a4b3Y005OhL1QWrDX8RDcaaykA0Kw1+D+2E8ENHTxcZr
Na04ioTRgN0IV9tQspMS1VwEFfjQ39i6KrNPxZwJlCbEgo/j+1R14UF1f+7haBrE
+m/30u383pFyN0IsKCG+qejzm6vEawVrkcD1wGfDrPwU9DNJTzv/FFLkwy1kgNWq
HQVRadOoOENJbmJQgjAfYlgo3oIOl/D1kICUt4o3OGQkEW0ktMWndQWTtMVoyqML
tu4uMq4RNuELC9DUKmpAJlTAUKhK03MXNlW1gMvbldHVMBJT6WpKDb7BSA9yQPrK
Tqb++6316qjGi+/uWdLDltrN1wFj0eespF69v+l4c+NHEUm7ABeJnIJm+b9bXEn9
yXn+07nqh6F/rNsOlk+4obVxTREeDIAr3ZUc5dXW4lUYEYA0Jdpuhjjg53SQWuEJ
5Og04m13IfLjPt1U55zXgD6JfzWqWGOvSgUntYcttdiCb5aVSeT13wznJ+JpoFYy
i3EYV/9yQn2u/PC9k/+dhcikknOn/LoKAmqHgXpaGmmI4ySbnXGitzMj6aRM0iqO
qr7ej72KxXvreNgl2txUAIGfPO37GFHGEIjPHkNvj5/qfCIrqQMSLe0ibiMga1ry
nWgCbkOvpZHlSnI4ABM5p9so+oy7kY9qMONtMnUPPlGwb4tXeTs/o5ZoKuOkSNNn
M73QoqpWKZYUTsyk7AqkWpGtVvtNKwCmxQnd6C8Kr3Mq5qyOjf8LLlaWyBLWHykP
3xeIThUFy6aQcAj7FFwjUkrDv0FPKSbycTC+dxrmWOkqPTiBHT1Pq1LaUCzDd7/4
XMKdfq1JblABm98x6sEjFBlBfvmnx6huLYm9dpsmfBKHchfB1xWOvjL+khrDMndE
gezHskT9dfpY53iNtD4r4DBmLmpikhmjkumWtvOeFJllfvZIhTgvaAHXnyudGYIF
1a+1SH6s0xbM9ecUdibv5nMyBCNQE25GjpHISJaJjXOufoNaEztiEVsaTTlGCYU/
Dmn2PduAJcGz5kjKue9u9XIdp479SgFg1SOZ7BcqcThFft5CvtEYCa3KeE14nf8g
aOa4q/DIP05gzaKJ83L0PJAvYLof52XNNg1i/NsHhvSRbQWCmtZO2EOLPE2tfbde
fhQsJMqSf8FQh1A8Ajugcc/zjjvgTTe7StOXGtSTPQzztlX8dKcXoGv0YqAlJjm0
fnb2J/7+GSiWDIn1jy68vavObI7k1V2DkGqdIe61FD4iPqOkG6Vohyjv/GXoKi7q
Agj+Xr/kmUhYN8tTUHYegkcZAGLKR+IBeqpxZ23AC3xfcqthkKI0kdFUyQIVlSTT
IHfnObAz3C2/EyAYCIbPnEyTrclCUxs3nw2IqagbSb7cIGKzZZeYl3FOkH9XTGFd
YMncUgSLq8RUiYzl98X7hjvhQygrY5rs2KoAFKHDhOGDntCXiKxswwRo8hr5L+8E
svHhAXtA8tJuIt0IklLeAKshRjHTebI3mrTKyOzVwhgzu6tBLWKYb44dWBUGRqct
nBa+wGAW/rS2xvMN3wHTbba+9n+pSMocF4lx8zWadX0T2VyTh6fHpdY5rWonzL1k
7UZNM/HU6jp2SxLwNkF8hjzSUsV1QrXwyorjo7+pu6ejAB9PVEL+TiP2PC9AzmCG
wEweeEClX1XW81gF3XCNRpHxb5Vm8tV/g5xIsp9bSgt9+g58iAd/Xq+7TKb0tJ7v
LdFcO6hiABVmb0dqFg2hajzKE8HtnZk54EtFE4dsL6mKvu+pdiUbj4txdkChYDMe
I7BxUSHchiHX7o0tuE2U9hzS7M7ErmVvw4d4meNTChtrb0xb46sjy5Wt7rwJsek6
Cz+Rc1GjYd4548fQO3kQfj+DSv/1czIqxXQF1MNzjXGZxYgENUiszQ45AFjSQjHH
9r8/0+pZuHdyjYA4CAGEXt+Y1CNxfA0/OzlURHe5wJRNCfySAdh3rJgYbFzp0jlo
xQg/q4XwDaupouFPkGuuMWnHpIj4jZ/0zfS1JfoF6cpoxoa8BoO2z6nxGFyd2M7E
Sg2VXzyFq33kRARcb4Sb/ruFDEjfXp+YjjTSZ9S6paToUZRyKXcqE4bEuUUstBUF
fpstvbfmZN0x9sKLcDrKP2EXyHxj/kU7AAGnX9WoSSOp113Fwrr1RuQBAGfyFuUK
4PB5ZsgSCxsCC5NFSzW7VdHBGT6tGX2OFXazIstAMtE3n/D6igcqDk0do22gwDxj
ghausERMo0wPA0+nj1MFLMMssPIEHZJqH7Cqwo0rdllUobDUTuAnVUhECxAE3J4t
dKUMrK51PG/MgCqe/d2svYUsZT7kWSJCfmm5loRpYFaE4YM3LXX7dhx/zj5mPjsT
dq4sLW7oskPZvThmCTvKmig8Dii2GEWiul6wANOHRvekVhuCnJO+uzQZIcKmeWno
TiCBBnE+lmuqv3Ru7xhfOVeEbhf7IcM4wGntyuspffcfqQqbgYhMv9bphaaQC46d
mMHq1LCZIzJdbiHC+0FimetYIkRQjEzWZKz4MAohTwpyoAv4KZHDu2sEtnhSqKdS
m6JFRHjjik9ZAoGSTotoASPfpzn2zetX5QXCVlrq6IjGsnx9MUZ46X38QQ4G/oqb
n//sAatLuBGcvajU/CNwN7cv/hlH+ftug4tepYxqYIIZc8Vj/Tb+Nkls6UbLO8Of
8Sq4oXgEWn+/bLMDgz4rhbAfZvjqzCVdLnLDJQmmPyJbFAzWQPoXGDJuOR5Af96r
zPpUM9Yjkwwntn1WD6v717X0gTHTw1KOIDLkaRzOltrtV2Ef3N9iornzbgfCTR67
AterMFTyny9QCi/NCcy6B15YmIOwLhI1EPpAkBa00BYn3ERZvMcgOYXpM41+JHR1
ay6oKNYWxNFqNP3AZVzjNSHLVAf0aT6gMciUnx3ndiB6mMhpxeW5EyufLva6yzcc
V3JAGJnqCNS/TOMmb3CaI+FTfa9qU8h9Mr8vDbmxa0eBgUOZGNY02NoW9KNAX8+P
qro8m+VDTa3Jdt5oqk7xjnTXuPzF00BtiNqSZybB7jfp0o+hP23zkonWTb6k9mVK
G9G9q1LTWpn1YsyEGKcL2ps476l3hN/JiU82iWfbygB3OCPklrJYIn3A/fNk7JwZ
Ln52p9Ocb5nvHlHuq0w7QmfLUxQrRo3PSi4pw6Hyrd8W9JXX0Z5VARRtoPbzaQhi
oZRuu0Bc/4UZgrFJmOLn5luMJvqWTAiUlPxHY2M+rqk38rO05iQekWfVrHw+W6gW
SNie6UKFPdjHGuZFQg7qHMGDUgwh4rYB1fkgtzNfLRuYsG42acmDF2yv6zXgz3PM
Cv9ImWNvaFIicWWWH1cPsfw8BIy1ks46YlKvjH386Mp1VSFAB6+CSitHsjMxTKdT
1NWt8/kToeP0hlz37pydi2hKjDCPZOP+ZDyJR5yczG4lhwc9hHb/6UJncz9BI1zF
N0m9qzE1PYVX2K3GHMCU6OAGNw9qwCsPYP3rNlbx5XLdn4tmYoNcgts6UEPmqCBl
Yj2WhxWoOJVJWvLJeMiS7wqIZE/846WszJrmVXRYAjHzHtfZCOCORW/Ej52WEv8x
AI14aFo+Xzt5XpbuUR3H76vHhHSd3kYJyFfH5C5SAPmsy1uvAfXSDQkuLeALyH5h
pTV3hd7To1tkrtqoCB4v7Ul7k8ea9v5+wEXu09jse4c1VfK0OHe2R26Ui9Vfswj1
WBP5U+04zhsIxhUq5TPJ6lZZ4oqWraRmKB3z1eHdmVR2X4lb0PWfd1X8dx0Myc/O
yNoyZSLI9+earZh2Wb4nxTAR17McOAGf0So7zg5gBF/9SBE6f2HVXR8szdZvFKZS
vIqXdMQcUVEF+fxHi1r7cxFuwbA1LHgKRLs07Mnm4VrzC46GOTjwR0aa8fPJ61yJ
6T9JCRvzMsuC8lTXQToF8CnfmCBCzFef+t+zezooUXWTFfcDS8Cp9iKcQBzexRKB
uUuH05eBDKBcarxTNnKjC+wVlTan9IBYpimSk5vnSMNxzdyKxsqR10Zg/CLopXjT
J/18SWoyEtDkqlhkwJvCW3IB9kQTM88kbnXJtmO48h7jUEQZ1L+7VE0C+JJaGqK6
sxS2SvRHGQgHn62p5wsL77N5PBOVbYZ46WhmG7z+HUm9ayCJTrJkcXj/OkF1LhZB
qoL8/PVviXzzhYBKxKiMxhUQthK2TfbWYaG1UxkW/vwVrcXC7TLetpxIDYv8s8lH
X+DT+YxBfUQjY61mxhFeRWsXTk7LxmV9uryQZHFgWWHfgW84ObmLpat4yx9Wl+Sk
75jCDx3IWqYuSZrUn85ydk6+KjhU5RstJohSUeXttlOGDoKEz6kV815khxX2e7hM
h+5SAr59StRnEdAestZ5Kosxr16/IisgnIy/Q6V0MmQk80cyxCL+V5d6HDiDzuuv
Qz7zawWxZ2lPSTf9gM9dj27XpBVVtD7dBdqwXwfmbb9FCzV+EsDvFOhZ3SViUw9b
0h4LFamr6G7F0nTJBUy89VQeCzLrigWU8YMbdRpD+ySWgYiMDEhvu5uVseJnVIUY
kqRQ+zwRDBU4Xbu6EyhZA1TSjbNuOJ6KdWoMT3rSHRpezpRY+ACOXPqYhDSbEAEz
GW2f2NDIKVrurVir34YQMKlu1mEo2rUgO1+o4yBRi60luFqsTKWjNslElfRrBkWp
rzAmevLKtgu9OYsvwka337iSAXcDsHDQHYIOZwsmIf4CqoW0Gs6gjFTaNbOtpkag
U/XBt4IRCZW0LhgYu87BLjWrMy1an4LFoJ2Psc9Ias3qm6VFAa60iigIrGPLn+sZ
goWFlAAUI3SEqA9PLuUCeUxYn/SVKBcwG4gAFJ+cqgRfEjhhJbHo5hRvqx83a8sC
cwY3XHiLvX1g1Bfu+HYp9b92eYQg2JmE+zE7MtyczEt1EnLCNqyRAHvkjB6L/sy8
g++1sSSFMP9/3Ubo/8dN8f+VL2J4miFgpulGsqqGW1IY5whCR1yqEPuFJNlVLfJN
efyOexzzW/kuTHrcRARoqGfDDTp4qnJb5c56gQBYycJL7JfnFR6R6BtSAPpMhDb1
+ZkUYhBrJRkztmRUAZpjpGqHRpzBU43VKyDPe8/2dgcqSmQZVW6dUD3Ci7yhxhh8
trMPIdWUPstM3kJSOFdCLjDw2tPjhfAZ6dyjMGCqNT2Kjc/9IRCYh7uMJkQKDK8m
1QVqAvHclNAbCEao+cjkqm7B1GpSeK47bmfZkL7hKUYjB4UMalQdjaDHRjyQp0Am
m6VdEU1TclgmEzFzYzrfSwhwwqKt6l9Q7GNxIll6pA0aELczuiNHcMa/tOdtqCOz
hA+jLLvmqc/aq4aV7ForI619YskFQXpuBQe0Arvbd64UWIgWSWucWD16J8A2/hqP
zNYkEqIJbuLkdZ61HiUryFWikPu4DZgKR+xX6F394SX1CLR6dBmqCP+Ns6+g4QXi
WizdfFILl6BtilvzHZJUFSbkNodNMK7qgk19XgeoRfd+X2q5ee9pyC19SE0D1kbC
KZ19DOrv1sezODKwdyFoVXbTgcujdR9J+IN/c7eC5Ng9+M0P1csgXliZjmKqhfGX
kJMHAX04zJJDq6HfbDWhblRgrjzfRLaA+4D+VYcRVQPPSPH9QyPuxgx+7tiRwf92
z9g6fPuqjDnRoeu+AqC7/GBLXzmPJVNxgxuyLq12bmNMNfQf29UhaaAVtqKzED92
/erXINJh7cv/gFeP1pbmcxDf9nF1GPNVo9qgW0fTKgsLWCv4YvuNc1ZnN280S91w
rMHJSBFwXe8isZXNLTZceF9XN5qsY4QGWBwEzvBEdGuCAAj7KzkUkGYmWQb97oNi
revsXSmi9MTy4ZihgInDpeQh3XaRGN4qIhXkT65+0AlXbVKBtIFeZ8pW9lug8IgZ
1Uc23h3THjMaEePBJmLlzxq6ucoDmzsbCYBnkvsoB5LmAT/nCoyh0kcpYI7b0z4b
MvWsYpXKQZKMFtmEdJ0kIY//qEaoOWYIpG//JSJjdOKMEe9wBGfz62zzSIhZImsN
stlSyLjlNfAq/h6Id1NPKLyQwsyKMOe6YlFYcWyn3Cp6XKwljnkMnQzsYntWGoDy
cCda9MdRYod08RUHrqslyy3kUO3ECfri5q//Qs5ihVjxmGnm2EZnf2f+zF6FK25l
73pXMHYbEK3QRjInBKJBbVnksBml2jaek2AUCBL8HqbVb3mSpehcLLmfAhPOgxza
O4km4TC8p5G/zmKvguZL+kwO6oJKQBSq+w3oXkvw93yQVXGQyXMoul0sE1nbAR2Q
PdPU5HsbWBHoaTOYkj4ghN4nFmvMHed0MYfUVA9uhU2ZvF5grHsVxEhJevMjsdsr
3aEuRV7z+xC7qALuTgDLNJgAMnJ+ldoY+AX41fc8Nf5FKZp/ZdXubU9ZVg6s3Jxz
OUCkOz8fP6almut+MFX8r/gfLNiS/KlyB0T6wdFWbyEDEzl8hrKJNRCzc9pAidz2
5lUfdN5UETPpkUSKX5bgEylyQGoEWEmV9elxcRmqoyhvm/FoWwX9iRfnqhnJnLPj
dwJxUm1Dr6XB8RaxeOASecEbyuA40YXxKKYZq7OdAP0ahlE5ZFzQ4qHKi0WxriJF
ihSSeag+foS9wdxNdf1P9X+R7tZl3RA7rexVRyOHKJp/MKnAhUIYQX5A+7HMcsC0
KMsIHwkIEPFacAXc/fc1Jnx5oRfuwZaVG6GfEEa1yNQ3/WqmIqqRzlO8crEioqT3
E1NOZzdBapZ1IqVpCvA3jjC/w4mlj9GwK3V2tVz3KeCTUAJKd68y7hU1+q/28bYE
X4XtxhWsd3qx1SlzeHSERRKKRzGDFyxLNy5dYycl3nQVECo/tMCTl7VwYtBACe5R
FS2CPmqUeJ1vlM3d9B2ZARjbhtFHW+Y05hkUqwd01yMKGDVcogTZTzKiYZ9PqD6U
BhWZlx6MOUYOLK23sDNfr44LmyUyYc8pZx1/BNPC20I+Y+50fXp2fzK1LGQr++q7
OJKKInIyzixnrJtYQaHj+hSoL8HwbkX7x3WhYpo8znJpn+YVFtWUg7Hk/woEsU30
floJU9I5apGh6IfEFnfbF8FmkeKO/EG/4/G+XD2wBcNyefx8sEJXdUOz5l/0wpxt
xj/QjPiVhwc/slEFHPZFEkkHHHy1qIZTDgocR0IsNjbfvRJAcaY3BLzqSgOqetw/
eBWVENaFOo8yVqX3b0uY3GD+4Wbr5dU7ioo0nMukltGV6unbOAf6yOEEozkAMohS
T4tewrOGndy6veVim8pnY6t04Yo6/gr8NV7uYJ95nBkv6pNnGFj3vb6FHzKuXJaJ
2mUIu/8TL/1u108DZmfigiwWcnfghacbeZkm4oKl8V/WQ8InVzpjAOp5Sr8CUO4T
PsyOVwTbGMlbOx38wJsi5qi/yj8tqg37XMmq3k5YHkXCzMlCrYdM026zERiT/W2D
E6bXvhcV7RQvTV0vCk4El7YxGn4+T7XJN0otpAwfYXFF1arZxRKOk14qzvKMghEQ
AsZkp/+rRt8ggQihwsN9cdWXcAzC6WRbCuwsk6nilDTFvyTaAAXCw/fgm7OC3/2u
wMeT/BFRtfhtr/DcEr0M+CFBMK/dQTUaBfMFAsVfqQhooRVLsPBCYBqb3L9jB9MO
GEtOw5Jmyo+hIVwbOFN81t/lzwdPjb84wu+T4SeYOXlLW2NUD+3kygziPqlDLgFR
vMvs9VQoYdvRN4StaQu3g9THN3Xr3pLV8Zy8fTLCm/+0aYVcDHYd7x5uMxhk+9Vc
H6JQ/0VN+A01MwZ+Jecv8p+uPL9cZL5ELzLsvNFJdHPBZcfk4cK+AWVOmh2Dcns8
OeOhaVMzm1yhsciN1I3vAR2Ohta8iP2wS86tY2THOiUdhPCIC+xlujxZ94/M1qsz
ZJqJHMBj2/F4MTTZB++2bhN7QSviLUHicX8mKlmjwMH3u5T7ZKMdflal8Tpl6F00
Hk/eJ+lWtrclpBCyEkmRlWorZw2Qr7Cr/scR3tzUvCOWoN3V5yMm6zJ/1xUPVMd9
kHkbqYFumq5hbFHnUmv4Qjye7azVy0gemhxcU1Qw1R19GGaXTJO10PmUg9R521dk
M8bRp/9WjQXR5JOxju/4s78w05Q5WJqqbkg/d/wsgqNj25H8TlGs4Y2FmNCH7J6G
hfBgKZfy0Lb8Kac+VHFv3Drm01KULqd4kRGEeGIyN+ylwA3bQGJmyHSRchxkDw1J
5ym0H/ekgdp+Q1MtVF6SCvXj+jPXA8wu3g+CoG7gCfQR/npStlNtRmEiM2n2ugCR
pdej243x++CPHFB9/VDdos7D5nSMJNwD0K8syaSjOEJKdeRK5zesm6QGA7N2gqMh
trxWhgHjohL/a5paxbR2NHOzEz3x/j/ZQyeSpfd6hqXKW8JkPQguEkrHFgspWAya
laqDvD6Cpk+2eFVcEA9fod/WqtdwPlKkPsDzqgnBAEdh/2pOH/ZdhbtJKNWOsOE+
5j5nu6SDzCsIjxmURazNwBm1Xbe0Am6NXFcswb55VNXHwfuyyEeaoUxDky9VcCTV
SalYIvR0T6C7uO6xrcmYaSERpmD2A//O/HJDwOv6DcyZr7HAtdfaN/InhFh7g13M
u7NAO784wpuODrVTNVUXPe+km0zlFA7rfy9S3iaESfTUp8tpyBN3x+7Mah2WkYCD
txdeBHjLXx9L9kApYq/AO0KBhqXcse79HC/+yDxYDirZNOK9TqyGNJH5cngWFyuG
xdFyPvaH86Z7uge5b1LyuDPeVya5i4nfbjRJS5peG8sjQkGEV6hTlcHlOcs2VCiR
zGW9QtmKMGm5Ns/r4LQtJ/xOKwapnE9azT++4gMhFaHjCW9k8l0J5aLjnB8OJtiv
wRaCoW+syk3f+vu0NK7aYNyYP4X9qFTkIqHGKc+fHH95cPAtaU5UCHT+Y4bGzujf
AGKsNtqW9MMsN6pnH8BZ7avaZ5mDa3FekL7kk4rkNKknALNBD9zhrZ3b5Eq80cnB
kSQ1IUmV/UW2hHIAzLvuZRj86lYluDFH8JE4pgEnXTGui+jBfGd64G/v3wZBoUNF
yEWzNnRDlqX/cQJXrLXmmcJykzy8EW+ZT+m5iwW3NSL7HE46Xfas1uNdsIOWzcwH
08Zim0agGUztiE7diymwjSTKYRUhwb0burJzZhF1GvwQf8ffcxTGoyXT9+1XYUm1
VwTHGlEe8Auy61EQVUA2I/ia+xQuMVm1B9aLIFywEYHieYdvugPnGRAfvqhSmbPX
0iv948LJhQVLF0SwS3JSJE7qZXlIlG34Lh+oGF82K54dC6y7vDIc9Dd0yo6BdWxe
OrL3QmMi06ase3Gp78y9zCDlKbhtZOy4uqSLQ93Dnk9wb/X8gyZJFW60ZWoETUYf
7nmmN7DMh7eKMognJhcRR3xmEn25tUmNESFQU/d+js/6OrAOkOsV/26KMzIPj79l
wSF8wX8Avow2rC5rIT0XfDlgrsbyFJN4WHCQWs5NlZhom5Yu3T+dCNep3hq0Hr9w
W63mLBeaKBAAvosMzdmBrLvPbgbrgW1Jp8DEu1zIUDjlEcxSxsSGtfHroN8TocmD
IG2PBKFwJ7q9oqV3mD2kX8nbnDbHutp98rTxdlsjJiuFg7mJ4OIOUayR1Cx6QBeD
MmP2BtUjeQCxkwNvu/MOg/7HsoNPQW0w5qa5b2pQmQkp/69O1npfGGqs/GgT+wlM
PeJ5PB9KbOJMbUJdnUjaUFSquBWIP4QykPX9P4GsAAWI2MAf1OEaGNj/S0+57uxx
mHp6fF7OY1JYFAuebqRCnKtG0cnWnIpdxQTH4IT1uN0BfNIJT17DmqDqgElYsvHr
vv25bwYqLHesqw336Rgp9ka6F71CuATfHfcbNoLe8Fzuq2J4xT7LitTixrjscXpN
kCTkB9vVUujT9B/RPAzQk7P986E1093OIKUJruIvbaf3Ndb3+TswPruE7Qt36IuV
DytvgackdiD3qBBAHnKmLWmZ1h4G47NIYKnQc9HHwrVWcGvWjZpUopNceVD9FE5y
+YqLYsJdZQiJzp2T4vXWbhU/ml2cwjW2Gayee34FTjVq3KZdoLQ/3UEMAiWWvB0F
cGv077LRohDVY/sQUkzAwBwLnFW2Qq2cI0uFxS8pyRVEG25X0VasZWCJVk/afB9E
2oHnzLDYRn6pJF57kt3Qx0yHtwGTOypLC0I4qyi49aW/ojYEsiVZw4Gv4vUQ77T2
ZTBoVCtXkCYnbarcGdoJN5FJH3T89LlFA4NmPGEFpScAd9Lqkg/AsVYl8rIPaXuv
mizgrdXeoe4LGUAc+V8zTOKdR95wq60pokdzPIvTx5AL1dR4i/NIryImLofX2kf7
sUMc5sw4kzi2TVlItpiH+7rhJ2UiqS/YdfepGJo3RKthgMP2CrvBtrjBQYqRrLCH
JxIGHvZMr50EeWHOeoSgPbrOZEG/35IufLqFHc+3Lq5lXwMTZswOIDPjK/q0Nvcz
b7taAbIyzjZeCdv9iQ4GFnGNt8N+OGu/tcc+vLeWg9zayssRH3LWDVnGjKhLtRon
Cn/dnEkIS8o8YKu6Xabx3q94Wt/UJ5JBhe3OBFz0JFFkVZZPW3Ayzhm4GRM3Rs3E
tTZ8bj5Jz0rb22XnMWS1uvBvvbc9ACwFqlER1uheC1Qm3p+n9HYZUld0Pjk9Cyd3
ccKhcSY0bUyBMI4E1D2tHwquk2D0sQSDD7NjIYULIGqnCS3DAKO59FCA8l4tuOA/
HUqGjhGTlTAiTYIRKlwhV6O4nqXsnVcJAY1YwfxJIRXZEtYkO8lyIJAnsg7cIRMI
pkq5X5G55teBr1ffNRnf5GqSP491p96HGTYTGEYLXK7OIn7mcPpUahYFZWx2tlCJ
xWg2V457B0KV6FYf/PKonqlYkYwSRVQVZfENbwB2p78ntlxfStRYSlYaZjhF29gl
TpWkKSHUi8th2CRnvJ3X/hnod76dK/C7ZVRee2690Zf0sCuKX3oRB8xY0D7X9fxR
FAtc4JQU95d2EJRXElfQg+AnNFEg4NWwTFAHGdG/Sdi9eNvrAkufDt5mgnNx5YVI
SwBBYW6nRUJWuDIoVzvaE5M/PYCG/xqWiygVtoAHQSvgnq/zqG2fEXS3F2lkWuJU
sZJzbPfln7KpMzeFyUOOAGOAZ+aKd9L/50B0cdYI2Mtvnf0tiu5yanUw5YH2zTTR
GaJWj1wL5nNzwb15SKbEGpFe72WMe7Lk3ukpk7dBd0FAg1AHyBxEgXadHe5viFkw
pMr2CXfVinhU14GJ4lvUCzgSMBrhUIQZhrrS3+Rj0kJfC+Q38k/J0wcG5fYbYMGD
jC9DHk/fmJ5eF6fdHskn0MyNt6JonUmWfejO6T77uYx4YnEzofZ5aG5NXXNDE8au
t+a94Sw6jpggn7p3imkasGEP0HXCI+aRHnNYVJCbvjC+G40rLQHQvZ6eqdOalxr7
AdGc3Eue/3SsDiMyB/v60dxYpwEH7nC/SdZA4zKIeqGntzpoNLZr0LtaUs53qk4n
W8flCxUFDD6eEgqQDyDVk99UXTLQyYRlYBGZeBlJyXNeGwHeWBTv7is19MW2ZhsT
n7y8XrUENpH7Rwg/m9B2L3w198QLsMHt/Owd2D28r4ooQR1HPFl+VyfrJbblXIbj
tUBA9LPdWbSv/ma0HfCpCE8LRhLFAlQ8jBxgjJlZ6kjU3sZmSbEfboCRiywyBeh2
i1abgxPDLnmWL5gJmQCVTlFgJs7pz9XklzkU+WTeq/y/NP3w4t7I07CzuiZNHGGH
uUV/EV7HsJFkG8NYWRHwmp2n9n8ZUmEKm9Egh00oIjOhfRqH5OAXp1oRI3nUKbr0
waE4epEn0yUIlwnashTmkK3SPPa02syL6aT6wjDMlSTijkZXDILC2Os5cS6z/Ygg
z7KCFg3HLN8QBH214AHzgUNCYC9ajJHiplv7rR8vmD0gjEns2PXPFw3qknXwZMvV
xydBIty1ufjb5ZkFZUym6Ez26eNsbYnCi+wTu52t5tnR7W5rWvKrCwE3ZBhBGpo+
JzTvQ0nZ4XceI72+tsRYlyaOv4Lt5N7xnKe/s5K81vgsmFHijpVFlkp8zV5Gjqiz
/VQw3Vkhnmn1YekKClQ3HPWZi7Rxjt9lpJF+6FaC2XU1rVmq4XzInt/gEOmgINYT
hkFswdFzoCP5O6foBOPyyXPtOHrvsLauPXVM4BCH2ykijQ0C+CBZmjR65vZ76Vr2
L/azbqNbZM8ZSka/aKNRdt0RHUC3CIIzYs/YLb2T9ozHqCuqCkMjxDBm1OTAeh6r
FAU1kehet4b06N0I1sNPNLQ/wbPZDTlzaImNl3wj3Cw+ISUhnF0GKOdEXL+3xopc
hEV2f7UmEJovPfSxzqwuYkkeTWINMbLd83sBL1F0nCSOt/HjXOow28LYFcDU/iJx
YGBJJZC+qJckNKFq6sQcs0zx/OajMDjhTU1BGC5pdTLjBGxW9Bhi5EKVAd7xUIzh
96iGL6U63CA1xleCJ75LatURo5vsHEske/PLbGzRJQ/lY48mqEZlLGCt3W0T8N3g
5/yKKEVCzxH5cej4RmUa2lruDo3jT5B25d48GQ4ki9c6Dmjyj6d2bFHH5ZIzv12A
z3bN5ycBDDLTkywMJU7hcBaTLiQSnnY+WJbpxSlCRywk9XIJ8a70fdqnHQJWaFjU
TTxQdW3Dk69F1lXn3yPZDb50yk2LzL5bo/kO2xqR5iXFYp2XbdjTbWgDB0CfaTI0
+Tx2XAH8V31lL5yeoA85sLl0D9Zc5w/U8OkZGFYyyS9K6zNdvrU+UclQ4q1OyA4u
tvT7B3R6W1PjIXG9840EG3O6XFplUKFeYG8U4pInRjFpzpX4qp+liGr+MIy7gP1K
Vj/Lsh7boaVaGtVRiy1dhw==
`protect END_PROTECTED
