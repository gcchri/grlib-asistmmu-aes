`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3B2mmgYcV7bGIXOx3uYdV9yOAgF5M6zKj+hzgzjIR+e8H/Tokjac3EzznJINsHnB
7c0oVx56P2VHht/NCfmC1mco2WavWq6V2h4iWF1spYH/IroMduugba/65KLi6nIv
ClHGiXsGaBLkCFapWDIME/NvVsfmDm9a9N56KSh5ry8vWxkMf/PxBRKbnidfN+KY
P1FxAsso77LNsl9qYhjNKvIfWdtd66shquDolB1WZk7MPJRZmWfQNQSpXgMS6CKa
jV1RKNIX/++aP9IMIWlVfour3D1qgLzAjC2yTPeh+RV+/OF2+ObzLV6/KaaPRzah
//ArI+0niXvo8AcOnjKkDYDSLmN9SBf9gNSUQ2gitKRtMCYIQvsRKd1CdxXweiGI
epo5xFsFzJkE2dwOBAhfi0gq5AAUGpO8yf4+j5t3dkfinHfyn+4MDLWuqAQWXhzA
VBUIm2l4SNqb5ZTTCfON0f3OXniMPTb0gyWa8/QHKtt8fYjXT+4YOqltAIZ5T39C
RcFqy6e72zCMeRJKm8XQ0EB1WlpKd44Z5/79z/eE2yF4FSNEsaFfCoD3L04U10t9
1AxxX1OORjcv9iTxfSrl27DaOCewdm4I6UikN2XaYQJjBESloN0ACcgI9RbYwejs
joZdla1YZR0qNVlrQsXn+n+r35sZ2d6erp0g38sVWZexSJsAbgIMBBDIXMy9rAjG
zEEbVktDQKdiwwTontfTHhADn1BGtgnhXPpqo1M5wKFkLUvrzNS1fipG0Kuafb/t
IPO8IKvPXbWliQb1IAI4+O7WSKsNVvO79BIF4F1jG+tU4WXDsfd+Gb2PcHWT9G7Y
t3djmBT6FHTLeRxO9s8+OFCV8sKxe6bzWQHcbyQH/GFEPUvz4qnlD95LmoS3x37P
Xo2dRB6+3yh06NntVeLe8yMDciffkP77z13Nur533mR0L1OyQHOobRzT1DTjwuOK
rbWuwVP9OdpuPO/FqqExBxsVBY9K3HRjgiY2gaOdC3rz/6dA3oOrIuUw/CHOLSmm
1eacayjft/MQTqzNHtePAPDRZPtQ0hF3BsUvj2Tu/ZhS+uCkd6MQo9nqgC5fl1RO
T8dsO32CXPSAhugE112aBWQGL88gFMdOuaVoHcaaRMzVVl76I3juPp4KxHpb6Mmm
rnV9ww6PPtKoF9svx3zGwTtpBLFcTCRjRZ+S72L+Trad5Lu/9LyIz6KlDpUnERBS
05LaUiv9V9V6FDl6xgmY8KoXh+uSwMevYSBsriz7u+Z1KuXQKJj6UrdOqzZv8yrj
ChT2CFQz7aM663QGe1e4CxetG4zSNJ5Dm5i78eC5zIcB8yy0h/OQxTgDqedrJAmg
9KyiocWSEfChBg3RX5OV3kXY+ciJbkdS6+ZMe2dyGWO0fegQ7DLahQnk6m1e8zpo
/vHJzaTBqvhE6LRPFx+flFw5+OBOegqZuMjsp2GEnzIyUoUi6ZNMQOsuATx7T2sp
dtBC7jej6W0NM8aZCwNRqiHL62efgCAkCfYfROBUvcXBiprY+flhABM7aSqnEK/x
K+yyk3+R4SqgWcNDHAvXtPnnQlOewJhfzuA+YlTMO25OGSOV77EUaZ2gEB4neR+G
Qde/oGStMiGUdOi9NUDdng==
`protect END_PROTECTED
