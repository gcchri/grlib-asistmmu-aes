`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ty86l9sgDwfNtnis1AuDBMbUhSQULwvF1+jvo655qOOcXyKnnVrHlexq5hS8VOXf
/WOMmO9Vgt1l42+6TK/7qO+v8NTh+W8MTRwOM/PkBmYUJgAk4Omj0dKt9Aq7UTxe
LzNZDODBhG/TJHVAfDbO5HXgNRkbZP9dq0KFmMDY+m54DvTy2nHbArywUhj5W+I2
87KFG45slc/FGE8DR9FcGW6A3ATmrGKVb4h2lCX8STZ459HwD4+IEmerZFnfgzeH
xw/tbmdyzV5TfhiQmBs1pHix9cM3+pAM/cjarrc78rnOTtGre/m1y2v0WyEMKv0/
hxl/kBW634rvsEt6TNdigEutg7C6x92FA/NOkyY5PQi404FOOfTJ1+r9l2Th0rA3
my4y0NV895EhZExOImCE2KgmsiEIy3HiKExDHI06udvIfolSMOKw1125hnNTGwKm
Eb1Xa8kK+UfejRh/FXpqEnzz/H6OUj2M0aVvz116Nl0SAPViNwUsrHREv/B9OEqg
wJbtDjDD3/nOpdGtLDSpEZ+EKc2NbGSgEjlbUXuuLbwXSDnyqFlM/dnUZSNX37e9
58osjL9xNMu4a8OqXI5LXhZohoJZWtlgDVzQpnQFgzzHB4uJR3C2y6zaHiY33i2f
eiippMh3DlD+4uDsvykfrCdFw2FfmxL+xvY3CjX5fUJIVn2vfM73uLZ6Nb23NwTD
MduGQI4535fRVkNJpQ+kPplSUV14E7ye9ue/I3dt40GwAPaDajd60tDtNIjcoMAW
bWboqf8LkDVMq+sDpMS+kSfmiA8V8/xMpnP9N9VnsiuUgthk+K3laqVqEsx/RwZ+
AHn3JravUE4eBuVfZVa1DgJD3hFDakDOzrlgDQq0pVBHEQ6x0J6AZfQLB2izhVJm
ZmKahYVLx42nIm0H43gWuI+GIsgH18SYxxklYDbt5FGCqns3j0DqrfO3eqf7kBxy
tzwKGqf194zaOkAjKPW+Cka7w8aG0RV4vpwcXCHUAffId49ykSCbD+5vc6tsi0F6
/z+uIUGC9Ut301yKNqBP39dVyX+qqyae2K/Tq/WUGTTSCfgWSr10eOrUdspFYKZp
GpPEmk62xH1d+W5cY8mAjq0FCypxkTqWv+nusE1EizO9MnA568TQrKLL7KsAD6Pj
c0XpRSbmx9QSayYxJ4sQPI/BiDswHVV5HMFqBuB3g6RfxckCscyypcatiA192bsJ
lvotb8HZcudmKXjKUlPsuANSDog3PHtGHml2GcG8nRFw/dsrD1H1X/RuX8SatHaf
Qi5fpMUQgiax5KiQo7XmFtrq24HHsVCNd7IYHZNunKjdeU8zIF7ovB7msW0UjxqS
sLPGWpAEV4JoCC4YEkX5A0Mql1w5HOJLTKDRPvNy9V4LgoMxQPzHKVPP+M5nBN+k
d00hl2gejKnPh0cmB3Ilwwx+lzLazP2GnRfOo6CY8NQnIg5OCGuSElT+1Eu7UiE+
jjySy5gAdnyStqmn0nChJyNuJ/hboGu7a7n2gJC5suxcbuCnc9Agr0tKQAAxNO7t
lA4ySYI0O5D7vzuTaqOvREaW1FtutggFvQeqz73iMp8RK4FM78Tsq9Yr1oy1s4yf
PuGAM4Mw8YysiwFFdkE2JIe+f3c2Lccu0Wk0B+KkDAuqiZdal358UyeCdexUmsKO
E1gphDSIcZ9bcbOmCntN7qLSbxZLa5YMV5QLw/RJbNl7/m1NF44fwBJXRhyFzL3p
tdEjCuWqZY+wSHGvQNWgMTp5X7Nc111plBMUpKyZTlNUaXet2yfloqkNKw8PmXM4
fuf65r4mrjtCBxq6dxdXgJTvyDsLwahdJU2v8dq+PbF2eJBJAbXSIPtYpqk+XBTP
0elB/SucaZL20yfKlucQRWF8oUJtLY7QmDit8S0lAtUYIv/bVkdRlLUCC/wDnbIy
Of4IQRHX4Oo/uXdE9SofxXFlEeVxNFhWizePrzlwleDyHKvkhlRTcalHWU4YPVEs
iN7mo1FAB+hkY5KsUjomFV075pwVZpgCiDVBaNkiRz1fcpn7FkLiPLpwNnFOFjfX
PAxEHGxZvrYI0O41R6wiSZAUHrucli5YvEVBBXkkWExHooK31uiD1SUwFrlkHbSN
mKwhxONTHBAvWBOvtmAfVkIZsFzBJCBONVXmVG02wk70aJZ65DXvlvUO1JQtv/Oq
X0ZZ6YPJivnPC2777gzFwt61qWtHZTQggL22EmTBditDgD6Cm8SVaob/zMXEpYmU
V+yM8WqFx0S8JZjAIHyMHrEcGpX4zMguTk0k3oVF/enhNwoY0rZlUxHf6++cMfy8
2BN2YiCcVVhl/JtPW/mUqul38bkYqPrVZ/caPLT7h0DqhdrDR55dtQhybNI9s8C+
45r8YggUYWMUIRzPgZ83t/om+Jv2yvXU81ow3LKxz8duBsNSXmR8KCgXCHK5UeNP
bibn6rB0VEPjgNE7qMNjy8e++y8CHethBD85kMn88zLwDd5HbDITyNmKpxNujwf9
Rt6VCCGxN1wVPn2y1E+DOTb+mQihBPv5H2usQVpub+C26M4gPHIwkmx/nGMZvlJn
DhF+5OwMy+8oTfpgNkrnce4DpRMbMF5qotUurWoy44KbKnwoL7siR9vR0fhAwruE
8C+QvWPNUs8L3tHJMkJISCsW7mbJTy2W3EDOC4h6GQN3RvbwD8J8rDOEBADeWcKF
1MgyqhJyRtiQvRmkxl0u27qo+UNVNoDKpwmBh7Bw3jgMh7DEs+0pWeLav8tSZFrm
ZFwDrsUxFIGmVX3x/m1gtCTW2Ie+wATQy2DtLLt4lWu0uiE01cgGc/HlPLEFa3rR
EIU/Aivav2FiNdoT/WejiL52rTkIZPnaZsYEYFcy74ApWgNXsZiwzQHkuNqqWeCw
f+1VzMddEjGWPSTsgrIZiVRVOvM1fhkqLzeyPsJscfX3ndGahUy8ioleZgQttTeR
tF5yod7T7Ps0VsmvlAG6WY39hRTXqZrXtcc/IHWM+zsnJ//fQr6gDJ8dpgy/XA5b
D+uUJ2wEEnBU9k3Z9FzPHAlMsjEHP4yOsLdHQ3FqTrn91+5EvlhyaBIb7z1mVf9k
V/llZWgFNY8V9tDwYdz/jmmtB85ru0w2wnLDBhrLjYzL2BsAzTfh10HazP+TB7sA
00dtZ1eRo6H54X4DqJgfiR3OHJBgc4nMfMpaM15Op5/gD/oEM2oXM/Uq0FhZywUk
bk4X0tqiaKCn51Ok48uJyQZTwYhMpk8e+y9x5GHaCEOkz5zb7eTPwcEg8fakBwjG
KGnj70KdAVPd/IS8h08X1lBv1clgiap+vodfaFxrxmA8BtVixBz+6HFK1B2rWn4v
nUjfVlAwbXK8nfdnqZGw+eILd3fIZUOaUvjwjX7I5cA24751RDSk2Y+f0DtEIuTd
SaBolVMXUOVcbA8U2X8qmuZLDUMMA7N2YHfWpxqnZhKgRr2RL11eAjgkyVZNktpi
i/J/SItLTQ8QX/WOgH/iVuU2iK67dWJiTSSe4nYUHaiebd7y2oLXigNmHRe5jdNL
TzmD/Qv92iNzhKP079w81A5pqyb6jBEfKNlAvPIx1hdaVzggNLeh6oKjmNGFYV84
ic0QA0OBxL3/bsgnjHjdpYY8gIZwIphOBCzI0QV3LzUePYN+zY0pVaZTRLdOTxph
EPZW65ybtqwBPFA5vLDKV9YyTKmS36vSQuuEXNhT10T4fIxjd0KK+46Ko8ykLKGq
rTNx74+o+G+345qOKeO+sglaVbq0MEqdYsHB8WVSmh4z0eNzgw91gdjSe+T4mtWN
KjGddTcbhMTIO6mKqbgzMqqorfRPXSIc6IMWtjkUtZvHIQ58NahDjR6wQS8ViBG4
JW4JncIgjkfYpfu3Ko0SXqpUZXU02da6jK5LLikU9s4f1PghSRBC4asExdDQZOIs
ewfL7ys2LwU/VuLqKqw7CMojLnhhTIdoX/UpfQaJkWX5DoExYY/8wJIEf4FAozeP
QJ07M6p4FiOiNtEWXPnvGagxNF6IIjf8pzEUZgvpXWLsOfXMjnwQkEIfSsrq7THX
ruE1Gxo1lOFySsH8LPPWv+4yxZeA5/Ba73i9ci+AMLJDSsb/jsoFjuQyO61xvTuo
2h5lYk/EXpZ0jtNM+gB5dszUReGfMLRq5r1o1caip62LCrdeu0JP2dsnb7j7CjpW
5RqnBu+rYq3w3BgCfF6vaFTRi0ZeKN4J9Ph+p0GXr9GO+tbSq9fdc3+ZFXuQpP1/
FPnDW0rnAzLsFwtYqQNVQa1cqtvb/aOWUiawNudHtssynp4/aF3tB0vVtoeKrosH
wouSx/oVbLylWcs1246TbG8WzcV+3+vtIzPhVVuUowLzBLXlqZ/efXRPhNFT5KaE
XP3FRgu3BnNP3BsEuedy1n1qlNz5hPSTPf3uz7u/OMEF4jBhvSse2LoLrK6nlC0m
XvpzCCMo29BRc2DlXBWsbEvrwa7HodqYdBoa5kqROpDS+X1xtQHIphXGg5ZFHZp7
iYOMgptkpHprOCCP2MA4woZq6ctRKZTZw35jGZ1hb10pe2Tj5HfIqopEVohKq6fD
zl/O2o8Rgj+KmhR1WksV29E0nwXsvaNsQ+2e/lgq0e596xwlnas/TyKe1PyLPgfM
hXVcLWi1Qhng+zzwRD9NW+MpBIDyVuSzrnZ5ZRyRKHlY+lwYshVc0ditA9+lyEIr
rvTROLnz03fYZB35XvEkEw==
`protect END_PROTECTED
