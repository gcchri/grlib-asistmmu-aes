`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EYHj2z/UQtnIFsv5oSyvLLjXaBteaXvBsMD4DP8RbyqDgxilrvEYLyj5H/41HvZ6
4UyDH2uHvi1pVqPOWGW6K76YmlZK2LaX/P/ct2X5+8d/aEFo2hKT0JAXNnI+US8i
zUDVVEmsHzM88BzLnk9tbf0epuLd3Z7+A/pO0lUZe39HvgsCsxudQclc7clghoj1
vYnERpyTgbtBGhezv11JfZ+dOcvgb+ME+u9sTraTk4IQ2b7kfoTgwcIVNEgFI1s9
cJlL+f+qAZ2NayfCAiz565Beap8jGrS6B++APww6zN8AnGrXX/yZobQFeQWXOaxM
yG+VNLtpBinpVBktsLS61gZIhZGCKHZUU0FMqMBzpsEshVFy6veQRDA2fJSXNo4/
Tlhzqss8xDqKVRA6s0hZINynGcnkQ1HQVqv5XVtwuJyADcmG9nwqpCwp2S+n2Lux
rrcog8vBuiWd/Xia1ywg7BJF+cm1IMl2xn7TN/omiy7CQ7UMqqkdZ9EQETz3LIeS
`protect END_PROTECTED
