`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
16VadTRL0qLwHrxkswZ+FemH3Xn2HiRKPReMBwcyAL0HQiHYWGrHamNpLRmKndfw
wWXzxk8W78zgkCua0PZmV51cEmyB8X4FLzmg6wJXKrPq3U5FnWvpInr/v2aGy/lu
Va2O4fnU4bK2r/iMqezGsRsOfnYnnygl7KzaiYk7ZKBCKt55r9oCRnGWa3CXyzgJ
f86GuvSIxOGMcq7heINfDbSQyAABsTOq+/Z6lve7lLmm+zMvI02tkEytdm7JINcw
6pk5Riq3U4o9xG7I8dWyah0Kz09Ket779A3lISVJBGR8LR5W05lqNc6MKwEk4omL
0GdYUOSIjj9qtWcs748Jtmr4N3mToVVbryUbI/5aL5l+s+Y50IT9czBiQC4cjuu8
3imVCRvXXTFmc7cE/0t3tF4cXELirsYFVjJdaM3FOg3kNdm5pH/XxDRrvT3G5Ppe
YQ34OCpSo4FMcLZIm+/aON6lcDXdygxg9Vg9eHn3izqZ2/T83INroktM43P1D1RJ
fJXovBgYTU8NCj6WmG84cM8ecSUackN9zUfRktBJ2xRvn9vVPpeC5FDQVz7IbmKj
`protect END_PROTECTED
