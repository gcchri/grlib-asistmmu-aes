`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
69LGoM/Km1+35KnBgyG3GsvBWRZt+fcyn0j7I5FsKjiP3orbcIlXHF4D3viIedfd
tsCmzQYedttWoqH91CClq8+N2jvA57INIrgbO71Iu7o5cj+nB9ScJjQ9HZXwS7xT
0kB9oCAMaFr4ydGexuhWss0ZMTpdinNcXkrmI5pLf7kMU1kN1BYMCh5Rlmn3i18W
eBUY6jChkUWVUBs0J1OM/I+O+mIFaBYx5jxuEhHTm2+scf74yXPVF7nQDVaB7TYY
o60BxSxb2TJ3dNXZryvPAGO89dEaUJI+DdOt23HcVGQ=
`protect END_PROTECTED
