`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
koX4jRKKC7Tc/CO2ijhG7wS471PB2qsoha0ngmlkZV9CBVFcYQ6pQzivIiAmy0MD
dJioRKUIubMb+mMSoa4AhOrP8n/mFgdd+5Y1yMeZ7h2pOX9SRRNF1lczBR9CukYb
ft9P84pdtAMA/za0rCtvBHaHXRON6MPSiwssEIxt2NAt3JuMkahv66QbGO5BydjE
gZ8t2kT5T+HMRM3aqawclyKfAIdmUMPZ9EQ7QLCnJ2Uma45ErQ+KLuZ1gZ321O/B
jtekINAd/DxAFypK7vuKye/iPvYIAdzBK1xNn6WUYQ3sULei3JSqlBVWoZouZrsJ
`protect END_PROTECTED
