`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JUbczb04RzXHBYwE3ZoDNW1ijT9w7L6NnengSyZT++X9AQwgqHlwcQ8QAF0pASJN
Mncdd8UDlarvs5a+rbojl4PQuwiiyl6fMN6u6Y/yLKbfuqZLfni1pYHge6hLmLTN
GqSqCdYb0FZ9YhMfaspSzrozlkkX+yxMMVWFWe4xbj5s3zGl9DyDADjOwEnuhS+Y
8ISOmokBQBNtrAHaS34oRVqI4OHqEXkyS6Q0IMdu5Ef4BBPmcxEkybj0NDjOkdgT
rrtNBDHZoBBO3IBgSqQp9TYi+uXRsYHL2qyeuBn128zVtU6dhYdbHqdpU6AFWyNb
PRW4XEsunrEekeLJMxY1tScJKJJOwANyfjFcMDWk1zvx2e3o9wjXdDwE+33gGGc6
yGMQdCdU6SVrMfGfNJtZIps9kL+rkEKgXT95Gn/FoL4IIGeW+0KwidVcxVTgpYO5
OXBFHCf1sXBjSmPFzZev5nWJPVHhkPty+abpfz4u/bM4DaCerim3DNQo8g8S+YeE
DRRUoMoog8GkXtAufYKyUy9wT7846eXi6bfXwpIRMOXQtM8GJ53Ip+0VJ6NQgcr3
m8a48MHqcAwc3jQkKCPDzQ==
`protect END_PROTECTED
