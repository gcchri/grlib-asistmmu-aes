`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UEx72Fv6i6OdNXYsApezcJOkY90n5GZArEzcrLEYUhUrUSKa8XDtRzkWBwVmF083
VCB3diaxH7irazXICM0JDcGXPgmopcdlfRIH9Mrpg9e3PpfPZbSK6PEbbcvMvxJX
kVdHpR7I2W9ojSukh6xO6t6FL+IebXQwlxoiuJoT6EnraPXGMw6kB3kY8PtL+tnN
MMKX21YxcAc8t8GW0zNiRcw42g3mWHS01yakRGkxw46JDbDTw+92CscAeS5MgCFz
0XWr122Kfk03ipIGrArx74bQXqXVJSzhtk26NjgAJI1/dWCHufXVf3x9UtdHiOx3
t2uFuPqLTerkidHZUvitTGNpL6QBD4aMYW7guc0t6c17PdBdaqCGL3n1Yp9Fr22L
fsnNa8lIUYG8oXuVHUMBNHPwqg99TdwpK1jHbTF6RqCJjJKST0jrcThj+dQtwBEe
`protect END_PROTECTED
