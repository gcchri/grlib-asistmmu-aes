`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8v0QbOHghDvdPt1JBaIArOSpsQqTyVpSJmOE8poez2OTmqhAIm8aYRz4RYWzEPLy
DytVYb7n9kr11mCA1phoCyJQ7D8jgNX0/qy4judVfvjjOZu3hm2C3NFYW3th7jWd
r311zqqmtlPGXPHr3YGU4VZUnLqtPzNR3UUdHmU63/nMDWzsh6mY1jH2oVoU2qaf
m9HS8RzpESh+nRRB2Y3eFN7cWhSxlxSLyDptMLGSqydry1B0dcHSLSRGUw83pHKY
+2K/GpCJo7r/LMkXY+80UOKnZyKq9Vo4Mriz6Q0tlNCausWR6A2BNxOrDrcEVa4C
fbNniuxpYSNo067PRynlVRItAfaFqkKn/X7YbQsRPyoTTqLscFNz/ez9pm8ZTFcv
Ez2zpwDvYfuhKBymr/M5hDyg7TitDM3gb3YC9tCae4zC6XlgZlA+/CyCFkYry3b4
dVr6CUgOMMwMPN6Xn30vHVnk+p1A43KzzPBQcJOby3YRJJmui+Iu/jUuef9+gnVe
CtKF0dt039MPcd3w4VheJ/qt/zVKp9ofbXOxOtaoqCPxUrEmq8Jk+nE+J6Qet6yA
`protect END_PROTECTED
