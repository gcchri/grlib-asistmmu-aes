`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OwxE8a2Qpkuz/Q9ZddA5iZ96IS3SFfSBEgiQtOjgkmrdJ/hdZBjnCDhDiWUR/OIv
rsc7c5JzkVx4SlsFxHMQHPJIH/IsbSO1HcM3bvPDH0ujAd0dVIvQIVzsh2Q5LxPr
flJU+jvzc20r3qyLS/o02fmdKDZjDs13SryDyQIkHnbPK5lzeYE7PuiKKH6zw5DB
u2vLkEnz4jcmHeAmEFULYRBOOwwGpfkSbenA9/EGmY+J4lKn4tmyvRI5ThcbPHtf
ocoT6yfWGJwAGSLoT1sXSS5m/xMFr2WhvUg7AORWI5OGbxJa3QxYMvt6gwjpYZUy
bRx59R3DvNTAStyxK+BLsg==
`protect END_PROTECTED
