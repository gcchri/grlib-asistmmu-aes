`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vw5zhTUcNgWGLf/w62QNHw5S3lhQq6fVSFc4XTGXu70fDKHMP6i5+/I+M3nzQ+RV
2/KFSs3chQJ98TH/PJRasaycH4P3F3JjtwDbU6DYzAMsk9B4mhAR6HkvHMDUovCg
PrWXnNFXDmr0zgCEQQJXb088CPDl0HP3hpbd8mMc4mFCmD8I7I8wDrevtTDbrY/h
2JmkJmOyGkKG4bR685V69daVmuLFv1ze7nFYeQuoY4RLJ8sdyZwUc3fpo5oIQC/U
TGmyIm4mqTr0NysFyadMPNyelukdqCtYAhTe6D7J4T55RpG/ySqGT3deqgosUud/
s/VBxzVNYYxwRWykYZXsQ9v7uY+ne8yy6x2zi8bAbp8HLKIAsUBxLbdTqzFbO1bd
UPj7Gzu1THdiuUbHUW9HTXfX9l0cWeGzZnRtRZEzbHfMwuvDL9+Dl8b1o5kUTWWX
MWeaNLF5njywqvjAFfTxujg7TILw34CMbQSKYzcBh9FKkWJE2h0Ns5MKGY1FnyHn
zwlDFaMSfz2c4UvFvBws9OYNGQKQSElGg01XDI3ZMPHOfYAiWtUqKDaiJK8Um2Ca
GscXVL29AOQpUlEZ4qP8oxfWnrFriY9Rgo1XYRt0F7vK+9sog2lrdF/xhOPCHtXT
VjPLln03qysKB2HAbhiWECokGyCyHwlTOoLxq4dg9ccOTyZ1wXBJMCFAeKRMlcd6
j1F1HRH/WTKPJ1Db8y1CIdELOeJ4xJAGYCUYPK08QAoEnXSFoeC76NW0XtvJGGLk
tfblDsbaArOVJ9ktSxwBssXV0PW60Hxz1XiZclMswLjB4Ii/VSMS8xZzao+KYWss
7czqOGFDR7zwdNosSbLPKmmydfF5oENxDxPX2SAlQ/lJrcbMGQNhemo2DJ9ZlhWU
cjnvBDejy0unBognL6R+BL5nPvhdXaoQE9deDiLfs38k5aIHJUa+vMzdNWKirbwV
`protect END_PROTECTED
