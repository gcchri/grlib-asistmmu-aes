`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CgmziIjEE3jcPdv7KJ8twHHZBUk1WRVpgfvmbKmGkTKLf6BNhgGXaFR1hMQh5cql
J8WeInpofWLbTIyge+rMdNJ3XGfmN5udspN3Dd6HTO9P51OkuO+PiqzYgc4l6dfC
EckALe5R9maF0lTnOxKkkXxwZ5RA9GY4eK92jWNS3HR03RYrAMRr/M20WXlUymXL
bg+0r/c5G0J6AFBCkc5oJ/jq2V/Oe8Z4fliiNq/+fV7yd/30LrxNNK2KWV/JjNBq
9iiqNxFUvzTuL9/vLeBdCxXalWfeUiY9XUeyeGkkLjg=
`protect END_PROTECTED
