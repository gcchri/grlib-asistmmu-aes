`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ym21hPMTtsdRwS8X71xOZ+/GF/v8S6ZdiQdt0R/mtPiJvMXa8b2qbAzCslKZCs7
8+SvdI51taovOlMVikulRj0gjsyhFgLftPt3iFIYq/MzNLpB8+XB8KQLxdLg4OVG
MlhxmPHTpODNsMOJs0f6GWxNQM7/TMBPAUxdfupiBstImx+6Qn4YkNXimIzx6OAK
7ZXsHfhVsDW/Pz5PsIIz15LXu9Fz5BQG++R2XL91pe9pLPapIVCpwqdH/FEtcd3e
dbWBwAzQ45J8ZVXMFO9ccYLfWnUNZjgU2OW8oWjq41bE7YQ5HtkJolJsQhYptVni
vshBf5aT+dnzDNI2ssIMo9lMF1cBwG3rOpqGOQYagUlsG7CckkXpPDOXiznacbVb
I74EwUmgLdoxZ66vsIFBEccGwxVKuVxXBYfpX8ZmXc4unU1IaDu94F3ztfPebaPL
LSXqOiKEfruEr01CiGod5FUnOW9LxwVzlsetF5PQQq8MqIOnTBPQPsYUDWko2WLZ
kTayfRgAvppU/QxIr0mo2riNrNNZieLbJt/t+Bu8BCzT9pHgvAbQiVKjR3+KcAy9
nROWp9eTw0CwXqVgFdfrAEgGyz0y+LMMhU/7hoW+67zEhlgoumdCrJHeFmsWLL50
/Jo4ZgwvzL6OXCvdrnPBwA==
`protect END_PROTECTED
