`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q+z3qptKayvHib5TyFhhUPhf74ZPB+lHA0P9+jwZ64KFn8/xdsbbz2JCy7JY8wYE
XM88L5DZ462WW+5X5JMciAhPddhrXcNXo5nj+kEZBlwVOdTaY6h8JhWa/gQDXm7u
ZYV5nvq4VuJACzwWFQdOsoMtCT2CumXKNASG/evVcpn5hICafRr0UiEhuGpmJbEz
ts4qpjgGmYlzlqFL/SRwjg0o/pui381D44NPzcd1oGMOrYrZlpFdz0F2NnY1HAdD
Ez7Mdbq7j+IvtJBZ+Ptxe4Hd87k44kGBsj3GUOir5oTC42MrwhEzixmoo3fj8357
8azfAk4nVQ50yEI+k52ekWPF9yBRRy22Ja8/Ilx0lGLphMgEYCgDoiB9OdAGya2+
5sU3ZXjnFWHt58EIoamzvx/ZbmX5XB4sfquWZ0hEP2me4agjG2ljxPKDcxnj3ZDZ
9d97vxjmPbhmSDKkKNfIkeBGTd07gqHudl3YghpGIvkE4o8z+dcsYiNJ+kaPIONJ
GYmxn1dNEChiD6mvP2D3JGThJ9N8QkPSWV2K+H7nqS+D3EAqgh99BXVXkUhYAY9l
MDFU7g2S1Px+HpzXYLw+PIx5bkWIQh2vwOtpeKYx+7G68l9OQWl6KDC2m+eTRf/A
jL5GzHEGC6EMe8WIeEJ4SnY3Ad+GmOds3UFT69p6DhLHnsrNrUl86cWduzYEV3/M
x981cUeYUXLXwCa6rS8snaYeJ3ZRe5q9dGrqjAS5cUNfZ7z9rGE5zaccsn1qIrt1
b/MZajjmtQtTELR5Z5Cjusn7pC8Q7RxUXqQWWMKZEAkpnrQ9mlOyjqx57jSeVyic
FImlz3N8zQGO/sdssmIxc8ayHDHj0v3d12APJElS00KmLHM5nBoM9BZ5MWfoTzVw
CVZhKLjPrv+i5vGtCR0FvVBKtCSoBUu5D70XIgXEuvOpEE5Cyy6IrwzEqLUPH9VL
nVWTZnIJnf6fYk0XtuqkARTubEi8loJo087tu1/lpM1k3O3EZ16m9/H0VngLi0sj
Y45SmmX9jZ6urUqDH2ww/B9cvwn62rX/plX1ITEuUhqQ65omDJSIJpvydlSF0ivg
kGi0RKRVCdt4cZi7yNqWAAETG7PjnYGE2j75GQtOg7KmFol7/j0cdTsWlesO44iS
2sMmHBO9AZyH7MxtFF5cnzXeRAxB8mHjRW0Z8VHDggat2gcyuwHAfKGSxfMcCBuC
x49EwFqRoYC+WGwsqLuBIEMtzjmlQh8thuzKF+MEVt4xl920ccUOElaY+fCjD4lr
aSksBoKZgHl7SLrCJamwi7b03s7fhEbv3r3THQ9lxys=
`protect END_PROTECTED
