`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hp2HzZ+3AqXmoJPJMog1ePeuKnpERKhkCEB1KyzNGnMPoTJeOcaJ/7Asry9D14bF
foXwy+Oc/uP4MVCKh0rj349JOW7vJEfTP1/m5NF8TUVFLUIU9Qm/Cu/Ztlduznqk
cW6Izp4YBe3QWeFCAtrtefFpwMEQ293iHqEJ65Zvd4h5RJovaf54oxbEhr4YHxHi
4ZxvleJDPXaZXBTgnpwtGTzoJwUYOGscLpklE7yDNsm+RzMHhyU2LTzj0Bz16HtD
3kKKyl8vvJNxQKZCq1zPSUa4bALJh4zGzjxck1FCTyhINi3tqfA78bLTGElgEyCu
xWxaTNj9y2y0aJGCxvGalr8J0fHblCMT4PJ6eCflj/fFlqfDNdNPRoyTsofJZiH8
cib2CyPhNPPxhaAWTzCek1Z9cL4sYhrK/VLlMUlpEdwoi/XR0buT2czTwK+58T8B
PX92WZNPiHXuZ4NwMap5oRNfk7KtESuHPt27Da9mYJfUpqJaRGlA7nhIpSTgu+Ug
Lae2TH7DkugV8KzmULNrsPwEsH/hVY4zncAWQtxVIKvKbazMfsTu4ewPlYZCNzPG
qHHC/RdDct/GXUfl5J+PaHL62MUYCXezViZTj2Tw1C56fvhpokpkf3olAvM3jFJX
jz/hUe6TZ2dGkDCPBwJ93MnBOtiv259XAKr/06GkXb95kSwKOFUaveHdD40en7DS
djPV8dj/jRt3he4Oa1IYEHyoX5/5Pz79HvKAgTl2kbyH/+gKja/Fq9WodXtuG8OY
iHvLgOPDaFcENbxErKnVgUU63rkRcpDbNhAJiCZQ5mRT/it/bkJpYmv7xZz2+KnY
UqZ3mzYMd1JBPdon/AX37luWWSpA59pVmJTJMaqZ6oFVubxRRu5TMWMCosAWJ18L
UI8bwPzNYNTF/DSel20Vb5cnJfheLCK4euWbpIaR/Ez2xBB55qnRJYuNMn1rPH4E
c0m1zmJpE61+JR0tI4iY6DPHyR2/TyLgYJayP6lu25EINUmj4pE2aQHgZMccOlHD
Y5DrLfqQjsMHOLlbG62bggbxkrzgxdxWPU9HW3mvmdYGtX/K8OaDXciL+UVIsQdh
ZVOcgp8WmmnAbb9SZpWe2vLCkBcrlqz/mbBwCDuvphDturuPR6XhYsBmzQmu5MmP
kVNTSTyXJ+MBKJEwOpjFPSo8xw8vbuJaS/rQXwSS+gIoiYZhK/MNBe29ByoEju6e
c7QhDkDbl0yMnDtsbsD299/N6DSnWh780A6UuxrhF8ks7FWd+LKtYALWxgugTU56
qy7d8dEAxIv7wygDqP90DcHrY49MgogAzEqQdHQWp78rBL7Afd0iNzL83y7qVXCL
uGCtkZM6vTYZzUAA2HRO10qrU+AfJbbH6u6Lf8XnL+d3katdtpbbIiH/54b2Y99f
e+pLMVwKIhU+4NCbBSKUmQ==
`protect END_PROTECTED
