`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G8Pzcbc8dKDBDi9rRbrkavZqiDm2Bdtof9y3OfVq1Ov/hzxEn8Qc4ie4mz7JkjJv
LVYUI30mUGhqmP2eXo1PQuCUeXgJ6hg6vKn0ck2ATQX5w8YXw+mzr+MX9/nTAakC
bWUVkUFDrM9Zu0CUy0LtUL2ohEll3MzjcAbcAfwff6kwFZBD2FXLh/1XUz3JUqzn
z0eesm1qIp5iPnrbQzMtJBvM4vHRk8GuEqXWs61p7u3K7D3Ijx/KIg/P60nBx61K
QC/pz8JQUDl+lpx8uWtDd2JfMQUOsyi0kAFHfaMfxCdncSsne2e00cGTbZQDjgfE
oPIoC334svM7BVBNC7GGoukbvX8knrjmMXcjQ5a1fe0BUgYvSb5WbJBo9HsvzSDz
ZXlFwmeFcjSLeJ+UzL2iVg==
`protect END_PROTECTED
