`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XXy0tv8NGLD0ngkh2m12SqjytqR7jZMecCnOBm6RbBAA9vS9lQ64VUYkhVXUJwVd
1qOO47JsoV65f6Rp0sAdd49OkFNHp63bjQr/LGUMrLLC5fKgPlavDjor6vCp2/4O
OJ1SJ/coLej+NHFdcQtWuNcg/8I81fmW5DTXchANRvSnyxPN2zqy7mBn+RfnwUWz
BM6v2hjVS2In58sdMjwvmdXAg1nkQTRL8Z0mhAnV3o/xN81VuFrVSmZHe8k3q9kI
r387qnJspKok0TZKSHROVtSzi78Me0lTnJNarIy3CzfsmxverCJd1wHfXtRpUAO3
aU03DoSbzv1EcMk1HVXfydRyuTVUw+WarHguzcgZRCtDVq2Zhix66aWvgbWzovII
veJ2FNTdsX8Q4cIhCf1slFvWogqNI0Ma1vufJaKY2OhTgO+KplIdcLbH03awojbB
`protect END_PROTECTED
