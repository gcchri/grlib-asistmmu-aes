`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M0eNHgcLPzk78puyWl5b4l9ORIf6Ceu7/Cd8lawduCC9huI/EWgzohtU1Vwvyv1J
SSRhvCuRnCP38NRKmY+TUmpQkdTtQ/BTqdII7kOSKyOEdF9rZnmYcaRN3aGCaBin
ozlxVV9L3WjSXcSqWimgMkcGmsx9k1HCE3L+kO3gLvms7QKREQi6A4XIxwFmyWr/
GSq8Ca59vgLyS254wmXwK+5AY3wiLYYXbTIaFNQpGVa9WYeqSxKGVUXt94AaYh5q
kMpRrkI4ggM/uqzJFWHnJb5jYQxkokRT5ba/ZWOTFWpngMClxSNQnAC+Lk+RQQm1
NODV1YZD7TMsZlQuL5H6axMiFwdiQThVj2/isyvgaSKS9TWwRG8rIUZJ4+tCoKM0
TaIBV0nArrrgFVXJ7l1c7vo/dfYadDpajP9oGW0jMLUjhcDx4UlFjDdQrTR4E4+3
f2qk6zENGQTFNOM5lWuWyJzFTeKPSMNDnO6OqeSP4nSrrH1hmVAvTGWZLBsdFc18
i/H8o7TEzAsYlPgbETqPuDF/xa9Dz5tW85yyr7XCsbA=
`protect END_PROTECTED
