`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s0aZvBI/YRQRuk/AxWB34OScSJHZdGcYP6mCbnZE5PznEqMoC4BiuU+voEUxTanV
iW84rT6kGihGAAhi6A9HXB+pbviHbf4TKwZQ0wUL+VHWN700y+O5Leoy0SjYGN8Z
ejpO5Kj7Etr6gefq71qw+wRBDAEhpzwI2bPRuU+i/6wr5RUiENUhFvs+fwVUNO4u
hrnkrd5aU+MOw3/KEnRf2NV+IYE8boZP59eJwvgbDtOIg7rcunPMXcEBd06i/nG2
rYXm+dfDMUshlN1Lc80cKOaSVldchltf//GlcmEajxv377Kpa3KmykEKKnwtxX/c
M1gzSAfG28QHnIh/29lKCPc3/iXGFJGS9DU4B36PMbiagoW486MPs2Cam6jqWiqz
qUXUYswOfzFwb1dfOXlCCxCn0AYKCY+3tW/sc02ShceIHcyTJokBRLgUXVp4Q7H7
AmUQSWKQc7/uxd2pdMcTTEBKDwZDWTrwScqhYCtRTFTrK6dEGrZb6H2UgUldlZ53
`protect END_PROTECTED
