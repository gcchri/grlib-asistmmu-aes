`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jjkO1L+6itXnJDNjlHODhUrGvyvF8Jl6yPMmVfblqNn3VRBCWB7O44OHtx1EuWUT
QgZO0VFN5AgCnZrnuMUl+zWr8U7bngQEy+5/SiOvl9EHf2mCeOEpxGIwdYzaDv6Y
Jqt01w5NXjhZY+Sjp/+ghjjq0V03oDTMWfOL2WbVtdntiUlKMy2mDp1hS9k634gp
t8JJimRGvoWfMUf7tNssb7vhwGJn7iLY09T9qG+9RVn2w6Fhin7INMxM04TGfulm
JuyM+/ra9CuPTgOoiLdeLQ9Xcg83tJ9JputX19PAoJF/QXsIHvIJzXEjJCZ6ibFp
zGt5eeHegnPOa6DrFRY+JMJ+uynJfuwoGUmmMYJHFbHdQcna6XgNc+EezHadOyPo
C+HeIp/r2SGzqfUj6uJzVhEktHx9Y/lAmBSlEQd6DmnnJwTgt51xpgJ7n9jrLuwU
PHkvwqYs+BXtqpuSSbLECPJjkN7SMAwOU3+9dDbNOFcRGNqirdQhCm3t4Wsmxilp
h9DgDXu33MBjveIvFoa3Nz4wsS0ZuGST2wASKUn6Q1qJxLPwmQF6E5iHyjiDNt/f
ulAAN9Bs8+reGI53pKJ1SoZaTLRlgCw/NARLbypYfEUIVCFyFEaw5YZ9LwQ37iGc
sqPHECUO+FnwoRORglxrjJv4iZ+VvbbmOTVtSTYb1RxEqyTt52A8Hskta9+wGu5u
MNlvUnFuFI09G0aw3nqCg0BSnF0UIsc3VSTuFhZP+m+OwEHl8LEtg5p0syIQPdaX
WrwJkxcR5WVa9xxPRYIfb1EFwRv/wWDK07+QiMNFt7g5bFY5DX2njZKbSWUUxDVa
3Xb4BMDlgr5fnwW8xZUFtyzwAJ3c7aW91dgXFULcg/HIDzWKmwVO2OHhlEvxVLFT
KXtl/Ggt7SsgzFAwpa6FXzFOPq+mVE5YvEYvY6cagl9XU0WStBS4wQ0qkc+BbLpw
IEs3AsHsJmNtOn3Efqrqzyuus1iTP1TXePv28DobrRtiffRAhwkJHiG0sOMmGB24
nfrfLIOWLF1N+NQATde1dNWZb9R+O2HaDc3hFl4uXbcw4fzvaocw+Acxd9q0lGSW
Aimji81KVeqcLuKqIDJkfc2HR/BWiDB9i3qwswINxq0I1uJEAFVQ6mblUNSMFEfY
l7a1rVXhRpA+iXGopDqFx/Pkg6WE9HU5kvunjbR+fPc/Vi3sO3kpaDrdl2sCc5+L
Vdekzdjhluvyo75UYW23IhJ4yp5NcDYjRCQYK6fgZCPd97hdgofp0/xhqbEa5CM6
MelvcNUaBSX1O/mCVxOL3sxt0v/GATZHWtFWKwHz8j1zwWbS65M0hrsQBkhDzHCu
wSa0TtDb4tc20vaAWiPW16Wkrj5/NoiNz6AyRsC5H/+fYoDAkeV5cNyC7XVIpW1z
Ni3QvoeW3X1b9RiSkkiFtcN96mtRPFOb2vXYToECM3Ntw549KArSunx2E5FELGOP
V1RVyK6UcJoPaR/6M4FokhBIYVH0TvFmjp9/iJQZ+FXTz3bspLk0MaiGQhsTnEkR
lYht2Y87OXXy14G8g3I+BLGbru6RMQCOxCnSdeNnIg0oWhLSTT/DoClwbwLV6MPQ
Y24gKuwHoZiN1KfShQqvKjIPlQj9uGYF1adoZM/Eup/0ks7+w/1KigzheEDu0Pf6
mH7hBUVx0LabL3fqqXxrNa/Nu5XAEPY8LTCyLaUESH42n0r476/cezVNgPFbqucA
gbyJF8PUd6cvJPDhDb9Ed9uX9J4GIiuUIgEY3JSFDEgE4Wep5Qq3kBr3+8qKBQX5
7c+bAZFIPaGBtO0fMMup77aaym5XFVgqNpXzc+YcLk/lO6CNZVSyfh4OHpgx2LRR
+JFpmxhEaI/jlJNSJudh8QFIcQJ/FNoUm1dEL3iiI4KSacfutMBGbww5T69ee2R/
ufVMIEVVRjJCyrfJJSyVuyTPqlWMcDHxHZq+ZYMsmOpTgSibEzMEao0dsu4rJ/n8
YUfKBQJNQufZlDoWT2a4X4JQpRx8KtbOehFDxH7lM7nlKNXzwXbxnSwAfuJV0O8r
Z68W9K6Uh4vSR4N/divlmEKCTI5XXd/8Sb3CqhiEv2d2sNfeiv4x9eu/DPLl8kAb
Rn3uy+1uQ0wNnZ2EDO0hnrTW9uBX7zhUyqBu9wUFYdAtJghOapOLDXaGRQUPqBfz
3NIEmkLV2DwFE4632U/cDRtZ5v0+OiZVRVZiCVlAZeKxTJvbZi2mtxD2rZI8ps8e
i2vsWn+I9Hjpux3ycZImgfRuZ5HlRkCoiOwU2ZKb8Ko7Nqg5uMbfLxmTGlNWN45S
2J2eOfqmIoM5c9H2wFGqfPhEdNpDyHYvZU/DR586Mfw1GlDgWJC+Uu+afYQ5ytNq
1cjSPp1o1ZeBgMriiFAw7c8kdcvSYUSPG+o0E7mg8URD+jflDKE0QCA+ZQmXsFph
UJc0aUH7YnpwPxkjLrmbYOEGuhrEHlllLl075t0F/14kqYPpt/XTvt+TDvg2KxDA
fWCYeu2/+NVrXlsNdKcZuSQpIIszIotokHcpET63sxMTHqcUTkkI8EAlyNEJExCg
ca317loeaqU0rgIUawuAkNJw/t+roE3ZWQrApsM+OjVsUGhNJ0ogTSMxyAEgblWp
SIg0CaXlK5HMO337tjrBvKZfOBeYy7rUHVFRmjcFGJ5y6TDkv542+8tOKAsDaOg7
3LT6djU6SJDtwu8dnlKUpZc4SouMD5WhKoq3slpdC1mtz/UGoXenhEMIFRAnp051
/vZwIrGMm5P8/wntRq29QQwCYPHHPdth6tmdTlJd5tc=
`protect END_PROTECTED
