`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qK+ewQP89YZUC576x7F9tP7v2jR1ko/HaVMa2esPbFO6jscMz3cCzJ5GbLSI002u
MclsSyGmAViSrKRPyja+xQkC9J5FeKFvSjaevz5hd0Mpd13LVSIqCK1gDKCyRM6k
oPjMvZScqnsy8BKk66y0NViDhhCxBb5TXLArgiPkQrjOdtKCFbqligrrYb+Crz6K
OGHrr1z/wU59aRywbb4QsKEj/wkQNJRoya7Iuwhb0dQen83bFtKGWBQ2LqvQXmnW
Ckxb+Esw6FK18NN8W14ak8vxwLD3KoCYvIyyWsMuBtFirle7QRuB9BqWwGzii1Au
nJOWjtC3g7XT/FettU4OxJtqWg0Uitu/LeA30jm+2m/B+eGqB+s7DsNBO/ZmlyPB
1ejh5qqxAvjiLCuExf0JseQCjGDnW5Nhw/NMINocst458G+RM6pFi/+i08mvt0fN
DUFwJz0Nuh/gz9SGwkSzc5vDtRIR9xREjVLikdu3SxIfoRyJeqahcGp4BHDSUNf+
JIh/sW9Y/RZQP8waMRGvlX8YsnXtdqIv82jh3dxHHPSCdhd1avhAxPziYHyHcIqr
EkwScaTh4+YYznjA8KiGAovFf+3yHft/dgq4Cy+SC/mdj5JAVcNC0XVSR/xGDUv1
39JfJ/dzwbXTqNkL8Ei1oWo8BMvEd8ts0xjDEUKw5c7zQVm7eEHcltf3d/QWEj5S
jb9cQax+IiI68s0WTsRbIUpu7ULBFmiSs7CcwxwHcp1Oww+UT8tteMfkH7ChqsuC
VNiqFgp1s7RYuf5MHZWq9+UrKZn6mnQyS8GNk+d7s+86nt4fUPLgc6W+e9DEAQjw
mevv9qGLICJFszZjj7qPHubkN+WFxtH654JZRds83uhRMI+PwPYaQTe0BEMQUjl0
wFx5YDEkXJcmJq1aq2W7YpipBXzqevCqB7sWh4bDoIz8vfpRiBr8eYKxGsebTlfg
EhJzkxvtjbm0iCdFegVevTUT0AYOXhWDcNOkrp7Rhof5LsVT23ZWbY1X51PmQpTw
/94586eKWctc4Ac62XyMkax7A9d4+Swm2iFG6GAmcY+U/P8Ah3/MpU7Rey51kDIK
RqteF5RcBYb5kxMWwkAOmSfJ76EByxOv0auNSQiUwURGgn5I0nOtKyMlotcFAfQX
`protect END_PROTECTED
