`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SrjhWUgjy8qg3Ub29tfuz3chdWyuRj222l3FL6Qv/BGbALNYCZ7CddN0ajYr0zQg
JpOp2GE3HNb+JK6RIKP91RwFhxG2l71UA43cy7H9Dhghh79LPgJTQQVLsWJT33FU
QveYK3xfdHz3Rj6CfhauLlIfWzHXnCsXRA7xZeV7dr/eaRlFk7sYVpj7JFdmQDZs
xajxfjIHC+/TkXeexHAfxU6eYnKXn48BUuI9u+JgeVjhB8xLe6YjyFrRh4zW3uDh
`protect END_PROTECTED
