`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uKkXYXcfU+74AJKeprda5svm1njcQUkSUFLzuBhFjn2tAj7I+9ngnI/plI6r1R4N
he96hykdM1aWfgkd/Q5r7au2+ZZSNeacC5DthQnqkVtRwIrPvBvDKQyTMQLZ4WOJ
lYV7lt21jrrmrWLi2c+QEkjjWmBfc3Oj1Zym0zHllHSxpJuaLIniQfAxFUsW3Leo
CUAiON9nqoBAXsAhzSdpRgUhlkxWqBTq//60jBNSwElnrEgjaOVF/5vx+ia6Y93Y
SkKDUnuB8TpM6R378sFl12LQY53Vh8h8fIWUIxlHW3pXAUsW9shg8X/09cm9KyKv
NtVk1wylXnl9uMtNK2X7fbcpe8FJSwxQfC5k60AP+4g17YN+bQa2vTT//6RyvZ0V
fYfSIERE6UNQ6u0evZ1SHQHK2culN50r1CRrdkIst3g=
`protect END_PROTECTED
