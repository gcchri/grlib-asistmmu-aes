`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fEMGQquCsl9VSnHwKbdvE/cSqQxEpqaKoPhc9hPN66F8h57G8NY4T+F6RZ/w1L67
2AV6wyKLgySF7X3wDKw2mSZ2MgyN/9vWvJEqu0Qs8ceRPWt7IHxZRmy95Q//GGn6
iHryge1ZHAYasIjUC5CM6YTiMvnKv2XafWrSfKD12lfQrsMFhTBt+GAYPar5twcg
ID93QDhhrx/Uq+bsKE0ndP2CtMcrWVwz4T0itKjkDYiokPRA4bl5coK1dstH8Qhy
/L6B6hJQg0OeuDBCI0Ytkav7v64so315fdHYExppRr4x+muXBaOouMiO66iVTsQQ
XeXqxR5f3Q4BLqsPFblVvWV5jqYHYSR3VX42rEQ8Di+DN1pQ3zl5wysEYW1pqinF
XzUdzMckRGvfvu23At2+guniGRgkrRxlgokiBceTAZk=
`protect END_PROTECTED
