`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BfhLsLD+4fiQwl88EHQ4KZgXza7UKdaNcEBG9lyZM47kdlKffL59PQHi9Mm6Su0S
dl8YH6q8gHal8tbtnICxhqIMROZLak1FQLNwVOierIr3C+e2vNtu16wU50Wk4EB5
lmYIqJMKgvsmKMZAKpcLBpRnTd3D8kMDANiXr4WmogpaL7MQymtrzMs/0xJ24OYJ
prX0+ZsN2OgfpQmsoOM7Em+KlYdh2siMmzaXH4KnnMazmGNrdIPhJwVcbcOLhzlY
nSDYm1c3kZ9vHZPrBC1Nuvm9scHRU61Spwq3Oq3i7quLsoUOJs6vFVLioKZNDTRP
hZJKs0vi8KofeYw//R7RviYGtbv8Kbgt5OvHYEwUMvpE6qr3LnFGSfSfx8EezS06
QXVitPCf5i/MdmjtJEfCOu7a1m8IuIgOfxX3m+hV693nCKOodLq87YFJrixgkzmC
WsFKs3e7a96mR/Rwy7VqI1t2YY1IT6lVv2yPMZy6+U6k6MYtXDKq8tdir2cgZ1hq
6/8bjBzZvK1wpFJqbsHZJ/ZFDZ4jAMmEBWuAOq2RWpJNIYNYynzNsgkmAWSsvtJ+
hn4iUmUjaBARKKVjjo1nZ+x37+ffKkbOzkWUgUHl/YSMAxMR/eUYKNNW2bYOwX02
EfDbJyVjDwPQRmkVzt0lDKpqpOLS/ndQ6kjbqHTNcHmUEk4uhLTexWd/eoB4zvVP
ZmJXFHU5wcP4/H8Xcl8b1ABLwrlzd4W619zgLkfa8Ah50vpjUwaqZ6+8tYSLhgEo
cLFpA82jxhvmM0DFf0CQAFEmogNE1/cCfvZ+oohCQXvJFUOou/2lpuFOGfk6wXqr
xmFO/jopPfZkFw+3wbp1zKIgnrlt5fdM9zmNDSkRgwrqWvTdMm09EltqjlVvxZMF
PurKgOLOTchb/ofv2/tJ7zPcusfNOMmLfO0rS+n+xqbNlr3ox3X3bMJp4/UsaTDa
OpS2ACl/lNnaysTeLNH9ZSYFGU50IiFpDSR/OuY/mD+NSu+/EMREEh1dvswpi+ob
lFhT+ogaSV0z23vqotZzlC8IhKF08WINa7q8dRQWegP30PbDtxQ8goR3Ybfi1MJh
ZvsX+p3n30lCI1CmKSllzFMHJcMZxVD2POUkyXuLtU4wguKxQ0gq2bOQ+JZIHtiX
pOIG17hg22EwBN+zNNE0Qvm+XXxq4sxh2triGscWQDNU1BRZL4xKfv2oObcpMuey
EVKfzyTA70vD1l54JDpcTrbEN4frty0HvhPKXoE0Vhp6nhQt9XpApMDFQJqHw1O+
winqguUcNQpIbsmpZsK6PoeSQRHf3FmXWAkTT/HUu9vKgeCz1uSFCNLLerNw1Jfn
hGs5O2zHvXQut6z8TN65CXqlVvDlCp6EAx0HxJ6tZFPhpbqhwOOFknjgPziuZ2VM
fqHmOJPBaA/IH1zEe7FT1Kl/LkmP+AOPgwk+eZU3hwqWp/9Q8uIoEN3g4fBaiIo9
jUpzCo/XP82keK700xa1FA9MowaGN1sv/3p+Igc+cZk5p9sXVcnczfIdYvOvoKfm
0EbyTztGJMEoH/vdydIbI0BVbFX+Qr+hxp/LNsosmos5knLW8jVStoJ9vZnxJJtR
ncHe3Ja1Tp5w7kmNNFJd+1rGdhxoWPLCkudL70NJrlAQqAsJ32XMRnJuXR8xMsFV
FsWYMLwljx0UJdvMiyCNOBvr9mplIrMRBDFSKS88Hp2fp7mvRo8RzhMqibzdURzE
TlVOQa6Br6FOdZYaxQW4tfeDAFhvJESZqsn/ktLeURA+yMCr+HdYcKB/JJRBD7x8
N9wg1EgJ7uYXhC1WNuct9iJ9mUErgvV1QSNsdLya6zwU77ER6kPb1N3O6i2tKirk
kLCc7nqWGhytFKhgOBFxCSP5poVJvP7/VvyG/RxpNxWulb4n5HPW+3mJs0urvdlk
UWhYykO6m8rLK4wuoDW7dtxOPDBvlw0Rs+fDdKTXmSp9rkSJKY71KEReAHa91uzL
VjPMGxmkyTLJXnDN4ROaUIPIALV+6L+N2MGvfYqf+CgF5lNfG5jalAnP3GUvKu3+
pu+3YHfKZw7kjsBFKC0ASP2ZS+FHGVOrv1rTVj91nWFabONY7PaXOi6Hl78IB7Ax
vTLazbhT5IPwOIWQtQq9rQnsMfbEuiq4L2OQW1dgp/LcERsieMMIHs7ZIg9LNOPZ
U783xb6BvAUJFwHEC4WjGg==
`protect END_PROTECTED
