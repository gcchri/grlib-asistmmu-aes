`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C5xLjy1OT6bJwP9smGa+NYaiw/SVViETYXBrNbTMGkc8OFPw0xyNSP/p35j3IMYG
0mxd9WahBBdJ4P5gJI6nI0tdOESgz/LkauuCTLUbZWHBWAe1f2Jvy8rClb1O7cgD
W05WZT3MOP8Z8W/iEIdvsbUHKT7yd3ki5YgW8r6GnGiGdpL0x2qvEUEHo84Wlqzo
xQ/6lmYgw5pxf+b5CGrD0drG1W9wU4ne/rVE70UZNE5Si2nfwaPw2o3UDxCCcnHV
MSMu0GKaElO2bLA+UyAx7xPel4MN7mPmBCko5/oXCvFcnaMILT4hHxlOxhKpNlLE
YVgEKUoAAsS8ITPC3bfeV/hgZ8TqREc1Z+aRVIjfsSSe5/NT0uH0BuMcF7UYp29l
V7gO5HN3geT5MGnWcBweptc/wggxS/zy6K2MOkk3t2Vx8jLPa5+d/GG5ckImaROg
UXT0Njoz+4CLgVDsMqKdqdQtWWBDGUctOQl55KoTKaksftc9X37e+YtfcY8yFRTQ
braL9+rNCnd6NjI+iN0aLbUn3UUM6x5Uh8mDpPjoP8TCcPxSf0Ylip98X7IAgmRr
GVTIAYZY9ZOoHSSqqPOaVqWJxRZgUv/n3ceCbPyK+hR859TMDjlXs7BiyEa0j3U+
KSnxjyijCXJ6S49EJ7ZE/C/6LguYZd8Lfz0nmDB9dHE=
`protect END_PROTECTED
