`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GB+Py28R93hflroGWk89vn7eraHm/NSxqO3LUrjuff2dCpdlgW/AahT7t2x/mq8x
2ItMesy69jereTUnnfKG2JH5GW2z580tr9CPYaeHVzD6IO2SkoyZzCqiAEswaw8/
14fgOkzllhaCmARofp11ybCUJ+2cKd38cp3yKCe4h54ypIAXQtfSkY6erJkjMjvB
3u1vMHdNMOp9GzPYJuWNOXTX9OrJFiorS/vSEooDdS0e5j1VkSuXNo/J0JZsmZUK
VkYZLzRzKdXbFYJUVKeyagZzYNfzLVCFPkBcROlmy5TyOYhjnWcCAwErM9ekJs7q
sj4xd1POLs6Y00fn3EeNQFyScWYADY6bDqcH76O5hxRrHwnB4zrctS+nBf1BfycM
AQRxOe2/oQIAYAZnRVSvP1yBKTHbA+kCM8PcmolbibmtbGzM9LZUsd3mU1oaAOsc
`protect END_PROTECTED
