`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mIWNDQwaZEc8S0xng7aiZ1Io5DC3xPEr3vDajKxuJAN+rl7TPFy4Nkae442iWnCE
29LtbwsxOxBpYWQKdT2YOyv72jNs7LxWS+TEHok7LkIHdCMaHdfhDlkqLhimfUks
kCk7lykxJ0CTJUExpOcDBNH62KHmGlELNqdoPctPe7d+AOWdpsA+KVJGdA2SP3rD
hDHOvBKeIxj23tFKpD9vUaN91fsxTH2a/BtTfQWjGw7jyDzrjJfNBpdMAepT6s5w
DGvgpEj/PVueJI4m1XvM+r1LxCg5WpgcXEXbiEWod6T4/tJCZECLZbfKYd2KkNrB
0sszj0Qu1sjEsW5nxXUM3TznDfYRQIs9nuZhqQ0HxRqYUq1AbQfmzObUtWD6Sele
tD4NG2gL4fh6yYze4zm5PHNVoW7MRSUN1mlA1mHbbO/ij8hyMKypEku8yG0kk83K
ezBDM0yzAsah214rG73uH2TkBvFq6Lkn+D5u74QBytZ/e3EZaNeQ3LSVfLzF9Uao
`protect END_PROTECTED
