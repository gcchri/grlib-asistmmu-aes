`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xBgSxHURez6Jp8/Fh+W+GJvUHsbUC0zBwMWbDZADxpgx9ZDhj2rCyA339Bt9Cxas
9AokabeIy7eMXtmNjw0oMwKnEK2m3f9XxlysC8TdY21X8wb/DyfXP3HI8n06lVqR
5KOJCDyPddYQhw7YS2Hs1p8ro4eCReXMpc0KA9+CyJu4QP2oLfrLGjQxKghuk02w
LEdrX6XvAR8pj6fIvjEhg1RYPIJmNnv0sF8XDLrSucHCie60YtQNizbMgR6cIrAO
aVf9lOO4AEwv0LEasO+YqT8usTZRFXWdckCuet3AZVF4JMK7yN8kM6MMsBmd+Tt4
fC3yVw6aZB2XLXA08bCc3I0wN4aKwsai1iWWjVDkja1PIzNZ/gZaj8zu2msIxo+3
Xnc8og5IMkilegoOA4Cx1Icgb9JLCJIdfi009SOSaZxMVcJUTzfXNBrNSrWlRhD7
Tizft1HsqPYgZcDXhqMG7hu6PFQ8gqMED0nsN3kgtf8XugEWoG7yLsuPwkTLB8cm
`protect END_PROTECTED
