`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vGbM4EqyldjA4XPNthUJzkKUXYGV6vvyvxqVEsHE2HiGiT9aUj5aL/ZcOPFKuheZ
8YNwV2ExFxVGsZSwbn+X2VNy1sZHO0sLEN15SO4vLqBFmB2Z8++0wf9HikTdiFoz
GXi8FXGt9saKXW3Xhf6UNqj5VnX1hoPLqQRl8szabgG61a9vh2dBY6R2bK4+IgM0
q+2o3vQ55z0rqpl5AwRaclkpOKWxIhqT8v+/LkqKeeguTrBrdvaPfHKh9R3SiRpd
HuS21Pc5Mj/+97wGPcCQc8MvEr81Jw5kEX6lIcKXw7QIfTyTBEpTkQlbinSuVH2q
VpURwppNZglPDRXjffDKauSeOJan3YAqE7kMePrKYLdWy1Mupmj9dE4ffiZYNpOY
QOxNmJR7Zhi3mhtW2hwtJdarkSfOed4iW5tUzhwLE4+UkSn3syhEtLd10fDcNavN
W9PgWpW2wR1jcjkXf+CNhRjJRW+U1HHVB2PHxKd16r50bix5t0QspvUVAaTLnzOS
Vhf3ZeFmYEuadB4rvsRT21S+mBhZ04Ea/MLhpzp+pYkk4Qge4778kcTX5KILYE2N
Ud0Vj+F42sEr+KvQTYgDdH1AaTznc16Od764cVLlQSUtksxBPufAggl/os0f5IA+
`protect END_PROTECTED
