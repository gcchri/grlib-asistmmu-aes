`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QtBH7Y4NnUoXeBs4tDFHstV+5UrGEFUsS5vcLG1BgJBxDQiUHjYw0oCeprMZusav
33q2jVwodAiLK1VSfQY54M3N9ewBgNgS0aXoTn4f/dos+X1bJlF2Ad7FRpJFVYbO
V+M4au1w/3DTVq1Pxyxz8LEywd1xlGLyyCe7HoumXl/RIt8TaTKYgLjpBMaYHZrn
qHx1/EAg3ByEZDzZ8bW7cQotyjWf6pdMBMUihFpRoXZNAPgUh9nRlfk80owGLhEr
JC+JPjcnDtKDIgNYI8tQyPk66VIw7R81XKoHU04rxuTA+/dYVYTJ7ecU3jKqsawH
96djyaVePXKiAvhGUXyuqiIiVJiotuKFyqZooMMxieyDbD6z14p8tRha7F3t719w
/xxfeq5gsro7p6Sjxm9OwO4PUrVXEdNt54s5c23UvoUxB/n64ZNnpvT/FYjmFPvf
lGqv9h9gxMlbiNbFAQhYTcCqLyOUsU8CPvITj6tzQUP9INlbOYolnJSEjoS8piQv
3R5RhXvf08pe2prcTz8Sd4jH7EfCSOVcgtxUcaFoyX1fBERvHRQdmssQ+RAdjg9K
CYjPc2Bkd+PS0Nl27RXufTfYg1qni5EbGPfUcw+C9ZSw6Ka36n3ecVzEXt+MTxp+
yRDxSaE4zr47zW5XOpgWD63fwEOxBI78ekFYGAFlAzLUBHRgs1CJXvAgvspTsbjO
XOerxY5iyGEhLL//LZnz3OZxErcMi7Kw5kUBIKTnRheJkUQaE3X44DPmxBqtFWIl
Txe/5d6L9/UAM2qhpGpopAv0zs+g/nGeW81BZS1YRU1DWvwZ0ZxkcPo9Ozlqdvi1
5+KGjFbwek7GZCpUbmYO8+NSOLaQY+JN1c8qFFah7hOixv6N2/zXcEj/pK+0nwg0
eTB4cqkfAFBQ3KQJ5Hk6sEu4nD7aBRsoMiDwlcHauiZxU863+XKz5DConpDWnuIl
`protect END_PROTECTED
