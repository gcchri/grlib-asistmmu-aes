`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9dBh7mcDs3XgB3fHtwUP6wt5Nr1XEaAaem8pgC4itNBaxv/xDXlaNvKQMmFFMcN1
bFJMl5kNUikRJd1zObxi1Zckj11/v5JI9P19FznPfnVBfjgZox/ntX3IdECJVCsY
rVy/fobz3JMRa5+sDXed4uZ1MO/Gfx0Dy3h1b1ic08dAvCc84hpe9D2h0CgKGxiv
O1BMx93qH7a8D5qgqLeKZCRcWasRYCiLUPEEuNLaKfhllNY9Tx3pMC76oypLXp3y
6PifxTHVEZg++e1Kmb/8a4TBcaY0xWzYNzlKyIRO4xcVYoo1dveddSJyHh9pl0O9
MfjkASb5ttETfHcPDhy5INa4uY46RZPj8wyDH/1u7U+voG9btz0VKa633N59P2ga
SC2W8K+tAc/44qzRA9oDyIqw+rs33NVa5dv+QBNAZkYE98RSv2Sq7g+CfNZ2CHaZ
oCz45uSSSU33SFDMNS7GStrl41qq9UjZA+yIeCG6v2n6cSiQVTcurMxSpblYFIpZ
L8NCGrsKK4hnD+oDvW7MLYMuUVjEXr12xarAl/bWgZWoyuUrDhzQvJORp09yyWTr
g70R8RhchWYsKk8uXLE2e8lkd9RzxzrEPr8NyLAUMGt9cNJ9x1F2KKj1WQx3DML/
6ApKEOcN8LXE+HdGg3Rn2jMjLY+PCcUmbZN8rG+Duaod0Q/PzkpKYHSlsXHmnmn8
aapaXdX4DEcoWEE5u/b4okWWwpEr2pmamLMBD7UUaSdLCceUyhXpuGE6QAbJ43Ux
B4T0RsUDGjyuWIteQ8449qHzwY3I3QZATLCt3xMWyyjpxncRD0aDS01AQ2AUz5m7
ySjJ8/qilzIp80itTPTWZBD4Ubu/GiY7FHe0XibtmJJgTxB5WBCzt+54J3HsFxQO
I0DdKc0xnXXH9bGJXmvkQr+gLjhTzIHH2nMAAMqIV8DJIFgP1rCwhukkdgyg9EyL
YQPay/PpZO9ufCAImip8ya+54W3BOl8VtWCk7ubqpP9msOOUXW3q9V1uBNAqnwMc
nshkBnUBtTyaIjMTCop4TlWCV5xeW/xJMQ1Sb83kTmmHtwLp9mZkPvN1S7K+5J85
WcuWJG0JEIFkKq4eWybhxA==
`protect END_PROTECTED
