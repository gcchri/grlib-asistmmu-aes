`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aaowIvmXPzbHH80bSANgRqhcq9Eyrob4r2WAYbPI41QSoljqUx46NzYUhmBpk/Cy
M0kp9MWqwxjmhRbDi0IeD2qpH6/bxW81nXE4see97N5pyKPt8tm6ga94baXIGoN8
IPRN2+8RivbZMyoFCTKWABd0VSSVh70NsE1D3lwdACSQsCUMKPkUamVsXEAGoUXE
yxa9Ek6rBfLuqEaZ+pkqsLC0SGqHOe+1EwpNYVvq032LXf3a0lNENV02qvFf4uX7
95drXNM5QsgODuWYe1RTAPLvoNrFy6jH8wjpotU1QppJb6jbj/df9FMCxOsGQb1h
siwQWAemXq5Q+OYeF98lkhsL0MHvc/PiMuL81hfVhTDCFulAM1ofHW+8x2JjpUAk
pyACZb8dNrC4RfyXPbgrZYVKhft6Ol34UAbFkR+O2XXhSZCyM87oybkUI0fatatz
txnKU9AU6ibN7n5UaTtXOW6MoZArTvjVLbuZNZIl20YO70UquGFtL/NzCbFHXac/
5UYxwf4uXADo9T3Tux4VKdt22cQzioCDVHX7zRtdD3Yt/giCbx0LgQyGZ8Wfd8im
0sYNOVIU+P13nT+sBgI9ygnRZYsJRAwbB/AYbPAXb+ns3ufXFqyoVcnpma3Z8aSE
OkQ2w9EKCwUMNQ+xxctN7AwerhRkHwUvwQ+TTjvz3RJWLlNdeJ5iC3yYsx6OtI/x
pnL+/5fS0OlW9UPvakmcoNAHaaugyUZZd2ZAOvm6kFMW1W0TtIQfTyGB8TAohf3o
uv4nrI8Bgn5mKcnHjwJMw7y8zY8Ddruiu1EumTn/1kjxUZ7gI3EHAAC8kD0TPX/M
XuIyLOQZT3UShjmRGo8tD02IVJce4pwXuIFGSvRAL/F1hVBSpwNdpe0zzvPTavs1
/9HkeIzOyooalN62AucTyz3QkrBU+9IHGjSYi800SXKUou6CTCVNYd/7TPuEfdjh
`protect END_PROTECTED
