`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rWAIEFI3GOv1iUkIEEGdfYQSHc2T8Siq6ks3MzfjnkRDulgHVtFGDTAN9NHUfd9V
nDfifV3BL25YB6X/dpjwEjlEm0EWt23ilHu0TbaQXfDhWHXKZvdSP226pUbw+dF6
rR7H3D5Yogn8EBC+vZIrvHoKuov1BJIkM8kNvjeygK64BmKPKGZ8xiyztnuNlr0t
3zBQcjGYoEl90zeroYgY6x9j0RUui/8hfavnv1d1bN4PYxwNm7L+FIdDMn1DuPoJ
wr5ajRyW5DYQjWhhnrPC8U7AI0OTk1Qpxt29189UXjTbco/wLw/tZF3OKvUifR31
7WcLU3FSqT5maT4nTSOvwWu2CRo0DCRBCAkd/1HyrOF9yARmNEX5k6COa+PxNeBt
2gw8jfOX+29TW9HVY7sPsbzYOoChg62x8++L2gAkcu4k+v/pcDfOlofW72ot0sHm
91Qd/fvRfc+fKKSNHyxQ3g==
`protect END_PROTECTED
