`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CSS4vKRoGPRzQuG+unTXXd9IGhYY1t60PID8a2QnZq3Lu4Hfrlqu0p5nLQJpLvcV
HLOT1JcErYmtDfeev7mQfDITHXQG7Ix7lnnHHnG24WPPOqGtvHk5I5gYNmm/j7wQ
npM9wMV2iDWsVO1jiwKTnoCBAPYiOBY1hujyJ2VnSr2aOUXAvWhyK9UVyQcpBV6j
t1N1QIXpwk514Ly51VbWGpKLbEMRrZ9MqNDhIW/tiNXht32g5owHx5lowfCUWQ1Y
o+YGmYVYTOhHIJuDZubJ9yeM/mgwu6wPbK5HprVw4DjAAg4yjK13WUSr4mHvPZ1t
y+AtkncnGT/ntdj9awTxQx9KGVXQmdtz+0O132faLvCDy8tCPN0cc1OTdn0BbKLA
HKeGjKG1yO2BGggRFFrsHAk3r/sVU5qiwpJtu2sx/Cxw6BHF+K5oDLXrWE3aPiR5
MiuB8ew6Lm75J/h44lEqg/MD2NmjYloJZCFDFWFFJ3HIlqT3Pxj8Z/0ehW+wBvTG
rl+b6hq95I1MrXqi+DcJZiKJuDx/yhmB0e6LtZElsW+djp9Dr5ZztzEjZOlASH+t
iis4ruK7DRm4Mr+9Xu2IeccOW7aG3cWCqnDMCdUhhqjI8qzRo4tKYl9UCa+7VzfI
/zRkePkh2GRTZOR7O0lDXFX2De7/hnbh8q5Va4R86JVLFXUIy/C3OHc7wPGJcVPB
8P9HAwIF1Bqq7XnpRlAQQxKCXjjTXYwo2HuKvZWoDf43ZkK8zv4BJm+UQ2hG6yNl
YgNjOl2PVYhyugVU6ZJkBz3WiWQ9AuoFOSSArGs3UPq2ztu8y367H95GHdQn3oXp
7yR5kTCfTTcSEvIomS+nF7nQ4bVLY/vVC24xI/LitAbEgugHY1FATB/6yC8kPvr0
4330tIMKZmBd9g1uo4U3NuUHH+ckRi23pad1FqfVQpfKAvHs/xfpWHOFD6W8C9wv
qCIFE9/f4i+A0k4BTOS2AKLVX4hRN5JtOTvevo2Xf8B2CPyvkqdukYb1UlcNBQ1p
PJ0KhB6Ct9FKMVSrPjsQXGT/TPzPb2ICRlGvk+ty9n8sRAimP3tiDkBBF1odmjNc
pjqn0+HDEsoRgQPqB6VMKwvcSgzIq8r8OoB7eXBkEtbPlY/WxilOv4ueQ2AOhBo8
h01tfSdJ1eRD56ejS1K8b/X5Dq6RT2tru1RYuErbYBgY1+ZS8L5Nk5AB4hBV+/hl
S9uZbHnagocYct0MBsNoePd8mXHvCyj5AV81kx9FFAukozHhFYTpX4iqeEuevWDu
pnLhWUpnVVSjYx1+0MvwfKaX9AeKri6AYfYcsveRzdiu8IvC5nYwbDhJ2lKUk5GH
nbc2xHrrNRibZ7boSWqiCg8n8pwJMs7zfV9fX9s0ODDsoJ0DK+a37fhHQ4DuiMW8
MhWaGIirCM35KGYeGbk8wxNiKB3YEz4KBXnnGNswKx3eeWyt98mwPxceZK3/pdSu
pVkMVvKvuFuRJkFLuGW35NFA8TFk6a8VhzcbJQRbldPWIzqHiXDWznrFeNMEkr5U
Vej+TpWQJLc77ZPD+TvxY5/3jQazQmKb8r7Ab/6oL4M/y4CIaOiVfnoLpYwuFacl
OUL6jEHCtTnj/B2DIi9587E/7YjuWkP7NhmIsgvgg0qf/9cuAK98skIUea5RPDyr
mnh/RoncysJNQcP+sZ8zMEUpagWoZz2saOZgikG9VkUSl+imA6z4JWjkViPrE0L9
fLEQbDoJBt9UpNEZUQ6izbQKyJYU5a+Hi3mCsqQwoTSMFAqxz3SQXYvxWr8pBQ+P
3CkAnDD6xDXpr0Ubk7OATdawXzP1JXr0WU/Pbhxju69vWQ/RWy6tUZ3dcO7P/5wf
S3oEGlclI3uXqVXPSeQNOGqIUXJ0oRSJQxrEtRL8kJ5kTHZBGX+0mIVXvyhJBF4a
5dZiFVuHtmafa4+FlgeimD+shO4gvB+K+QPECCe8aWINJHg/wIezwLrv31Ape2ES
rApyo804pXwyIvv6/k9wMj5OB1e8Z+BWSXT6MP6gsNIKDGueTJjyoBAOMap4ngiY
XDFFb4riP8liPlYiCGvpC5EyuIUlWVuIjuwwoAdho6aUolVHGpA2WqM7O1FSKKjE
GjDRmfQU5EZIwl2wbELHhN/piXdX+tMsl0Vxujuo8fZeyTwmc1xkW4sfIbiTcUwZ
hLqcKXZ1qd69NYqzQt62nLkxu//1DzeJ4Y/0b+Lf98DVaOIBpRrqPePlG/6OxrGA
M/OUi7iqoeBtv5u4kbMEsG+iQCxkXGZEDRmVbZKZaFaW7VC7GFsnaHBa2oyj6O1t
9dPcOzAKXfeeCaELL0wiM2e13uz9YX6Gsi3NNEUlPAxeRIekNfq6WbbETFHHVMua
pe2bLA5S1kBtTy4FuDn4OczaC/YpyRHmiB2TARktpQvW9aUd5COXzOBEweScm2nY
oa6WAWBeeBqhSUqr0epeqribggudmx64E2bR49zUJsYubo5MZVzUKNOQyfXSucm8
jpvjdwYnz5vJyyafMWmm4n780bCTMh4Daiy+jlds2MhvaA3X9kARnmpzH5u9UCHN
trxeSmquePBpABBV9scsZ+ucQHUT2EDXKZ+M8gPSeHa48MvraJ/OU9tbs8wdPlmg
oAWfbmJ9WK2Lh/AN38oF6zBCX/8puNRfdGIIX/2fN8ZTy+oPFpvtwsTt4huv1bRw
qS8XGLrTYpp7VLXdAl+MHfwt0GYT6WvxFwgO/OMEEcPkfeQnTXYSwQO/XjmckVNp
DXYh8EHD7Wk3TaXCRG52f90kHi0q44Y9Q2JCkQWnxzgILeWZy1wgZxpI4v1h+rjt
UbH99Sz3OWrhd7xwf5eoe51TYp/9gWyX1EiLnXE9a3xK7Rz/qfZk2Qn0RH2tkMgO
abVkqKJ4sOYpyNiiWCeDRH1WIupcueCXT1wohwSHWfuZ+WkfAUkqYT9gxQ1iHHbj
`protect END_PROTECTED
