`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jkmMLrqk73FA0O4+m6TNK2F0TWSLYjwXW2qt3mdcGKY/vyjzIVF+ZYIXj6olwKIi
DczCMQHxCgk8ZL2NqnMmUyIQ1D7nCXKGjRQO1jdVDXj+DAxZ7sN28NYUDWSgqxOp
wNZBtnbrh6ZGV9HvOY1TSO8CPx6LNL26H9dD5+ObmgkDrPAJc66CXzKzHA7mEfT+
swdHmKwqKbP/y4ik75aeawyRWz4yYYOhvbKejsWQKbm49SQ38RYSdFqA7dHAXlgc
gGIN07z9MIESV9uEZ9zLy4ecGMIU7c9wg09lrEgX3G2wiapJVS55XCWlkrHRvb66
be6o3BFGezLZEgIH47faN1EUgfdzbg5lDk6GHXieeagCYETEcdXjNwZN8HzwWuZH
CDU9/ZUWPQTlDMY2iU9nhjuLT5kx8igbjFxSzd3b/mX42bTcBDb5gQ/qEBw1Y4z5
`protect END_PROTECTED
