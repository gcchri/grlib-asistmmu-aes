`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aPmHXTxKgQ/qr69IAJF5W/c50rmM4nw8YJ8D5a2Orc+tQ1ErITgplKF5BTZrwyoT
7sihqxtojboFUeD8xTYtQ8rgqJxFwr3hTlC3YtmhEyXRo8b/aS9hrJGbsGif9Fdg
V4V3g8Ublm3robfZjZmxZ7bAjFrHiF+ekFkEKs5KxaoavDcXGCVnY8QCugY0tFtV
aw3VBiTrkEkJUEsEjulGt3xV839CTauK/LPeb83QXsUJqWkANVr9akR6MoxVBi+/
5X0a1Yw5sWL6t2GaktpedTmf0pdDQrTV8tyFNy9ybSi32fLQQ3FeGabnS2AOXEis
XnjNsBiyxAaxf+i+h0C8pB+N3BNECwRqxro0bIO63LKl6HEt8C/1oAI9lOIx6Yj7
n5SHqgM0ogywvHo+y6/cM7HqbBAERxGp2iRXkE6QoY1vVQiqiByYLespy5mEDYtr
HtfNVl937vGKRyNln4uCoBWT1AkJW8tU7DWlEFEFA4m5wUvWKqt/JrYKVB5kZoW2
t+2/9ihpwbdya0xUOeMDs2buiRpxwfv0Ed6ZbcrB7mg7KYarhO2Vvl9O+6wfEU+q
8EWcp3rP8DJxIzubdx4/NPE2jqY6OT3G9TgSGkgugVK3aS12jV4S8AN5KnmdlhUN
7lsklrdKQRDdIoR8ID4ZeOEMtECphPFzOfAFyFxysCVnEiT/cfQpQyBS/EfFpfIV
qCE8NrdhJ3wJR8jOpvcnwQ2SCZ/2g0KdtMYy6e67wQXyEyfv3ff1QQFgO4jVdy2G
EIUAnXSK/REAJdYK1i4j1FlOAeb+49m/u9mimppU4by1v+9EIwWCLfzGLkMfkUB+
z+xIM+hLvXMmPaSUV/YZMQOnzJzVqHj0LYAX8CycammdQSrLxxRLOLDJu0yYSO65
hcqXtScZNCxrctvpykSXTVlpYKIsbzjdnWCMn/x5KxIO4f2zn4SVlKGe6fgrtF08
mFgcw1J5uUWSMtoGZ3ktKYQX4TBj0aiNy4QffRKD5P4I3dpGK1PyuSdST+hqPR49
pyY8qPJAQrG831qOf2TDuuXpXZY1V8dpEXGYiZDquQZ3BezASKETU0cHDRN34ZBj
wlVu5XOHzNyIl5Y1a98M8QGD9sWjWfZVtXL3Iv8NU3YV8U+yVY7WxRGLbEpOd3Fx
6JKXh7TNQhDbO1jaaxKkoWaVBtOI+n9QKvlBOEXUGhNyalPB3WjxxPgrAUg2p9ji
C+jCqoT8+r8ju7ZLFo4FFFZCcvj88tKQuKS80FAfhtccxPqnkg2vp9DgvDAKfUWG
OKduypqkSH7akNc3HSshLHlgumsoHbcWDKe2oLw6ECgeIy5TooSpSBXF781opZ46
b15BadWwE0E/ZpyiTrb5ptK2e4W7B+Mo4U7OGgkQlP6sU/b8LC0YmNXJdZlo0PcK
51mI89otlftZrUdLF2MjDw==
`protect END_PROTECTED
