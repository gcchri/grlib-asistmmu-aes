`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gE8LprAeGjwZcD9DkSDu81QmlNekWkWFvVVUQLPPjnPiTW9I8WWqkcWbrEhbtQeM
tJC6XuE/zI83Z1jtsRC+A4T4QKcimQMnTWIB+5Xrj7vm3Dt+pMtKbOxkLPpUNU8g
s6jQCp/vSktXIwzFKbWjuK8MF/406gC/qG2efbIOdDEXH1x7SVlKOq+XU+i+iQYH
dgcPVRk6IDm9ZbhmoVTt23Jxg/xOS7DvnjcR+k1JZTmGgG9pagPOHVNTmdTysPmn
9CKoVNKr07+Pph2x0fYj2S1KmgYIXiE7x+xDHNIxbkjkmaq1wal3G7g1QjDEoQ/3
23JCMWGUhi0RI1R8wXvxVikU+/qacqoFpGTT2irMfPGipvrJLkgWNFa1xP0rePLK
84YGXxiZZnAVK2jl0SrxwNH+h3Avz0NA/6i+ginAzKE=
`protect END_PROTECTED
