`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6NjwLaDAdUWFwjXXUEqc6/K/9BMGl7DLt73qlQgpuo7iTTyxOZIkpTZoHcTlu7PX
5BXncbDZruLPG5G4L8vW6aFkMwJqE0/sGfiyEjtZpyVbeAU7r6q/UxsAYLSWde6u
SVoy8ZNfavaFumKhPrhv2Eh04PSZChL4yH02MjTRd4AtOg39dgC+S546WlM+y4s2
g5uVxayLBbFghZbMmYeWd1nUvCXM+oOmjhvlOLq5/5EaCKp/uDzWmScz+YfwFCKx
BUiv2cT2CnrdtSVCCHSjzQ==
`protect END_PROTECTED
