`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ErPM9z0h/jvGUn6PgDDL5fAH3gNvMyAGzcAELFaPkUtnGs9/4GeEDpZehJIGabsY
lrK7GmaZ2TRegCCXhvIvR+eqwiQ2rfiB/ItSl+wlQZbIdMA4hK8T/bvRGOku7VcT
Pfa6Q2EShNG2pE9WwX243Kk4stqt6RVNOa1FEqc7qHttE3Ja5ZD90TO7LP5y+jN0
I2hJH+JMRv1Ehbxjq/vPc19xcsnj0FfqXM2MiQ8oXEAXWHt8LtoTB/iOgwSn7yfQ
A9fV6qddYLu+C8QMgWYn46n/lHzBIZnDVkj/URcGQyJS6MBsjxqYk0AN7f6gW9B4
fnkvYIA4DL7XDwTppXKh8PI4dk4tUcUy3LTxgGI4CMq6pktWQhOujlZF4jYNY35C
R999boe5wvHyqBf/pqwYWTJa6svovgHWxfDm4RPpnGonmK+tNxUCh6TVmGS5L7XX
lGDLQKDBiiuFxy9PItSqviY2FwHdcNUZFDtQEC2pexJ7C9CdsaNGEXfThSUaF8Xd
r3gnXTsyGxplqJ2MaByuoas5ErJEmuei3A4rLQpejrYNDJwpwbggleHaw3jxhVZn
IvMk5Xo6BEOg5DHsr6BppxUstU6UYvMN8+SWTJ3jT0H2OEj9grCQ4eAnT6ehHtxv
SQBSJqtOGICoYDsQ640KeI3CmDUJP66kZnXEA3//M7aChItY3E/9R9w6bqgqJnsH
4VogIIxy86C9/iF6olmxXFmQW2JH4pbgHvmCeXJ4PZ9KLIM9hW6tOYLx9erSCDh1
u6ZLtu4LU9uBIp0q5yDwC9sIxfUf8NAy/EUqQbhBdsO8InTl8Wz4rfWQxChAOEIS
Z1sfZ+WUBJDLaWIpS4YhJdzYpWMLdKUt7cwG5BQWJX2BCS+4L+gi6VV0oOZtfhYR
HS7gJHSChEIYcO3QPrQjcMdDfgTs2TTNDo4PR5YahAgrAEtZErS87JxxEnif+RDs
W3fXGkxJd9gYd7ih4wmaPupVAO2bUIIOwDwqI4PzZSYXbElJ14YhjpvkyTZxMGdC
GbjT4MI9tH03vaGEdJMAwVGf0RvqdcGKrif3MxaPCRFZnkoGplRmc2tpTs8Wpz2t
PYqHW7PXIEUUIkTyugSwWu6BRFszvkxHVlZxStNw3RqHwzf9IU+luZCCV8QGg5bP
0FtRXSUEb8uTWcC0IWABnTlMc+IJi3CkiFMpiHVoZRdPLya0YW1bmRrhF/B4F/sx
oF3Qvop2vQ+W5arGep0D9FU5fhFV4KGEUbVjBC8AZ99oa2XlbUV39PAtbo8q47GX
IY0Cq4oBYh5yHEjIcf4YCSL6c1k+7lHPJlVKt2LmstDu2RqvroJjp0+zolAB0TcF
5+kqBzswyQdxTITtaVz2OdHeyg/3a+8kJ/VIodTfeu1MWmDM7X4Nm/OkUqABHMWj
3Naz6Z3z6qFfzddOOEngiT79o/2ufLeJTKoyIKt+2qqhHVro3pL9ilSuIRrJVhSE
Qp4twuSt4TGV8ae19GPHzp81yGGlbbhAQaf8vECWG5agUAjEi85zQn5A1oHk9fjY
I+97ocQUG3/KO5wAO43cQA69zw6l2LXo+7K7/bWE2sFzqaUtZcM+3AP+gfAjdlrT
ijIZPv4+bUG0QPyGgvYD1GfOwVjs1wb5Fd9yLFOWiSOM5pPiXSHNv9+uF4Qow2Xa
qH2XuABDd9qbotbaXPR8wJRBzEhZKmIEHZGLmuhwQ8CdWKiKl5o3jOTdfbvrzOHm
JhQjLGrQqbTSQg+uG1RX+yQMo+8H374AYJ5WVtCdkoIdC7I5cvGa1NDDILOF3Zpz
P6q5LvpvHeGdxrG3h7CA6HpmcWweM9zy5Qk/9kupSVX33XV1BFN7RXmUowyEpffo
76gr2+D+WCoTwtVFaP4IoRi9JQJcje3qWzdEKDb7VdwIam2Ch3bTTJYE3Zx2K5u2
fxHhLa0etIwXd+KMInOXpf2TA7LZlPDH3240jPfoq3d1UPO7tSfmWKRUhP3xSvyH
WriLF/1zWYerbHqTdT5oe2D+ZH488y81law5ZJexHgxkistTg88Jv4FWkpUzXiVn
3psFBbn4/SL5R45lTrRb6ALHEDy1ezrToYfJEVX6K2ObRZ6klFuQfrDH4Ro0CPV8
Nvm2S+D35uV/W0hZ8esfATz8acjinjvaU8y+0yImz5s74TTot95gTMk5KwS6cqRd
R3mQcUqyCM4fhevTNqJT91HMjWwBiUCwUrrlT0TaWv5/LMSOjJAw17GQP2mfmoT/
wzlt/A8dego/Jdt02ggqnQFzyiif9BKvAkUKQ6iDtUikuDlguC2vkCGcYJGelc4M
GB1Ox4xK3O4Mv83wBAQClFdumWVF4OzagGCaIPohiWEBLwV5LIA/2w5dFJD+zSEx
VkAwJeY5LHq8VU6Xu/tjIW+KL/hHQRBzUh5Cnl0i3Mf+lQdKD6Za7FrCcStF9iLv
L3E3BTATN/Gw94kmbjPUK3h1StTAAciU1fiFwa8ynLiSmFdBphq1JsFIwfy4O48D
0aYfIRQ8fq0O7Vl8cGgMjKUGZ5EvCZ5waOZiB3pXKv8g33so9oBpFdnuz4BkCvhP
3Gop7CT+Vw11jG+1F6Ja5eHoq9wYHdt7GRETiF6yPlJvhV/z4KvosF7YM8XIM8JW
wqEi4aDm7gIdf6xey5TbaZIpumD1+KUhz/u6G287tLSnPQ3L3R+coB8Ce7njAhso
yt72BFH+adq2C5RNrXXpIumYBM9N9aNHI1F4mhMeC0O70H8zCjskfEy89YdMmUvd
JW4pz/nN2nJQr7A9VPE6RURa6wLUxD496ctQ3XenFFB+/qldGPQEmvM0MpLHAKOS
EB3HJMz8Ruj5b7UcPyXMdXN1GGstGeQnqwh8gJ98AF7rBCX9Y0YbXFCANbwjpVnk
4n5CoAwMjKO3VJgLufC/M1WRQW3XORnQVX1a1l4eoxnDSlZFqSM5Tx08BR3qQ/o4
DWLFgJQqFw2iaRWWGwrSlhAUKBQdTRnKw801+6wQJ66O4Q8+6XaFcKzceqWXD4PK
EeH4TWsNUc0z4O0ZGZNeByaEsR3eiJWyDtpgEAk6utshIAUEbDnv7jb0LlxGma+d
IyAyvn+FfuR+dnfPDO8LKIOvW7zh7ttxLcVA071c70o=
`protect END_PROTECTED
