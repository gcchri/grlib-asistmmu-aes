`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MiP/fopxaPnRry8os7miS0cKcer+sIcwXsJwPGLAPT9tY56cqO7aHyaRM1LEHjDP
pOWvrxa4aS7GjNbC2RtkuYkhOMf9s7zQs/GEDH/luXRrNqMge6q96ikZ9esgTMyW
jBEQEsVALebtSCzrN2aHXDrkWyVn0Lll5Eaov5uI7l0Ay5Qzq2BPptdY77vGTY19
eXN26RQVXA1sXVZh2hrKpVBi2FrsDNFFpjJQ0SMGXbTb+Fe4tY60kSvQETqkxsa3
elGnAoy6wgf4n4QQYo1S3+pQe33CvxLdzIDwz+mGeFJaKEO25OyiPKLVhuNZow/Y
E0WIRmaFAi9LVXrYkaJtFBUovTgA0pgjFIgUNJE9y8fWu952J76BgzWH36tcGMXZ
YTDDY+ysMv09Y1M3WvgEScNXyST+oXsSipfa/w+U7xAN18rvBtbhiQQV3BIMQ49O
cwz6XNjfnqvHG5T0KU4L3WCnKqMURY9QFHu1NK5YwnnoWC0AeKT2tAM3Aet8cx26
`protect END_PROTECTED
