`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hdw2GIZ+Lrd+F9qHjn7g6ly/4T6kij7chQmd+Cl8VDeOQ8Sb9VFTOSrJtBBTkz66
w4pkF9r/cnRkTLVw176z5NRdQze1fkvKvFZUMyiZwt+CfYNN2e+hse38EUj1jkxK
hdvCrmSA5LiCgaeGR02lwvIq46WDPiGNtjx4XW6dL5t2dUrsU1YDydb3Bnm/mBrG
rh3E8BqWJhcJyFsGZ4+ocQ5P/hbql3ugzEDwE0oWSg3vRSOD9PO5WuHSXM4x2L9Y
QulwFnplcSEeOrGlPPveB2cecg/49h+eDHiy+KbuB9uWag85BECNzNgBbxiktudj
K1fN8hh3bJLY9ntrbPW7rVk19fdQJF951XtuPnoetJjfSdBC8YIZgdLKERbJNggc
Mv58bDuepv21DO8hDUpZyZgRTrE00pp14Aoh8V8CTpXs8yJUxf5ZTPrASaEZQTGO
/C5Kbt/iokNuAAYQwmOC868ifca3I9t9zCndR/s6hJbD/7HqLfaZ96vAAd+6l5Hn
uNlcbk2AEOcrdmO2vTcwyQ==
`protect END_PROTECTED
