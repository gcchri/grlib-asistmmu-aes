`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d5N9VXeVG07KbCSkyVj/zQ4R/ClNWvqsiY9Dq1UbVuaunNM9ADubeCoEeG1cEk8X
1uEiDWUviOFuuRz3jLU3RKQTWzSmOHCYZIlzxvgflDw87uqhlCQ3Q1u6w5PS2Ctr
XIckbOhOekga8eVvExmWiw661sbNLRv56ghgnbsM8EhoPAEDQ35Ol4E0HWWhQPsj
bM7tJk0kDBBCsJomyVwhFkXhOVNaVa0DRXQvbcqePeCZ1fPepbAs4BY7YT4wG0J6
RzIkqFcL2JM3xDbORnFtZ3Ct37MMzFdb8UkfTrztAtEyoit4tuJkqd/YHt8WkKJD
A/Q1CRQa/EjOll7qxoAtdr+SQNpu3WLwawpwcr7u0In+ntP5zDqaeKuUqCweviZw
L8NxiNCwTJcyUZWWNxZb1Tka7CtaA1RnY4Rn292Xfd8hQWWbJM4VHPtHgWkSBGv4
jgbsgpkulIOy2FO1BUiw4r9QMAZMyvdzo2wctXcPjd0wOTUnFQdzpf8kGDZEZzyC
eqsj/FJKzlD6AY2zLx7G1YmCfJcsIfmKF0S0Pv8lLguN8fl4RQIAaV2L4H5dnOp5
hTUM7MgUGAqJn6ioZAVgUc1LJ9V1QOtgd7aC5Hz0/idRQts+G6k2hJQ8IJPWW5XI
HeXXmKi82jOeKEVp/PI5XHqwKJCm8BA8WhtJCQOTlLq+YIm0/jwiNeV9PNJ3PPJo
hMtiZk/mqS4umoNSoo5awyyJx9R9vHibmBLscyRQDWH3h0HRvJOf6tngyoOQPgWP
lreGxloTYeUCXjokLVC0U/T+0us8SYJblZ70VXP80PvJXOEKzevbHgvWlV4JfV4h
81BQ2cnYc162n+M9k78RMlr2mKG5S1jMQ5zjHPe3SiA=
`protect END_PROTECTED
