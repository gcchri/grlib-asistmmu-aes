`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EiGK5ll7WuNz6ds2xIl+x0OTnzaJqqFJ1DdRiXnwMwEC1es7c00igxJKaw1X3CxJ
S4sU91bN9zXIiwX+buL5jH+pBq/ae3hZwrj0/3mCsbUWHfSmJrnRQJGNUXw6/mLZ
7fM9UM/L21OrSn2kkxW/kOQQWCV8IWIS71Zej6o+oXxlrobXRUNL5PjI20r222W8
WeVt8lJeOCUyVEhV7fUL98QCxHf+0zQ/eHkjXkctPCOoYffa4kiGu4nj8C8yZN3D
9HmmCfsSFqFTo+i2pfpzli7GudTG2ue/ZsYV/KDVy1Q=
`protect END_PROTECTED
