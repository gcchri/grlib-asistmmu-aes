`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DjVPwDHv4WoHBN1VPfKTUa77bRpfw3BCQ3JGwqUEqYH+PVrGg/GU17br9UajkEdg
QFDb/rXWRLs/IIK6hn9wuCHehyJEDdqQj6LHCjSN7OSakbJ/+YldkyGKiNH6CQf9
KVwI4Rmcu/KbCuGqkJgmAaaUaWXtxAGdWu2/WTKOMDwbzyPQoaqAe5BPrTM7nepo
5/tYFtv93bLrq4U3pFDghavDNF4SAaaIDlHgJxXzJWLuZOncFnjrnbg8A4NTMOed
OFOuVa0Ea+IMGIwNoN/F7wycJlhSsEtJ07xbqY7ruXRlORWLS4i8EaH13P1cYN7e
RzRwRiMHxc7r/T1GYTxD1927VwvWobT3J0smCcjWRGcr8SkWwfMSfprqfo7KyWbT
3SVdMp9oFjEbLRzm6lplNnox7RDUSgfN+C6WzlkK9bJDa5A3S/OEbZoKjnKfTVOP
g99LpTEwP6jO5MYBIES7+ezVcfqUO4tuv4JFfFEiOIryb+Rk2K1eET+v4x/Weqze
Rcp05yNISbNNdCdu5Xzr2qpRlavvlOSG1jrLOrbVycMbFQY6MeY6YV5jWq5Yp/Dk
//yCNJi+soH2wW3YcL5r02u42SPJ/F4RE0FBWE1CC0WR7VnO7Yd+pWCNCtkfAU+4
wzCpFFYOZgqhVjmoj9oMxLLwK1UfQu3A2U9+DQVbbQ4rJd8tgvVXuOKFRCG1Rhac
vekg4xwzfRmct1XJ7O8zvdupOcVfSSLcRz5ggbcF5uzAQoF3GfluTaDHUBjLMjUX
y3VBZwvANEI8jq7XjzeW3LoPn6mbvgV2sXtuNLG8SMyx/PPdyNWmiS+UlZh3Hvo5
2xR3g0I//sIFGsWzqkdU5cueJ2n14EQStMSpd+yYiuTBVqU1Gb2kjZkdA9+OM/9Y
ZnpJWoPNd3RxWGpI33tzSORhgWqyUU0uap5E/1nJisDFz37G7q7vyEotttQ+kMOV
O06uluLg7AxJeQNzYLaV+Mivh4mtMn4RWOtSKY8FJ69d7wVQnjJOkbjjwRnJlls1
zWDdShigIraibe1vJ0FtRDM7ZbQBANyFoKDt04ufJQGosOtjvw8thO2oUP0gFecS
KTv/yh7Smb6oKmD9UrQ8ILp8NkmjIaq4137ax4sKEqy2GxI/kUPdGfYNvVf2JMQp
ymrUV1R1qakg0ofF0ACT7rspYSPy1lUBkIVWhGHaqWpkDdOGknq4fzKoWN6Oh+v7
qQsCgQ7jvTMUL6yj4RioWr/2MtCNmHfd62YrA8UP3oOelpChUMCadRCfoyn1LCwE
0cWDqW7GVuAQN15XyslDUZYlop7lWFliTTB3dwJpBS4ESDt+jX4VCGaRU4lP5GOQ
7Dc7nDWARcqMMjXiYq268+PXan9V8VvGQi9BvYMVX8LNYQWB0C1ZijXbNgthLK88
yXdOopA4J7zFFRPMaMErPwUmc4ymVQf6UpRtX4DLA9BROV1eQW7j/QhS46ZBWpHz
4+mCyspuEEpKQl7GBdT5am+Z9LHLfF5Vy2yiDuLGJwQDMCc0JG9vAbKHtPXKjNoP
NWikTQ9J8QBAqaVl7JDraBtuMfn8UItD/2kyzkQxwjsD/MkEdPdUSkfh+63oyxEY
1sy5HvV+I8Tdt/ooxIpRMj1WhQXk/yqzLeXytmQS2lBNMkSZBjxLyY0nUDLnk30k
mkeG4EFI36JtlcERHwmwjGJCQJ+lQMoed9EwEc6AsYc=
`protect END_PROTECTED
