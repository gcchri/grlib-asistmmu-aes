`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1tdL9YyPwJrj3138cf1C9b/zZmZevKGUsmVJ62p3WtdV80CdjZxdihhxKKbPic5Y
OaykBILpk+XNZIcD0UsG6TZ5BRY/TmltcqUaR+eL74GGgz9uCIPGqzWm0rbu8W85
zBmKM0rcjhNatRgIsfMQ/KnLfjIXfPpAf8QZxoiNXsDiGFQrxMVm6WP67mxly1Ms
FqmrEV+XNS9vBa33ka4xYnT59QNZFgCbSf5f7238aj3DvrhjGJzqxzgC0nZ0eCrE
oL0fJczpELLprIOCT3hloqSQnMsZbob/SjvodgwkMB0ipMAu6Q09Ct8b7XYnvD86
btAQ7woQcpm3bv8obN4sV/VkFEv+zmqkk9JB3xUtOEyCuTeSlEttArcGIeRc+f50
gqGedssRHGGOkBS4NW2Hy6XXs4+fkESzlrWlvyWCHB0cKVZHnwRELxVH7tMNnm1P
VtClvy7eqik37yDALTxBorEA3dlOgwe2VJSxNppma/W1R/KzFrG1Yo3YsF3ojK8a
`protect END_PROTECTED
