`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G3ro9rofFaXkw3UY4EuAhqk++aQxkNbKiQpzX0XV5KDMWxnzXvP2ComohZxLHc9d
BZ4tjwHaFpA/c8jLG+gMpNw0094OOd/BlVXzUhTGx8/OxddW4Pvg+sAV1itjgdL7
89KDrHB9Ixtvr4YljylZxg9xbjaHMapGYJyqRKJy4rFamt2we0L6znb1xUVyToLg
vQv6Y6vxrsNOy3HUFBfShV7MRrEaMaTqCoF4cMrF8sf4nUOLtW+pTlTrmvrI8LWA
FgUo87sOuK4Z0mT2lisKX4nxUgoOc2btqxZTZ2uHtYtLnmzLINEPaRLc9oaO8AZP
aKkh3ERXW8OpyY6SpX9zdAsRSIycww3ovbNGSlXXUaD7z46xgdIMZb2Q7YmRGmlN
L8Pio1MjYs4lqQm9x2qTadKmx0pWbmIz5GTlPJBpJEYDVqeLYMod+W7nqoNNLT+2
`protect END_PROTECTED
