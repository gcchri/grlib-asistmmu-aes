`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oy6fiPEkkBH4DINdq16KIP+/KatNk4gNGaRbEwTRCg8EAvhOgGw2bDwT0FrnAw4K
d7X2b4fUbHjD/7yaW0BA2ubEH6gts3PNtR6iao3p+Uiym10HNkm4p/9e42JdAYXC
RB//AodtQBr+gYi6MDNG9pQjEUWd3firrpkJIokbisF9YsPM9Y0iZPSJdnlHdBxC
58OjRtHCsDrO6okdrFgqDaDId5LtTF70tBLgaNrBeA6wKwVW+kp73gn/Brv3VTjN
8d/3wWJa0eXbI6CmTWBa0ONiW3cRWeQeueh1xSR6KFAGp6EAZOanf1qYQ7qAAF0j
G2ZMIJO4MgYx13e/K9NOdn72iU1zZZMa4cNuIXj1ufztMMHV0g+vbVHeCZqvC1Am
g/zqj8iiN5/m5TcWR565vgp+bB2KPqNN5ZwHQdUF3egTCHSTRLHuPHlEz84/EUq8
VFIQuySfOVdYvuh9zvqSKA5D5Pn4+AkL8M8s+FYObucsCqyKDFSJdQTVVWulu2Oo
ORuyGcSApGWpkO/nXcdo2tGLsEYaVbOjA1+ywe7cz9bsEi31XIhxzU2d3Rvlgase
WQNETl+SIZzGDHVDh28AqsfWB/Ev/pzJLJfDaqnSvS6JdPX0Lq0chTPBM0/loof5
z77BmE6slowWIyAjZqeMbmszvn7KItoXJmiBLwIaF5h/yufnJxJFDlQlUlQbHrVK
q6LG9P47L8IqErsBoZvn3BrzYgQ+AH/XCHjLQWlmxwNFq0cisdzAz8TILH4g62M+
V2DAtLh52JBdwi/1pDkzJnZSyEhf0BtK94AIj+wogspOFFDi0Iy4vyOhdKxbQah+
Gx1M/Qhe0d0wMSPxnPecTHzsKLEoJAB6lL4FP6LcvP5FpKFOUTsp9yTk1MaDD55u
RPBV6BOq1wr8J2qkYOI5F2cJdeWZqBJT8TTefov6dpeFBpvp4RTi9xbdec5Us9KX
nOT7jkUUbPc6Le96UM1f5wcwy8seAbKg18/nDqP79XdbC/sVBGWX8bwLQL95FiNf
jf239RCO81oNlWaNlkvrIiYnkfHEdoLs1larZvIdQOxCWybikWaHfpRJSZ1LJ1kp
Cje1B3E8CDKGiEZcQ5kIW+F/A9PUBkyPpVXFkkAGnu1ywKOv3Qu6+uKnhJsTLbt7
qnFKziVzJrDGB2BocJS0kRQGP/lXZXP0JY66niqplwmwEzQFSLFEDdOPXbMSCC+y
j7ZTLYmq+034idNeLpBrnq0HvtfizesyQp5qeNibxXRcwAqDd4nLiW5d6o9s3vKS
2f/IF1ZARbnaHf2IauDI7kfG6nscbJJ/qDmeEVQqBPAS1UT41fcvFnEyxtOhgXB+
h2hfnOLLwyaumFProJGJU/0pgvXEBE/hq2rj2JuKo8WDGcfAR9d10sHGscUDetS3
qOLCCQEtuTKvMjsVIiOdrEdVf1uAxLnvSByHK8DqApLMrCox0wpdGZyyMQoZcySH
L2pi445uSPpw+IHLD0PvujH6pkzqG90XBV702K2kVkyBbgC2CO1YaMtMIfbi+ndH
+o7MHItvGyvn0Ql8o32P+GcavxNruGi4/7wYRuHwFyBzI/QHmPLMIf1gg3Chp0tP
fY+aThPRjZ8sR9Ll0seLjsELlv9pcAqvZOA56bsQbtp2FmWVz+ziTiiiGMkp/Cwv
8NhXAetiGxIZHwQwQ2qebwGYFUN5Fv1oJ4L3QX7d6Ub368lrJL9tdXmU4JB+T8iK
qFxP2Owmy9J94gkj3GmIGNLlbj6GoX5vCtGbtvBG1JaGANkOuL6XdQ8D49ehh/4t
K+BSn+HMI9Sr5bD7Iv810wWgsVR+Z0UDy9fRGzTmrkA0oWlIHa3YIaVYgWdKy1MI
5RpkzlPPJH913LA1AKYf+c3GCQmWrj4GLbhdTpKeN9qQwQYi96oBmTzIj3rjKArS
JGaH5q7JjXRH5IWbO32Fb+3BPJFDAu9PjAqOy/dhxkFAC1t26Dqxz2oo4scsW04A
VVXzulsJ0fJQjtXLOf+Os8cCKZvXGPbUjdU+QmezYDvMPryx6YvQa78nqQZYwuaH
VCCN+1A3us37jlnQJdb4BFYPKQbY/187ic3GJi4A355n43lnIIa3cKktsp8RvNTs
VpIPWU7e4s96biPGPBfscycWYbZtQPBCIr7/BDVTVdIwKco2EvBlPChwgoiis4yl
/8uAbmusgr1FmJQyhc42n6O932YpRqOo/aQtBpHx0zHzCg+7PvRzW3T1N6S8NPUH
txIRfsAEQ2wLYH74gimykZ6Ws4GgorZfvJ8fmOFGPwqTEVIUIDQHgdmY0M/b6HZs
N2XUunkFWzy39aFbz/s9eqzdptMjnXJ2bjqdputttPQkpObP6Bsg+9uTiWFvtisj
sMouelnQ0SHRXmeA27DMDcJEoMOUo21RiM6YpipYqC+SCaQPdfyby7D8SDekMRSX
uFNkkxWmdwrM6ONh86VFN/e0cHmUUMKk8Z8jNbFm9fpUIRyJ6UDz46ucTKv86/Zu
vacTWJDGpve2nJENzUau9qC9HMwSajsP3GQRZQYnJeg=
`protect END_PROTECTED
