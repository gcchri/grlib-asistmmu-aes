`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4zGtRl+FsI/1FmImzFUcPWUsVdpELKYpibXAkff2XqObinCLjN41xiQffCLQHCN3
z0RFjC7mLgh9VoQLEV0wcS2jlP7j8ZPa2JwkS/aAc/pl8PiNFApj8fNunHJWz3NU
KtlIZrgT1eYO3Oo9xrNqya8l0UPMOz3grgw6nh7Hz4QWRSyyBuvghRzh4nOuORM2
VGCF0CDodvOZ0TNzLWjIp9mo7hxsiywMQS3TO2zZEGQqvvXmgv5C1JlsfRSunYhM
3aUQ/g2fkP5f6mlgirW1uZ5OmNMQsBV+fMh9mUak38VgSWvTARptr6xZWXqVSVah
IZycnJDg40t9AG/qecq4MaUsuxvZWqjGQXAZRcGyDTZTb0Rb2sdCB3jJDrsITMVt
EM3lb+XeXxFpCt0ChYGHKrrnhjWutHNGYB+/Q09QBCkDuaebcxDSywIrFBuDyHO4
+b7B/JK7BWc1EU4PNH6FTdYwOEnGR+3xcs3BiE3mqRJLemHtI3ziYHrOeafec/C5
K0pYeMLc4Ao1ru/H91eSdquAAabdhW+aTsMcZ7ONlMX/JOr1Ge5JON7/8H5mEEh/
A7h/cvbJvWguzmVY9Uy2RCHqJKojW3eXFge/D8L6Difs3RSRSy9MYeCzEIco6T5o
j7vIUNwf30Dn1nkjicx77WOsmDEoTNnO/SnjcY/PyI3ow0sAM4r8PKA/PiPP4hTx
0rKIBW8ukC4XYE6cJL729RzKN7UxF2sOvLj8+jEnjJnosGvRI4zxGK0z0M+kWljV
DQc3lTkbgMxOAotpjqpZakXNpODGWrPeVyiYqhl5O+WYav58Sv76cFzEmG8JrL8b
HaOsyB7pqGglav4uKLnjacFMNVuH8EGJtwHloUb27uK2iBxXJqdOm68Os+SnLcza
92ib8yd9hzadzqp2qRzxtDMp1k6KOP+6hy7Xt7B1/1aekDgYOM5yzD5DymAdaslq
qCuUI6QGOPFHMDRbwJi7XLu2a3v812wo7AM9PH9aQHwtApyWxEqjSKAZ60C/f6Xw
ikd4XeOh7WMVtWrkrJyBGzobv+dOd1UKicwp2hOE0OzvCP8mon8674DHFPAXeGDY
M+CCjjHLFArLyp1ff819BEpFeXC7FTGHXsFSxUoJX5DM4rK/fwJe8HdDwsFKaY0+
4U5ZVOyP3rbGp+ic/dg8mjUa2dsVPpmquYb8J4Y8txj6OtvX5BmZYuQAZWZmGhRq
HvQqu12FEjzUpB44fU80Ww6ClxkClPU2VtP2qwfMjnmzLNRxLn0jmLFiMu5kZMvi
`protect END_PROTECTED
