`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lt8j0fxfGlyUqiNrbL57Pys8Dp0/8btYbkYHz0CQFFk7nd87snVzdONc4T57ohga
o6aXqWPpRKoGmtrKA/qp2Py02yJTWmHaqohxR2/h+23BAKoZBVv/+pqjuSg02iDi
SdQ5m+HgZAhOCy4ynkPa8emMZFtBH9R31gMGSky4hcMTSzkhNou83+dGR2MxwXBJ
Es0dc1N6Vimk70/1Pjw8g4SxSg0FChkC4qFWJo9DKsElP5J+DTRohpzyeyXe4yR+
6BVXQnd0TRZUkvUlt0mjPRu5xXcsglVWJ3KxWNNoH6etieZ0FkbTa4AK9uUgRbQd
lspIbjC3Fbalf823MWYnw4UvWOJrCRQblE2fCzNiT6wYZL6ws6vzfufmrGi8TJbp
v7akhB5HznOS8nPsWRKo5F0kgu8NkNgFMg/1VqDxeIygKQ1nWZMVoqDJu/b/opZS
l3ad/TfDfScCS6SxClNqwA==
`protect END_PROTECTED
