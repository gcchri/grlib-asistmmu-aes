`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zYMlKcaa3PvbTNfqLDOdWizoYEf7oSQd8vOr7VMogm6/AxpUM1Z0HoRCssWx5Okp
faefi9NCOwOtI/F7ah8ak8ehHW+dRUeSPqeC+uiZ2mzI7vcx1ca+uTJTlmaBaSMS
68RJXFcgJjv/KSKY5CqizLF0gMx/bvf0NuOlh5vxLdBn9aSqMF3M9HNeRVRRU3iy
VTgo2uerTEYVDB08SrZ3d1Vs7YbdiB4e0EA6F8G7S0CjAA1G5+3NCbJMr8m+3/z+
e4DJY7q372WfFnFGE8kY7JwZAWWR2JAVSS0oGuOsI0RUvhWKQIxzXiLOYDFtwwbQ
61sOKP5i9KlMG6BIVy7hw/3Qm66/Tr8sVWXh8z0MredGqzdeIBizayK3Fk/aR2Xd
qEQlfRVyczt/f/O8JuuY8qA21c07G+2tPD3WtB/TwHeFa8CMF3UYqIiS2fZFiXr4
N0LfOqSJwF5MnfMashkiN9W8H02GxbYo++IDpNKKiYRH7sgrCRDI/E+f3rFyxL1z
iVWANySGDGBRuSXsccOZO/LUKgY+9pqle1UEIVsth9YCfxqOqiQ1eaTQVpq6Q2DB
r06gYI/p/dKMWygnK3SW9NlmjXosDFDICM+RDsX8okKl5mVxFlkxqzhXgrwk4DFp
vbnVZvjoA2/kjFOjc6T7ecPhkIk9vg83JfXiTnipuxmK3ryvmZl8w5TQLXiq5tzq
uiXGPAVkcMdHIFhDTgLPaF/q8GUWOEekUi2vaNYCVrdcFH5MU1ALBth1QR/Fkpo3
MTEYtEYopsqwdA+xtzexXm0780bGwEHRerlFdOwAZVxU4KftTb4H8UYUVuFS8B7H
K0jr9ItOYv0r5Zn+xpFOHxeSEnq5EZs6ODNh+C3fp7z4AWKBt4UtjCa/RwTJiadH
75DqCQzUPCOBZiJuMru8yEDCqIiuEdEHffNglyRyM2jpLVYQd3SuU9WDUlFCJQvg
seXc7185J5EhGFa2cCUYfJ8C48/dce1dPUm/XQdI6X0bFxeB4FcbLXWC9einLOS7
B7K/s5BXxZdTJhXqgaYDAPqQSwplsgQHa4xX3p1K0xASZ9Ymvtvcdf0AsBSARq3W
56PRdxoe8sxEQ+kleC+yPXPNUlSq5pQLDx9S/Fw3eLYnbfGo3E7Avju0vlXnqlr9
a5ouLh92LKPAZaq4ouDb9bJJdjFwKC6I2Swer03S4USZRUibhFRclNq1h60rjwQ7
yWiqug0e4IaV2W1UuH2kbFxbZfnAPnXcoRBC3GrqRixqJ+jkHXNJNR+ihr5sfyqD
LqPXZQd3ekfH5fnXElW6kWFcqGb1eGglMSqFT2hyjcMGzhzB1QthseBKLdYtT8Kj
dJfwdHXB8HiOfTF6S0rhHSSvbyKRqonm8zmhs18o3+N3o1u8Y/LQjjYPa54AOzIX
rbhGZ6f4RarPQWPclrmILES4CFD1lKA2iDBZpmE0k84GtSjcg2OVRyvmjDMY4mCn
A2waRi+OeCr3SpvvWIaieRn1AgH6Iuz7jHhRir1iGp3jEQvHisOi87TEP6Fjo8ff
JmICCAaUVGUgeVAZjLyzwlMsI/cTWgBl3PQs8i1yiiRSwR9T5jHjF9scGf/Uc9FQ
a9BrIFkb6dWE2Kr+yiP3MUpDuNZ1fZI5zBg7ov2ejMlO6oneyy96UONWV8iwW7D+
/7Z6cSKLI+Rgd6M+RklEjWGYYdhhX10eNJggIv9EClm/V0XRX8VqKJfmhXg2UJFh
w6gp2ybqL6NpNRzy9hJCDF/QE8rKDrs7CpSL22/vhvFkgsbzCS+qAP/CD6fHmujM
iLhCoXWoNDKNBxQ7lg9UUQ/tdvt1UmZN6lQgbtY0M1nxSXXdbE30zKaj2D0oO7p6
UnDYOqkOYfKCpyQhKmguNZeIGz6BoZHNMdrO43ODXkrhkK3VIGsyWuv6k8VA0aNk
SoE0pdIHhmyLIOQFSP7kch2A5pPxmWAtolrtH7vadfp1fL+WPW5YcM+JIRP/4UQi
7MnEEV+lY98zDEkCrf2q0qEseSmSSpM27E5obOeM98OK6H5y6FC5RCypI5N0GOY4
1/R+rW4Nk/0/U6wo6wJQ+gV/IoJKLlzCN0o1K/gTUJoNcN6yEBEMR0PpKav5L/IS
NCisDXlscSzAAZSBvkOrcBYlq1Cjo6r5IosXZC6D1MPurOK9zLEWZGYnhSoVFxGS
4w+LMtJeribfK5WA37QWC0myaZMo5x+Svre90M6K9iHPHZtMa/uoNd4R++Ix8i3K
gDq10OdccNo3B09eoNylTbk1V71EVGrZcKSw7OCenJzKtHtUdckB3zQOdd8X9f4g
ugPO/42B9WU5VXRtB97jsWM1y0TEwEJ/L4FRjOaniVru10e6/kCucqi19BjDt/lb
QiTU6S1fc9sWwOQWaAY9ZQRRuokqyv2Nat8Sd/+PSnnaMMlM3i6cL62KeOZG+S7g
28SIrI4tIUi0pLhyx3pFUkzSIYY7m3f+w0ylyIHLmFmDnDbuKhOP+0GNwcUY/UD+
jd7QjXKH3LZNG4F9ziNJF4uAJjVp9PJKkW0Llak/0d/pPSzbW+vvCUwGuk0JStvp
sZIrRMnlYo02IyAqZ/ZYdjRyGqH4J5PMXPXewDGeNi5Qn5XPh6YaU7Wu/AKW1+3C
ut4tx0IVihAMp/mThmns3rrLwPlval8RjFiDKmHZjiNMBXw9qaJqgG9eGy3oZBe2
HFwtWTCQyjUrmYbF+jIhmZV96IqFsxcmMWFwtiPwoQdST+F66j0roOjfaSK5tlWA
3If3sLL2j4eUJNerXUz4QUHigs3GGMbzKHUT10XEPUt+9foAlC3LXdLChCq+7eo/
R/5oh6SEtqL801p3fMa9VyOwDs+JaePUeF0VTD+StqsZkV10BM6H2+aj+NObSzIg
ZKP0GEfbjdUrWRjTbn+89ZxBmFBVq3G3hCUJFHMFadm3NWT9j9B7PvgzKJr+ZcKa
s9okrlSC/4HgnghclFCLUTWJRjBo9X387sUJWsUSA0ilIY/BbeZPevVQsZt01y3a
SPfe5eheMjKQPmo4w+MGpIbht2nWmJ/PAzRbNssqa3tVJJoNUIP+CXqcrCnT3Z0k
k28QpRBdH83E4y4q6nkKYV2oMIsQpcPS13ZxGGkJQU0qxJkz3UYtAlyvCVDPeUA2
aNCvOsXK2DpvL8s2DH7rENz/INygUQlL1R1VCPy3PhaTCutVLd+Fh8g/P801t0i/
+d0Ph8qlYfk6sUHqAQtVNF73x4uarTO5ZI9kuO/H2QAmDfQjscowq+PTN31Nfp/v
1ZiDU3IeKkFgkYK9mV70RICPqP2YTY9rM2F+8rFvyhxmIoQqleorRDeG/UtLM9SU
bkNoyazrv0LHm3q+jds+g0I/qLt/01ZosCwJugzCs/k8K5PIG/WcFZTsjZ3dj33g
OSb9cmcWUbHtY25E8wYZfY+kIznARO4vC4s5FyCgSLGQHiZyhsm3qg0A9e7Xr8Sb
RTd/nDAJ+nOTKcu4o+fOfRagzkKVLGUDMGbH7H5ZpqFM9Nu1B9aaEp4w2m2Cm5vD
yzJC4z2quK5HmVDTxunBTvyiUezZIQ8GnHEQ+Cxs4fP7iXc4XSArn7H6oXIJefXS
P+7KD4Bge3LXcWnTFj5wmlnTAaWV47zmJnlUQVbupPrr7hibRAdvz3DL4QefA+X8
dOL8d3LTlUavPIOnDqwpHIDJFR7TUyaPrIBzEA78IytLuQOu5nGUDj1mwHMGSC61
S/TltOEu638DXIlWItjI48Fs3ROqwF0nOS3Ww7+ltRujf3wsWdmZ8XO2Yl1F8mcT
8gU4vC5B/2ptnmPp0V70DnWG8W/BAYJt6OZN+bBgKIegQ3vaOn2uaTRQjSVb6bo/
F/ECs+VppkwrowrvojfNmhtEjfe/KpEbXVTtxUcu+RGCJZAzgAe/hrn71i2Mc4ER
wbNRURSFwVfRiHN300Lws21MNKhTkHICFXtjNqL3wpVfvnBWm3x7Qpnz5Nh83MCo
vTpyLL/0gAb7m+f21/ILu+/Uyd+JfnURhyvM3hrVeBCIeKnfRWBJuG3p+YMCyGLW
pkC2v0XKvPg3bBidbT0DFiyXPfiB0KI43tTL4EBqIEGsmX3pQCQwmImUU1VC8f6j
TqVo60ys2Gf0kkCzTdO6nWU6HhPXsUwKml49ybeX/EWgIZsTCecwyn3INyOqGkQT
JnytlZs7lHw8rm+l4OEbYSXLzBScuRwsswVxUL2ao+EJt2oqJmzd9yUv/5F65lGS
3eESat/NxAAgUP06CBC5gxqT429aXrjv8gzlMgRzbMRo660OmiW3rStjucByTDAw
tFeYx21WYhQcVXBBnIdmgWe3QtU+xH1K8kOjxWhuapacSIuaUq4JXDX+a6fjN9rR
cn0JQptzbgiHFK1v8mLyZZqUJJ0rbFRrgnuHcUU29Sav4AXUTGgTXAd2fH8mJ6Wy
g+Qr0AXcOksrKQHkDK/Igfo2wCvRSoPKCeUaYbefoeyai8QrP4JTEIUSpNxMq+xI
NiCdnCrDBHbgb6UBUPdirm33aRGaJ8613nAoG0FWR41APsS8/l8s9rW6hjY3n8yG
UsRf9cW5HJOPrjQ85IoTQHPJcYy78yO9BIg5xkusGyFoC8+c3cN8ytCBW3JUxMnK
XL+n+o7uQEtpOKnh4ocFDK+8mli+llW9m8kQQ7TwiClbfqR/Qhqx+hrRGLEh2VbZ
SK5J5ztARKSh9qQLGm0msba6gXXuyjwOzz4QoulRKlPHNpf91Pbp3mu6WyxBTlAi
8uRlu3r2022Eeb4Ud9DReOmHX0dkc0K80vOOZMn8q5Uh6+cHUW7TEBHxfxZVSOKn
pGdqr3Ycd30yK1tqoqAwqkh3Ek5y1297iEU8DPU87Pw9TaMPwC49ooc+rcd9TjG/
cdMsF4FoTzOGfjHDlI/ekfi/NGvweibCRhGDZsvF/X5d2ok3nrdCdLMpIOZtzJCx
wCiqXkO9z4LJpbBab4rcDFNGJ9hMF6BWnsLW/Xb8KGbbdFrbAGuadxNV/LNPAJvJ
pZeHPpGoSwtADCs2ifZtNYSVT2zEKvMClsN90I52cuYu60UBdJBv7y01XYeH4pgX
94hOSX3gjCCt9/rz3p2iasTU0Cr/ICxhVsh7B5VQnqb+M7Bzkc89ZtXvkKWKXEgD
BiafhL+WwQ/CaCDWSi/JHF6QIEowKStJKqGnNsuiEffBpf9AwPDMzVGQ6BBOYcXu
9osTf3m+2EjqCbI9Z/hozA/h5VJ48j3KsFGNilNJT2FbUJODQMShmAzDf3rV2Bht
tpvsmyhAM3yMAuJ6VLYRP3fUrNRa5kdODla/0SOCbRjBoj2bwy0Ut8TOmr/iBI6D
vRLPhC4W7+ct0ViqU78QwkMrDIZ7m5CAC8P9a7+xoo2VUc7VJ0dhHCifh8Q048ce
q0QRcVTfhmjvoZSCIA89Sdp/qF6X0UFsbq0e50FEAbsaID0DBggYBWySxBeDx5eO
TW2FLPKMbtIFg8r5Lfkqca2s8AsrnM7MF4z2oCDYFyl2Lc+HRPkJgXhpA3Ta9AZv
DwWgm5EeXY8IEGn2G5wMW5q57abh8e7YLZrY7MBx3dIG1TaxSzc3NZa3ch69q0zi
dyuwc3wUDedyqUZJ/4ddaYaoAnlj1+4KswJB3URRuxx3QJc02mhHQnvKuHpPrvhN
42swij7cKXo4PjCxm/hLA0tqc+76HcebRimUQ0IvgOgOZRNxuKKS/zCtoLn5Izua
k4ht3j7DhJe0P8xcuH55I6fYAGs8lZpCDpAwoqHjR9nEpdv/TmyU3Kxlg2LbSDpx
RbWis8EsM04Oo0vT6ZG9Q12eDGj0sYJfw9RsB4tqcotBWsvxw3AEgk0rQi2J/Rfv
BDdSK9FMbITLkJevFPp01xM4ZevzWs59XvE8nNIyiLeySWQ2qadeZaoSTaJMC0pb
P9UjACbiuJTmSKFAmDuNE4221ytnYkwNTw6Zvkzo/w3jJrC2Z2Cfe8dw0sRpjAix
EPt3d9+SY2cFB0V9/xEyJiQcdSbGytS6SczJpZ7VChZ7Iuy3z6GoN1j5gJJ+70mj
KoG74N1F/lCSu6J3Ab7jnRO2r4huioYNgBdeEaFE4SvpxpOw5wz8WRdLM9Ubosem
E2+tWWWE0xuyouGkrzUQV2DbzDOTHFujz4ltBrsKNz5k2qIRDCd6+UOYOtPY6Osz
nEQGZ427daa2lyDOG8zbz7oC9bk72ic9PcVgLLALFvEbVsbbXXDKKVu3/bu6GY65
DnShin/1PxtoLIgWkBbx1FqbiFsFnjI7wf7m824XH/Bs0yHoZS7U984MMCOP/TRk
S0Kn6bu93mabOJQql11YQA/gTtnzMpPW6FDDiNILTRKO6VvyDx1o7xdQ2EviUeBh
i+1XwEJFGScRxEcvi/tql5gg9atgCM+3W615/BwppiRafniXQUpEynaQEdkyy+q2
LZUJv5fRVvVQahbi79Nynq3xARzom0rnEf55doZ+asJFD1V7nik4vGNfCVqDr8sf
jB3cN+TpH9bYHefmeGPqWIznJ6yXZcUjmuyEQR+9OXfLB03rNEV+BtQm6FFh9lZy
mAGYKgpxVqwzaD/OkBu4iMCDjioGHSvmeridkH/RDluXFJrR0JTZ58a7PlLQlcRu
U2cVig1BlFYCFTmd9Taon+9gC3wdJUyh80pSts3ey3/aYddX7p5K0AqIJdapSA4o
WhI2F+CrZrOhgRu+B/AjnsxLe5Wdm5AoJTjwNs6Zr7c2nc/sJPhdbkQwdecWMlyt
QwrzhH1Bv0DkQdqXwdEj9vhm0WYfoDq5FAWOWoP4kLjF96GK6IL8NRL/ev3sItUp
vcAgTumkTL54zJlTeo5oWr83Till5edzxe8WrNIY+Zi2NxGMGF1KhrBNGbxCZzgq
3W0mCzcKgQRb7YYkAzb9YddJXDJfPB8J72oTkNOQXAnMU4fdAWpD4ERP8hJQtR6C
nBp6OzEeypn9JvFtgLbcfkk4MeJYdF1Km1hrzRF8I/Ja6RX/xjBuKV4I+toKsUmv
rP1mdiT5dcsho2xnWdZw+AL6q0yTMd8sqWYtdj7wIrXJRBcdyHHvgZWAVHNcfBJM
jxdcXs/QGJQCdkXq5L8epGLksx85zMp5VACsddG01wf1ggzCESBkOfJZUiHbV1Kj
3OWu01Hyw3xW98uhGiUdqcRC59HEc1lGHbfEP/5YWGuslzZTsNUVgaXhPPtiKYUg
Po8SuOwx523AfLDTdMKQa7C0cPxId5/LS4g9s1YRTtA1yZio8OG+epIOhUiIaB58
2bk07D4TvefzqbY5Rvefm4Ed7Lo7A+FXnkH8LYD0a9Ha9EiimECu5mD5ZZZVXxyt
ishCNY66+EiccvUYKsblG8lnsKPphQG5I5RM51/LLCYcwYif9ylvlyNaJ2Mv5jEA
yzoLWUVhSLPBQtAvSGmqUDOPNYVRh8G/Ej1Q1pdmCSVBuAFh+Zo+APW5/IhVmQGZ
owvyGAN+/UENEz1IrJW9T10eGn4chfDOKslOtQ4QwrVTW7c8hnfD+7tsLHZHMalI
ExBnQtpOewTNelyThtBb3mHwuIlWs043sXKDq4OYqzCuiN+AKbd+xylXfDj+8J9v
PwryL8tvDW8ZVgp60mbBtUhjEKOJ5AeUu7/1gpvcBJhgEmRiKCLbvuygdFDUswYQ
xWTVtO32dxBlJ+29BQou9H8GuYRu4n4pn5Ab/R+dIgwWM2V6gxqfM2fobtz8klfH
D3XpMma/2wTfJaM/TMkuTI5jxvXHXrKkaGJ2ZnvjTr9fNl77VU3KENVmLAv1EEx7
1XOvYMQ1NmQk7udCWtc23LTrmWj9XwMwETKSa4FpDhVbTW8g2zkYuDHyBv/xsp93
Gu+yW5/XXq6Ps+hC5J3GYU+u3CGB+wZI2Ykgpx2HavUzxcmvd+kj/gBxHbomX6GX
qJuJ+u0KFc24inu5+iScYn7xlQjNMWhJsJfsQMq3NecdA0De3DePYbgUqRROlN6E
iwuCpn3lqnQ98ksQ7F4BjPACPBYk+lhKwlgcV1nvUhJZVztNPPxfBX518DuS1kHk
LDOIy2WUCg0imWZLkBrkz61LouqPDj+RkmHlWGshP6BPCOElpNkVurYj2iqFnHRO
SmQXNPy7g/hb939hg8Fwvz8iq/ichL2jd6cektVtS9Nv/4PoWzFmIWb9A5PgtLLv
+SMs6VDjHTxOfetLIltyVTPyEl5s31VGGyW+afS9pavIKtYm9ERfjGdAeLvugwoe
tEHpeHJl7q8VTztq/ec2a3XYkwschSXW4kX3w61mLt6EOxmuEZvKo2hqew71F+Kk
JkAwljWckxXiSVvZCbmYPI4lmhGJFYHQbBwPUi4UBwQ2+BtfPeoLiA7ANo672usW
eWz+FWPAk+bZPsJhT6N4E+0axFpbHljiW2AS+Yf2onIYwW48ZANQwwjTuXP4OjjD
DUz/zmKDSEU7AMHy0fe07zpJ7gpbR4iylLtkK8KEWOGFtz0UVPAnXohTt7GF5wLd
qgdfRVFWUxFTKGv+MctcrhtSGOZRJh9hL4gpMs028Sj3j/Lvv6s13SQzVfUdxTX5
6l3G19WcXsaSQ9NN0cIz8mG0DszEPj9sez345exkBs1iugGaP8F5FybSQwT6awDB
TXl6kRM/AYAWyKlfTiq20VF8Ed6+FJMTZ0aQ6ycl/ux2I9/zjSZgM+uU7L4g9nhT
YxfY9v7iRkDyR1hYrxWqd43Qz6520f1mpa+GscJQzU8ll9kXa9d0Avbc6caNC0I5
18LxR9KdY7gepUTypgd74YJI0GwYQ7r4uz3NXpLN0BQbOlrWkNLOUm7Oqngn4RrW
/j0kwZR5/HSr3pamZ7ZWOaLsd/mecSmaJeRpFTVnChTAuIA3xjZpRlp64Q6VTWnD
xjm1l0IllpW/vx7sYTqpGTaSIwB59UA2wBhcnb8trxzs3Daocyd41GCXB/ZtU1HY
qnQ2DNGJ/MWAiJiVEkJRrTXRITMvdoKWjwuGgjN7th3zaACT+Fq6HrlSxlLVlhOT
M1NZHCaMwcLNzqH1VT2KF7aaTwGGA1HJx+/gMFtwv2pPS2sXvno2E4RiGH7bGdsW
1OhxFWKU9gjNHLzINcUkDGbmtUr3pW9rlqqjgXUndXCS6hXl0NLb498VFK/eFc83
KH0CHsrFYubphh5JWCbUnJGWIrlyceKHdRctUXKJrgwjJT7mYjR9mpbCB2erAGqB
kYhcCGU4EPRhF/E9sFoVwDMdAOdEKWuBfwUsLkrZ5KvLNVp5zXotgFmspk+DIaXx
A3lh6wppMkOjthMTCuKfyrkHcwmUOiWFlQMgYOBzxLfTN3kwjQxmMWF1OyDFuuga
zKroi49fzGtO3dlqulV54XqtRFbMbE32mVqgWCzZS0RtX3FptjHj8uJDPdY0svBq
fxpYHlrOKKvd6Rbg06Du0CYh8baYZ8Fb9gbgAVEEoibe4IU95LTFh5OaIXGzWV36
tQq+UYsqrzdvAnQ23IdW+/v3FnDD2AYD/qICqXnmCN02SA9do8os4nue6b3nGqFg
uSgTGT7c1MAYjn9PtkHBXo1+XTKsSB5PgzxPMrQa16Ok/PuXJ3FplcDqfcphehl6
5v3bCEPWKlkFkuNVBfEoTCWRkEE1S+HQSSXkNESO5SgG+8NznxB2NSe2O+v9Ql2J
HqXS9xL4PPK4sA4joduYyv0+F43j9D1owywtHpoWvhR4W7P+5sk7bwvDySRgQvOM
k4h4uYlAtSfRfdTlCFE6XzjGDNAT1nrvlnSBZN+EydABF1hB5/Z9smtEMPJ6mSmz
xAhfxHerCvxbma1+c7j3Aa6NtSi16awCwz5Tz8PeI2ZFk+lHqPqSCcsvwrvHm3IL
Jz9GCVwc3UEQRX3rZZkPa2mzM4jYNWskU7DzJ2J7Ws0qzVZxBfmMb6mwJpQjROoQ
hONorWdLYiBpU9U+OPWeQWfFIq2MHZlHuQCUsouSZFyTDyoAZvrWosaYUy6ZlQCu
MAkVt1ofdE4mxUbtbYwvNysdflUJqGKanyX3tNhfrFq6VOrkIJiYX4lRKRKbMkIj
d7m44mn9qhxA+Fa0dMApVR0ra6xH6hE9LLjUQblXRUcKbgAu9Fyshi+zykr9ShRb
a14DtVo1PC4tg9m9LabPy9D/dZ6Uq7U233VmcyhEC3Ee7uHQSj0AtqbdoJW2Bg1S
ZzPueKrEk4f0mrGRTt3qf2fjlwy3ra7ZHd7FTlXnreZEusngUAfg5BdngaBcIGBZ
lBtQZmP+dixxmjx2uT+2ZfuYcWJYrrGMjrklOiqkxnl0Hd2seLK5cjGu58uZiuwF
T+FTeBpCyZFjsYn8gLhZ812L6CbbzUC0Pu7I0wDkXuimEKSnA3vU+QVtIhfL9Jbb
8tETkoMS8ZTGm9gWHsyhimedprY84EnACW1a+Lglz1MP1BU5aHdq0HRVjLnofk3O
/W8znLpSUZG99jOWXq0GkJOIlBAC+12lk0QAn9GmxzsAXfXP2ckCeVYV2IIZsaD6
dyJ7ERS31xVnHL3tQP5RczC84C9xaAeFhXkUJgsbLAHyTd3/i0kU2vy8i4neYB5B
0iBldNEH6uvBFc7bOTwMCNXk6TCHEqQ43pFIXQdf9pDFY9wHCa1VCBLjEOAGJUMK
/BUJAU5wVVGfpBMLDoUosVg3uLoZWewJCoJhtsUvv3PFJg3RwVxzuHRZej1hbtxa
jXyPCL5mkaz+RYA67lu+JxF8wokTyscE3Uc1LAzrsp3SWp+X8jv2ot+60E8GeR9B
JtGOIhyyHkHBnrehnnM8+yXluDsSR9dqfRTmf/KqLPksRH96lncvnMNhLdJsDN5Q
agKBLkWt3F9X4XKH/n8NZuUzMsqj6LDdX4RLzxJ+vy2Z60lzp66wu7YylSH8Fq2w
ewphyFIi6v4/+8xlQDASGZEMnok5EWusTOnFjAfqPtXPNRiihk3PYndvLU6BkqAJ
USzc3NqTvN+JKV4k2f6Q24jEPcbRACo9pm+exgH/uUg2ckKpUY8G3JDRzNFPAEMR
ZzG37CMV6PA+kCpXUiZcz4t93qDAn28TG9vOgfPFASoxd0odhH4Nyv9y56yNelT+
l8+lJP+hLC6FaDARmfQWR4AYk4sL47O7Sh2l7HvAE9f87djNBut7kdYxlHxWsWEK
i3HOwN3KOAjTWjTL4HnFK2HLjvVLTOXk+gfCUusASeREl1wv3Wg/lp6VCf0+V2AT
9XVuvNa0TU7wjphwfyXHWpCKX6+rFRGs6z0m2MjeFPg2bJl+HnaLyJjeHvTLildN
tcAsVftmhEIzx3nZxU77v8aHwDU+WxXLaSBRM/J+6yg8T7AqsazdHqlvX78We0FX
M6GkWZi2P62NLupoa+RFXG0qSoGlCTKhQ/a6qqViAmHzmlhPdgQwHRy4xfjUZeqI
0fTQfUaVwPeityMcOHwnZT0ctnm64SikByidx58RzBMssDszVPhTBEGGITdkWihS
qLWNL018WC+e5BAqWKTPLjc14PVfV2LRnxUkhNWbA41RjByLlUnZZWazBPTe4Vom
+vymuU9QuV8bGpgFa+hfDt1OwwtsrqP4QJLqxfv5UY4jQhXTBswRC+y5frmT2Pn7
qCjVSr78DizrZbtWFz2xGErWLO+og5rO7XZOuxxiwngZTcgQKwVUxcXgZQfDWaTT
z19eXc/3LmIPw+SYcjtSyEfnHL7/GOuiTG1ut3R6lfDQx751DoHpA2MXrli6dT9L
HADzwQi3Vox6mfBysPU7C3G1GdDNs2B36s1HOmeAvZRaXq0vyKqji5iaxWPeHCle
nqeeHQASYf3Axncdd1yfS3R3LvYhfFJAIJy4xil73hf/g1QiY3nYefawc6Lgqqbc
1BAmsZDhCk4nXJGvcyz8n+LJDjmqvaBO2ENbJcctKt1Z8Hf4bONdSkcdsFUHwUxg
5T79TZisQru1sMNe4YPqXLU/Af5A42yNlXhOchGfhpKRgwWaUWGqOljHcg4bObpM
IDc7S5+IPKFCKWrlYJa5Q8WTAalnoeJp8wqv4X41kISPywbrrAgmVQDKPJemsDGW
BuWD7coSP5NO3Gb76c0TFfjf2psP7egr0VyZb6luQiWC2JnJGCtBEf+49wKU0vnQ
U3AWMbYt58bBYYE3hhSS+As+Ebi68On8MMcUUJ5VgQoDUTj8PdZ6Qy1dlcX4o1jJ
ooaPYz/DSC+OFo2Im1wFNeh5Ph5VYlDPSl/0pDRojCQI6koTKalQGZsN5ku78tjp
MP8AV8PuQqVfid5U1jqeHnyNyem80N0bHSA/f8WrchNRMP6cuh0X+c1YFsyKpgF7
jS69aq4dIlmgW+L0gyjBKLrISMpi1EQhC996U2TeGbTYjbJO7nZWT1nm7SQIlK6L
9TFaP75jyWZsjikbFBLf0LJGfxyRdv6bRw07yg62eQpZSfJmOOUl/iQNLRxrUaoj
fF66bjkBNbBVv9lk8H07FbbjkrHdprjgFyT6EVFIFR8CnqGOb9nQ09Z2BiOzfPD2
BS8PdjDN4BgJEWnqoUjY7NkEbrLaUTaJpb9pPor6cobS/djJUASaivoGo2o57Flv
VJOi2dqK3Cl1ymlQEfBURq6+xIRC515WmaV8hjijD8u25SH3zwIXtvZxFEDco0Fj
EfKLqlzbb2q/ZVRl7Cm+ELPGATYEQEgQiluxQqA/OXamtzQOIvrM3lEV0M1FPtHx
3EScHu060H0NSR9gZJHWrmrNw3Ni0zjRLg2u/oKBeyI=
`protect END_PROTECTED
