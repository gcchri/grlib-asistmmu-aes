`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lOKe75DZ6zCgFDFm1+ZFmACInNnvZdXMf+Oiimj2mrIy2tfuoODs1Qsl3vo/a32m
kH5v++WMmqLV2yDW4g9YLzdLrmKmJnY3yNbvAJs8kzVO1PFqGNs9vO8JI504+sRY
plfjKP9sQ1ikmtOUgjqKTt5W/xM0ZR49emhSQUwimSTV5qr5iuspdmhjn6ZWoOqV
oWY3JNBwrMq1GXJxTHqZW3EKs1JnQgH844AWro0iElCk0r/kO0V+eZ8W612JW0Qv
CRVx+Ax6138MNa1Ii3aasujo7K0wW/SWAHxTG2jSNldF5mS21ZccB/Z1tzup2sJ+
L/uQVlhXIBAtFs9PjQ2e+GxnC71kjjhVs8ugkRkreRyNF288fRVVLIJ/uNSfkscW
x4XOSymJyPynPufq5ifpzS+L5uyggR22gRrje8ios8UBNaeOrTX+U14E/TFSLkeg
qbmTXQOEHLj80dyVF8O44HbokShIThPOZB91Nd2flXcRhHeq6cj1psWn7wSC73+c
yJiVTbqs27qAnz/DT0334MxEguxujtnVSYx+p5/CPpLfEe6IIazc8OoVXsYB76lt
JWZ6oy/SA6q4xKtELuTmGuH4TXc8hgU5+xS2yuDhpzwIM9yJzMe83mcG/vcHRolw
+IwKfCiNNtSFzzaepw/U4DFA1qzsNlflc6yJbIBY8sFAQ0rZeTRh9nvT0RAs8ct1
xM7DxUzngwolgccpaCN6pcnH7QOYAoV32XS5DL/v68VG2eEf8MVxn5rh5K72QDXv
g3AVypmb53CtLeHtkfcSeUIFXvom2V7izsRQHOPMses2Y5Z6TbKwTaq0NmvuBLnV
6rKOWkpKPpHkLRvgOhDZ5DuZnPYk416Mm0C3xShIX3jIF3GEpFiNeSZI9RSDvwJM
s7nmztNYMZ5ob3ncUY2LYF2h/QPYno3u9qpzMFOSbUWRDdwJTQXqUTBxMp82cGqG
q4GtPCDoQnWqlsTNhhZq0lE+NmBINwtUF2BvPf/iksZVear9CLCvqRD9Uolp9ReN
ebBreSUkYhlhht60zdaFxWmgK2L4guIvI8PG0tBHJ7X/fdRdd0hGgop1cjiOu5Ya
SKYyAd1b3j34cCcEds6/amXcjTBc6UOCFjfl1gMOTPOArCVsDs5+6Rz6rrKfkL/5
qJt68P3MnDoVb4ZjNQFG2LK4eplmaGIumK+RKqOpARsaZgdLwZEhcV6nketMUDUH
qvv4DGx8Ml1LkNafmLjZuHjW1sVp1zditJdTuaIwth5P7wgF+RjivKhcDHzJYTmZ
MuoR2TFX6zfTfg4e7Q4iEcFa5TXuMTtDhRHjaIAOVzWB6SHrh7L2ITKqVO0NgnkW
1NlWj1gB6WYVwqRVXAijWel92Ce6TmHtfreYiFCyF0krw+3BRg6RsMQl3QVEKCnS
RiBeI6bo/Ni76/Q10zQScaBsef54Jje7VfFkHwv67ptrqSaEZKtAV5b19hFS0i2j
ilnSbjIbl9TXJlef+TZb7NeIhspBNi52aAkdwnCoTu8TGTOsr5Iq+9pg6bIDuYU7
MQHsV6iSaEqi9hZ3EKaQPBtZORApnDwpgfBG91gkIWTKtja14nILu+I1W/hpx0m2
BgqoTwlZsVWWbf0g9Wc3xOzVT+3LE//+XJwF7YphTVvLxEQQ3QdfyO6WyDJ8XxKJ
nRLlox8/03tBVo5IpRlKUp+RcxmapOJe/3Y+TjulwRni8NXLOcyY0qwlB6zmxH7f
lbd811V1eBFmuzZUbqOTyNcU8GePFCtcocXEdwyo84httGhXmTqk9Ze9JlqT/Jde
qulhtXRh6c+41tJ+t+3F6I6viqfaImTKCItVSi9TNtkZCY5yl+ZlMs5JZiyjIJ3o
cQON8bMVfC8jS6gxpAU70z3Xqyl1xrewk5yTjg2qPbU8GSLveSnxTbdt0Rhf/Fnx
nKO8Db1Qcm4lvRxXhWhjfBz3sxqf2SiB9+U71iARoPUmPQK3MED6LyEVBtohRqEG
ugQvs4/Fv4qQ0EWF3UiU4IbxmgvBCMzvStQ1gqDirBa+Uptu/Kvrv1eMLVckkUo4
3t8o3H920TldF62896u4QvxJutnjRmTewHDHvjzgN0JEsiVhFDd+fclO9UCyUwTw
0BKIIMoA8TVqRr2gDg5L/eFMA+3LNHIUnhdLvtp0mfmUz037oXK86GpjR8U7y0Oq
GcfMD6pb3xpw72Nh9Ak4asFVzoviXdLn7GJp5zK/xAK39iNRVOI0VfJLPcJj7amY
xgeH8AErN973zqqj2mPZYFTCenZsx65gwiz8xsLDEeD1xdeP8scv3lPUdanW8M4C
DzxooAxh/yrsRKOcNnJQyrdHwfxZq+YDqVR+cB/ndBdg1C4x/gxAPWxnGUpPYU34
j/qay1xst59Forgh6hfXYpNZdMlEtyEOwH1ghd/mDHyOhBv5OEWXMvuFfeRFzpVO
ScqvLwwIxn5gfoWGtMfQEZoVOIdXKnMZrljiqnsSWGD48Q2PgfPrLzr+PH6J5IF2
5SJTqu1umVrufaXh/rxRd5mgOBAmI7lu0q2t7FwotkWdV5CHCHwtVHrwvH96D1k+
wbuWRuSGom//9Xq3g94F3hX/EdRWXS3HqgoZ9SozmOzJaZeJ1zwq3VknPjsVmpl6
pS+a4c/1X0AjzvvMG/GhPB/VemdvuUF2eKMkTLmF8LMuOJRPQUA81EVwevZ4r4oO
4+f9WsIQrM6LDSCgGZ5ezNb7LOZONouNCseRuE3qUk/W9O/1zV9bcbsO8t1T0IDF
JaIUez5UtJKfU1OjtC7aEdYsw162VIkL6YFDnrdc6VS0MSrNSKFrRCzeUcRVnpU1
9CNXFLkrell+l1UGpkf7js0zcIngA781QAGk3SxdUGZKMqS4/8S5/z8DfGmfaTRn
R/iyCAvbKQLMOLmFCd3oExCa0c6txOLnv8EvCLKNIErNXb083HKSOYW2d78gItod
k8Yo+tDHOWD3i20tFbt6bfQnw/SFMhonYZ6mBKFG7EIY2c0sKeyc0P8eNzqwoL5r
LPbhow1PDqKf/YuM0OPJ5k9rxCZ9h9S5tMIPwgJnKUY6v03mR5z5PZDI+p30nWfg
A774hqdb43EDicaPjcsbeBB7tKfaS0MZHMRUgM0AzxfO3gmlwq6LWf/aOqKaFkbC
dcPUP5Xucd8tYnJK5pPMxP9e8Q/9sV2Cqah57EB7vb7EFYKiaeB5JRa/EWrGoxyh
1y8D8Cam3TqbuchnNa4UQZlxz4k9UlHa2B2Dctyk0xD+F6XBljxzZK7yF3QABnPq
Ha1AtB/gsb/DUlVNyXno2l7JulOpFHWoB4XXMVZNObMiW+r+Q8B96DhFGCDkaoAi
OYddoJ5qyuItcFkl1WxOqhrkXoNjTVEfkYl0o6DCixyIPtagOBW5wBclqBwa3TEH
m0ZJbqelEDtYGE3AjrPmherj7K+UAzJSfUfAE+tMLw9CQP4mzIFNsmuxfcnxVteo
kCgrZC16dnLVAB7dkhiLeSg35hyGKk0y9C2M8XoZpQxRrlBhbJ426ikYDenLbhP0
dwZPC563oSO17mpL55LqkjkyjWS6ZPBtHEa6YpvmBHJa+jCeoHlqM4wiNpqtsauu
Bw7nXrMjoVCl2LP85S3cGyYBQqHimfc7ixR3TWDv681Zl7fViPkY2mKJk9tvrmIl
OHjwKWoQcSNdi90eme7IGSH1X7ZSi6ZhscZoT14poxxYeaSd31SfGc386SSPCsG8
aBDCRejp/lYr2Z6GXTrZJujsSRaNFe+EIRGQ7OH9WOwn51ibegRqI/GYgZJVQC/B
TMnmd3teqAiZ6XovhhTPK4q2HVxMNWiHbhc+y3Em6Sk8vuHg/m4upRciqv79eunM
gYQ7iTtAZyArco9m6MqtfCVFmbyQuWIz+EAd5Uji0NEOYoGcdGISuQ2Q0FmUDORi
gK8mb5Hrn5Ud9Qpd2bipgqv3RmQS0ao4MstgTycFUIex7Sr1oTGbMrCqoshsyKVA
OCHFF5X6+iRQrwRZSzQXtLSQNOYI2p+i5MnZ6oFizYFYOaGX5JavpuJrC8QBdY15
3FR2ptKM/UGVSXzgKT5gsEXQeToBkJYzf6iq3KCsMVtwguBuCx4b9fOkftVzctpB
7rY/xKdmD3St/yU1lbWWlakHchsQjY7Cigv/MtMZebDR0YiQYWlVoPDXsCIk1e+6
V5KwYAeDJou6hD3noDIeMWTfJSNayMUBhhyMvuq5S5/0X6wNskrFnDjoSdUBkvmI
pHh6t/p+EYKCzBlPwhtkaAKPsbVfOVrmV1C7C6ktSjQFwTDk/EvAeQmkrlS08035
hrtjskUtyENIvjqroDmpx0XgtOFzCktrZ04VqXbwLxAsAWeUVyF+7B6uFrfZ6LwX
X11/UmWoYRLFevFogOYC+Z+V0UipbUFv+AXXOicicd7oMNDeNqefkZfLoGY8Xauk
V4R71dsEXgHIiiXZ2C29Rf/x3OH0SILBsy7vz6ig6Wp75a1h9BTbfopCVub/Owoc
SU8mBLAWUYgrEAeVsNT57T3P8tfpO+znUR0/DHeuZ02BVyIuHjA+PUP7DnLHJa+q
CLcSjtDOfK1XEUhj93PuLfOflgLUht7hntAYcCxUj7IXCFRGsvxdYu3GzzU4Em7j
hYFOKEmBECxY0ovXiDNXZ9oqWqr2mPHByU++55ynqksq1pt4d/MgrQ14ocgwBX7x
x7ltI7aRiBknLcQzyEprhDj8//eFabu5ffDRppztjalccBYKVWp94ScllOetkWru
U/PU/tFjqGktUGvdKKktKxCJyQdqMJ1gP/RoUGFwx8qULAMwhIGeaBel041vThet
`protect END_PROTECTED
