`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y7eo64Ca2zDUDrXdg6xlzhNkw83EvqcPPFUurpAS0ty5cOgiqemeDNNszMnz85U2
ciEQEa9HYOV6y7EzN46lDlQc9J4v8lluFC9/r7gMADt/Scd2oxS594BMS0TVbMmv
uL/Y/OdCg7hp/kKIue5n+QUHxvS4thwG55GK0xCEyaczBELwEcNElNjuad8ZNRzs
QQG5mFiomkjKwifqmS6G6MD6z4kjEc7cMnpJ/OoWVISawCgMbtJtAND3UgfFCDH7
HWO7/6xZ6DFvprsFpZmRf4bD72CUghmu8T0vN/hmvEzqSbQuh6+WbOHqG/DdqoLh
fi8UmaGJFvz2vbqezpLSfiYmUxsyBWXAea3VbLVcB25YgePWR7/Lg3GPuT7ZGns5
yz4jyfHVTH6dEtRZTLu5O0tLCR2A+4FkxtPKRgNO6lBtso/Wl0qlpNnrYDGWH28V
OuH8FIWU3Sab8wBbraFP6yphvhkmkRvbgZCtqnJx+Kvh/IIO/Cd7Z5y+ba79i7re
sAW28dRcIRlj8BkHVWDDtFCsKrpU8bTGVQFkGbwkkuxC5s0bcYtCUNP+Ux5Yc+UD
CMm30tdp+2eHllMuxPYPmXmg2zKYRnhWE6vZuCJy/8SCmLZXZzXMQZaxays3F28P
utwY+XxsGhpLh04Tlo4WfayFkpriKcvVzRCsxofMh9+kF7q/Yl7s/GGOJUXlo08G
TulO8ybceeT76aNlRDoiCw==
`protect END_PROTECTED
