`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kmHdl6hcyMJ6T25454fR+c9OhMewP6wNBgNChfOkKy7n3wgQT8/6Vw5tVnwzqDO/
CZVVXb6lAUYDFfRPz8v1l9QI/MoJ+YcwjtClvu3jjs7zxATpHQAjlrI5GfdSHYzt
tGabswuRn6V81qkyRdPQ4x93WycRra3+9DfyIhdydRyyd46/1vxuoftiQ82LgKTV
LV+nY8YPK+Y8HuKTtkPLNe75HEgx975ARUw3O4VgWQRjtYnakcomVpR2O27MMa7k
IR2Hy8GkiL0mtbYFztRHcrJkxb4/l2UC9KNW+V1Vkda8wPuy0lfDzso79uFcLtFr
tVy9/qRq/4EMK1LpJCVodTPWpQQphQXltMuaAPnXg4A+E6obRIkz1lxHX3lowSkL
r639A03GAqtbSusQTwW7LgHweCzEWYjwKeEcOte1saSn+nY2chzZJ/q52IcYjP35
JlMnNSmSSJcgRrnmHrEHE9hDZRZ7DE8eiZ5rKGpPmn8GCXRq+n4rY0EUQhHA2oga
4TzVYS3PziysEwmsYgqQ+Ce4hpSz7x4B6AHUq6cu0Gp7IiIhosCu1/BbjM50g/G+
`protect END_PROTECTED
