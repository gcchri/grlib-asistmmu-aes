`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D7xERQjTjfdGGi4O6RipHWgYeQRHcEzytgUnaAwyg6XxiSkvPw7pn5vcgbVC1WYN
e2k2CJnSVnai1xmqdmnFoght/K46bDWZgMk5Mf46eElEMOHMfv57OXFRo7oH2mfP
3RlbtnQBxmqHPHYVfVZMfpXihORk/SPjbvqowrrKwu/EkDGtasrhtPWgn8Dso6+/
ZFiYDVBYpr8seuWGwuZSxYXWyXMhCZrWEad4UG99YJcdY/M8+5NTH4vy4B0/t3f+
dHj0y/fCx7dipCHRmEJE8WqqBIWcBWz4C5MJcBsxlc2x/yzofFl5Wyx6kR4swwvG
97osUU/A5vDQ/zfAAbjgKVfBc8VcIWrFs4OyX7TNsr3lsSYV/gYR9NO9DU/3lMFu
3KnuTPU+epOK+L8SZNLo7C9hkG7vN9ybRZFADtU9N42XusWmS50tGcRj+X8680Fr
Ehqztib1Oyev7Na4MyoQ/w==
`protect END_PROTECTED
