`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KTi7zlXNZad0fLZSm2n/m4tSwJFB4WpfQstzhMPTSD/tFZec4RtywLGcw1zaDkXM
A+g+wCy/zHugaeiip+4cUJofKS4E+qrT0uYljq+ck3tB/400udcSpCd2sbcmEJRs
dwM3vXweU09+2cfITB4lZ5OqjsUoctt66jVY+zUtjLY2LwZbFXUNP1SHJQM/wqOg
VHFmhly+UYcC7mwaEUhWyMRWkeokGaHobpIWPqh9m7a8Pse6iqiaiq0LYM6LD6c8
YIvEFOW42MKKvHsOFY/UMnIjUna+hKGdUfQXOXLNlGxCkg3IDc9lCJyAsXqCd7yH
hboEp/YkteRy2frJ8qUvgSQends5BKyUrgfAuHuySKIJN/u9h/nTnQl2HxwJ8Qj+
OMhJAJzKzy3bbSaWfBRY16f9+y5v5TljLMqg3I51ipzn3yzDUfab/7k5ucUfcGfF
EGkklY04KKn0QmPSNNyw8J5LsW7pkyumTyiNpT/KxSQ=
`protect END_PROTECTED
