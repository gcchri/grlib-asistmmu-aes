`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X3SGwlgFt4ejhJW9OtFAgBejhDL9MBeJ/pXAHZyeC6aWPGgWUefMijQqBbdwXD/m
MKPaYgob89ovFupY9fr0WYiAN7KBLzZyWQKRMO0rIEXgAo5JdXSVBFHjtjADfDoM
zL+Q1ZsbCupz0yMsh1CCFR4+nZZxXZmf9/oj+nhb538FPIl8IwhWlHGxObr+I7YM
6ieTl+sgQcZaDyOFRfejn4Pprij22moYrwYDKFfrdIQTFfQuaZY3mJraURVP5kGr
FKwO7m5zw9rixOGg9/4vR2Kacf1/uIOOKbL8qDLBbh0M5VxIA6zW7idyfxgh5wXZ
4Jb0ZSE7kQea1XTmk1kC7A==
`protect END_PROTECTED
