`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gJNnlw4YbsIDfgG7vbTG17bHt03g8VGYz71gO3wk4Nm7GMZyd7drQuwexyAuJLDc
s1Tb8i00RkyQxHIdZuw9IN6uSgSgBOS7+WeB1h0U9yoVtt19GqqjVVnvxdXOMEsP
V8GRa/LImitdHkFhUO48/rXDlq6EPTAN4xA/MH7zcfTMCGrOgwVQH3q5uiPiIQkH
rX86LX93367D18MCCmZdDLhxlgEqOJKcCfiXTIQCn9fjikxDPjb8zL0zmONUJWV0
B4rd2BKlgqgfDR1TKRZygJkrXIm0/4o/y3XHBmzSc3kXP39rYE+ohjp38HX92zzt
CFj1Tetz1cagLqZ7il71DdPPkmUMzzXJc9oksWxpJ5/QZC32gtW83ftE317dw0kN
O4JGZYO5NdAoqsOOPd/0YaXbraNnwpLS4wbAVP5w0c/6JeiVKYxCGLAZ9pLgUySl
vHetH8qBDoF0HKmsD9umUkB4yCp4dH5XefVqh6rsIG7b9/dtTfpdPv0aHpGFjvuJ
cujTdiuNT4fm9MFziblyIZCUOk+DLCwKUn6Wfub/V3ITDJb2hjCp2Hh8QfFD/bCB
42dbx65aUYgxEvVivOmiFjm8d84vP879bW4IzAJhqi6+7bhd6GjZJzUH2y3iEN4C
iV8+ClkVpN1o7tNmMuxHgSEUbM6GafPdOzCgE6N4Z5cMFbXNi86FEmIbaG8/3vyQ
`protect END_PROTECTED
