`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XtoCNsKSQcBCSJ26NQPPk/o+M65RilblVEIk8B6l6BVfalvAM4GTj0pfNMlIqBy2
XwPSyqIMgIlg7yuHQ1EZ5lfVDBmpY0KaiclIVlJ7hgOQAHTUKm08o3zc256GKfwm
z9RV83OyCziAOFaagG9XErEMOdTtFx9/qQKvTrY/Bzq38GoQ4RNSAEFKapImEDw6
w8Efz+D5bp9e1Q3N52wBYO2DJ4mgYvBJqLEzqmpRS665b+4AGeireC3bKccpdM2J
oV6Hj23XUnuqacqW3EYVK/ruZokYVOp9B5UPEPl3CEk=
`protect END_PROTECTED
