`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xWZccIh+QAKYihqJ+CA/DqyOyLWd1mocXYDVWw5ggByd76X4kW+znL88ptdSyUGP
Dljhn6s7CykUW9ZpaApKuWoXdZr9YYoO+Tp953/EcBikCUf3yUtGW5ZWO6GlzWnJ
Z2+GpgCj0aMmVU+lpheYNAx/fMXj32AxVqG0wkk/YaE5WCvKqJdbSKInYh767F57
9VI96Uqmv4bu8OkONoHqM/eHDFLp/eryxnphL2nLbOckbC5UqVkZaQngqrQW2ll9
kC3zdYs19iP7LqERzzafOFFBc+HCrFupEqvZbpI7Al6Gv035oNNJDPaez9fcA7Me
LlgIEiuWsMF5pMqCI3JH0DffHX+8SiOMyxcecz1/eNays++9ofw7KWuutcOMa5a5
baNqF6pMUnqLw6nvKUkJfsEcJRL9C42yK7UfDWYAkN/C6vIiqHBZ1697NirsEqhA
zuNSzdIe3tpkFrDy/nJ7TCQlZiadn8MBvkk38ny0uKXFoCLLMEIUbB6f2VQKZqA/
wZYAcn7zOsW+dIrP5/dTX+aBOrQ1dO3v32KSBpakfEFxfPrK208P77uCAII2DtpZ
fYOak44WyQO3H7bWfy8rIxCZUNVnMlwGGM1YjFXLUBq4ibAyL4/TDQ2XGkXYmpAl
14Iq2XlTvYepOiO4rx1C/59Il8StVfyFj8RjnmI45Fk=
`protect END_PROTECTED
