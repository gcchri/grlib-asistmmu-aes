`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6vGgLJxWP9toP+oqR0+iEgLCvpCGKesmJI2TKtmqFS2IKbdmjKp8kvh6KNbufB8M
ANeIzWgN4CSWAsPErXddOSy/GwUOCIDWTdkxQwMnLY91ClVRUcceo1AUhJjlHVN5
XpwkqA4Q7kf8AtEMQBYRXQzEcTuTJIct1HTZi2lhRLqbn7w4MQKK9W9i2qvpaTnp
C7s2JK+DNFVOuvFLQRKfvuyXKZwyG1D5vSPVQqPyiXifMPdzwO2k+LM7rPWcGZ98
jCrCccfQXL2PZ4ZXkTiqmpMh2QiuKv75LQA1HdHMTncC/xjQ627iPNcQcYFi55+2
bV6vzEqwFlldeGCW3DMZWcIbskNUOeyXd4ZC3znXBJ1tNwQ1Ml+qNQe/epO8SmtD
NzaPc43wq/t+0z/TfiDsZ7u+aARkBzUJq6TIjiMaKBQVMcN2MyutQx+8E6oPCPc3
esni2+pJKFHKw/qIhUEYa20cEdCc6GquGJt5hVBRe7jPBRNvBfYZ5NE+gOFlNgdS
KJ5NIbxlqG9j5Z6RG3IitY/WDS2Ns+m9VpKpJRIKqQwhZzx5RgQs6kFB47GeRzRw
EFjauyHcbGuxI0bs/O1Z8A==
`protect END_PROTECTED
