`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oe662zbf/AcBbRfthshEBBMDKGWSEpVuQwwOWHA7UKkcFqS+o8g2Yy/OdZy/hF35
c4lCIRS0A7gjyfeaMQqCOnC7eL5Z9R13Yp0FMatC0pkve0aFjQAsJETaZu8FPTZw
01EOwMbUVjMIGxX26ha7YNmaHo+yIVT9PVUf+mZ0TY2V+Ltq/sR9QQ4jvtgkxqhp
eccOTPXP3Q5l0L+VJNAWfrumVFtKScJZjAgS7rVnSP24/mDXx3rYnE4rUg/NUNcM
9HaBAFMiII/2j02Ap7+nQHO/5KtaiNcTTFX+CHahZsmhD6Ux8AR8NDTbQvrryjV6
Lj+LzGHDllWJLbk5eCNohV+laN+lid/rEJQ0UDJdTmwODJX/zwbYDlaOWRv7d/1J
P7YcgmsUqimfRKFMPZrxmUx0QMQYqUUxHksRoiE0GksYsSqVF/a0hBXa3iECt7YV
nJ3d3tiuSTA949X8nIkMfQnn75ekYZOLlpfk7dVYrLXzdmRHmOjI2jalefco+8mt
INGutYCIdZQlAT/6apJoWnjQlFqrV621uo0S4Pk5grkvH2Q7X8y5KHQ34ri2l5+9
hi2wxdiR6l6QusmXcEYk/NgNFJuR06ce9TrxNXDOjJUFphmSm1NsDRd+lgnWpp6h
TVAAY5RuL5rkmHrw92+MJ/dBs6WPU09RR/Ziuxseh2MdaV6XU80JzYKimxjsfLFp
zwbbgvHg5SBeJ9+JUUxjuNzfkeu4hSOVflz3iF8Fj+ze3vgZqcDuCt9t7czZBiuY
3HlFVtOvdnCHspDMV/oqCkQp9/P7KW1E6NTFvSLQ1NkDkx+g54G5CtX0MOx6Y91B
+k4wqz9Dso1OJGddbvS4maukgxV4kl4J/pJN3OLRJrLBflKTr1jsC5TYNPW5mJl3
BBSZNFVRJzwnmFmIPZ/2bimUZGBL+5cQStgsw5Elywg1DQD5tFw/NSsI1XBngXf0
annOavV2opoFqOZEpk8xMlImygA+MSX6S1XqOVItKQnitgDLXkQ2BZpshlp5Tihn
Ig1B4JuW0BWsnjllNp36nsXiRYELVA7XYZo+3QawHl3fneMctrOFPI/5gjmri8o5
+Uqh7nubHunKtFht7iwsKjh+ngmgKj+hKBt5JWVXED0g4zvd6SbkV3Bdwka/meYk
T0TDhbLr4Nj6orRtgFM1UIYKKa3o7zF42lLZ2dxPgMmaga6RQG2cHgw5tGcB/EJf
x48hxcBMro8DmrgZ+pADDwCwKhRfAcnEYEfiZoQsopxUNt1oeBMEWINPBrUtQDiK
9IZp+19H++kVUxxJbwB2z3C8XS7cmR9TjUE+94OQD2gGH+rDuHzCR+z5A3EE8ZOe
fHW729gfK1S26ppMKCivYA==
`protect END_PROTECTED
