`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GCC/yk5ic6a53DtQCgMr71tiZAD7dePzDiddrO7s8lyB+yZ2OlDfHwyHrpNHKu9D
U2LoDjcLKc4IfawANc8TWsP5OyQdao2tsuPekugFS4VPEgG5eviAClyzKAv/84tg
2eX21NYEOvCEKtDuvNHSjEr+hbdJ9dl68adpZM7mWxgugNvIizr3Kr62ci0/lUDU
KObjN/YD7DxO4Rmm6MSjG80tfgZ0PqSEy6sGQoCbNJ1lLJ+kcUY0Enuu/byupxEq
s1WjTiVwmcm/2NZQYl3tCRZ6L1Xamux7bNFiaL9/EETRJtEU1CTNNpdXDyuxb9gT
h3jBSW6aBPIvDVaS6bvM8DSrBQkQ/JlpXuZJ92Oj7E0NBdxGdT7svnuln918W7fi
XPxjJZrGoRLhqZa2re3PK2GqdAFBdVMyT0AQZiExmCQ=
`protect END_PROTECTED
