`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rO6g1JrEN0SaBprk3KQNzBrj7yUKgKuBD7e+qvMQ8Kv1OMAmBCs/eb8u/aYTA8jO
r3q+PxixXw42OEikA2yirThSzfkNkZp5G0SqiQI+MpAMBF5x3wvoMk0+ExIvmtfg
k9jXZ27kt+QPQPmq37HoVCL2bMGxoEzFnYreW2oQXAGdWejngITQTzjKNsBP9NYs
0+RzhrT7NYdRkMT4OaNdR0S97GOjlkK4vDneTzG2nuV3qtpbYBQeRdmlW0KV9wrG
eoIkSKemeZqWGFXt3nN9JSJX/OrlFjf2FrutKVTK1MY9PNX9vyMXzPIGgSU5LuGG
xULVYGTPqq6t7TBPJ354SkDpMtSy+AdwbSa2cfSXUf4hbtHjWQ6AnZubol2FpoZF
HI/5H15wyzIQAoH4I09oe+R/6+tyRBforeKMsbuieMyfde+iQuj4p6tlcFfBQcY2
3bLYfx1aIYWgzCAMuOE7tuIMfbzKxhT2PGG65oBu2prjYeguu1yqvFM97qsP4C8I
dS2WztTK4Fpi/O48Lzao7/GfnkKIO1Rgiq1Ob79//VFGbkQcpPM5sip0P0mYAV7p
koJz+8i218HrZQ8oHjW+HQvKWFs0gLuyz4Qcca5wf9D0GwhSKUTBPSEFFdmhahMF
D4N7jwWaImpjbU8R7Qa3QtgsbKCXj2uIrUgL7gTroFUc6r/YngzCHe2+t9Q18t8b
qnT5pJklrck4Dpf76Gd9PDsu8dMVymbgQw/nPpBdIy6W6bFhbztgsMPcER9AWQij
en1+uIwjWfCWWz89F+1N3xtO6ur5NsW2kku58p0GMUsECTCpHo0ESQsrOb07F5vD
2mHG8IW0SJfumBL0ZmCXPhM6Lui6vJZXC5Gyvg8x7e5w90rgFYQMVmZGw9vGSfhw
MhgKFd3r21+JoM46TSp5O88mlm6T2gd7s+ZS6lWcpLB3f1RD00RXIIgIO5ql5ikR
rppEmc8AIDuYbQLMVDf6Z33lMgSdm3Gha7TznOVQFQ83SW9QoBNKtIyh1NS+1l5s
nDF592cwLimZgLtb2Muna+v9RPitEzQQ+IQONIdlRz7K16eaX9GzOdhz8F4+PvsV
mL02R3uHLtg4YHhT+sM7XaXRy0n1Ta0rHIEEarmLYhFxUPeQSHbAxtc0w1+1KYpp
jbRGg/vcVltLjfWioiWHR8NYnrfa3CFNmIFSc0Pocer19RxrLBohpKPDwzQrzoIP
Hh8DJzPLXvGlfuF7iX7ztAjZ0D+AWsQSDFfFoHqMxzUs4/N4jVWMkuHP19YvB7g9
Zag69/Ql7hoQNuDK8Id0HRUbDcZrcRqzhHOPg6WtDC1Gq+FDQfjZ/yzIfbk0Tv1S
uhIs2D3+T6kO8vCFAxDU3jpa291AYK1xIFwDYHsIjDIJTMsytkaIWfVqxx/TvU46
iCWi+g4CoBjAvSprd0TI7bY157f0IlfNxGhgB4wY/obxy51/EjvMA0mgTYAYVpZM
NNVQoqFoN7u1A5LB2x8iGMNjPuG+G7Jknr1YcWw/ljvG/7v2RxlQnFuXqOBvi45F
G8cgap51xnIP0meC5MLZRGnhdd9MikhlJ/k5+gIg1CqSs8CxSICiqXkdJUpaDinS
sWHF2v3gRYj204R5lIQLyK1ckm3gqql5uWcYGgaSIK9UNvKffWvoyDA4EOAn/CQQ
S2YpUP5g4WTjWUxa2sDDaY0USPw0G6GfydVFHZGsNa+1EeoquJCK7EhY/bMaSKL2
Hmh3ETXrL5eQTQfJ+l5H0te8ypdt6NaMFbjCGPyv59C7aOaVLgAsoqF3XWt1Hp4p
fAGuGYlGkLnAhZxg9CcPgDqrVBmWzQp70QNAVXWUyGaGjHzpf74YkWzR2Tmc5iv1
oSXnt6tdAZf/LbiiD6GKxC5CZpePd46JFPJNydVBT9puYIHv+X/BFI8ghRtFChhM
KR0e7SOPI2GwKi5ENnoGZtXyhrxq3RMfEzncS6eTAbOoJkUJWrJKhSixWGHNd2CD
JfcTq5AN5upOe7wougAgapQqDn60J8U1vSyCIdG1dYsCizt/eTrT6hNqZmQ+amuN
pcww0UOUgdfAyTVAQvTVmu9XUarxskVG0REovm8aH3rpj5EqRAzvJEvSU5NrWoa2
hHApXKB9I4Ky5ZsXIsh3yLWcXy0AIEYhChXrE1P+0LnT5r6hX4Lqv50Z26KCDpcc
UfUyj6Lf7cwkT4DKk/UG686XiAHIsFVPuTHEKhnJQZl5PV3galhNHL9KkkgYGxgD
/+xAjk5e095rN9cKr3bMHAHISmyQuEr7l9b/tiQgBPYC4fJ1EV8eRl3AkOC2n99J
TQjmp2ldLtE6UwosiacbcQSXWW+8DVUkoYGBEUX4CbkAF7EO5gcrni1O6S4HJRcG
SHs7aRASB7b40s9IxHEIAThBx4C+nixQIz4hqkCnTl+MIpQOGCWFmwmGXO3Qpt++
ceK6gCnrCRK53AxphTGCAohNQgWvLzAtOJueff0MAwuKxPz3R90jFUiBymILOMQZ
QXh7/Kg4aF/TGgZIdvu/dLU6rLs+wZcmaTulZ/4sH7i4CeyXPMbdmq9NbL1I8tI4
shNKcFgxrpvUpSXOHe7bvgEbC+1MCzRdtaeAPTNGlDk5CzhlpMgrOgnemo3uBmh4
TVtlIf75VTe69hrfF+9FJWB3EyN9PT46s4AIDbmAhnaep1LpaWDaJIpn9Pl8xlnb
9Fx95ircQ8NMMLryIBGp+/EfTANZ/I2rbNARWS649rZ5pHEryaCgvpgcG2d+q3iR
BpGONynSFCJ7BMkxLv7wOTT5PC6AJPs/vUqGUlAFPTNkhbikj5hB9enyDahu7BeY
oNYH2qKVXxhzBnV1QHzKdOasuPDzjcoXWqkg6oeetJCiZAe78J+T1JprL+gUrG5A
/7+uLCyC/gnD8Ifi0TFUFPeZOAv21oEShxgvTqdBl1fth5HPqa68fDQpTFFPesE4
AdZPzZ7VRw0hhTF4vXRq0a71QtEN4xzEu29fwjteHzofwgriikZ6r3O5L+cIVg/B
YlOTR8NAu0i6Rlk23siLeADJa9+V1QGtaW7UFZSHcug96NQndhH1ucX1UINvF6OT
Y35Fhu3xXZu0CEF7SHvaivRaRNjV4+bhIDKqikfhysadGdnL0ooHrWRE35f/hv7v
Bf9xmO+wiXaKPkJPCjGZnk9OD1dlPyuepAMo5dBnnftdmnsZZMCpweW49l5bUte6
zjFQL+xnuHj2+njMgXy7cBqt1iY7DwCRKdWbPvJed3xx/tp2U6XsUpREGm0QpwqF
A5ssrOGTsyLWX6JUXk9VN+7CQEq+NVEqJjzWMJ8w6D5KnUp96OyzRIWHRx5eGngc
iQcOsPepvoR9d3k7XME/Ij8fGRVPpvaTdlBmAxVJo7OoO/SZH+lwHLJFXLHtb3X4
dFBJV/Bs7oBAH250LH5oFFemLEgKJFnb+BjsZHAlWM4iTyTHui6llgWXZnK59OsJ
acnoiwLZeFEHT7096tWa2I/lb2pWquF0isydJQaXo9YX/qgOXXXVRyY8+8gnpfjt
H8jOqw8Pzdzz1ie7SXmgPVvGHTYAnLXEc+6WR3rsL7CyG9h9VfTB7WrBgABx8P2M
6rilsLO2ZTs6U3u40Y/zeAkUrR6lv12rIZvYFDCnqJkHytC0fsfI8U4I/WP1blLO
nUtRnBJgFWerCgRPyo5NBdlfcm0uwCIC8Y0NfuPdvumxTJhI57pJPz4FzyNx1RuX
XeTC1o94t1pFuS+6wmzrxcrfPB3yIn2kT6ByDwVRRbLAujgpRlksSnPtagy0kgAn
4v+r+Dv0AQDb8DGodXBOqnsONXPjtmfDHpxKlHlAuebHOYojzeqDa0iMuE1uwjR0
WD1wTW4CPcYJ12LvxknNOWI08gLs7OepgvJA7mnijan3Nad4tmzIBb6YZaMJtGZ/
UH4pyOJXKwmkCCv6ZxSGtnKBD3z7u0CkxorQzeiL2Deou3GLrqoIKf4a/0kE5sQI
+nDgWcC/wSiMc1w6lt15HWqj2BFSo7apkZoqeBJc9HJB89sc7rhAhoe79wSJTysQ
BxRTHzHcfwtBnlSWTCrX+GQySRbwUbCkjLquKWimHAqrUzQ36n9gRLPXqUhiXXqe
G/thrGMD5otHkuqTh1tRN3ltRUaHK/ddQ0CoFx8qCbgzILrHd2IAQStuNwdjqDRP
/s3HKVruzwIldP/YhZFjnEP+TxQPv2Y80iHNSTucz1lXpAIGIan7+Yd7PET7DAVv
4kdbczJ3Rj75hNV/kuzkl6RYdaCtkQAJp3ahscJ8GPi28ymF8m5TUS1gmZO3bTDl
f1ecw8PK2eDLA+foPAhn+dB7oTXr87YnhXQbtveq5tamPlxdbHco7cVgl6HlJNAa
7WZg9KR1PtKrirbybRoGIrLDDoGHKKGdU9AqNkWF6I7GGf8oQKxR1MkAiwmz8Tq8
VYvRaTnU4jQW8eOj6x0JQktqkzhUjhUJbQ/o+2qFA/RS+3pkz36wTO0iPebyn1er
RRYyCE0mZ+VPBasghFrquDDEuQ/zn9P/HeGjNFrTRRNp/abx1nrI6xyzWhuUBqZa
yzOVzUSd/pZUln87iP/HfKLGqQcld0wQtoiWmU/z3bqm2DQ5xCAwNg9XmCA0+ru3
SSiB9sSDxzfMkfxVtybKzn5xwKtvcj2EJvCrJHTOhJGopXta44UhqlGvK6N5a74A
hMFYWSBphEljay8vxFPbKHypLOhJBWPEguWdTdNdc6xxhy97BMsJKRL7p38SvlBB
lgakN/WHQijq/o0l5oNC6UYzqeuCvT9pVf1P0McNfDtaHBiA55BMa8SveFRRVjPK
r9//4DYnfHykiKv/iZ6QvVwwvibeKNP9O7Q09jHogEtzTVjm/2lBfryAUcChxTRI
b5t/GxDwr6yp15r+LObodE+Xp6VDrWq46Owa39Jonff8Rt+B0H/86F232sxXoOqE
3su8iXlB5W0P9mxMRxtQbeiMRgTumTFPDdxVaRL+yQF5HSUCcHVZAWnct84/Mu/L
i5j3SW3h62DL8Dv5KfLLJimAQPz1fIf8o3KOmFBGoegfnWUlqDW12R2EJG1WbNe4
uFH3m/jYqbg5FVopFuBjLR2ooacOMCevoHq3Camq91XMLq1pe5VTEwAMX+0Iz4lv
WU3drfbIX9kYZbuVi0oHQrd/OToHQULb169o/PhFmSl7m6FA2YtVRJ6xJN5U7uPt
We1Kh/xRU5myofFqVMddvH3q/dlCOBTJdQ1EY/Afi2CEBw/1eqskQd0czgWAzlko
4iaaFmTk6s+aN0L7BPgYRiyNlrcPPNaWY65NBosbM2UPk9sVhLQfPt26vuhlKdQW
Zpq6mOxCjSmm7u5eEQ3deOuvSbZqMskeNIDYys0EQzYUQ6yIxqQqncZeRxlR08E3
a24hXbtj+EOoQL8PCJwYQA==
`protect END_PROTECTED
