`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NQxktprXB7qZa/e5K8zrywwthRrszRtd7ASXcB16D3/PedvWQ59/20NcNEQvKqqk
AUdkMNGWMLvrCzQaeEgtguud0oyUJSeM6kfRrDZB318ZYnug54DgqG+XuGI9J4tf
6J0heSMuQJ6lWhvbnlQQV47YSgoqHPrdcNF2H3/hB+Y/2DF5enKRRzwYVsM0r/x1
YMpSMDCBd2acUz/lgk5kYjkkQak4k8FprwBn4SBorLYEwmD+KnTp2G2C8q9kfyJG
JxE90/TyWQFuqg/SVKsSXkAlhkAa3ywdVBH+wCCnpkuqNVCsGtdlzlq4LRy3PNib
+gJ7HbKLTi1qMBgrdEj+Ara/zmVlnu+9Uxz0kTF+koeZW8QdawjCccAvgRePa56A
E7P/CW9IV79Hgfc5XwPA0dEuk9jgfLFGXs+JyU1NYdzmtHTHOqXmQ5OQNY+DZkEs
UELXybvbNm8QxtL3sgZIaa6h6RdYqvKy8EaI2i/nRvy/ifi9GAWhHefzsvnT+UGX
Iu8lSovBzWd/cXAFBLOXhOUoWFiPwLturxF9LOp1oGGeccV2l2s04kE9KBqxuBOr
R0pMpR4b0fsdgKo26NQVB64VfXyYkhmN9NxXGrYT2RJgDC5YBZnc+2u6A6+JKVZ2
gZvnnECQAFE8OvZAZ85FlurWITPv2rJBSwdwfFb6FmE8P5OmSA49jYJ+yUOPQJcT
0g2ATCHRTD4VPbUqGWsE9sem7xwoVKxkD4c6l5C3kkcbsfvjUPxOrMgp9T0BNXjk
/mrifvG1vaJ1buUus2wmzi9l5pYlpH9jB7ggXeeayvFwXdas040qynrsNt8ilDdH
rzVh5+z+DouINIGnYxBl8Sga/OIkSH0k9t9InwMN67ciU2baS5Jisxhu594mQ/KV
h4NG6qUSXEkaewv4vs2B8sImS792I2bgYMEZHGk6WEuPPYpIa2V1UP5RDKqkhvxf
`protect END_PROTECTED
