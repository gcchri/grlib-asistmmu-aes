`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lsvBoKf5Cjq/GkojplVidp3TAPMCDrGHr3fFBcw4OAaNiN+HiGk5lQ3rFSle0oGV
PXqAcSCJv40HJ3pn+a2MTKV1YF70XW+i39YZ7j0tuGyJrM+yMyzXVVMvFCDP70zQ
Z3KyaQlmDUlK4ZkHXG8zaJ6Yyfa6rLawlyR569j+Udy2JYxY96emezYnUlspvy/n
MkC3KbMb+JDrpmbCEQ3MdCl5I+b4mKizzLVHEOFMpdC4xvyUW+gV5fPId7coxpg7
6OmN1ki+TxWdh27y4BQ6g4DldkPyI6tFogCPiHMuK1859nuTkWLy0D2fwZEFI0bv
PglSawXCQjdE3TpK7Hvy0L1MtM8BixObuO1MkGR0dOtM/giMK1n0y0rZcVWhHijf
VmSyMM46jgpAnMSFLDMrOfXo4rYhoNH3fyWToxQPm1Wp6z6GCITjkvjgobOjofRP
QXumns5Lrv5kiXrsnQI6OBhuRoivKrsZdB4pGmXd63qylQrhcAb7D0RGW+wcbVRh
1U3BnCgPV+ozl8URklTGr1AHYhWVIN7VhphtFjqnCgcZ3GyW6KWEruBZgMj/m2s2
FyahsS7jagGDjO0kQzZJUeyStrl7UiEqqf51APMwD/qsJQJ4PKCgd74YpfV+vKKP
Sg1Sm9mljeqf2ZHh9ZHyktKEoCO8pLwvDY1OQlS0jxGM+XeaErlDQrgeGwT1fbSM
gdMrmntQ8/uBJoGAlq2un2mKchtNWdfMlNnmZRfi/zv4KDPXhe1UVDop2mzi/q4a
CZPREpHLR8eFlzc8++QozvesLs7iNz8GhMfvNd4CNqMF2DkE/7MX1MYsPzVXMOn6
ZdA3b0yvWzooNROsBUVmmr96o+3WG4fbwE1SIrO3YMYW2k8CMJb+w7HDloGXXqFq
ytNhE782cxCgX4lPx1qravbMhmznWYi0IGZ12aVjJTNY8U2xpfcztOLFH8JOA7yh
HoW2hshKrfMKnD1Dwgi92bhQrCoFyxlo2ZDUcChoLKkK/SUtrO/fy8fhQ+Pi9bdb
fMxhpHkGo9B+SeJdDGZuCzr1sFFUxe90Yk2ZoIfX7Jr+Rp1Ez4ydzeALXppzGk0I
ri6Oh83U0ma+JoVXH+fJhLA7LZeI+F9wcvcTDaE6SWxDeJs9ztEd6MS+TcsHLdif
//Wiz/SBl7S4HVKOaJBrMcdxXaSpoJohEMz0vbKKMGlSQ80UR+XISAt2B0p/phB1
dxPd3JDK0REbTqtuSchOboa4NZkn0YsMnyDx4ty9KWjb8qXT9GjkIDJL1F5nhIoF
pozEBrCUiDIGtn1mgnrwCmiAAUYMqYaW0R4EyLMuo3sscet1Nl3UPtjWDa1nxtTD
dPruSnpRNFPWJEiUBjIA2+0YQBt+PkuKGORa0SJ8ayjS7bj/JqP5V8VEWUDylQjm
`protect END_PROTECTED
