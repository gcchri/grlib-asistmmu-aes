`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O+Seq2CxiYEup3rsvJfqfcEfksU7HpdzD6+apnktM8In/96d6m5dDjthZFkpomSb
IfdhtYZ3YhbzlpvqElduo9/5yb8F3CJFf07D1hW+risPOcysUlsSJIXWptjpUhqM
YnbmefwORkoG+DpsIVYTWuF0EmEzi+RriTZqhqX2CoI07Bx0zqIGbs1aRww2JGVe
MVP/NW+m8krjbWZO0X8rhfP1XGl6vw1aQ1VQZS1oNDFtZ6b+RIxEdQdoUhJ3xa3S
SVU/C/+CilRQWj/3iT5gr2U35wAEalYewL8sUHVnd0UjytEqY99s5uRwxQoohW38
HWGLQX2eFXYjzZtn7OxFWr0gC4cz/RLyWAyFT3FIkibAQJCEhLIJOdwHeBFTHKMz
BltC/h7RoMp5SRTc7Jl5vJy1IVtVNI98bSUGPRmwerurwbLxIUnIdpe5ua+ENbbO
G55PiIt8dn9R66azutT5JYLVn0AH/jKh0+qw8a7KLmpeBrIopIlb1UaNvX8CTrrC
KS81L2j/lkFTRd3hwSX0yMWYi3qE7gLty8U9ZxcBp75fxt4zjzHKH7EKO394r6n7
9UD1oQ7SK6+IQZzhpGYo+8xdLg8nSKiSdSSsA7hOLHk6GTJ0dKDViB+p1pBV8fNZ
dP/iQzZyWv5IyUY3HLAqhFYmTfr5aDe6Eg8ehUWV0K/i1yp9nEGlrdNjjx4B6EsI
`protect END_PROTECTED
