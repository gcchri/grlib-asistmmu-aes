`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IT9nOo3u1Q61K6zd3xOzQWuByQEvo99/vLQ1fa8gTEeIYEySG7yNAhyluzX50HZF
VK0wY1/MW9CeJzbcoowhrcnGK6jtCKDuUzRpbQIGqU6JVr9OzgST65TWIVDNYpWE
T1ZlBgV1h8PAzK+VkpHhy4+bCVjpJ9lvXhyW3JtPnMAqwqZ8VlRBnmIwCFu2JmqM
egGXvDBcteCl9eX5hcwNeA2Y93wlRUrDS8A5pps3imRbOo4mcLLz98Wo9zTiWNLa
jVAdazOulAzPxUsUvukIGkIbt8Dq4z2Tsj9LbdZOFTtpiHTw+dxC2ny0GXtgb5Zj
kQ4RqptvvaI8KjQqyjmoxuHlD8Y7rqDoMIE1Y1bIoen1AH9BAgnTMqM8pTdW5bGE
TgNOeFd6k9ket4jGntnXQcVogH6UG6i0/L6jrMeZ18aY6wQz1l2KNH2lX5KFQV7K
XR3rINWO0V79VGW6HeabSpCTa0lvAWSM68/KG7rG+Suu3Y737RcvJHJWmi9u0G8t
NJtr3C9QucK4HFofBCnwh9lfjgMV02lyzQZzKTWrI786LtcBpIMpdlAFSS8VVGvE
eF5pqXulOyP7gymIXCov2vMc9qdL82Bko7e4Zw8hP/uGYYIQwANe4Ru/Qb2qV2L2
ngH0U68vH088l71kJBkFhEZUsm0lYO7xeceFuLK249Ncl+ytUQFMJ7WFKVBWfEL1
wp0+xPwZTwxYdsWgZE4st41iCHIEprqxJpL6xaompOkEqZAEbR9mRoozqfoVGhDc
dkpm8ecfvm0c+x5TvsPdfCu4KxlM+JtI+IMrw2fxQwWWJCS/by9ukOgAn1QdKKPU
ZDIi/Y2GcbbKnwEJEZ0W+Zin/E2QInVIghNFYsr4iyc1ddjtHrqw3u3Ya5CyP+TV
bwbqx1/b1N+rWcrzki3wo9oLRzrW1hMRGUAyU//AVqcBgxlLeTfEmBtfe+wv+EQo
xsi3I0iLpvOBnSw03UokOxcnTK+lPPe9xHybVHWSE46msTa/FWHAs/yvVJqNjWa2
QEQlw88SuQlIFnIBM7XvSIZi9N/j5Y8Uqxd80U4Omsde9VhPd4Svu9iOiKvj/WrG
vd3dXhIdoQD0dWW1boHYthXX3G/3L5pUg7yGjIjE+f1Q7Jv+bP9K8p0y5quY5oeE
MHo4aYdHToo4laIjsKFckK5NZTJtBWK9+GDEje4qTARbU0NT6DDLxb05Wfee+gEL
uV+ivFdt7peecr8SYHpb2ePDY/q1sybAtvGnBveC+wq8Z9gR1ld359hzm1d8WT3l
qPeJO7I9CwN0SjVYt30/3OP5aDOlx/iSKCbPuBlFKERtvJ8WIAL1Lc8dFzGNDPO0
diZ8kD1+9fSieiRJu0tOFpsVVOI0ojYKCrEqxWyZ/wBURjJlPq+I77VaqeVuahbt
4penIi5iaQExMCp+7vOPDO2hCkH9h5mfv/lDadk2GA+UufxVwx/rfJuCyvl7a1nq
umhjAvsBWritblwyUT/rZwC1MfGSns8Y5vzTO9Gq6vXI68mmD/DSY/RyeHTqVYd8
4bpzcvA8zmJ7Io2sQdGa0UWUYXPHTUU5UaVrDBpwVuS5vOqOTvYvO5U2NOVYWcjw
KlrVE76GokzsJ6ncQKkkmiRa/s/IWs6iN4cZMCHZQydG9lGRZJn525gy8Go+5VTm
bdVbySL5u4Wdm++YevJiihISxFFOcTdA+8UX4MQddjYQ2W4yvRBsLjGQYAl8v6s3
c2qi/KyRga9KaJ/Jv3SJ3ZdZms20tmwW0DoqaE9HfQgCw0WJuTfOEGlWun5PreoC
aEmZJvkzZGXUKG7hzAyetep0bqljbT5wX5Pb/L1tL5b06sxWkmrwMfRQFelYiRZH
67XNv+optbfYVcDqsfscQ4tFs1ZidSj61uMeZcMapCUL7/Y+wuR0LiE/llMZixeh
ZXMV4FdN667nkv1rimnLEM/I1TWDJN9XSaMdmgGbcv2dbQ38pWcZa0Oodem8ePq3
t+mYpzo8fZecYZcHxauV8cJN60WxZ7eZflaue7aiVF5zoeu19NZJwNP69qjNeEkO
WPd7BG7PEK+oINu34ddMrmbu/YXqJ7oOi8qSk7t0fjeY3VdtSz6w66f51sz1ebM1
HIhfDfXL4qrl3HqdmU5oiVKAsFB2T22Xst5FSC6f0W40uIDgxZoUwIp0rWbe+ViE
xxzcXTz82+Qvtda7G4saqCObvmW88lgf5Eezr9LW5gdWIqkTFdC7N4mwBNLpbkXv
QFwlSa7BRoZpAph6D77L+pHcglTU3IQo3I3S6i2GdD4Dsob5ejkOs3E69IwevZXU
EOAYffWsXWHE2abIxxBDkDWpS80fDf0ILWv8QrrvONDDe0ONr3W4Z9Ol0aqOebl3
3bWLKZP1iPWxrVq89PmFYnglX8k/ylYIIT4QlYfuApudQ1q4rkdSvn2DcdHmTTGP
KeCZ9G92Y0OAN+SMpStWbCc2BsYGCqrBQqMFmHk9YX73KLDTUB4Hnb0RBk13dfA/
EPr7peeBzZN6DSF6c6Px48zcAyW30i+y2FVGltOVln/mehiXS+kStoviCGXejym7
zXAm7eOOykGc7UGt2Wn13lbHx1qy5dVMslKBm++cPttS0JZG+Lr9mqTDK0Oqixuy
YSgRY4rrqPF4DU3aghxJsWypAzBGHy36GLcbtY92MgI5eKhpiRsiNbfA+nD//7U3
OPpHN9eIBwCLJsDxp1Bd23p+ukJW8AGS/wZCLcQgcP0q58pg3dZ/Vib2z+IWAFkt
+GqvAR+9OFcmUhjUAWZmA6MuArxPvAiHPLvdm7pYdz4yYss/Y1LlFZJs5Ja3aDj5
7wPUbJQRjHWEkPaz0Ckgc1zEyWqNQGTIUH5skwnAIS7/6OyvbCshNkAQXFdo5o4t
37aisRKk02djZZ5BlbePArHADESShsrCe11wHYr2HTUZWpVS84LbfdH6TWZYDPZc
63dH9802guNXLR1UI4iJkVqG/AZ8wcxTvvyXdGZyPyEa5OuSjfDxIWLoocx5bshx
`protect END_PROTECTED
