`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S/pWdqSyNoH7E6+7b7772qi+OWhxknmJpzUuBfqQ5bO5gxEvmwcN5FeQwN1qbuFm
qPrfRHyXSFidcLhyKpl8fC6YXwzctsUsYENnIWK9vnjwTo6plXy2mJl3nTrK2O1w
w56APiQe5ROzVuNgGhtFUo9iHYjd8Yp+KxiNmwSwhKkNMYyrjzzw1LDns1DGeG/r
Yc2ADFZBnJOQ23wsSq0EUh1n8RJ0odcQu2BLpEGyd/rcjpDaQDP7uqAE6YHQY4Mm
GRz9OM9ejVKFS820pZ3EdZURIYrRu0/lP1EqfzK5szbKOXc3r08thm4sJjp1AeUu
0DcYHjhem3v2Tx7URmSlBbzk0DO1pcYdSpzbQHe5z+Czh8DC/bDeO/BZki6sLpaU
3KoCUW7hRrYWgBOdq4KehO4mK3qZ704s9ND8sJRh/pxjluywWcZoG7IqLLUjuAP3
L6fD/VJKD697Q84XloAOlSunzydOLqLKCMvm6vzxXOj0+mvAXM3EFHjjwg+ZfUCs
6ADAKAQbD7lHZKF3yF2hrc+c8nyCr2eoMKYkYyIoxwrFQMjA8ook67H5NWd/rKiZ
zW/noFDNCaAS6AfSFI2nFLAwUTYmzw9VaDp2FxJdDkA3cP6dyEuXtiof8ChcpKvY
RXfTNbEPsNh3M7yFDbQ3C1Mef6C950wSSlhUSDDZxz9q4sQxNwzlBg/c1k5rHRiW
y4qdl270AJw6j74ZHX60z/GWRzhlCI5CN1wlC8hGGYlzU2/tzHyr+HMO8zaWCsyI
ujaX5YT9I+qZFlyUR/Kfiid1Q0MNBEllaziQgNraPxQCl1M/DLsbIjcMlUVleeff
6POfcHSm2CYdms6BILajPez1Q+3D9Qixzgfzke0RCmqTpCHSsBKPRmJfU3uqnCm0
7I6m2vt6vr0lM6r28iu87JASqIA4A6K7EVAxQfeh9gBebCxoHam+/u6TTHWzKYEW
L/2JjI7phcOkIM69jCV5aCAK74XJ7MNmke82Tkf9uDkXh5P6lJbaCkAJUoZ0MHZx
jZP+p0neiyY8HYxLhKKap5rAhf69SyKr1Te+pzkCon95T01tR4QAMF09kbtxs8wv
EyCXb0lOTeZKzPXtsMXWc8kDhVkD4r7LF2wHR66indNMOxshieJMcQpqYNHcV1wV
XkXrShJ2wQHjaROaZfecp5FToo8ZSVZHTlyx+D7WkL5LzYfQSW3JL4/OSqX1IKj1
aCcQkuDTtjLjg5B04rSbAtzqeGgQAYCC/UwMn5G1LpadwUCHefV4FeFFiUHPEMTd
+8V0WoRZHYZYZFGiYIqqdyb2GnM4EZVBfAIhwnIgX7VkToa1LQhtm+CnbkWJgvl+
TGSXLme6JEz/69HkyNlPlH2DHjv0cOMisoLc3+jaIIFnb0Tiy+oLYCOefbtIoo9Y
a4jOK/tsdBHVTQ6Ygz9ogzwXq6BdjdJxD8UBmU7mknBPVJUorT07moh9VS3HlOB1
mEBJRh2B8hAcvK0k8isowliHGe5Jly5Wl7hOGPo253uiJk26U8D3Ys/MeqKHAZta
q9aRLyG+SCvbfFYqBfuy3jKPwvg3Cr5Vo/+p1ApAmwd/sowK5/q5gekDcUJuMx36
lsF3dNXzi4szqGOqaN1ZdorEsSaovoVMoNhPu6QPio8t8R8Rdvnwu5etB09VBf6S
u+aZRQqHddQJHKMGguW32TO1gQxqs0ryglF3aGNNeW/fu8sRtvohDh0gKQ60iRB8
0XLyH25cWeYUUBl0aym6k3hYVCrvFfm911okQ5FaiTjRfM1fP3drfB7BN/O0QZ3R
FzKoGJs2XtMYJVNxaPDXnVE9xTVqg1/mpnRpz5vaxrRkuOl5J7z+0L8ccxbMJ/Pj
07v9L2oTVnKTHkX1qRggVmbr8vemT5XaE2B5+Zqje70Vf/+VccGOkMUlx5N4nrmx
+szSjeFpjjxQHYY/PML5JriFSpiYpw6pSeg+kUiB/HzL7JIYViThd4ZMf/T42OLr
vK4WXn0UMWfp8v+zJpp4MpR3L0kY0XTwC9Bf4CZSqo+d7hIH+9mIvh2MhoRpgwDx
laF5EH0VrHzuqIwvqOe8ZtnBZGPSYVphY/23KQHXoPWbCA9X44kAahSZLRWyJSf1
T3sNTtEIr8tAadvz5zSc7BMOC0/NVd+SVZDayl8gX0GlLdyEbue90m9LiyUtDaSU
xVwi1ERc7bVhsQ6x5J9MbRDcgWatC9/aZGNR5lSUzusPk5+LfZllIQqbV3rkNi39
jaiIaCtVTo1HdCxzPhRweS1c3fwv6QIc3/TaMWZnEwNJk+/gqcg9N1DbfcK1g7iZ
HADPW6caL8qJT16VRNakydfLSbs+F41s7vk7GrHRU7m1v2C/64C6XG3xGYCzJdv6
zC13l7I9BTYq218DjrW0JljdDzFnRbw6n9+ekkV7D2+XbonbJxq766G2WpCL6/pL
/9qOug75QLx6mx3cS/lCAQGQtdDpPP7qeeceWVhQYPppYxbctdeKZCKdp5lfyC+p
yeJpsAbk7F2av/PPuP4u1Q0zFo3zAOBgLodPpoNF/U4wBc0lGrqQw4DU9Z6nqUCm
DQpHxVBp2gCrva9njwGrs/J/PRzAKl8uT93FeLaQ+5+2WC7cKTuNcd2jHEZexUf9
+YMy/0EentNaREPo6M1hFMp4Te+XVQFN6pGJqdBGqqE0U0coQG6u+sy8bLl/ZHsB
NHWWZLQlNnhg73u5MkyezhiWRtvsuKHbYLN4uMkNQjWSbGwOFzsPwAQ1LGksIbQ/
TbFHMKYth+OBf46nCxzdyxFFiAanV5iEbau7sJUPPd5nUlDrWSG9USsSsyNiBw9W
Ntf+FYG9d1PWL2biamRJggG4as0PjcmXKcrQm0APSJ8+0RmhLoigQUceJ8J9wCxv
UlivG1CBjoYqindQIQw6TNkowi7MIUuBBvaf0/pVMxJSqCmIU99CRx9sJTeh2u48
Y9BSrhPBcG1X3cIkk1qmny7CJ8ODQUT92il0SR6HyzwrDDB2NBL3ihwEll6WuB06
lm3zLkR8LD6FQwF70Imz2xCV8vjLaHiM4aEvQGIU4R4iE44IEcTp6vAHdCr5CU8y
MjGI2/WgyEK+WvvjBuzLkjhuwcnxM8U5hbnSVlHY61FwLgBYrE2cw3/Tghwlg0+W
WwYLzu1isZoNoRK4OXRbmixKOPrqR3lZL8QQXOF/wbIxKzdD0toq4+rAQ73OR+Im
yZpXyi21AqnYdDs/YT+XWWqKL95sI8pZMALYouJZWJYFoyCQiawrQ6RS+HXZsK2U
vllMCntRoQD0o9SOtyMJBVLZsIADpLFXHuSdlLfUU+dhcD9PUfmyEstCGKUt9/du
oZpdtP+SKsP+9T87B4AbFFTAH4zqsHLIGB/V7yxlbFkGPjgzrzydZg9O+zFqbsZF
7VPm0Y+/vzgVda4HpQCLkcv5eETbOa3qVSwUdt4U+Uou2tUrK9IOxqMPPDEAxqqi
+fcrz9Wy/cg+VfcH0smiUC30TVajdi76fNEtMF9UMaB6Dym+D7COOUU5VOcP4/wI
UtKjjr4RNQ/zNAq5lxlK9sT8So5M9XBv2PtAT49OJRKG5gdIX3U84HSHS7qpR/7i
NCa/p7fEjgKz0qhXMHtMqUKeQ9Bp1QdYzWaheiC3RYP8vFu7jWrMqONtq8tlY+lH
YytSgjrzg9CcWs6ZL75wLwDmd8dZvjImiTBgmAbv0wbwpb+eYLCeBINl3fYvUi2x
U6sifjYWNVedtzRG6tqLsL4uaxit1f6qDgfJeqLWkFQAUP7n8QKLvh/ArCeAokpv
tBlw81ZwwqHOmexGGo0orwIt5cKghCEl20WRv2+xyqEMxTK3TwZQc9MSy58+fYVm
pjh+Ig4cX6YEpBYozxYyXdt/vIs0CfKFt0Tka7Rd5m5/nZ8euQhgraSALnBXn5I9
6yQ6gOqvW/IWybEdpMe9e39+KWex1YtRNrPecb/UXr6RCK/m95e8sBhVhEt0+x6A
DvPLBHyopDI7j8/O0BVobgb/ZUgiJQrtQALoklZvt431dEJOlACiLO1lbeAzp+MY
j1G6CObHiwX3V8EQAJq/YPSLeAOTZwi+qwuPA3kaGace4OocG6oiUe9YC2TC5qrV
tex0yw+HL2TxDruneVHwV4VPuD44mOx+gz0yvwBlQchwGyaET9MmN35z8TSS3tIn
xUp0BxA9gWkzIKxd37JMygjq8douL4V3+eEwcJEhfWdDuiD8Fy6iRAeQySankdxg
+zjOEqtPSbFiSXGciXnBUu3lEr0CnQZzzo1cX1d3U5tXWItgZDFUOImSwns2A0Px
n5bF4XsPhRLEYxupJKp9ids2KLFn8DzqCXsGZsGy0HdlelUsKdu3SPR2jdYVr5xP
I6abIlXwUH0Vrh75BlF2tlQkul7xsF/JMxi1Ew6UKDxApr0jXdYrpYybD0a1sZix
GwAyTsBSSTAIfI1LEl1ODolw4WstyZMFMuOT0O35jKVkgNlaTKc+2vjMytTJCrSY
XgzO3vE7SRdZCBtF9o3JVTVUZsad9YpMRuK3zyZpaTxqXF18OsrnzCsD4Q1QLuZq
/y4aum8TzYEthl2hLiG/rcs9sMqgilL2DB01OH0kwTpFxBimvJ9A6FM1eZ0bJY7X
2kx4OW75vR9VNnrb09qJbeUCdUsVPWicKjd+NdMMeTBIUrYQ1FWhFx/RRZJN+3fv
i5ydKNwvheUO9l23lZdgYxuE8RWjOMvChdH+iUDsnI0BWQfZW7aZXkbAoIAyBF4/
1PGFF00wi9EZzqlC1kxt6GabsNR744Vu8EWDRYR2u86+7QIdB6W8bVp8KmcUBxs9
o/iA554zCM+LBJ3MHj8bwwqUjCqIQ+2x+AsIkqKW3P2qrRYau6ulkoTpx9tsEZRV
CIwNFZYvLUba/nZVPnsBD99Bwaau+c35KKOr+/wkmeP6L8hka4LH31/saHbGcGDx
KW16m3dQapMGAafOK7SoMdA+4WSzC6hzoiM56CMs3Ehh0OxLaBVWOEBn5iI4tfd/
CCC4mMYQMWRt5CbwgNtL6zA+sy8ksZorJarVZPn53W/LEX0597rvCpUYgNvwQq6q
rHS4dP8QL9iQO5cE1M/gr2kdzFvsrdYZ1lASgHCkpWZayateLkQzHCxwPBgR70wx
mUXBJ12w5Pc3wkLXPdv2+uS/lB0ZwhK4/VIqdrJ4q5t/ABISxDJwsl+q+FGB2ALG
V80oQ7rFfFAQIZVy2A4Qs72+Jjpvk4tkM1/kt8QdBlgfE6VAOBJYzkgXtbNk+0d0
jfSo0k42CYxTyV4a0VA5i1UTxPq4BJIcKWi3djEgrCIIQ84PiizhCShYHQcS28L4
tduxoeafufoR5BfPL0SOcwOx9NJNSHf3opQRb0THgJ1i1boAFQ451OEQFu5nZzh9
BZo0lPsfN5XEsCF51lMslgkEzbPlLYFvYvPZ6wdAsAYVJIRUc97I2HW5Y8dX9pAU
AZVT6I2uV3d+ldn1ejM9oNLhSH2pvWZX6/9F8v2b1ymLKj3usWG6a4fZZh5SaogO
upOHspoAtvr4hgcJvolU6hoINLrO+JHB9xMZJ97Ir9kcd66tZaGghyCkXvO/O8Us
MmYBfc8lTsdaVgdWWPGx31UcTMtOTGB6uevhEVtS8Bd/niZDj5MSryS1oboy8z/Y
uXeJg1Wni6UWX0RRBEgugjqc7KAPdMy7x+x+nXEg7ji7W9Sc8DXc8cdZjuTFIDiM
jYyZ9Jk/RRCD7pWfBrz2dLrWRoy1hMaIgY7u3NO8IWSqLHdfenjBoDrqioSmRTSU
vJ0zn5aTS/LS/veDuTOo53ZPTyX0wAzHZJQzdMBkKudx8QRsnXPR2LyPwgg6uKch
GsKddOT9WkkCxeTdj9PSpfKy8ZcbwZS3qKTjcfsz64VmVjNQ/ifOLaFIMyGyyq17
ijrD/6eqzE8dvp2HPOdRXgakqMqhh2sZVHjf8MMeKq9lXch9jCJrdkD9yXC/MOOX
w0yaKIk8JBSW4f5GwnIcJa7+LUGpjt3hJpdXTjCfA+AODgllhqAoaQziEcuIJKvz
uhybmsIsIl7M/PIcYhWW18KaLS0659gQV96G4bE410KymHKnzLfkhTMtLODllAz5
5Av2C+TuMjASasWGGQcowoE3VuLwH0DuHnwwRMD3/BAvXtPaMxSepiCO6STggru/
QdWF0IrcIwIGsujq02jPlN5Ma7SkRGYrYIhUnJ3xabrqEfxT63UpHtrTvygWpctf
w52pwppO3CgXWJFTYKOi4sXGqLDrXj9/hH1aSx1I8Bste2f+IKK7uLZ4SihcrW2G
UiotiG3MNonM+oLeqEIQzq4gcJkrY2BtjBh8TciYzi3jvHSPM4Vo846tUJZ0assn
YVkp/7coYYZI2Qm1ntzs7Q+RiOfL0gl6sKCuG1LB0LNyy93wGhGAETTDROF3sNi4
OYgbCLlub4H4o4oLdLCJpbH8eZRJ4uTXs7aEPCrbKtF/BSiUyizUjVmWm8OFt5Oe
XOtjRIi+5ifo85MMXGC9G+yo5JDioZRSfcI44jtoSlBAiH6AsQj74nmrDpzfKtwp
KNskk41LQzBlo0SAqAZD316EsZXSD3F03JHiQ1MOXvqmC8HqTvvCi8jYLYi3y5Ob
/F0jZ6MALhHhP1/d79Vfm8mo10tmiC1siYBZsgMe+LXBNWaQIhNotY0IHlRQuurD
xLOmNsby20Uf+xnr1BxFnlWfxS9+5ugKgCs/u1mJbQNW6WFpFro4qC3n7c80RZT+
H/Qmq6hCfnwUC5l0p+aohPZjFqmDIsPxQjCnfGidLtfltxb+5ZpRPc96XZdl8+/V
n1HU0ynEmclfmn/o9p5NVOwAXxE1sAD2uPApDKa6mYudHLwwT3rf2sbkRERjEzwX
LyxnHTLYCoNzFvk7wa4xu8pTdggCBkjeS2MHMiTBQWDkfVnYOSN75SknsqhOQSFD
x88JfSjy4xwT2fvcOsJRKJ6286Sk+CdecmGdH2gkUy8gLHlB5FP6+BuObhHjEP0N
PNNvzrN8r+8KXyMZsCHD2BOUHa8AV31M33WnG+QIG5Y4PEP9y5z6zPm1KUgfjVb9
3CHYNqeiJiFBQsySXXyD/JR1CXWZRS6krHv/LtD9RXB8uOEO0DlWJRHZ9fdONTSj
tCcGlcVeG5nOVFsM5lgsc8ip+leTFOODKR+bPVf23IXXkhnvsYicZtUmMJGx48gu
EaVGkW4I7O5zPObzHsokakbOfDEGQ/761308FvZjoZLbLgyUq8zip/j6mosqfIi3
puGFjSo6Ra9fQwTEc5kd3k0q9T9tqmUGUTWqZkzbw+Itqniz4VGD7iwe1jjekmj4
ps/PjgIZBIRiLL8MqqUoulGMxb1n64Fv7Uy0bhm37oOQ69h8v1gYJhsGnnRDE2LH
w7/zEBRDowgb8btNXwAE/eG/yCJ5Po0sov0Ak/Gm1yV1m3s/gEBcpOX4XjwXZs6i
8pSpKTabzHhU1FSNZRqGQiHzo9vHkyZ4KcJEqDMKFKysb6UbL+TbQ7xBhBoCHR1w
xg/Tw/n+xuEZ46eVmIaK4WRDEGxrwwyk/dKOsbYdLZRaiYHDwvLHAXQEIbCrWwT7
YmCnmLdTAl8JsNXwj1RWwXqd78o1bS/mxk7png/R2S+LHkpNbM+jFlFfSKhPXgHM
jgSiOxB4RKecp7KHfbjtSrOUoC/5fKBk1MXlJR0FuF3SKweBAKclredE7maXbPfV
H/HgYHMiDHpxPz2UPYKmxz7PNpLfJqeGQKZaG2b5lOfcPsE9KkYMpXFGjFvd+uXO
yZMdGcrP9SbQCqiajcdZwqBF5tP3pNYtm6l2Vb9mZeZlsLN3LUeYNj51t11YydQD
VjcRfQlDckB14JuQGOG+iwbFmrTmfFkcIS04hn9Qi0UrE8E0JXAirHGf8kjvJf2/
ao17+E3P+5hrzAxAH8/zFW778eb6kt7dmvQC4VK3ksTkwPjingbXjIam1ydCpqbi
naWZdbiOvx6PP9Qz2Y66AR1HkY6igHBy16ed0wLFz5gchJzSMqX1bPeIVChFgZfy
YHddTdWxO1swhdSyl9TdLEqlaTiGVk6dw0XSUNl774yk8COwqdlIixDeRvY08MDH
GwQS93XtqumWy7+dCcLW40+GAz84wGTbstaEp2X5K4slsFIAPTukTUujvAREZKW7
PYH7RKribisZj2z1TC/Ha3lriz4r1ELUEDLShkjHqQ4ZNw2NWikbpFwQd+M/IeTM
ACoQBZj98Hn4IUr0TxLp+Y6cJeMhyj7Jb/2j3uGSm2wcYpA3DE1Neaxc9d2fKNyp
Z5AjycHGOfum5taEfl84pQ7VRvSRa010ZjHtM2pYOpnm4dkaB8+MWk/gIu1jMr9D
DjI1tJwY96iJupmvGZ/sQbWBYYU7lObPcHrOnB8DdbDHqke/WtB59Xf4q0GwXHMn
aBAIsfTdH2TYM8dNCT89jSAY4hbDQPY6s0okoOVFAkMDNyedAHg9lyCtp+2OiKyA
ochu4D5keqhvlajQMT3+y3R5MTf/drVrL1rtfiXF8p1fMY3RXf+co+qFjUe5rnfu
YuwCaIpwQIEkl6jG6Etp507KZVRjxSAb0nFeF48HxRgIzlnXY+gKudBvA0VzfwGs
NYkkZJpABu6wDFkZ7mHloKaeHqWig8W4bfK5VcugZcD27Nh9yV1opVKvAu4us8Nn
KjyfrQoVXYf3zOEOWG93o8wlsMGwQgkP134u/zL9+raIqbI1W/2BgJVlI/1NS+RL
4EuQdz064nPGtZ5EZHPgrJyZhDjt1Y1ngJA8vn0suPS80/HvVED2YsA7S/WB1+Ct
kdn/5C1mp6DNz2a9/JQJGhgohQQza0jskvoafJXbtfHAqCg0YAy+/0+WrdkJXYno
YcVNwtjMk9VplPym0tNZGaCCAzn6xTUiL9UNcCAcPg7BWO6/FFbhf9U7cX9PY3ck
dW6mknhWvLKhiI60Lx2ltJKgsQy5/Ta2umNi7ue3RcOYxetZLWktyvf6CV+Po9Vj
bbkZfjOViLu7ZyjHeuMuI8Ak+EwsB5wc785nuXqaRiW5qw1HE1kfGYDIVUNTYazb
8TA51LjNJ9v4MEgI9pPcAXYdwrF+ISrnMYHcrzOiOiEE+oE18aJLpGRYUq30Y1T6
MTXk+pPxixgziIP58fm/h2nlIyvIOkqb3Gycv9iYm2QvH/1FvRd/XQZpCWXb/GUK
Eey1tQOlE3j9o8snjRks1GyR62kssqyiO4Hz/iwCSMcRDZAjS0awiMTUFUlxyqgW
K21DKgDo+TrM3/FM94V6zWY7oZ6ghHni4yg4H7zh20KO7/z5hRxbZGBDTriDxSA5
Xdna6SUeBZgTGGq1g5l1rO4Y1P1ZQUCICaQAV5gnerE6YWWNRFdGBwr6zHNr1gAp
kJ4YD6a/TltFY8j6vcHz8uUX4Ymvq7F+HKL7ovBZ7RHZS+aDGjyNUzWjwEZrtsVv
wyGy4+9OntPNuRqkNx+diFIZaHLzhhOffCdLStaPalgCEC7vwNKp7YRrdeiDsYtX
CumV0TwVopZDsMoJ6tGET3tJi/mme86A/WYgVvXC9z0oCU4qcKIt5mU1VtRkLvie
78WIzD87/QateLHtx5iIUgeQDaySau/X7IL228Qb64rSRQevKX2itnYdKofjBsJb
jetRYMSBeUQ831rWEX9Kx9uUFrKoVzmkapXJatbIKFXVyAqYyJt167fmMY2UOUWq
1nqYDFzc2n4m5QFdXZjYVIMNp3R1jRgFeznRgC9fVPhfdHIFZ9GgW7atBnPrPRuM
QEUEVLOwzQJue4Yhun7MmrfSUlScbN1eoA9CcKKdQJKV41K0ykVXzPchQqFeHiDn
SzJkaBy05imlHawseoLqsEEs2WrFxfYFHbkwUBpDHUjiLrHi1gNSUaol/uVfEpSR
xAp9FwfuIuk4TQtg1Q0I9XrsoNovxGXGNl9smUEK/kb7IUIYPXtaE7OzFjUVCD6N
uBU0Gjc77hYJDjEQW4wB4tYYtas7ouztjYaUL0OEPyfAPwubel7nkws/IhiQvbno
IY3tb7WYmYTUiGdGxKetWfx8ZpWepogYwXNZZKEBlcZEhaBC7IuUsGMc2dy45IBN
SRJppSKGFJOQrMCRvDIu3DWLEeCPCvvMG5H7RXKihqc+vraPDRjaYnxI3oMEgXEz
hvcQe8N/0jS6XhfFKWW1FDntkm65/wlxSXEEZkIFd8UGrQJK1Yr9zz8v391d6aIN
armKXiUDm0/2cSPd3M4EaDM14m08C2y7vdwFtdFtnDZutTL42o9yD6OnuGIdEab2
ffiJSk7aM0xXQ8v9/evFJltmDrPUyYEkYKH2TEX47aUHqA6oTufUyK4m/EYEK+99
t8WMTH76Fhv5cVkHJBb+KpMe3BWvhMGx7UDHnmPIZzfF/vUmxemXxrDkgINTUClB
kkuv+FDhxlH+Zxg1y3n7TqTV/agGDDOU7TqpyAJwmufDTrcDml5z8Khe7dMe+HpJ
qB8FEhbF/v8q1WnCTXFRn7LaHLR1TIA/uLacBxAGkOGvchw7276tj6w2xp8JEZQ+
W9ZrME7zZ90xTn8/UJ+ja4SVTZvMRxEAsB+RoQvKchso559rwTofDchv20Zn7JpU
zbpIWzpEz9PsxBUh7cuJBzL2XxWQf3TwxmmTWSKdRwxpYXIaiUUsiuER2HFDeoiz
WRG0Kf1WkDhCskToheY1LmrIo5W4S+JMwIb00xNEclYoOiTGHScV39H2VohESBDs
OYmAnvHH6YWcCiCBneCPXV5bAYhRxytQJtTP15sg5YFXBVeweDn4xS8MWPDcFemQ
EfWLYEIwHH0aVw8o9B6nELtR9Cqsym/dmzGcBnDrOpp7ox1xflnYjBtyVSyI2tSK
0gjKIbR+nRBdQH5iM+vP+QmAxsXsKZVhFBGY+8S3uvugY6J3FFcH1aK9wVo7dr2z
UIb6cs0tMtJTxfYUwnhvO25J8fHB7sEZ6mPYszpD61Cg77uFQaWwu/yKFlMuh+m3
TzA9/Ivbols72qkMGadmQGghpjB0Kdcdki1oyFeDL9RwWB6OxnpfZ0jfGGrPWJdn
fMjMFj6S71gjeW27rR9XjsHtteW+zdGe3tcs9JeK5WkNP4hyxe1VYa4koVjJWw2f
IhyR7Omq+4ybjdzbluEIIdalHglVScDWA05bcwY5RcXvELa3V6s+4bwbZqt665MX
klJmGdwJyxwaQRZpyyeuESmdJiiXvpguMh5hxuhpcdm8FurV86HqR3thhWc5uN7R
/VoU8xL12kJTyc9y8kZV2Q2DM0YljXp59jejKWBGHflUPCy+1YnJQADf/NaHv0zR
9IbGI/1UjCE0IG4Cw2JL/WaaxZQHXu6Lp7aEU4yKpEnqGNGOcdCUdjrbGcqudUQA
nf/THB24jDQZyLxfdj10FV3KI6XucZOiE97JGD25rjSF41aN7xw+tT5jKP7S+Oi+
rqapp4Yj6kHRK44q8o6B3O8jQJqWY+RhfnVm2PImmVaZ7kZhpd3nr8bwC0AmMv9l
j6qiP8z5p4oESmaq7P3HIG0qxKROmexEvewd41kQSyRm6giFnJlupBTbaqIegjZD
QQJhD6bqfZP9fv4KYtqpY0HEDHuEWyUt9xJq6KD56fotmmoFI3sdjbp2uty8jAqU
RYrYTYdVSJbrqN301GGGNWQLeOiIbLJ3Z/nOj+8BDCJCNTVG/P1PgdsajuyakK23
M+MkeZH4W5cIJtarPqbaN3GJmo+zLWzANAJMhuTnOmbvI2Iemz+BhCLZuRadOP8s
k/XcjmcK0slg0rCQ5Tb957eQ/mp7dIyR2Sj7Mmuqims+Sk2prfj8iDQAlgN9q6pm
Gv1AGpdg0w7BZ/cCLWWMpmzvncg6vIzO5F4dTDP/QLgxgNFavAf8kU8toGJEojM3
ZCEfO3QvZ1RS82sbnGJVBktsSg1RLoFc72UYX6PWuLDOTLkjSy60cBJTZoRupXON
NjiuRGWvRDucP+xoSxjqTLE+cUpFboWxyQbLGnUA03MeH982QBLLX9M/R75EQJU0
m5z0jJODCB2/QNltqjc1vsNHSG75durx6kOzonAbvSB/aoczNUrY8U01B3oxa21/
rY0EpVXrTgQbuuNhIGJ54xepl6iLqvbNbPbkMSoZ81bGkxMh0R4U4dRE0gmBC9dM
gIlvAHHgKjv+GAn30Zkfcxwtc7TtnFPdyoB8kuFcxXB8fzAg9GdTgDgP53sT3h5o
0xQKmRlqds5Mz4js36wFfDG3mwuqkPYtdmF/v7ivMkGUVg98/3+5j7Pvz10ib/TS
Bc4XvC8G+Q4H+zxIKjFE1JtOPOwp1ZjeZ76CMTmJ8YAsTEi6I1zk97huCIi3bPut
YJM4gg2/CTGZ5OneBz/+m9parCFGDKWAP+6EUieQAEa082BFwCDj1VP7y7k2/x0W
DNqMDpqbyANwuBQndl9szUS0cL6wDAdSaR5qu4a8uMKVHE0WS8JtF933IV2k0gvS
KlpprAkcnMX9aIYNd0VrXgDprEZhcigmcUb+sBltlL5I+cIjcdCsYVikqYsmOzhG
AhB4a3fE1M5+hhbYI8Dxe9WCW5+s3y60JibFeIbWI3KA1sWlvPua1sWybjgkUE1X
erCERqdCMbPu9l9h3V+zsfMn4rCoW5g0NM17ko4+ay9nJ7LsUstvk6UHvIz3Lfgx
ElWaqVmkLZ7R65XNWxvpUdwoTt1SoBSdOfA56Z3k/EFFMp3WNcGVr97MvimfaC9w
E8ogCZd+f6L8v9O9c8qQM3Cq3doIEv8H7ruuz6tLSINAhJZTzTKpfYhxyIjbzlX7
vFtWlm3lDGzahinriNq11aiLz6XMtI0lFT7E17pToiY4fcWBeaObODMB3/7EEyU+
YQtkkG3QOdtuwRjpV3k48IcwWfSmrjEnb2LSO1wxvK8oWL5E2zl762yVJrzgwFBe
CZpU4thm3i3hLHLELwT5fIO5J80pvwcLqQLuoPHsbnBoRolYMI+Aw7lH8Z9nbsQ7
QrZGV72cVzx5AcyrKzh0qw3SAzoo0WBCJiDrXLBbjrm+Q2hjgi68koLWGBh0VfLS
HLT0yMt3pfUSYew80p+SHOzjIAALIG5PgMi6Xi5PZ0uBXpnsNzMkInwb7G7V83iq
KIRDRpm/srXNx/Tb0J3ffQZG4K67lTjgh7L72Ta52jOOUCqi6aVSGr47zjsirSEG
29Xb5qJSBR+YG1L3WSQYWWM0W+JyBQiJF4skjFgePWR4rm5GqABUEsVth0L5w+Y3
X5KEOA9FVR6Q2Db/uBjCPjECzPMuhW4SRxGsNTxU/hlzn2g1eAaA1rq6EkX/a3mO
8nkptOSAvd/jiv0H1wd7OJQmwURJZtIIehvw+hG1XjjjdNZbBTqNWK9r47fh6H/h
kAw6PHi6trX66nskqlHCh6DP87iAp3durwtwoaYEg4y4w5xnN5BhY/wSiq2jhM48
J6aaG/WZHk+SAkq1fRr1t9GpxdZS18xZ2ryjEVR3+SUJfPDpfzhl0u2Et+sw2Xws
9SBD7jKquz+1f6nDnt5U2w2lj7XLzcrIhal4EFKLqhnhNm1aw8BFgFd8q1GUu5FC
pCXLS1gALk0KYhxkNonRA41joyAtDo9fbdnCu+5sdDyL/mUlqJNVBq3qCcQ7pez3
v62jlLbpthd0AA+hzHfAqCYOzGeU8/c+gaykQxn46ZyuVXwWrBeYhPMWPCM8/sDG
ZIkHqzt+lfskM7xUD+9ukzxzG/TjvWJydItKRjP7ZRaKFWSXL9o6z+pDQPnfEB0s
7SE2lXtiw4y4Oa/V9A9+jr/yqGcnNGx6duSMuwhhbewM8vx3jZn7iPLCRY6i2YXp
nhNY3HlHqmsudWlefjwo/1uRQetDe30SbjpHG6PjnEu9oWRxsIZrCK3X/eyKY5BM
kfTmi4Dl4DeLEbhmO9CF5idHOLM2PtmqxuOFwRDb46B+d5IbexefnJ/EPuiY3M43
pvV/I/939rawwZfb7YYPG1jBGFz/jXLEcfmEPkrIBEUmXH+SRN+Qk1A8MTfnlFaF
1g4TVtbuyylmLfR+V4t6wtiiScxPg724LwqDJzp4sZIp27cPcAHSLUmrJiezY+N1
g3X2a7ws0ylYi17jC7iwTA0K18xV1anxWMEvPfAIGMx9BGm7g/HZH/k1euToiKbj
kjjeVceMvLkg7GcwtOUC0BVgQ22G+JezHi7z0/1YSdCdAwWtSzVP8vjx8TaRVOGD
0OiUDxiYa5LJt+rDukdKEaKLN7Ht415FOWELh5v5SK7R+b92Qc1NU5fi2MbEb4Gx
XHQuHcyR0HqxXtruVKceV9hWeBvn8VZQTCF324wPEc9qvk3s58EIsv53Y/A5RtFA
pb5H6aGUVjkJQpKCv3tW305mdwd87IZaIZs2gMSJLbnWxbP3VjwcCwChIRx5lIvU
yGHcdtaHbrdpzFbquhow+DcOYIgBVC+FUvSPTisy7ZsmSyhg36nygEyGUz4mGcVk
aqdE9KIldj/SqadZlFpzTBJO4pkEvKbN/Rs+AlL55z7SWlz+SnolBXuQ9P/7WGsv
uwmEGKLiJvz3Bbqo2XeI6kL3JkxgsiPxVAAGxppDTVc1M6ODKmrEWsdxiQvMidnD
Cwq/oHqGJzxXDXfgzI2HJ7J8L1wIcqd3Y+OODY+Hdk5B182QX6MjtXw8t1rRKbbc
LKcIU6xcU5Sp2ybJxr/x/GY4/x4vV4RRL8FbxMRvUvTurPsofWI7ywc0CPbHABqM
4QUJmiRlrjK1ZBJU1hrwwMAqZ/SMOJqhNQSK8yfGJoa78Lvim/iZoqDDB+jBMaKj
pLGh4IN7jFEoEVcsIptTzD1UbSf9SjdPGdP+qA4IMfMAgOrgByNHkBrvALtIvjFB
U0oEJ+DUtt5U+CvcaSrD8FjRQPipSpITfglhWBJaaHlc5VIhfZPegFfPe4zavJ1c
kap+P27+9mm8jHxoMbEc4SH68Fwi8Xz2V7WBjeIFiGteJE5Iy+9TsCJiQ/PcsOvj
vGxq2FN0O7CaFnfxlg/BYMhk4ETr9CsUivEGb6cq3xC/K8eepNPzDj3tkPD31JV3
GwCeTrcyNRPOwVopzeD21U+VlsLBd6u85RV/z1FaVbm6S5XNrhmNojE0UfGuXUq6
lDzOaCdS4LxAxu3VPbMeoTJBikQ+uAsEXTrXCMXZFR0DRa8GSnNC9xsWH+a5un06
mMEawtPZ9bvdNY8A9pFsDBbb+CjmuEOxE3RxAeE+iSMXS0rSgvPA2DW8JYn93KRx
GShP65HsvPYhTevFCyIGVDnutRhhaUasq5MqG7WK490PjxgLUWCksDfV2j4axQwx
+eAVibWIig9SYeIt6WYjFMUfGSxDihrNGJK5dQrcZyG3OZ7A1XyGUTNV3tFbHHBs
2IRbjxxa4ARVkDy2ny8TrrLB5MnbWYB6tqY87mPJmxl+45bl9wHasUQV+P4BJjAM
Hki/3xZ962FeAvlGFugdHKmKU+5Q5rIQAbx2U+eVDjoGWX3KWokyYydg+CV0l6vr
D2AAMTTSOK/T9CpXZYKbIvJ0T5eI5DiLkof7r4/gl9F3jBKWW0/ioWUq+41mOVDH
yXGRTpvvAeHs1b2hZyXYxefzsJOFjoMk2RpsJMQMWwnDsHXUvEEBQdovObftrGOy
a0SCesTnBwBEhgS62K2LAtokI1zw+w/qa3Cpy7uFzIsFJ6QvjQby7OnlsByi57JJ
j2Pkr5zdl3BThCiL4H79dPDPRaXEUEl7POIgJK0+vwavNV3uv0YhbMIresEumCAJ
WN2PiwNz5NnMGMxi8T3mWfQoupT5fWdGLz55YV8aUs8j9cyciW9qc+wJRc1A1hB7
tXW32vKqLXJkqEH3sCVYGKvPev7OACZL/un5xQJdj5h+0ivICLtyXkNl8mdGwbqx
6Axpzq4Qc40hHu2FqkFCROkTPLZAIc+uraqBvm3QyULl1luzppvvlBLtIH0UbtCE
VDdOKSaxwYV1OQxKM8yb1f4gu4lS3XLp1+u37S9d0oF7ytmKnl+XhukthEU+5qYh
YFSkVK9sxdUDHTj7l0Ui4pASRPuLymYiu/bS+KPcOy1/U52XDz3poCr6kMdq8KFO
Q0LUiratwELv8JEKwx8IZhVrm/v6zOejtKDGnFVBrg4u5COqLA+/i1xzJAvv2kMa
uzo/qU32sAKGLo9FIeG89Zr93hl/YuI1/MUXBc6K9W3oNAnZzj/q6dZ+xzDmcOB8
BOsdXChR7z05uGHj0/aM5ro0EWxVtTiE0U7/aExevZ4fSRSQIiGbRWB9YdiqINzq
oGW2ek83jhgwtgcEKOu0MKJUfzZWvfa/bChuglzxkSawbLl8Lj5wNevbnmIBgxJr
k7XVUFMsshOuCjP8SpLbuX+rgEspINHK64QFap5W4Ey4kagB00jtur6KovRvMbsi
1oWpSYn838u7gVaBHv4DVPoNDCbHjLN05UcIh43I9PDkYmZ2XDCHf2l+xZ+1KTPu
NcG9Bedb0dnKQLapZwj9JannkcfgJac94ElfLCQoxw5rNkKXoADJdAgG+dL5wu34
z7Z4HvL8Sw4SjbjMyQUNQ6E19U4pYHPHo69///J84W9U4H0uFECFZ5cMysLGQvmm
a1jIkTSAHVecwDn6NGGgxhQfPFMKZo4THD8moygCI3xueQr6MAtBT2B4kXN3szKP
7l8wKZ0oMbF4Z6C675ZvUeBMqaEnnuvzryVn57jkwPUGLzzKhKGL+WXjhb6uBoA1
cv/gppI7ob5sQvG8/aLR4WtaVFO4nR9b9LfFUE/MS5SnfU/dk4SRIeOTkBIZJDTN
QVTkEQqK95Sig5ezzsgcdPZvZ7Yl21T3cXocVDqjSbojW9nCUqC7IlB/b67bNa3C
cD3/z80Ft7Gxf86ohL6YolQhJtG47FhusoW6R/tmi0oqP8KhI2jfOifD4y8rlIRc
nTWOing5rOTVUosM5XTg2ptPxZLcO9PXKvMQJdsRk/Dar9l+QdQ90Xn1Kl+78//r
CJ0oEqBQCCYKksWS2lRs0EXKT+FWie/FIWRLcG66wO3Wj1RXPmlEH10jfFEGV0Gv
uMYuloziuN2dybAPBzisZhSViMuFWeheM02ileCtLulKujJahbDydqlKKjCBndRh
AYTqYpCsUmrWajf8HXPWJP1KHxf+I3W9DK+n4vnrO1vorE6lt+SBjZA5/UcIsEF0
3vq+lzS0eeftuMKku6sxx7EzI3IMZ76IUSKGHwUk26hVXfq+kk9ldkCRCcSUMXRu
sBo8Mtu9vWM22HdzGaOiTHa9WWpAWo20YymCDzW4j+aYqhE0pVUJdqVVp1J7ZFkg
cEAA1gI57BVW7i74mfolsiiidHafet+7zsXTzpBR6EqF6cR2VWuZPYA6ttQo1jqz
FSav3t67Sa0BtTi0ZPRtB5dRCXU2YBaxAUJWTNUlkEsFHscifYJovZrpmKULr9Oh
BaZiEr95S9UXreO1zQvPt1ntSJVIVIpIKW3mCEScLWPba2qgq2pHH2ZP0lL26rix
10WpaDH7KUDY3L3z1DMPXQ6il8Ovs0rPH/Y+dq/C4WPnpm5Enz0tJfCce3bijuFh
GSS/NJz9mVNqIltjKIX11/LeIeXRl4H2XW00X70QvEEtDqRT85oeA3VSV4GPtQKX
KXVWmSsg6zKEwEGFDJ/yUcmVB+20221hs407909TiYtKlY28zBNF5uexCLvz35Yb
mLRiOljHlYBwJ5I7OMwn8efb9B8WH6sMGdma7v2M/+JcTv/qjI0q7TkJ+91nor9m
oJlwk+Yb5XAOV6IVwArXhPQP9zjJSkTLfZTvvNy3fbloAXg3FyMH/LeCFTUTwfkF
62K5d2wdbZuwrWkNEhg55RS+GfuMUgJjUoHnolQ1luAiEAgJETYZuYd0UO//jtSy
RaGpsH/oQcaSM8oMLhGCOZdqrBubwbnbM4rFCroSIfmEGcpdwqCjlV0J1J0AIcQQ
51K80QcrEaoUwGMGB+rfneqqjqhMUJhnFfMJvshXQk4L4vAQ/M0Y1tjxVF4tDC8H
1vul/CFswNTOT8/WMz+l4DEIb9WccutuRHrIileAjWF/bb0QpGdtb6j8J14I2uc9
y56GWolA2ZEozr90eEW92KViExCIauu/gXwjRgBvUpyCNJSkjOgu8zvHy0wW8YGq
8hVAakqo0JgL6kyr9AnJ7Lx3bHmwa0VZ9m1eiqQyvHDW/Nelc/yK3iVt1PFQyIMM
MtwVgYr0KnyztPTpQvaAYc/aLmaSb1VaXWc+4Idni/Nf20OGB67RjdWb0SS5RROt
lREM9w4gqB+MiFIHJ0Smz1JNXvb6Z3gc2G7saM5tmL/GLU61A9cYURcbDN9ijmXz
fwygd+79p6duXG3dP+cvBZPftp3EG+ovTIFqWrtUHgWWgQrrpv66ZRYVX0h+oOSu
bzZ7KPb1NRUBvG2njEUHgOoNiCIvQl0DYiB1bcL09XeiQwDg0V9owmtyT4eaOzg5
l1ZKKk9YM/JRMO4UPwkO1AhC/CCTpcjJSPNg0QdD5GqkhjVdo5qT1JAA4HxxDvz0
KYbT7qotV23kbIeVZPlHWTr6UQANnOk0a/rcJdcrrw84fNyOWk72GJHvc5s+fhGR
kdFURyMAEDvdccm7BBdXcvWckUJdyiftB1bKNTIQyy6OGm2c2DstgKqmXfVFCz4D
mov49tXB6pYiD0a6NKc0mtTUYcyocw0Ks9Z2+IvZ4xYIta2Et1eyxSc/2lvl/O43
UCKiwAs38PO5W0J3oMGp8iTY405mNgN5ooGHEaa+Jx1L432QE9MPDntrzcCJEbMN
1BHKc3qK/jt6D0RRyKwIaFazpnogfxn6b/Z3BNoYnpnxkuSYP6V1TL4QonoQnkpP
X5xwYgLVSaSIBQsuYN8l5jj5RH20XesxwDKvzU7D5lmlsM9WToJX4p1UkeS8qOEm
+wyfIUKh7iEKRLAZLE5hf+n9QsWOsfceEW4KjL8LzhM8cWPz5ZDkqcBHqzr5uCe7
6GvA6dCNLzyUfQtSf5QdF6eT//cQZpg5oqbMC3vzofXxz2Sj+mzT/GHfPEz5vSNH
+bc0yy3Spa/GYAlGb50kIY7YwLlo95qNSUrVQinSPKy5mVO+NyumaW3cYvdG3nRR
FGfVZk2HWIe0veNfWKmmTdRoXYGQhJCJNBJfXDGJywGLsXzYRUuwbTDspPgzHA8e
8C8uZMl7TjweTbQ3MyWnGkYacEYT9q08GT+7bxf3Vit32iVGk4cK1yaThGPOzl/0
je9Ufg7rphumn4vI6wFoZGhU/MmyI25bYT7IsxWG98jgQjDfjcIhJOerOEBxpdcG
6oejNz3SjBVSlyj+FFsz/NuqMx+KvPj/TWoyDsUL37hUQ8UxCVi11391QbtT7mfq
DYBy+GvpFWgXzhgD3vdzUBIMq0U3fDid/gk2fLWIe3RQGk+SSWtEZaY9bxE2Mm95
766E3Hb3vKgkRSrm6evhR+jkr5wpnHge2e8Gu4mejuO1fPz98NM/pMSIfpEYTtY4
/a7J+XrhL26fu7Ctx2UOaShmsN5fL4+IJtK4tEIyIxPLJHZlZpwhD8J1FutB8tTg
xIuRI1Ll0b6GGFgh6zYqu2LgyIwH3nm4MZYoa/9L767QRR0un1mKiGg+tRQ6AWVj
fgKyHRHyIxXi8Y2hIRnyWB6haPps7HEWirUIw3pEgT2hhSeq5Bc5KLxVss00HdgL
V/w8Qhd+mXL2MVVHV5I5OiPGWC0PLhJhdJRDAcFMHbevj27Mrg7HFi0EhnUtJv6A
cqtHtQyv+5zuXm2for0gv/zKdwRGQ+5I1354fAgBNbhsoSsAlNcYbaCIfSz17ZOM
KwRWpLz2Q1ufS+0uXO+HhlghmU3ECmIYaQPl4aDFkFwgHa+KgzuJ5sQn11dtbznc
s61m7eoko6kzPkgzSbzz+i5shaKlv6fWQVEKdmpuHPiq/J/5Ycb1Od7f/8KKy2A9
jtytiR6GVTvPlvIBqM6wAVX2iIWnMLbI1il7qAh/oIjIIkbuHdMq/hDvBTMk+Q9s
Uh7+Jk0bjoXOzdkSHzkb0pMkzaujHWOMIqm8t/PbxSP8b8VEDJIMHTtKyba7M1OF
wTJnjrJawtRcNBOM4CmK7LgU0mNphbjcfB8h9wfoKKLjKeQXBJcIpzmb7ckoyyrc
9xZYOWDj0D8YwU31OR2Yey2O3MTixHORY3wgqDCs7fP2UrKKxSZnzc0cjMw9LkKa
V4zCPrT6nVLMKiyegzLsquvPDtsA+bDFgYSYRCpmwIQMsmOHTzhOPASK1MNGRENw
JjgRIO1zjMiuhfMyohRVSh/lM3QP72auvA5BYtw8zC3gZx4RsCnXriW3oVh1oAT6
DHIRgq1LZD2kjIkLbCmuKiMsdOOnK6a21gQdGY2WvSOXKrXERDhbrLhtQP5BzTCV
txrSxkntLJal1TWvX8+YV6DSU3FV25jK/RQo+c70JSUJ1g7lYpL3FreUDC39KAzG
ty4Nymt2xXTyJ4tl+BWasAkiA/id9t+yd5NqGWVqLt7iFcKFo5qtkePJEqA66g0T
q+0bAd09WBXjWVvHY4x92VsxwDYtj5IfuVlsOm4V1iOMowfkwucVoFn6sdqyMLxH
vKEH2MUNh4rXSYRlaKLOQUV7sOM4oGicOvtFXrFSwj9VLTBcI5KaCOtEGJ5Td+fH
98U3yRBb0G62wmAUhluwDxnxyl2K6lHZ0VV1y1f9uSHgJH9lW53fwOuwJWvnGw6A
KCZ55ox6Qli+zJVBR72TiK/MMhZ2xhBXJdbcC3xvQW1i+CwWbvq3GRJAEQh0QfqB
SDXuBLJeS61iZ1xwVOvxhBbMRAHixH3xFZpfU08Q47nT5/bAWvjaCEHJcCcdIYzN
zyhEIOJNrIZaPqc/XZ/+qKjWX6YFJBvffdwrqE9/6G7/peCjg6xe/35QiUE15IUD
Y7MiDW1yXihHqIJohLmnVl52VEZpL2tUDFfWvoPx49mvFeD8ynkCYRjMJH/MVZw8
/ycN9Riof6ppYepGWOqgEVPX/fD7qdVzD3k9IaXWk8PEP23Wy/Sqx+x/c4SsuJm3
qfRMCzy7WBb5Z9dQMpQsRcPSSqmJNKrT+P/cDEn+h47JCY/awuWN295ayNin1IS+
CUIK27w/Pt8byKZUAfcS4CuZ54RWyBw5Ae3FD8opIJdxZBiuYz3AWQH/w5K/f6YH
U+zId9YzeTmZ8OnXD3ySAgme2a9YpDQMOwifSr0uz3C7okvxLTA8Q43laDMtYrpe
Q/6/GGX5kStdje8e7v0eLUQIdShbHIzBr/ht6XeNcfWdHrYvtMHSdAIZqiQQzUD7
MIPj2mo/WGkAdHrcnmTB0k21MvdDdIkHzWE1S1DizcHLfU2CzOChRxrSyuFNsLYC
72SXghHEZDHfBl5w/AQPuTWTqfPjw3ZtKEFoYGNmxUPJZKxCv0o4JJtPBRXnKgSD
MK9g956PHo4HQ8rixFoV8f4NKECzTPCfHlxzdPe4vkd7y/LVGKM1k7N/SYprWw8L
F4+LH6xP404HyBGsm/RN7RryFUOyqXOJo791V1wPHCRr3tC0BaIz7kYNwFqFwuKc
1HkMhfx6m7kZEL7EwFlFfAYtS2lVfzkjuCcnAnDHk0ZNfTFeeVAWriKT06iFRLfk
R5uaEXzp6ec8iwoRtoa3Wmxz9ymBxHj0zTd7Fa6YyBsusNO2jI76XHsam5kepl1E
tR7oo8oR0F9Wet8z2p14KXFQTt9W+NXrrZOQyxxabVjrcU6p0kH88Y4EjJn0/SK9
VdDu9R7jsNe73ErmK3oh0UheUl+MMz6FO4Z6WZfcEJr8hbtWMHhXdbN5eopn9SpL
Lq2HbHTgQSbE8ckj7jdB/A3QCmFGT+vwFJlTE9DKs2aWGC4LtI2lGpOHVuAEx3Dx
4zZFnB4dJRePteJdh676a5Bc/LgFb+KLK6SjNxsZXga4sjtY7bzTKMNifSrjzNgh
WZ8ETH1vALHrMScdyXHksa+V7RUBfWZTZZWopxYjoLc3v5NOf7Ox50aOkRIkL0Us
azQeO9XEm4gJNMxDoiiqwHSY2YPUgYDCAEJTxCOCIDlh8AIgXxTm0zW0HCvnEujs
F+9ItcM3vRDI8XwvhtgJPgeenm8Q0jYh2aNQqiAq2KF29yFMxo558u6LQ7hs8TFL
l6Ynr80/AFou4SJJYCGyu37gUUSy0+zKjUHi8D6zy438jWwF9z8f8Qluk7zu7/NU
PrNY6baWGJX9yhzLTBTQQk/J9gdEVi/l9vcciahijopoOQvGisZpKHzGQ61N+h+M
fG3ltSMcugJdCxXtRU1/I8uZl9sYT2VSRbc2lENhOqQmnVbhujgDfSkZUR6/NeQY
Fni4aTuy5B5cY5ybZypFcEuc6zJWWuoTx4nYasIL00ptIUF16Jm+892frNiwy1Dd
y4CKrHh0FZzLFlZMPieFQFw90KhDNSevj8Lh4ubQyZrCPnCj3LLDnIQFdjPB2UNE
SmwaUlCEV4hkqu811e+iYshk1ix3rk3ikK/VbagI5USRyfx3HtH3/rpVBETvsE5K
QrM9l9skEK3k1oowQNd+6lO/KsIhPTk/LJEWP799pz3cQaHSd6smwn7Fg6WJ9hOZ
LVc2RCKbpiUruUg0B+ErbvnGk20dqQol45HYp9RGbJ9qteGanWJEpnZLGU6ijoR1
jzkC8/QRuD2GbFBY+MJsAxg6b1PeIHL87VtOEUITNKYiVMlSiUeQRu8qRbpZyvZ4
+crbpX2kZ0gqoE/aV+dI9cupf80eW8Eg78ApFVMf7QFsMyIUZQd4/VSmUuIVNfES
2l0Fng+cC6SOyz208SKwTyYRd9eAe4nuheJ6Zo4mTWks94UJewbcBS1ceiOGAQA7
iVu54SJvxsHl6mBi8MfJK1dpaBan6kpfgimg+5IKrGbD37MRLeTialLNpHePFSna
fUhE8adiwmafDEok1PwUgFtzyAcIxwanH10VfHRyhOLuGLdoYT2+jF1k0Z6O9xkN
vcVfDMYxiOE8ohpvz8XOHnh6qzmWS37HkakTT1T/EJBWDWmVU1JXu2nkfdVLHj61
Yf0HHr6D7R7qf80F+C1OLfoomaDCsrS6bH06+CKpzVuB05RrYBeEIB4RMw0lfc/i
bZCXPBR6v+mkYJipZlsKTqz/BMQVAQE37LycsJnkBOrU6XI2m4QkF2IyPrDZcBud
yrmP9EsqvZ0UN5aFdIm7imBmiLEppChqRG/ZhLRPc/bItfnJdQUS+hH0NGXiaD09
3TVziu3OF33El3XenxqV3Ksu4v2XdH9DcQRpFsvMzsEN7M4Fp6MHF76CE1S80FZE
0EyisB+rcRyDliVAyqiKc+GWDVQwS6NDZSU3T1UU8aM20cQBGZj4HdQM9zchV9cP
sLX2oyAnDxhnNQDQcOKAuOZdciKGdAD9CRgb0tPPCXRKs3sVcxNhLlMMWIqwKQtO
DvEROlZM/8OFS3W/IM1y4gOeoYw3Oh8Ljv4O/dqr4J0DJOJ4gZnDjLdy2nv3bHQD
7pnkU8kI+VC8EycVn1jSA3FHvV4K9cfDuXPR+KKFpsbf7XLsnOszclOwe7O/Q4fB
mUj9k2N/90FW4gMPiw8D39shPz1T32qob+Qx61obK6zW25sWh0a5LV/wwaIxaDVo
I8/9BNq3HmWWge7eppgT8j+qfBSkskCFtsrotMnnEF1xLJ3K38Dovwo5BA5z8fH4
8raewGzJHyy3g+N911HE2Q6O5x2NC686kXXCGJYxkhlyBvNwH/VIbWSCaKiV2HjF
L5f79/2xeOGZ6q/q1KP6rKHHWve4QmyfBNsVjXNUo9qcaU5BIvNk5pqG4aFc1Wpj
8lMG8nJ16cftRd9nCJSI1WbwKADPEhJnwyWKDC8R5ZA8/0/WA6kuDDpLF5OHivPQ
IKZZyp0esE+Ib5z9NnJD22BPq8cOgiyV/2Zrgg14k00os7xPm90ASqv57gFmRZB7
Nm67UWYgnBUPuUK6CDxtrMYUvl+u0tvUAR0GJJYssNkBHQx1tAnxg1RW0GsHlFvX
P5OJ5VJCHgAwfoddE0+sCEbXFt6MUQziTdBYD2mGF0iV6wmq85VoG2mbmnGrNslC
khoemhvuSbwlvp5V1MQG/QWuDWB3jVLByguiuTbEXZMNlRUfpGe5R/8zVTMqRAoh
GUZGQ+pL2RuzofvQ0fhxJbsue3twrH/eUNwT9qTjjlnLJey3IO0dybhOLaK0i7Ba
nVD5ZBi5U5scGZ90UZpLt3A49Ok8HE9sgkaAb5YOJk4XQvKAZxXlSG2ZgibUj/2N
yL72jOcSr6fvZv/OeJ1xcsZs9+qZ+dpugq7MXqcH0vLbjCNNpKz1aq1XBxOiocuG
C2YwXwdrPFDCMjk/ICBB8FCO+/x9VqugMPWpUF8EOowAYUo8NwMsxgo7fnJNwL1C
YgeY5EgN4xOIdYwKV9oJHzC2r2sgEg4Rzx7jve9ZH4P7K+K8QTVH5tUff4upLvUy
ixEgAdvLs6MSSxp+EQxeFRCki3v8h8ob3RUA7r3J7c/2LEiJOTWXSJ9yspd2MEDR
l8e5CqyWtOXWXjLWvTogkuNavtUtwfNAQ/lv6Fekx/Qx0yKwVGPKrJJipJraRcnr
3lnSNU9YSOz11oTij4rzRqJG6MoUbMSCd1lnR7GlxhVzOrrY0GwgqsoTyYmaaCVi
31IK4GXOe4Do5fIDxx/wMH+ddisvZX9gnF1Gj1W0qB82wOyu2FotNi13SKVxlIKO
PLvxCEyyjG1sNpTzgG4+il+4lmxMhb/Mm5M/N/dFXhNFrqk/SrwkAEFFHk8QoF6A
gx+5cc/sFbKaHbeykofc7z7vbhnJ6bXHDA8bHPQgmgp065IXniOeBGY6VEmn/X0J
bXTSfgXbnMZxJPeg25NkT2R0gt6p7KiUdLHPvLzBsE9+N8TB6S4s1x5jOfl/Hudm
p5+wunXf8KvSocIP1eEKDCdEV4CahPyUxvLs8r1e5L1rqJkfmrJrFH+tSY2x9xNo
ZzraS+E0SCUmCdvQRLVr8XxUaje/cBB0Az/FfV41knonjZ6H8mY9mXONowQLpxZ+
CSDKhaR6GFfGtyALKUQl9CPv21YdweDLjGQJaCP0YzF8darV54cMLDQ1WQRTfdwT
7Q1WXxTxZCN7f/2jSKKqdp3fhKCQUZOeBqoC4bgLiSIrF3jRGjetSb1lUiMNhkLK
LnxBTDVuA0GwQVqOPRz0BAN+L66IjcsARZdlZxyvXFkCActUftWVQguJDgn0jWAR
0RNzxw0MkLhpi1eDHhGAkHTyKoeKJbaetiLgrJhnWYTJNRMSfZNRQWJN7AraTtKx
ohcq2oWm/VnJCaMVbjZ8Yv6Dbgc/R/NzEtdZpqaTb0HbEHXKHtWvFTxRrasr6AZF
OvFkYmZmU/S582smByNP8rM4d/C4GdW0XwVXhuj1/JgATQQ0ck1qwbT24imuSfkQ
80/iF78nxS7/jcW5X2ULhfwA558q/iWPgCrncMTZFJDNxpleUN/1OcXIlVqoSt97
imHMVDjarn7cbqHJmZ3bsLnQsCFpzlXIB8At/IqAKj+wGOxeZ/8IicZdTTaXd/OX
soNeGvyuGBqJBYpZolGVvhAdwKMbyXHpBTHLFl9IfRQeMR5M7oqVmUZDUqm7uvx2
r9860efh4ONv+URjee4TYoxLaDXnL2LLPSsfS/UbZIdk5t1Dam4HkV1nzOgC6da3
IoPA8EoR+7w4FCaqJNVwxBEi+dsfqA/W9Znw37POugdsXkQAeK7URMb5/2vlyQVb
z7TS0N/Rax81dtMo1joZk0MR6X5rxhkemRdL0EV8uECQX8f4dLTpaYhbWc/lCOlv
PYgrV8DV7IW5Jxw8IiA8zj72Tt1I0qyGskDB0/IFBTIyxlsvUqKfRbE0C9H3OztX
bR9K/vWL/m5ydKDxD2TeRCqG0XMFkR7Ut9vIk2yeMnv2ktpFijeykfunHSW6ke+Q
9bn5LHhFSbYlkdXFHmiLf2ZqDIkPyOOGnChFUjoPho74/g6ZIDYG4QLLlBnmbukr
JvRdfQy7W4doUi6VPbShX1JbKOnW7cSIE7AhwCgpK0p5PQRSG785s3IeqrQxxZbS
w960SVHFupXj7SEnkPV6IGs/pxatsHiHFOHrZORxoScIK5sNzd08DlWEdHOPOxXz
g01W4jFZqpItKOAJ2FT5vPKYZH9xM89hy60tAzgbnVCI32LOv7WR1knRDoI7b53l
xYVmIYBwzn1UmTR3YMoUd65LwgpatVXmSMnu4gRJy0TlYNAflW1h0vrEdxaWLvEX
24dTQ5hGY9zMyIrGblnGCyhXQbdEaqFKOk6hEFPqMrtMVHp+KAjseY5Fg8bcI24f
xCYvjX801791TKDAbU4EskEBXsddR5S4iQ4KK9m1Rh9knrbijpt0+LFIdKrmBTmx
HLqokVkn21oVNEyOWeyzcYn0pxWZsozumuxhzfS1p1RacVOhGRmQlA3yhnJDftvR
1ZWZKY1Be+3ETRKssLHEHLdf75dJXi6Z12GinjKpu6S5FcEKJkQ/0TiSWW4fOIUp
GKqFSJmEXmGwkDyL0b95XuFgaO39Vr1YRMpxO2etsFkV9gXaBW9VP5EzMqOCv+L0
VjqBtxIieZLixmZKp+UpheCweUYXIrqKwcdo7zaW96XrX287c9X6y0OsEVUcX1I4
2Eo4lnWuGwrTQHot8D3gsYsu/I/F5Ko7IHqxG9guM3A6foDYww6CDQdReRjjpgRa
6W5gJUCpJ6LhDhvvLZ7AQh2U8vxEORrzrrzG3JDL0ptf/OLNJPDiefvlgOLfpoKu
2lAHeOYaJMK5TBM8aGTBi4eUfIkZvFEJHZ51BwwlgEE6gOZurRG8o7xX1pLSd5d6
3HzffRKbvJBmX/bokNxjG+YVKA0yNIJRgZhoLrK2eGVQ65+5XXgWQU4/ZotyvTIq
2juccErnmJqwfP+v4a9W/RRL/Pp9fsLYmtsYKuFg992f5L9H21U6cQq2TSSsQ53X
aEXwSZL4zs7RVfLmb3zVY4GL2QfEsrwh8B0PZOgd8ga5fn3k7zJe/fdVnOao5WMz
dbanCHoaPrbijzVKnXzDJP6MO+C0hJOfLwfIYOLJ932PwH6AAZKD0LZ/k/o+yx/G
kwMVZ2AJq1fB/YoD7wXoz5fEOAq3Xf5GuFdSGU7cWO6WAfCYAHKlj0mckzUONveC
VZsnRGY+6aNXSkbgQGGXmrJSCJ4JvcZtNTk+Mar13u101J7Oeekps0ybBnWHSurY
+DfPoiXNIM1+Kd0YojVAmCjSmyHAhA6axaoeTyJpHgKlq6Xar4wbPvkHJOvc+HUP
hQLQ7ZHMSpWpgmToY5Zvi5nH1K1l+UoFAzbtDPcu0f8u/59B/8yoeSdabbvGf0sK
6BebhPuTlIV26rXGBrD+zLp8Cy5gPlvNp+AunVuOa1cEt4dyzPTpotIiT8gMru5L
srWFpkYknvSgz3VPakQndxC4WsQP04OOVKqJJBnMHTIfjHabE9R25koeDcPWAAm3
ot7umJPShcrjAr/+wRNpkGMH1zd8f54ztT9y+YA6Hb2vJUwL4IyC5AAZWPS8z5wM
VERUTvVU3+mRr8yPm1XegL+8R4dzv2ZoZSU8NWfvld0spFTzEorn5HBUYdxIyU2V
6YJkVgqn3Vbcj0n224cJstBY0D34pRe/12iLTYF1xNbeQ4vO+AD5zW/DhYsUIjzw
8rEluQNOJOGaVEH43yw2Wevxsp83X6FZpD4HcWVmLp4sGGrUnVZjaNSoZpzc4L1u
FqYLwe8zfAGRUQ8BA33lfsKT3R51EJea5lNQLF++/wPvD/neEmAR9KOKLFIWRnRV
KZMYRyoBNtdv05sFjhK3qfhLQsdm7LYq+Wp8PbvJoyK3JQ2aVQGNuz8YGCmUgfPj
8kiEqnx1ocWxN7LbFLRYn6wJEjuTv+ZryCk6LhmnBiiKGkRRnPEGWJhrSvK+tbCq
kdxHEh56kUTi85YxTNpMYNWSEzmoyQXTRBfnFrm42tFIxIrHqHE+FHTmnptHN67f
QcGMCySzhRGhjKscsLP/OP0xuKI8Xn3VqbykzfQFIGSZUz3FaEDZaN0ZaRWD9ccG
2xpi5eyb9sEWrWynaPq1PR8PsGBVnleTS8mdAJf56gs2zUbqzJxmALTaZrrnTewu
L4x0kml+bDgq4knOinUHgKDQYyG74eR5q0DSXjBn/2OZJTaWe8/HyF6g2vpbRmIW
wQcGGbr5tXcMiW1AzihkJETUmOT89yA1vDah4NEuEPyHZA9zWYVd188q1HIZ68NM
IK7HUZY6FO79wFF6uajDOzHQEVPzKx6Ce5tg1j2xe8ubfoNiA7ctWCJ2CgKgOx1L
HsX8FIo8ekIIUIsb2XBg357PnhmatFJDp6meDTkM0prhKdQ+GKQyInyHmoiYmo9a
1tlAWPcBSYxeadO9QbTuErL3dtG+7wPFz8Dr4bK3LBog33TyqkPx80PSGmhWdXvv
0BaDL0SU6fCU1IK5EXbpbaiCG/hLNIgmVaalnlgGRZ6agsupTUzOx4kNl+22ohej
wNaMZwDQlnGhhLGnVBcpFz4Rufg4UNjoyaiSXknsnPKpzLqpbCvZbcW3bzKiGA4p
TB8enWQnBMqXxy2bRnPGWlHSxAg6R/XycjnRXHmYHoWPLbb6yYUbcwns3ez70Qc3
9/SiVCNIBJWmavVO5VQv8qLrtt3NGJq6uGr45o8nvb8CGfOR+e5opjlrrB2+IdXe
w+U8y7hi0jph9FQGp1Y0IITt8VwrGa/KypnLlyWQ8N7WgBmSUMxdZVrV5FJWf2lX
UnyRjDmM3zdLZfFZyni/RsAOfJhX6oq/gyEwMf6jdhjPxKt7pFV6aBCt5O++1cfL
JJ7aBkbSuQq+C+jxjvEYQcZ8/k6poPQMNJ+Cefh1YMZT7Kp9cCmc3jaoz8vxjtFp
w/JdR4ief7OPUZ1LBdc9s3KeuLHc3us+NZeozdK9jgP0c+sMvlyzf+sgH/LO/IzP
mfkRNFxHbyqtrq3xfm2H32Ok7r9ZbzWjdH5v4GhwyX/mjTsbeSut4Af5eWMgVH66
ORSIYYk8n9KDt98ayK+j4WfTEjfNUNdbGQQP1G9RrR5ENmHPS1gmM2tvYt5H9vDo
2WPgAaTdNyygSQW5H2fmNuaclQaMLoro+VmUKZ+lyUWwoQgCFY90meNrLrCqJY5Z
+fXIsJx9O5AbWNSd58N9ghmx2CPtRJmC1cGJYJcOmexLtMCeusxbcDtozdXHhc4q
T5nAxKFPqKDqWAs5oK8Knw+uBDNnyB7xxuBla/EthhIz3I+/R+MYqzpcfVOgcHZN
q2B+9I5hQc5DwTsdLGRsBp9a+d5mQUN+5TypYagIxav57igxaihzUVDHm9nZC6WQ
k9mKULkrp/ItFzWBBUDpTUKtX5eMSBcmJtuvzg74XTHoxAcwESfiyP58LDlWjCgh
zgq+F6A45iqMDI+WtTVVPynKLmBVc1+/UqAc9Gr/NN+hfE+SqPwB7g+JCkcbpPWc
rq+6ALtPaS0K/WftpGqDQXh1+OqOieeroHJKcbx4hJKUQSeJ2b13ptksSq9UJU8K
UxLpbK2sVlPa2PCWVbMTv1/dh1As0NYTLo1EPUA3Dxt4Qvrh724Nsce81Nf5rer1
dQsei4jbM+HFDxFymrKzxVjRM4MYaOQ2+7LBQnSCWXLrwisp+usG0z1P0YUd6igE
QMOVYGv+yaDHo5SgcRBXju5aKWk16DczHmpZ+I7EMmCgzcnTYbCeAo2l7citmi7L
B0pTLAz6L2j6nH4D+wS45FOSjqetSIxu8jCXmQSn2T5vblfbY6jI2CHfme+aNEMZ
QilZBtIQEFv1uXk6nR967sBx2GuN6nsiq4/qmfVKNOg9HLWYC6bxonOA6anANWaG
mxiiHQZT67Ib/Tmr7QzvDNhSrsySi3sZRYFVsqUiAT8Rk8vriQDs2FxqeItUV2Hi
mzaqPs4j0ZVU+sl0IDU2F6Ve66MyMqkwHEwsi1iBlKnkeo/95lWC1/9P/mD8d2zX
lJlwpWHFtgm4NLrc6XjGjhHVelsFmMxqFmOnRtDKgrfK8jNvjUfvMYYaLPuwiMwI
oFlRe6SnOlLv7LKZWzxFqO8qmErpnfBGA1kC2Cwt3OtMgWHtNbTVkxl+n6COT9AL
mEozkNY4X8+6x1DxWtuIej/q80ozcs1R+4oa0sD9t113MkOjslyDxDtDONw/I7ln
66Pnb718c9k1g4z4yn8vRjcl4BKEDWuNuh1cfJuuhppbFP54bku64WdScqA1VFzV
cRgV3sfpDXGycPKL+2/Zi2xJ0e6n+8q83+/b4knKDDrJP+T2uY1oJjE5D36vrD/b
yGYfxYORAevcOmdurVAypCkmXydwRrcRQ4QB+4MxOrMxaadEFtCeLhFFtnsNnOBd
pYRJ677l+bT/tyuWkSDxD2QbsXBysu6O8A9lbsLqfHhlbfdOMO5dZFCUSgbgfTXP
Zm/BfbBFKXVz6JFqMNiQrbS5hFHsNnoQlH/cqVqfytdze0+FW63Qtf2kAv3W7eOT
Wwz3HWaYZaqVL+xg1JVfjtN1+IUwdNpdlXQ97PsoQkDjZk3KZI1LvFckIflSVFZr
Hh2LHe5qbzzI1Sk+drKStg+yhKL4uJv9wvWz7+MXk5TMwDixIX+T/GfMoRXHekyV
hILRD5+m2VmZXL0g3M9Ov08K1bXO1L2q6qmIwbJQHPfqLwJANshuE1D6vHZcy9N0
/8T+MCFvFD+/qtbobgFeo5ssLb82d+OfoRM231pbPiXj5/6I4cWVMe8a+uwD+4hy
1Q3/xk/FQo43Wu2VEqCGFx8/6NmaGrPYTTBTKcw2hA779u8sD4kaq3Mq803tK3rR
CiZ0qPxRVbsGEXNeT3ifKQNtMkOpZGcFE4haK1rH9zSWNm7xeTbYDFXBEElry2+S
7lFkXBiYQ65zp+7MLnNvQwypQX7I7/XcaNKk4nIUe3wW+ccT/PAOSdhA3CCSzh8I
KsK3rDLZZl9o8gdclgC8rY/lb8OiTfKOAqC2apl1v/EY7uFypEpGE3EDrm58MHRG
w5s4cpVnMMowJix4DrkZJSgHn2A54ZY+iznCnM9aE3chttNWquByuzgmCdYKqp6/
zmZrHjvexQOrPpwFex9BtFbg1OVpeYS8cn90UbnDW6QeC/B/HCW/TGkQXxX4h63B
EbO46eM2sEtsycxe5b3WE7pjq9Xjg0q/OxR7oKyMUZVB0mWqqxa/KGWL3pShe2Hm
808VAq73ExSz5PQyp3YUlOHVO8B4E/3boPB5BlYz2t3r4xrR4An7jvKGJCaczVZU
5rnMItQ1uYCngkqg27EuXZo2Ay5vcAVArqGVILAoSBbJ5CoKtDLdiCJRYoEDtaQ9
+6wjnU+RZ/LJSLk9fo0t/KEMHGx54hE241hE4hxPnNfKfZfZ8RAdkurqgmrf1OHr
OrjTWzRCXXJsCKBqPmnidS3/hLwzs8taDNz4J0ngU2e068oYtp0fFTRVsQBzhNv4
M6D1SP/yre3vd9VIw55bMLdA3aylisS+NP+lmrsBVKJohuXK99JCJcd91FTJr8Hq
muIgoDEJ7a+UF6Gr+xkdaUOhjAFAcGWgpg+3kmcsFEf8o5/5Su/uMqIjAsvDtGwH
f+5lax27tAzG+QNCCPHebw2J3pdp0pOBORSH9wygEaSKmijACc7+MIdoibMydSp6
0j/n+3bs97aUN9mufK1fRCOHavad7N0E6grGWUEWYJfdL3T/cKWRh/B1LajSP/2B
6zQouIBWOHiBAjkH3qZiIpGgIdnH9/0ivJugrJGyUNs1ZwWgTlJdQ23OyWJOnOYp
OiAIfritzr5KFafX4hEql1qZW39kCx73n3By7duw2iaoMlb2VisAxV3hGS+IYO2T
0DXBGM7gXKMmzlH5eUnuj7QIhtnMhrRtN1NKGsW1RqMZ8l375ZydShfE972ErzeR
p6xuy5Xnob8SFvxOeUVrtnMGoMiXO6MRuD818D94aVJYSpKo5XjPx9PTg00vN4R+
4bRrfmiLsA2grBdDvJ/9n+sU26rRp2VS2grvebAtPpJyNI1SNiY5u9ODg4Ak/ZmY
vx6ns/Q29XBeIFKqmiAcZ+PEb4JRMcYY4zcVx20KZnDwjzHHJXFY2//pQ7hLTmPH
W2XnuvkW4crC6F/aG7S8rWqek7VAyK+1t7W1kyPuKhqorNz6TJqQFbnRS8P50Zh7
KjxAJUaqIEzKeybnNJr5WmT1QFkDwgSAtlQ+JB/2iPT8O4c4RV6imRbMomFH0mM6
ySXptXeWYwHpRmzvWq9aSY6CAt9SdddrqQt5gv9PyZyCCgjzsb6gzIJMwwqtSNrG
xTnDOLWwaTPpCiGpRtLYuxZ7SnDTlR0S8KG6dMQp4APsa002GofcN6Vl+lGs34ZE
iLshtNBSXtyO0e7pBFIq0V4FQocYIzIgT9HhGCjq64zh8WPQTT9rdIOamY0Y5Qlr
Pelbprjy0kBJVjhgUvhzcijJzlwEUh/eBV8gtjp7xlk1ut2J0czcZfE0Wg+X9sGb
DxIRU2pGcPAbeJV8ZHEkBveuwZGIpzpvpRyMjb/Qbgr1dgA+RZ0AI64f8GwltGne
bFhRDDXr3d/qw2AmUoNCvjr8K0e5tNq0/Me1XtkTqJne1atekSZFZCxzcvD1slhf
w5CosfC2wI9TbSXKu/SCZlyhpgMj5++GETSCqPCUgEveqw/ik6VdMJU1RoBYex6b
tqEZgZlmczdH96JAk0AMHLNeRzEXEwdytOEpTtwscMiIce/xmbJ0O43QJybJA3Uu
Oxx+2HJA9zMR9YfCHzyHW+5uVP1f9UzzaZWHmdK33PVy+c3YUFUG200WHhrc9l1w
i7j6KsD8YXa41Rdme4ctMDt8/Sc07k0fnYXA67EhYJAMy6wSTvrdNAzqlu8RUdxp
AuTttweHuc73+khVLE9Fu9Fg4YJKznNcaTRfQniyz3qovYSJiUkNUnNck1zhj4rl
oFVS7EKLum48uvv+chGm7HahR3ez9HIu8op3CYs/0jB7OmnSVDKggnYNlayakT2E
Fo69SeomvSHt9sW2w50SPl89hxk9TNqF7GploXPOnZdRAmhOgzk2+VMZMWMF8KG7
2qkTQ+WCtkhzllbFXfNBvJMRWgKOHjdiCCozzls8v3wXbe/Q7FnDOuqNppGkOzEP
+NkJrN4VeuNWAkqLN3Yezc1HDoGK3wU/jAuxjLGeRZ6TrlBngRY3wlBKIgsbjpjJ
cffyT9dOO3bWJ8aZ3b3eRFnDhXCaSWtrjMk7JDqJWIKE6FnqFPYld/f2UfSTzUxz
UZJEpMeTzw5wSqkI7Qqn1SKXxWn48C1owhN4MyRplp4wXlHUTlVOv+N2jbFSK+Kz
umsXM9OUwKKtor8sk0WE5LFSFpKhTrz0Qg/sQzM66t35a/taDWr5YNYihnLLOeN4
DFO0Tt3aDDagMpIx80ghQKwoRoNWZMNk6BqX4pmPNnKtNSpPa7eXFN1t5Su0b3AZ
AIecIUgb4n7SbCzFggu1fyM2PdC+2y9Ia7d4jKbcdRo4PhWCrcF8x5OZx9eUm4Fb
H9u3HMiMjaHhqGM18tChIZKu+GHkeqAN8ipA7qAWYH/6Jnu3WQD1Y4ppIyk1W17/
VqBOk/JozL0UQt1xZ/ypP5z1hI5Ukt54c+AXckNeUsLMySH/brEI1GGXog24HwCC
4huRO6sO9kzDGVVbx9ixqmrESobwwqYvZUer/MdmjT2l+1UJyuxUFA/MVFGj7JRz
E7zoLnwH9W15zZXaI2zubw48ykSJZJaxZDefKYK/TvB/w21nW6JeR2zV5NNNR6wW
g0wQ9YmPJh51QE4qEIKMy7Sc2soPurcB0pEkYxTwFb8MwtGdbp4r4cTh9qiP72vt
x3EVMlmz2OwWE9suhGsb2ChUGVl0bWrAui/tPz59Jwy6hLSQ72DdZgTwmlF3up+i
UZ5loqJKVjsqCy3PCh7l+ydNxGawxJRnaVWFDs5+utwXXNHE5whZ5MAiRsWPoI6x
+KLs/1sLlQ3fHUsuRx9oMuJgK9Kf0+anxOuPM5OsHJ+PpRIiV8DQU3aQW4fWBRnw
0KzGaXebP1+7fWFeiTdZXFWrRPBpfB9YYyP+ZvbBhJS/rjIDh4C+IE1LwQ7lpXE8
g+vB73zakwOsLOepel0d3HqS6uKP4nGuqQTUpeg00z1mYJIaahTizYcHaTn7Neix
ZnkDkfogwSaKfmeEbOO12o4/0o8YQEyfdzCKL4TKyde8gR6nPekU3gjSt9ou6YMg
j+6xLQXBB861wPf7LQgIolIXZt+QyhMKO6cYCIcFSMRRor3cuTntUSlEFpDPiW/T
Qgqz6LfqqfFT1yeXakjsUTKdgp8KuyaMPzp9iFIFVIFW4JnX9UJzihPWq0rZ/aZQ
Emh8BgYpkk++Xs0LvtLrO+/4yRzJ/owf/9Njo97lKpf0Q4U527B3c/pzEJStxqua
2GbIsd07O4lvw2wo2NxXcBpugqcTe+TjUA1B0y5JUHt8kh7jSKDIoJbieWfc+lVj
ARh/ect7Cue0MS/+UKACzXUtw3X73f4zpldYP5ddwsGC8QsrJwDQFjJ6oLBlklDx
Brkw68d+TNxeaXav99Hw9m55kLngLZxtzrl49YoduD92j9YW/SWDJHSCPcGfgvSA
Db6FIaDW5qUqDWOCMXiJuFiQ/XENQO4/BRPjbIb2qnagM0/5fFrDmaKWYv007i4r
gA8ChyamNKWnbo7QSY/T4sS+B16Rf8gPWtBNcMKIiyDjrxA9HC458M1xOW7m5lgW
aiPKtJxGWiTXXmfh3PPcHAn9C8gsjBOv37yz7DbbpPznQtkeVSjmDIQs3ot5zyKW
hK1/zvSJj05moFf3h2Ex+G9sR1Cxz1FUlC6kNNI9hy6U/nopfw7yS+zYusoe4TVY
9q1zTEbCsUtmMLOcUwqK8QryPRQeFZPlxsI2IIuSV034/gBqhKNd3OksbuZjlZsb
3ICgP32XSfgRyWQ5S5D4SCB8Nzb8HqfS0h4Vwdlxw04gvIcT+48hXCICz+o0ZzFa
L+t+4dtYm/OqSAx01Dy/qd/0cyd3uTbVT4P+howhpLcpDofaZXcyHUzJb+rwqYVO
x6Mf5cdNilTlhyEUWkN93/4zbVRWOIs/GIMy0D1AyPEX2oOePgJfRwL2hxQbZqFG
qE2CAM7SYRCWOuDaVA1NGRF9zL3B+KTtooPREKzwbwIMKAC4FzipmSJypON6dTuX
Ko9VbXtSdKVs/urtepMLxw8zkld1EnapKHCBJvKLvMcB2Zi6o94jV8q5QIpbrjD6
osBh0C08MIX0n3VacKWT8petJ/LDZdN/JeNL1fdcdEhvsdZxJ4IQt99ZDyJdE1hz
Se/l3/k/1PklSS+dFJKm9cmzhUcPIUporxR8Z3A4C+Q0nNQGTaOcBhiQyS1wi23j
2bWk4Dhtm0hXrJ6NJCOM4m8ZBXiC6laXTjJg6uN6ddNXcNS4hRwlr/RbaZKgLVvJ
5TjYfuY7nagFIT19lzrwuXR53hUUScUzBCNaIQZ0qR3d0t6ilLv0qpEI5h5coUk4
QKRkwd6bmH1mBthAf5hBCtJz4BxihWqqCsle7JiNYOsH9oMMu5qQCjubm8IGVd2L
KgGveM7YfSINfXeUUlN6pGdM4mh1WAedwiLhEpHrD5a3jewgC1u+3BhLwnY6XEiz
ebLdWxLc8Ywr5/1jm+9UsHOff/LXcpOnooldbSE87dCT+zZ8OdoeRB1vUl0T5LQu
+QuLhsABnzrZZb96zCbCqRlkwxFWK+vyb3roz1a54XqChvDDzoywqDDAaGW9Tnt4
OrxQK7e/ZzL3UaiqpwlP6HnENk3mi92GvnpUKzwkNCcx/xgJPESTkmZMILlIk2Ck
2IiQGyLUcNCiSa9elwpFduqTMmDiMDM35NzMArhJSOHHJ58NOH25BtcgXEcupfdM
bVPZ0iS5CSAenwCAXs+tg0fL/8/+OSX7KxH0r0KUdII58mHd2hPZKbp0lbrr3Cw9
KYl+M/XvAMWfgGeY74xB572zt0Um5f7xpnZssgpFzYZrCh+lgI+0tkp7DwI6Z5QE
PzzGk4jSbaDhz/hfTyXTMS9iuDsgZamk64WWKTDWmP5P6+U/gS0Ak3PSHEvrWcB/
qY8iuTfaHbkWTKrlt5zx99lKSt0Q/kmFBJJpJyRwg/qmJJIOObLvsBiG70CjU38X
VdgYQJNIpc6Yyjz3k3WDZTHRz6ayxQK0jYeSzrFKE8fYR8YwEodh7NkLDMpLrTKZ
ZMjyREyT4KheYbEFI0I6J9yQExcYzYck+mHkBmXRdiB/2xho8hdwEV8ulafLX0Z3
mKvfE+8yQI2LHmi8lsKB/1IocfuUu2puNq4n19ZHMqKWdQzRQjPrsktKTgbEsKOF
zQaDZUCNw9gi49bU/TKrmcFTJjknk93go6+4NXcyjpy4vIo2Dj9HfUh+Y5CMdB1M
ChzNFiWXLPJleDR1sm6srwHWrLd9s6/RhZsXALnL/prrrJ6nb1C7q786G5CYXqxv
Mpi/aXIFIb6sRCxCvJppAosTKKRT0r4HO5l14VQcO01Sb/SIOx/O2+nUwZ4GnQmM
bYsMj13g/Dpght7jsYWHEGHD4dqhPm07kvfrZo9jlNRLym67sbO0X+qRyIYiDkuU
VVHaY2636ESRZkuIMcTYyvIwnpGckfCUlr/7FeGHxzogGq0pqTe77dBmZQFaOjeS
yFCZwupSJTrZxWd7RBvD2er9FWcjzF7COrX7Y7QUKI+hjdphCZs/uxFyaOGWBivp
n+w0tIMhqgUsK18iWYRlOZC6znrg+MBkrTRn/WtmDMk1xiw9aQvYdNBkmrKs1Rsn
KNG4x+ihkPGhIrYqksjZ5VE4EIID6He1dJBbq6XQhHeudScxT8MsAkgpjrVMDqUs
HsmLyJxaSIdZMPrbRRt+w6ymWBlSPwqdGotoy0L4EIzr8vL8dEToktDDbsvbbzmV
bgF1VX1kk18rPILnRjylrr583avdxDOCY/PC9LRza64LwTEZXaVhMM32b8c1N3bN
faRIgeaRz1vHz67yQAe21S0pffKAQCKgqjZEhfGVQf+iTcYQINUkYEEraotvFGZw
rN6zgiIYhNGURkBnY7xAjPbO0KL3UCz/GOFwKOAmmRbFXOgcKqB7Ube+asZ60Bqt
8AxHDTsrjwwNXSkwi9UjTkpPqv9PT590s0NPpnloDcHg7BVjx7/ySYgpXXeOk1dr
ynJhMGArjPSUnFrdT/t0tIu7MVzr6orcoEzDADtXRXHFUyemSq8/wjlFYZT1t0QZ
3pjCX23N8ar5bLAQwNjQu+pwXixlOaouUcbu3ZhURIhhdiJvGtahD2+04Ndx1gti
YugG3pd8W2TZOi2DyDmWLHEyNjUXuQo1+rRyJTZpmh0lH2M5U04y/A+pihF7UvLf
FzRN4SPQKiSMAJ8QlzdZeq88Gaz6rUGZ+mZM0XJmpzflvSxgZMzIbxQxVAZvh/ug
f+VwByGZJi9IeAeFwW3RxrZknDRo3mvTrv3p5dzY1/6aHW/S6boc42XlhXznMpIH
gY8psk4WctDuKIKvXaHvlILHq5c7qJ1FOMnlaxk5/1g/gWjUNvt6MSeuvSlY05dI
7wxGGbj1Q0vQQnQNRbMdBiB5MxPRbYHRcv8TOgx7Oz8JBfxfDM3LaVluCNqQWfkl
SCOC4DzmNqCxekppWI+tcRODk7R07nI6eA6iVmXjG3yzvMfhfbOdQFANWHELuJSO
QPSC+mRLepSkDYE8Q8rU/W2kc7Hq+bjgkkbcChIuH1wy3VNEh/p7NT6h9e4ln1Wz
TcS3yprFCMRCHaRW1z2cu8Pv2bhrRczUzkTI+Zayj3FaAJ3UDGT3dYek5R97x4jx
jEi2tVAmCTqLv7BuEuIWAyeqyHt/0Bdb4Sr3vjHs91scKSEMAhQY+wuggxiPiJmt
i1KECpVW9m9rtG06hRpftYKj9dNc7aFvnXMQdlSl6NepRWHrwAAlNSM/fl/nXNdT
tXuHJxF1xiXP80V1RUnDgrFcTnObxB2IH0vW1dhIxckRSMm/S8qDoqkiDwzeMNyH
TjDxEm96+e40McdpUHjF/nGdlLoXYLfeiOCAmUCPMLYA7Fx57EqTfHn5LREtIgJS
aUyOGVenO7y6sVPey1mLExSsD7HzmYiic2GC7UOtPHiYWUarSHmDD7Em8EZ3STLa
UWs2e979xL/cqr/pcyOpzuaAzAY1ux2k+fadV1fuAGt+vK8yKPHsU6q0oc3pP9XT
CivLfg9YBEFNO7+2A1AYC8tJ7/89BIYO8hMIFiFRjMHAcd+o0Hsu/B9sIA77WNOc
wYXb610QBIhjUVyLHHiQQGCNwRxDm3iHKXHWcfu2STQh0li+Eh7HBduaxRKm95p0
+7nMsGjRyhaKVnstNi/GQ6CmBX0HtgSXP7fG5ihI/l1cbG/nc5S4YS1hpicNaRXn
yxmoNPewIFn75H1yby4isTSroZ0gPnU+yAajlB7m+mwP8q/KR7E4n2XjFAN+dPuS
Vmo2Uuhc49RoWwc9WFbiL+ErkU2sBrOELgNf7Dyv/d6yI9yAoXvtLmgXFrrcRrym
YieDPqcjt3bV+77Ls4pEpD36hphjuyL8aiEJYY5/6mMIToef+kLPoCPaYk3AlI6j
BqRSMpuprsiu0yaFl9LJUZ4BUxOiOE6xCqHTXV7nxM+GGFAqBiVi8AvpZJl3gRnW
fSJNnhaY2Wb9Tlpmp1xDtId1xDeH8B75EIQMISJ2eON1wCAkYeD6bip9C7ZhpDpQ
Rc0QFuOFjFHIDb4f1EXcNSyBrPRu8XAKUJYdlXPWqCra45ny/WncGNnIk058wNad
K8mfv5lB3pe6M2q/jP0Vu8FA/H4Z0spm0DtJmALfgDYVxPSXqMr158+iBy4Z58Zv
r7dIoXhBUOthIVPQWjjSP4421RsJYW7eMGMXk7J68TLWMfStT1G4f7x5iEFJb5V8
oeOWQUYL0a2r9/a2F5UfSroNXQ7qM886mahhNRn/cUUDa7L/G4iieZVc/vw1ObCm
XCZHa2Syufx5oDWzMmtBSIYxkwj1jOMmuHen6eWu9Kel0PafJ3OaboyloypnwuAS
nZazZsu2SKK4ltbxWNitaXp6UjVa5caKukoqFGq2xp3ydOYwG9E8hlB8iEtv6MV/
QWKs6fnZ5bJtwcvKzvnLI4Cy18gtmW/mi0L3OhL4J/3n+QTzKibqjLRwJG6PiyGi
u9tdu0lkw8T1QUUC4NqnAJI9WB6cQFxNECqD/aP+2iB/zqpwLAV6lfFqNkl8Hj/w
1K+Czc+lpS86O6+sGuJTbw9GQ+w+6QmrbQP8bPcd0aCkBqubRfA4JHsc2fiwEORh
9tkk6IxMG2xym5EjBklk7X8ZM92B2ssIhZtiWODW1gsC+WRu06KD9Zv3nsK5RUl1
e0VYL/w0HxEtpKe9UcOvL/Pgpn8jWay68aaPtSoYZA/rkyLhMdWsYz4N3QuDSg2h
tPzRR8fyjkUYmLF7U8+OtAYHulkz+fQzzoIr+kjJrzZM2Kdv0pPuZmC94mSiTqsQ
DKU0qydChBvWmPePfLu1g6hiyxKUh7gtqi8jXBYtON6rwrB0rdK5SYUjRF9amtKM
4IOvbi3a10Du3XI+sCyABRaoJ3AXJgbHL3fRaFTgZ928sxJZ6SYJw336T0LU/CHy
PXGN1merbGeLEhJRbJCwu8xGvO0feofkWXkuQMetSsjZ7M1OI1bLW2IEAQxoUqW2
9KgMm0+2nzqsrQcTPPCRMa/nwpSMNJT51NCUHrkAzc6lmR/8PwU/xeUD3RabsWaW
iEmdD4CO8uCRb91AQSKJj9rbKmdrANz5UUHiyFLQDLXbT83WDs3Y7sy3/BM1cuSX
fsAcyV4+S4pXkf9uvxiQWL8FSKUTL9pRkkHup9N3LHuEjfI3wLPkptzK8UWvvpAS
ydsPeaVXorL9MdmAAE3qSO2Jzgq5HluKz+/65L7iP8jSJy8ylgzdeYTQFSczSkgc
UqbuoiEJcmCZk4OmX1EwR43REmtsnXBfsegeEH9zLQl58ulZ7iJ9C+scIzxddQhv
1MU2kyIjsBKT455EzHxeqdWasDfcHL+J0M7wDH5ZrpVn6sivBkqVRccbKayo9pvg
7HPF17xmcnS+DGVscnAZwY1dIt/WsNZfN2KrUiRFuLKkDgMAZGfM7j1Iuuo44uDD
XQ3IWvudOQBTVDVuZqStgFlqe0vlVltIlIJv+LGo1kveXlBc1jA1W5AEYm1HaXfB
dfiEdwBZkxI4I9zG+qOGqZD5rbCbKTJjJUKWBYVuncg0NWOaIui+mBcjjGT6LeFS
kCPNlJAlGdZVpD82x4IU94NgRHSPG3EG1wFJRPBmUzvliti/HIOZtJvWRbWVD9w2
RkWrcZdFAXEwt/rc6dXYNAjkAUxt37bVW7GccTKr//92JbFjxF8XCZ+MoEedLWxu
VvRl17Ap7RhcIvE+r5THq8Y18LkmVOM0ZsjLAbN8FNAN19cB9CLKBdlMlIX01nSF
tJDGIWFt4HqcgS43SG0byhHfuy9OUjF+8jvZimH1Wl4TRPk2X397qAYBjQixBZrJ
Vv55GSUuQ8CB5aPfiQsIfoGz2YJbcAt7Knw6ObkeR0txnfd1lav6t8UxZr/UXRu9
4OwjFFpV2N4Wr6ZvqhDwVxUnkj/4piY67O1CY5XIgT1q8OWg9vJt7huFb+P+IbPV
hYQuOA/QAz3XyUtiRAM1Ta+AbjRhyV8nSTVSdyVYkrhNxl+7gOXxMFi+K0glVfkV
5vpBmq5WTpU+8jhRllIE62vJSUb+jhfwC7wHkZ1tSllu9g4DWSwvgaAcj+x4+rNj
8qmOOGQKZuT5tkSM2V+IL0S2hM4Ppc9P7G6GSBseZRUg3Sqdn29SEqvBL4uVcVTa
/9UHL43RDVcA7Suu6WtgggBa6Z14g+4otxSCzaqbqJ94MA4P+2/xHVApfwtwde8G
ElIUFz0XZJYwcauK0aI3To1e9J7QwabC8N+HbTeFcdjomBRGmIbo4JSTd9DgWyDf
s+awn+W7SIAAilVz4dL7DI4W5xt1y8R3+I2RCth1jtTMfTDSZqKQqa5N9/pTCTXQ
9y1JBXpRAmfzmMQs5UHBwxdwsJcdfRX82gec3tpl0ym+aeFnnuEG+wpcLRKz0R5t
ZpPuxc/cUfPtfFBEynZq5c3aQCUvvnuKWmh89t0SxXzXjsG+xIVytNgArVtV7/Zf
XivKBmn4Bmw8Rccd/AnnapufSlGav/lPDXI+kKnOzOD6bD8IvzXi9pNciUepGuW3
iu5dRPVl4V22oHBXv2ppae8PPV2Ns0DPdM/+9fJIj4LZKflaE5VTEFh4y4O42PaY
tXcIt8c1YT4zFTTeSdB1Bt7jrG8xmmWMR4Sa+bGyt3xT+ZWY2pKSJ2y+rUzfuPt0
vACYE+87ZtA0IfGO6edhFlXdhnE9nbo9qllrmMxHFMjXaLtliN/W5ev76NLJHIV3
nFgkupAr6R+W6m7mctsy46t36xubFjNUyfhkhVyJv4wczsNE/sa/O9+2ENwXg2NV
FntTwe4lFdBSixMYg6F/5qEtx8EM1Oc/7ldwQt0jiAP3q4ucEdMiV0l0iMB+EeHk
jiq4bXtWuu5hU9EIEJ1LL1TGb19wdnhAlzvOnJCQ+zL5ukEc3eCMSFwvpKW0Cz9h
f7VDT4zdrsFHvWB+LNMjOwhuqkeBmVyHo0dhv+l9oV2LtCpKkQ/cnlvLVwYZL98X
HWWUsCLoRaRNGs6r1VJ6R3afOsz+2mcp9D0e6FpehdHXVBmPoL3+y3oV2Hna2pNz
im3IVv6UMeXi0QaYue/sa11cqh+BdS7gkxDG6aNQeG+DTZ6WDWNddDXOLTzmo3+o
VsGw2BLl3lEbBpz6dIJEuixLrVgvUY2vROVcq8+pLucwFPH7Cm/D3WwCDwz8c6pk
GcpaM9KfDAJMMVxwsgS+NcIgmaGU7hewMV1r11cqjcYnoexwrpt7rB2kv79nZzmq
BzOnYmB8qbgUsimzUqA+KxdnWUJG1ru2tAMTWrV8MYO2E5U9sbZxrlKIzCpmP+bm
JGY1CFzbLAdgqKMsl7U+Mc99G1ISjKlLHzhdg8XYvaZTDPyK/64fbh678AbpNYou
P8S3DJTSk7neKmAr9yAZO9f2vAXTYzafjXCUQ/zYZXAnKk2kdgZDqQugOL2aPvrB
D8rxSeggHEJpBO9WO1iQalxMqAWH3n9Vag7t+J7RsCOcvJBL/UKVmoFpbqpGnDQZ
CnplI4BDyRnoLQt/ghcRfYdjw8Xi67SDQ39J8OGpES/QLS+pGrP1NHxNAGIIOeu9
MWgRE80STdCshXsR1wV5W9dcsWSlpJZPQ7O/H6MIYakB+vvSZJR1Q/ft0rtynoQX
YcJ51/8qlFJIgtKUrpPimn44PGYErPnqucUw+GFxA8tEgt4KAZRKxYWjHs5qK8FP
V8dJMtEU4o3JG0CMc8vfqahalQhwV5L1IxZmr6JbIf9cv/pmVpRwWOQtsjxObY1j
m//GRDqMENNZusSz0NPxk7gq+DodlCV2x6Ofs6nhWXpSXyY8eh46s7w8Wk+e6QoF
n25zx5vXv9hkCufo5mk8bW2q8RfIqIojDTe5WOrnU83q//+fjCCWKo9st3Uiwit+
stQK0LzHjcMgyy9rrCYxGUIqirJ23+5brKAGzEULM4iUMvBCJQccGE42TxOAaUZa
0U5QsW01dlnfVACVj8GqgsTy2ey7AwFtso7fnSO3D4OE0tXAu8iojwJCROkBwBp3
UYmVanqTOsxPc9CXNTgw3G2CSxpHrr9l6hTDDXJY0lh6Y1jHURw5gSWPKDwT9Cs7
yQpUe4EXqgAepm9O27wPPjxno/Kbf+fMg0+N6g4q6SnfBB8U08JvBDvRVjdS0hox
aHpMbzztzXMI6qMe2oPQYZb//4wgHWWRwRsryMtXRKvbBB4Ss4yrw0GfvFQxet/z
sY3Yullryw+ZBKbsdGm49TPf/QKkbN7BxRXWiGF0n1Cb+1jCSfdXbtdRZVJxSoTR
DWKSt9LWL5upFnthawWVQIlLoZOUxGFg1KISMTZViP1oMGzpKT05dhV1Aeosm3IS
A2SbZEL+utii0NDZKLwfKsepPWBjIxAr4GU3gsCsOJL0OOZhtFA0qvrvyBbVbWqr
ru447jqxBAiptOjFDTk25e03SxpQ48yW3xn46h0uLxmm6ad8vVnz3W/znH2twYSs
/MJT4N5YKv8fu1MIGpIjPH0zBAMN3h0Yv/K3XVlYF6cOS1npH6ZxdXwMVmHp9b4i
i5QyGmbQgrx5Ismi3263pbHKG1nHZXnNnwOnBypfgWXgrMrHD1qnD/xxbF96+xTQ
iy6PjPFJuxPU1VGvtMLUGEaXXb81pEcT22iF/Oq0tqTWANQfNVhwsCl3BQWKt6FS
NxvdAMgaQ0qVzXfXzJd/55t+Io/oAD6+zFNTbJLKROJf6i5NBE7Way8HADLIV1NP
2frPVbUDDgBWfQIgqF6+ClD5QS4GyhyJ4J5rQ6vDBkBFjkcLDLsd8vKz2CfCCS6b
EJrtoPVytbnayur9NMIvsgJp1t1Il5qIgu7zWyjGb3mpxvYkhcMFYOMSf8M+iWz9
cUPQnqR+6nZD4Z0bZnCCAG+q7o9VdBSkUtZrreXXdxL6Zn5TuWZAlmJCsA2kF+Fr
yO1eajhFZ/qQOOrVNXdBWpzHXOvMfFZVXPl9KF3pA5giO3toHuxpY13TRARdiHw+
jYDmCTprOmxZi4DGGdhazadLRi6TNHTZplDVtWURU9FdKcpA3ussu2osV7ouPsTl
6lSnZZ7Ku9EtMZDTbXM5jqyPXWsMlJFeAfUAtOViNXATc+TxAV8bTdSS7fZZgWBw
9TehONg7gR0sh5ivqAoCpK6PFSpmvKwYKj3gGegGC2qo9HMgu6SEs861ksVPGG5R
/ukTq0iZ6QnbIa7T/CWT+JYQi/4bpkeiRsvWW1nyea0TEu4TzjrU115YLbhG3AKS
kyRFDqfeFxgZxq6vz4fvF+G8eZe0xuh4UKAXBPKz/+6cOTWq5VMGVC/qTso+9YVq
BzgI2GX/lVSnirK0BfTfwDjEWk+c57Ts662RgEo3DcpbZV/vQTXdFU67xI8+H0Jd
8eTF//kd5uixsJiP9HXgUUjk6Br8hJ2n2cPD9uLDDL42hsLGTfXFQctRNUfTiAYQ
P2+3qUHgsLvUmCX9fQW7ninxoRYguOMW63hBVFjldumJgjFNUEWKlGffUqkORrDh
L94BSwYKxJVJSsZKuKCs14TeDwDBPoAcxgINP5X7ajU6DDb+Mio8Oan+yvQz40wM
3Mer0V2UUOrGE4/aldtSIgYXWsHCy4HOLga44fp9JiERxlF5C6F2hKz6QLpvX00s
0uPhmpO7Bd2owIbWqwdW6BiRA+aCtR0zpwN1aUszqzgwH9b21HQ7RDrTAf2ceL4F
9D+osl6ezV+7U2HDBa+Xld6neGK9teNy0n+QnzkhEBhB0YXnqj2AkNIYtkxsdylb
av7t0Js5dTKGPm8El2yOitFvwfHmjoRH1CEkcfE1W7e1JfE8BfNCvucvPpFAlfeb
f4u7xiXuIZkBmxzh++UTYb+oLhrTMfnDsaveC9cV5a9ueedS+IjD9RuptzIc7hKF
WpubjFTgtmtMsKmPwAQr3viH/HIlUUfOnC7yjnlfW01A/2f69uSSrC0X7tWnKEER
MNLQxGXsNds5cqUERk9NONx3/MMBhOYbnW282tyuVfPHdLlEQA9lAkTm7TnzYt29
ju4Z+LhBLuvC5bXD4ROmQJEkfnKA8ffzhx0xhsb8gtFfVZp3ILnTxo1UHhR2ix1X
ol400NZ9zog36YAL0l+SucoA1aHsworYumbfo+5XnprpNV6KM1H3fzQzzYa1MmtT
Kvf48Klgbh0hI7bQ2oyNXh9NAA9kMm1MfdNiNYlFmO0676Ib9w3ZbW+tGNaxzlsj
HJwRJtgjzkvoICfkk0ScWIdW2Wl+qx7tH/tG30yxMEY7rgQflLHaFvWQKOa18Bij
3qXFLlRg319PivE+B2D2akJe9cSwp3D56foTdZSZDAVCv3csdoVdZv1qiZuGGms7
9lLEo3zgCBC/biKb1lZP4bnL2OGWEBkq5ZZz3kQwl4OriobGFVvaAPmxhNHqMWQo
X78Qb75ARvFuSzCGJg514UoExMrIZqsj4UPilItUy/3i7P5pZlE9HaR03mqeGRLf
/OAs28JRF0fht1F5uZfLT6oAoHmc+nuQrd57kYyhFEF+TfrD9H9fyZe2b5+zYZSm
Fq0PFihPYquXOdydOavQM4/0faiKw8LC2Ozh+1KAQm+IRu2BLAy+Y8JSTBaasNko
bAyz3TNeFmcqBy10pPiSK2+XZxJ52e38Ya6dLZj7kYth3yrp0iQcYWT7KCcgK5UA
TLe+Ig8//s+/QbfDqks9gWNvyXjmA1S/pbDnS/zuQJL7XUXRb2r7SL5NUyttUafm
G9LKVkDvV29/lGOeglofgCE30JAMhN2awpQDlEBUqSMOvLSZgDei8uFAGZOCapIz
t4NAQ8lZ1qI3qNFl4mGYvZ06ubpa+WSti/ybJN7ratT2xlDn933vmK1ZsQ7GCyi0
MLRIypEIwgxyBSfxWpqq2qzesr3QOyGjyFxaiaeFNHNYHOXUXaPh/nliEH7AfSgE
bDRMWmZ/XHxFfl6T8N6LIsiDxTVjZQFsFOv7Zua1yNAZZ/rXR3j1EawdyF5CldTz
xC2Zx4YI8IW0aaqc+D9kvHelPigBA6/FVXcxzSyqEsgl7z3o7FaMk95Ju6VLrOx5
gbwL47U6pQCqImJYEfKSnRs2unTOpdZg7YnhIV+XPLWNg4+YrB6cPx1J1z1ehx3F
zAwUNYupotmY61PVTFYwXICVqWdoCUF0oWPzIkYpZQ1l58H1Z/ShOpXWFqbMbcfu
OA76aVrm6tELunHoSbFTBFNRKMX1tW6SYTUiOhhsySd2ml6S7ogS6TvfOLsqI+CV
DuFNRD6ZpsfyJUUPLX/mntXTciCoaVo/bG//SBCg3JiwIvCr/q9ghRFCPPpn3ure
nAaKWFQXs0T7ssEsHTWAqJrq3jNIOCXpv3KZTIVgG3e2wi01frDwIKUPDj9jbZRu
4w9VYDnj0ZVH8f8F04f7Ra/Yi56bpkGnHrz8+CmFZNSIenYfVH21ZLosxTD6Q7zZ
0PgQJ3o5tF9rBgj9591Xo0EuxZaRSdmT8nj2j9NJqSv7aS6I4obGTcgVJ12YYfwg
4vsuyRPP+Cag17164MtN7Wj+5lzV7QTRx5AtmN5+tiawDzCbH+zZQDcWAdzqitB/
X1tSCoFidYEQcpYoGo10wxp5o5T1IKRgFOGEx0df3GCOLshTmDkhG8TyLXaHPFOx
DWuInFtRydn7RnN+N1ok7vxnEeUvLzAPJrfmLLSWpBGUfBEfW0OTN/JjmdwhLOt8
rtpysJbGpnCYMorrCeE2/slMzAS9fHAJ23frdV+fOWA/jPoSXvQE9w1aOu6eSzj5
tpE7GjMnNFv/PRmRZSQXsIQwQkmhV8dY28b7/mwQ+aK3LuatKu9wPV0X+Ta3fi8n
uxAJGc50sCHMfk0nOyG9kxPLc537RzFPPJMac1Q7hsLCQPz/r+oq6Xh830UzmGo9
fOkpid7YItA5DGM62cf/AYq/nIdrLTfnNHkjXdDnlL9a+z8vzET0Y82y9mFQVkHE
t5Hh6dkipjXz4rd0TX9dX+05gYHXMVaaHvJswgqG1vLgjaZCdKW2zQvkHfYjZjU9
9/fkU8yHJLV3mGs0eflwzhZQtePR728JyVc9zg/yYHG8tymIOzh2O00zszlVVDM1
zpH3q7pZe0FaxyHOpQRSk9AckqetVCCISs5cdPcA5fzNpEUCTshY3sJdFHyNCCq3
kQF4MQemyQ8MLeP0kEgwIAb/M6adaKogf6POAxElBD9uD/rxNZn/2GpT/65+eLLF
cRhpbk0IBeB1DytJU5DbxmgtNu/oCxuGJnWDaoUY9vmUv3rkIhPJx29zYNgldyzb
YhC4rKpPOugexHZCrxFiOTm18tnKkPTt0pUEa4P0rLSjgZ6mqrsnLJzz4D8fA7u/
Nb20K6fj3teHk8lA/0elf3CRhnBYbvAiOqdeEh7i4QYPrHeYh/iBZyS8ROjTxSf5
Cr/Q0L0irIRKsVLuHsqpCa1WACLuNJKxbFXFZUgkInU6jUKakyFTNgfcuWZqnUVu
rZUszjDNvrJPTFxwylXoJ6dfMaolAsOV/iNUE7cvoDJbPy8PvhRayyR+0ku9alHL
Wu6RUMgDl7VqSQpVMMfKw5ROHRwycetzU17ctmCHXKLtnPx8v/odmYmDIX/HUIi/
Ec6rMWLE8zwC7PC2OKh6TKGx75HmFwbmsqmcbejxq5AKMYcqcr0ycIq7GNXUIdrG
gbVNC/lOKg9jzN2ubb5FoBX5yNKfFWvgE/IApXIEyu/zn/c+Q4aMXU6XtA3OYQ2N
vy0owaRRT9WRm3Jr1GHuEt46Kwi9/F0A14+i8lAM9l/e8j0I/dsgvDD8Qujls01U
DADIUdkohWxnXa4PmHxfr05KLf8kmxZxTH3MGO7AvMLn8teErk0rCUbGim76pobG
KQd2XAHDdaZG5I18y76J/CQRFaUU4dt8Gs/aRwZtyuqt7A/1M+ZMW3ApjVR++Wf0
7Ot8TDAxIlw41wPxGoX/fljPTOAmyEoql3WhTvuO8snxuGrmM/aQbfdPxhIqff2Z
CU+ASAC/Pv/PAKu3w2CVB6whRMNvXAhKebHa7NPqGErApj61A6GjVVa11FwhM9OH
3e8Ah/aim+ju3Gs8eRrv145hUeuoWiMjwQepaPHL0LIhzN7XPDzXW99znoCnRNr3
h0kVy9lXoAWSp/Zr48E2BCcQQQn/EixpoVRzCjsfy/d1Cka50zClFfL1ANz43TAc
CP8ynImTsOS0WpJMGNv6JbNb+OvK5MduDT+2ZBzVb7S+ALOhqJekBf7VWggxO/0a
DC6Bidkz8aYq0tEmWINOspETCjk1iO9RtL8G9CjJElRM1WKS29T7oh8b8xiTievZ
eNdTtk2jpYGhqPMkmgp3N50sJr6GR/cA6auMgVCqImwtN72r/c/cTFhsClkGs+Kg
8fmsjQkChVVHihczdYAVbuBMpOvEl/NvOWlC7WpeUvJ2r+2gXl81kHSjhS+3Jsg1
96ayEQ3QZ/rw33FRSvznwegz6lxCvpl2ARJ+lxNRW4JNqbcbsVaylXPCAsmu7g2x
h9ieCUXV+ujFwp++f5hpF6in0rrhS3Jf7xC9EelhAf+mp7axD7TYtzkcOgo0f9I6
P8OTNIu4FqMmz5K2AUjtenr4X+yG+ySxPF/AfNYbpbkXFVdt+xUtftaBtv/rXRPI
Y7Pdk/T1qa59Nrh8zD2XrRPGk/hNT3gcvprSgBU9gnwGGRToMaefAFJHRibCsWzj
0UWWxpT4LSuAxuXISYPE8w0LtwsI8ILKX2ijjuFCx90o2pHD6noubnFcRKiMq31h
22yFNZEzkUh5gLTQ+C1b3lOohZB5lGRkoYcE9BMZVNVAfh6/qw95bkt3sT0nAE/z
CJdxLeDZCAmIL1oUv3hoE4BfsgrDoV4b7EHYMfBDo0Mmj2RffJtIYcLhLhtlpqql
KY/zxQT++mkrz+TP9Y2T5yLY6iJkbISZAnMbYRr+hKCAHhEV0JpRKaUll0GKFBy4
RfianANOFaTUh02vfO/GBVn/SWRqSKuOzk8BLJkQEa006scl3ymGcFjsQGu1XJHE
NosAmosQCAtSyLoThpOsyjOqczcfpRSCGPhPyyVAZ2da4F5vsziGHMaOTdtm+ruN
y1DgOwxrpAjQcbVwAM4Vg/G1obab8ZvcvVC4pJlU0zW0bu95Cy4+TJRIQ57HpR37
eHYn/KcBnaNsL8yPKMr9EE1NYCIBjzBjtKkiMf2FOBKYx/tS9vn3K47bFUIfeo/M
DxW/qZa7c61lNMlxue8dHKJI6Mv28KZuAHj3bTcoG10hh2v7GiMlfsViWplwwlbF
pXzEAGDgbhLiRvh9WFBLt/sOSLp3RVO7IZLoyaxGFAUklpi3HH4sFCY31CbcUJCN
XtsSV+BwhJnOmzJJCUbp3QvczScfzAvf0DiKTKJfUq6FawC8M8hztf/hJgqmV0Fe
xMFjWfA/zJS1Q5B9ETOAqqEOBjwhtkGurSqpcDz4t9RavuoHfeTKUuAfHNImvbrp
P7zLMOd/HY0NRvJO35ybN/QgZ3Owwxso5rYS8bU4vKlDQ/Gfg0NcdqHBwl+qnbWb
2XT4XL9OrBWTchPEpM2mFrytDGYTKx9pxe0ZgA3xsVNOPJotCmiNenHYnxrabJtM
rVTk6w9VFN1LbGPrDPJiOQnEWu4I6qViuU4YKI1MnIdOxF28O7O5OwOJLcxq4S8c
+EIuuDQ3Qa9RoeL3Y1Q3oPuQgnrWfjrpVsWStHvXP6GyqFGYj96oq+nwsJm16CCE
uc33eCCi4vj9hytecNgO34izmq82eoRFFwxwLBA0+dm6/uru+SiwD++ZzGXtwZZU
mGREnhkYbQ1+zqqrKnUMBbksfcSvCdlvRT/hWjpgYWbpMDO9Wik7CvOtqAKgCbf+
peysBlkY4lM3NjxgtQCDfD/FYorZMcOLzDlPpJtee/QC/APcOlGd+DtcYDhrVcq/
Qw0dZMol2DyXF6ga8IDZGj8dTaU471zUhu6Dci4XqY5DMiO2FE9xdOjCplYEjMRo
jUxd9mCKZe5aCvnybaarrShc6JxDX0wg3kOuJnBwqdbXiCJpgoBDvByc5xxeWRdb
yVblQKsbI67F5K35rr6/3F/HGGd9fTzw8RgfqiyYB/rnDhMB39KioG2tgWZ0Dx6L
1v1rp42Qh20s4+9eWKR50EIUZfoa6QCOUSnCr9S97ENZE3bobn7H0cUormkURtTr
B8pGdgKtZkV+dKk0J2MauSGfVe900DtrL1NnHeB7+EO9B0oM/zt4l04LBN8iWFvM
DyBFeUKV3YrWyDv6VkaQh9qpb8+3QcwBXlTRlvt4ZziExhnz+DblYhb3r6fJh0P9
8JmT03EMMb9elkovLcr7v7PRX1Hsk73hpQHsEIAXqxrTzUiEBoQxFxKTHHGMxICY
xqFbnq+AqaqjHbg8LmwaT7NXEzTcCKKn9xwPmgetHqE9p3cW2LSqDuerjnonLtRP
6MmCJ2BreM3FYYkzFDvFKoaAaU1V7sPmFGW3JKZk+KuupFq3VF5RwTx5QuaWpg+o
g2etyGSI4ZTOpwmkrbkCaJR57DthSDPJz2ldHLfpnaHzHNhSeNJlYx8BTsPq3RMG
GzSgxyUWDTYll9zfL1Pbb+eFcDmgC9Cnlzo7JE4/fE8jXfrqWYPlk8D6SQDBj+6H
sXmDrV6A0nTmBIF1D7M3Vd7OR63bXF7xq37Q7WWMXGGAxvf6mCSGd0Zwc/Cuzkdy
v0N6aSUNKXj6CJgTBMDpTNwvsH5KrVdTVjC3rgSBruzUF9SzsdndhawBiqZUwbVB
gtIFg1YvLvd4Ik6I7ono7x61RP9dLCm74/8Nawz3KHUAwkOkuRZ40GBiIuaot+/T
53PHAYQ02WYg/uitUDu3OVmZhm9pTAyhKcIIdsEwPWibCKOl0i5LuN1TQ3N0Mu3A
GyXPitsT+VKnZLlrRgTeEMwNvbAqtHWTTHgyJrAT5y03hIzf7nLBSb/YfWw00Cqk
hDgUtOfuff9voVoa8ZiNb32dMNciazxf6ojLRg5HdGIKvpnPfkaCA3i3YiHCYUrl
f3h4wVfqyfi/9eX6zYPOOdIq8iALPp4XaHP1lZ8iby39eodS9h445sipatQvC19n
NbGN4qnzcbCG02zNWEC6uywUTKWnwBDdFoWmSoETfBBK4k2yoBfUAx25nA4mOwFa
WDW638fluSBPDBx+2UBcuVU0n/GvmljLAHZwuBo7faW2XZz/k3cOPX6/Uz5uwi4u
R0wWHGYJYNUwTudI7rhGsfPXzozNJEoaqzOaecQ6PxsxGKiqZ99cM0Py0N+HP1Dp
bRHVKs7LCjeGI7xJXoiAhMg+w+N0p2hUsBNMc6qtQeOHvArkvIiVKy3rggQ8iIMU
Houw1lCAx20K8PyZNQ6SnZVZSrEhwiLXiQItS/uHWp310/FxCZA9Q94BJWMCQHb8
fUbH0LlZ/KiCB1PcOSS4PqcJd0YtMLgOMescTyCJp+rCvcWcTBnI/ZrUOqFBeZP5
UMIh3GkXBw8Ki6hCxwrDfj0f81mEClUtCqFzH6LbmS9/sR3jg4bs/DZJGmNCNn3S
tNOAebkuZlOt7Yn+BfcerqlZNPMdMcLJDw6fBBR3HmMXBO2siAMmG3Y1vmO1+2Zw
uTVAwwETXfrEfoUjQkmCQnzuMUSRpXZ1Haey7sF3bLfC948Jd1OzDUh5foYMAvC9
7I0Pm9UktgVxfFb0nLAfKhqlaQVaiT6dzINzef3ToQAzMb2PbG0g1gzjq/j0j/ho
CSBjep/FZpuLWbgLueHzeGpFJSX2TC9tnD0T9PXoPlORl+vdzUZKgBbwg6HVw+Lf
UzzA1JZ5lF66sacdiLfXe71QqtNga3qK/3tp5va7uksZPVKBRK+LTo1LSRxv8+Xc
MDmgvcpzm0Fh2Obsgw5XA6Er8Cw/0soYVLGiX9+XQWeXnxzMR+t8DHIAUqOft2Ea
uLA7ze3Ud0qJ7pb5EgElPYgqpmWME7MrW8dmQvUTJSKAcs+chubb+XRl5q7CM0Bn
lkEcMlgl04pCCTef+v4bQNiaS+eexx/7ookCgBpBxAtuvay8uFX7D6kcsC/PMHIv
WZcl1Yf6IzLPUnKyzEZEMb8fD1b8e2Arj0/RcYIDtC9DQRK4SWay+H+2dMs8sBjJ
5WOtioTxv6SZR2xLgl853jbIxAYq6XZp1oA6SiZ+HsD52ddP21UlceOvxfNtaBeW
MI9MKb63zy5+R5JPwM8S8OxO6dXd3U/o87KVV6NIzZxgTyNLoad6spybgBna8FU0
JA068KSz5LWXQdbYL8moCrHMEkgEDLTAszr46Gb4fGtnhIpwA41ZzjLHG7ZiZ6bI
Nlmm+8BdVRFIDxfd0z2mh3nrb9QPJi/KxnW7joEPrO+MDeqJ63Jam/zJM0PQlCPx
Br42MahyIMJLAARAHyewtFHM3KS90y/DXL00SsYvZsD5eY2bBbZ0fsP6R1/FdD6p
M0J+xqHKxRitXuXSulL11SbZNG0Zhk4Ix7gPITej5TBqdjhJGwpkG8bh6SsDNHvc
39goKQ/lve/a23pwKaWW7DVziQPz6gBqdK+YiZ5YCBFLoD5D+YCPwua4v+KbGLln
+BJ/WqEbeJkr7JzgV9RBSyOSoRPvzOcsZQednHdY7F1Xg1U2/fkaoWE2iJxUs/eq
gDb37bDrRcxqo3eRCO7vtXtDIlIwevC9txnhWXL9jzKt8jB0gYJ4g6lEzZqmho4h
St+hUXqNrHj+TmqB9h9RQympBYyVvZWe8FNH/CQ0iPTKV10Sm6PSsa+gL8o4wZQb
MGWNQIHmII0EwudwyJJS8T31sPiD4WBUIv9MEMLnwr08Px/ADI0dZBHXkuEoaKHb
Pz6ssovtFTI9H3hRHGuZ4+9KTGrObh/VTDyehcLVJXLNL91q/Fy65GZSwP5TWz+s
f0pWBv4TR7RkHrum9ouagMEGawPkzVVZUoaPm3pnclVfZ1VcjHkz+CvbkrqtBbX8
zDEkks4vvlS7zeBhzUul17tyWqacbPQ6zb1mtgRWN8qSdYtDTYRPqiK3hkb4Ywa/
zTNLlE4w0qaIjBE7DRKkk6EpZGaAVz4tWdJJUcyBFiHJnzDGXKilzjReen0Grqkt
tGmOW7H3MdlMJhk/c/NFTR40VqJ6zrHgxcc35r4KQ5bbDa/a8bGJLv6pumVShc+C
azA8YJwtf5FzA9wnbwMA0vWumfusb1HWjqoh0YxM5c8wZFksqSJ0qlJbcEQU1vdA
FslE0++W+/ha1UWsLhk7O2KCDDiHHhA1FnBSjR8SSBAxtyeyTyvXHvG8V8M1zW9E
ew4ulsao9EiyIG2sBt2BMtJjh+SZmJNEGqCJVW32hjvxXlz3dILoKNC/b93pCGhF
AnZwph4bIjoBb1Au9L7d+2A6RsJ/NXhWJcuJfP5w3NGAI5+37iUD/8FzGXEoKa9H
JCe6SxNYaROIO/ZWTdKa/8Er/ur/MnVffgPAEWhX5Q4qOb6gBpuksqLvq6CBqsoL
9Xv7IoXCHAH3NlpTgdJ9ZB+NVz37eTD0kwakMAbBJzs+YLQC60w1016J32BeV1rg
mIiBWqe+snGHJnxR/Cf0KNOy7u23Lo036wtYUrwfINGwD/hVl8cuMGMJdKdbzRwA
3taCB+WA64OrtIFBTraw/gDSacIKCVHqsXUjCwbmBgLziCUVbTzGX2R0svr6T3QE
xLkMKH0Dyt5t/0aZPQ+9eRg6DuWg7la7SaClb2AP7vjB1Lsq4AonJG7aChTrl/VO
K+pecjZgorwJuFw3N7aMN3WdLEBZO6FJp+g4KTDowfhYtiJxuBi3qXuI1V/BvE5b
rzfMrqvBLbdwIFg++ylwBUdkycGFq8Z66wgy+mmTUcVH3QQGQReLPMOOfL2oVaDt
uhYTLSRTjWl8A1xd+8leivak5pu4UVMX5jkmLCb7aVWGVVbVV5YXbnwCCGfAcnbI
EMcMPKKZKtQ2v3gIPEFokAcjNoazzO+UVmI+lLmQ01wl5sSv/9CNSTbZ5Oczn4lF
nqZhBCJwLWfReOGtwPOB5ug6Io5rR6AIl5HYeuDC7TQ0IvxbrstTGxuTL97MgoS7
aDy6tJZoViNFh7kGPEeBFK5EJf3K9FQwU9EWofjeDHmCZqzt+fVIOfX1VWFUKE6y
j3iyJ7LNfMvsGQR4hNQIv+6gc2zBVdvj6rFQpr0XVri5zGFMNIWxiyDA0dBv9kcu
7dB0s/YHrMWnsH6XjEO/Md+ArP++523ZBDR86iRvIa1AIDdDe7pedEVwqf7fpEwS
CsFw6k14oLysz+1UT3w/Sbs8JdVperVP4lEgmk/jRZdoLahB563sEkQ1yjnOaTDf
j20V1UqOS544sbGAlnw/H8ziGyPfE45EjWNQhOuDQLYomSMptJ9jB0PTrdDUtYJK
eOJXKvKPtZC/TaN2ddv9k39ahTGFaegbR5VZG4YH3HMYpoLhhZlQbppqHAbxVcop
GTxnUAyCDEgEr5IWkFixRB1BmJWOYhGtKqajzCdfoEeCuQ3hVTcV7Nkew78c3CSk
iV3p2fYbl0BE4DFL0s4d5H99uz8TTjm3PJvDRJbdvj7ruIxvhKcAVxIjUZ9AMuLi
Dfq908RXNblM+7V8h+YISG97SVOwBVYinsFAtbA/7zgDk1XgiqQsRGXvvhC02utG
Pyy+6YK3L/mj6xvo+/cKliw/csK3sXw70arVY0oOVz9VmC63M5K65sP//SajgpEC
wQKqopTPwNFbWnAZkk1cNemQkHKdCf43vipnTnDWUnTIyfyTFiCM4VAIVFB/z97R
OcDgN7tCKngP29psXEv8gUlfAnZjPoLulwG5r6sTSJu71um+kbY6nTFUT7Lg26ub
m7vjXzXD31ViF1uMvJHH//S5VeKnomnhIUZ7KnJ1DI2tDWlftzUzVHIKJN29R3Xa
s8S1e0aAnPWSjwtuil4YmAiUJCfhZHzE3khnYFufhhjqSRQI9NFDIAP16O86Gpzq
J15YjX34nirFOM5MpFWEmRumYGxSx/s/93sfz6fsv/+kM2qamHcq39LBIGeMx4dp
bChEQq/XW+P286xQ4Fx1QWAzuzssJa+fb9s4U/wgfLiHij/HigtNSe5/cC6K9U6v
97Y8/HPfXqfmcB/SZ5cuJ22LXJZNRzSNKrQxLvpDJyyUjzxchxfPkQYji+ydkDP8
iZ2FmHpEmKeg9EZit7YaLznYxWEtfdHBXQUaQdPORI5bxJ3pZL/uKi0QhHuBVRsv
xfc+RYRgb9x3EnrvB/gRj8+Fq5K6BEZiy2LDGfPo2v44K9/Y+A/NQWWUyz30djXl
xVbCNHutXUIjd5tGRmp79VW63opaCbnhOWRNrj2TyBbLZ/KJEudcZyK8uk4K/6fB
zkzQL2JsnfZpNjXyeifNCl8GcQZryNgwG1Kfp05MzsB8dLWsFWEJaaiXuy2xQa2L
4EJM2WDgaGtudLUQbN+tHrRWcUqyYCm5OJq5JYBgJ1CAFdvzmNBVpIZLmGlYdibv
Py4KEJ3PuhBAh4qGt7xJbQFqOyAsSZRX7tqcD9Bj418VdEERMWI18Aq2XVnnUvV8
KBgdP4dluZ5wlJTVxzGDkyjxuZUAez1PkU6ojSvwJoMiyJBTqRGBiiY3pBaTvu6c
8RaHfy6pUxBbeduYrGrMF3lpc5JFS7GkLBn5NLnP6Kjt7Zp6rdL4AQyVXunx3LIv
hhkY6tIJcYOfGuztH6RYSAIHqmOwJbInL7rCFpXjxzlLa69owQj6NM6S8+Cqhq2A
jyYSPh0SyVi1lnApAsUIepGdm8kkrOLcxgQDpl4d1rdoQoriFvVv3wQUpw/OkJQC
ItW/N0sUQHtnwM/KTBRG6nCV58MuvR0CkQF/elpIRnLsbO0KF8bP6iH8r5vus7ML
+YhMfRTJWANEjZAii99JsRFzSw/ixzbvi4498BJh5Gzu9+Kmii5GEMEspykWzVmF
8lM7cq2gOrQXJdHC2u10DNaqMiqg/AnbPik9F+xYtjB+ED1EN/8Amd1TQwcLaBWh
BfItERTbgSaF/vAorLiMbsoihCtjjsxYSGE95LT4nVXYoX5PhH5I0Axn6uUZ1bhz
79D48rW0tEdebNPoWNY3L9ON2hkPyRfqhprhisb8zZj76utWWsX/uhV+S0lddPxh
UJVq4RQwHE3Q6wwB6rH6RAe+t5F/jimhA9D/owxPCq1brl0JDF9C0JRMru+B1n83
9ymF2s661J8r5vo3AL4XMtfdF8RtNosgxdTyHIJbrtx7bt4N5qhQWe5piHnQ9B5D
JV7WnNqK3KW3irSBBrsxBt2p7In8sabNb9inQF9J1cYqUzfOAoF5aCl9p3NJXFn8
ePh5wkdU7ZNezum/RtZNGb5iC4lacxhbnfDAxHT66s0BxPsiSrGhmK95lEbVnzUQ
iGC4OoqZDWPrQSiybLjbaoLwiLoVDsDtTsizbPH6dwV3nIQ2MTpuuxXaHU5bEaId
KWtbboS9RZYKq+QPm3+BRBcJ7ZVJI+nBSg+OErG5Kfzyu8gTzlg86avXAOcrywEU
QusDvWUoddifYgyTQpvE9HpgVV0v3XMP9Nz5Vz7OeZ3GRwOxsZKOkAuwL8GOPdnm
vhHA0Y3PqScfZjfGiPFwbVIU+9kgFsznp2b1rO8uPFOGJT3YWCtIZphRSjNHfsHU
COyjow+n58MrD4Zwyv6jsDtAMWvBxFArUkcqcuZmEucx/vkTeb18PZzz7AjwAqps
+9Ti9hviFckRwXWqbV6dyLWr1+JHjrCkDij+dKT4ppBi7vAHxyIhX20BwrFT2eiM
hSALzZrMOSnhqiseoFM1pmJ6SUCQPb0HexOm3+CwSG41Oz4qDtzM29EpGlZAp5TR
tItBtw/qFy0gbI4DwUzHVZmQIcrX1ksroRx8m9fI2A0czWXTed3lImcKs+nbeKdZ
giWkh0lfW/OroBhXL27jmIskXBHUZMxCBvBC/dCjBkOjcFXNeBN9QxVpiekikchz
fLgJWa9x3UE/ww5GnhiLImeNeRrfF3SyRmbchi9XlenuVLpvnyzF800mGAPIyL8o
Sc2aEPK16JuBkcSv+vUwGhMO/efhZR4GKMExerO56lZDaYbI24pUbkifxioYPB+X
BQuU/rufNqDesnCiOvN3DNnZYPcvaXcfApdrryhPSP7MB4KmMALUG3+Ab/GMWJC5
JzJ3ckdZ2u/x1iySfr3btuXmy/7Mj+RqAG2x8Jq6NQcfNyU9QQU9OM30SvmBoVHV
QnkA1xdHxAhLG7hsZYEm4VIe/iWKdKTCf3MyAMypaShN5+GYDtJnjHN+3FNaj66E
wzPdxbOKG9EnB5tQxnsgLF6Ys6JUwPyDlF1Jkjcjge1tuXNtQmSP3VJ+OVH53Aa8
UPRh4EZN2wKTEQOuHXsg0PWclghYy4cSH59OwaEa1RLbJIEUdoocUen4lGg15b5G
fNIbs2iZ0CriZu8odVrIcCaI06itDbsJ0+ENqMBg01arpnsahPJ4BF0SXB9W8+6+
hbZRfDV7za90VsHktlN9lF9jSp0BUIZsPZofNdG39iWJslFB3VQR9K2DBEMEvlA7
f6eblC2BtRg4ar/6jyUeXq30hR1Jd6vXEUJzKKREyUDMAUbyNU+ki9Yn21Lekda2
fc9+zAu2eCREB6KLgM/8i7rhTN3bBqcIpeT3PnW0U79K1FKFiwPURKFYoZNoMHcB
HtCMGuAPY9b/aLNJhaYTxbR+CW9GOpugvkCAwWa5epCOqNAro7bgC1zyeaqhduo9
07zTI3cdje3HB2TzgQCtZG+SjU615aYo88RKZcfE4HH+j+9v8DOir8FmTRK5y4g5
ENks3iEhQVADl2nnvBkQTbQUkUi9ht9+ZChvd77qHkAc+xOoY87cYmVpQGqJWQZD
w6+x3O/k/wA1UZenpLwNEiSd9KTGguHZa46V361nyK+/yk2MH3mcDv8RlmmFViXD
1j52RuUrehN43bAOLt+9bClTckp1eb5nmt8R0FyVYISWk2OkgYK3wD2lRLpWDyvC
meQV+7YWS2vNFm2jFZD1Jtg+LmvSUFx0h3nZ5Z56+RojCBJpavIj5hD0XtVk8G6O
7PPGaduoe9sm1qcuptmnqYD3UDhrgAzSnMfJCyeDiCYSFwO6bMVWhvoFHeNVmPIT
W5VU2a5G0LOl1yS8iiL3ZRGsxuIocno2atRZepgHK8dQaDktSSEWgBy5QEgNlRPv
gj8HbXaMRfSSOUPo2u1VfHI6h/od+XRbAFMlm1fHEfLG+xDtpOU28R3g3kdH5W8Y
7nmMbq3jSZJqZ9dZcNf2JLZiLQK/f4KLbzb1NpS6/gXW1lUsCrS14QSfcUupdhsS
W/QpJBcRAMvRjxpqcVc+KBXS/K8gYGl3PyfZnyK4rZNAAmeWGCUxfF4xSpLA/Ram
oO5g669nmOLsdEJx9B0NryCiQ0R6YZjjFL+lSSv+xQMG0kC3NuSXgsrk0sKpcxQc
oKuDFQHNj1wGqquRiHddbFC2onmyRxwLlazr4ALEkggVg4r478MgiBxp45lRSU+h
34Vxeu9BlT2df51sFGcKnXpYHJNfuNXwp0JIQjuU9FipTcwZqhkG7Jebxofp99cA
pNjxlHHAhs5zL204gvuz+ONZd9XlCJBhaczomYw94eADnSkW3i3D3z0avq81wyQS
xtwqdzd51wW8y+5SJHKlRzw0tfUg1GPoNM3PKDfxhPk053ypTCkM7m/tKtvmF2qi
LumEupRtZakOOaQcoye0UN/3oFpX/JNWAYR0DKkeI+f2JZ+fdLz1Owgvk/jS2ug6
59mDHaOx+X6r6qK3Q2+TEJiTLukcJ5+X6jbFpiG8JEmkFAzgn31oTpzGaSGdJj8y
vQBckqWR11gIgycC5wv3Y7R6ggVEgKqe5xu+ki+lbOUZNkXtF6drm23SY4XTdTpc
KW6+jWbX25f2nUAFsfFJ0VFvhJbTwXXs5VNkKAqh+m8wFDAIp3TSEC1AuAzjsulE
LPwx2eYY87RaLxRAtO4cbE6aaBqLDa2q7Pi5S3UDbpDPnYU8GUXZYjd7af+Ef/ng
bzpzzdHaYn21n2ZgibQ1KsDYwD7i4otpkcV0JjCb22Wy54cLI6o+cIUB2veM8kV+
qMu21Vtqm2mfK8WLffWjZEKBR8l+spCbWJ/eSGF12gkN1i7XkYV+jROPcfO4OxXB
5KCKp2xPq1kzBk+ggjlwHsKYsGDa0R9vR5ltcvjem+1lAzC5S7nt5/qNN6X9Hlxn
wMnST+SXup/WpI5Rbn+URAQ7KPCvnlyD6pG74052Qtw+t8TFGnEHZSsd5sJpbqX0
YiCpU4azx0cpkrLYYXNW6uoYX5GxqIc2B5MUlDskN98mWtu+mcrvJZVHHiTLuoxx
YVopbAhHjZVCzAlN4OkrG+UYnaWQ/WV3cvISEJwfudNJNaE3WjVZ7k3VDMm52OUy
YFfdyjisRhP6eIDl7yS6flKl1UDY19Q9YENSwxa9IUQRNWUpG2osjtJOz9Ktri+s
n/gI00Anf+1YgtZ7DBDWYXCdZYDhSVYVRRqSIu9RjrAfgKuvmXtY3w7usFpHHtPJ
Jmi+B/pA9PqUa8QGgW+gT1F4H58xSmBgmvNOUe8QySOJ1sO8o2YIva7tFD1sSu5e
Yk2ecJyNMw+OdUeA0/gZZ2asXsTuIQ8fPvKqbfyT8OaR+kYdHeN3kpqWVaHyxQwh
qIBwqPJoa+POViy8x8dBrGLtJQUqppej2oDSZCNgK6kUWXXNMvV9ljuIb2ZsxG6Z
VpHxRP8n8+tRl9Z6d0kQqLbwUNTjceWN7OV6TiHKjgZSqgYtJLkBaIOnztAyr6sD
K/RGP1MowK/O+MbHRUIVTzhQJLkVIqyeIE6ckj8uaIsBAidIPGl1f/AiHFR0bKeM
KClEPVYMQmrjoYKw4PgSpT3L0FjB9ia/5y6jwIx7gKa4MiQf63Kms1FOgvqspvDq
G7kcEpSQYIcgkRWKgirV4CvuV5o1PT4/CgZ4a82oA81zZJRJwNrSbywTWQoqPgw+
ghxsIB2HCGpYTMg+vrbZ4Cc0l4R7a+hAZ+EBtn0MZEgGZ3Y802ZUIWVmJbYVlTU0
t5LYHw6gzpZNxv7YTMBaAE2JZHuIIvg70VrFE1EEzXZG9/NcyeTQyFr4BHaBKDT6
6NIp8GnCGgSlyVTBH8pw2wER1NIJBwTgInkqKBqVOC8d+DqYYg3gpqhv943gw8FV
wZPjllmY8Lea9uUBVecihDG3LszzY3kreD/zE2x2abhPCHQkrKIJ3UOOrClDnMZE
gU9KoWUAu6wTTdq4jZ/F0bckMbEFXJ8aLn25bF5qxOHP+xzX4uZF7Mv6IAShj9c5
W3frm9O6rsMmB75WOT934pRdwJn0FUStFQBqZ6p2Fo/wa3tMMnQcfdtR4OrX1ZKm
ezRnDLAFm9IYOxOG5bBowmOKSWbHWctrII92m6dd0snrMfGiyPoQgTiJMT2Ie4A7
w4YrDXgaQG0ebMPSfaKBLHSO7tzgF3AfMOhwxjeZ4FovVWNCA2bPZcvC5j6M9/vV
ReKsXkhz2rlZjv5cC/oQKsI62xeV0QPo5dGq35MdEobVvVlKZ4X+zOg4QWInr37G
Ru73uDAOsNRkZ5zm0cKB0QKypLwCWwqmNsb2e4k6uw72Z13BXwiEH2uQHe+HQZeM
UTePNrWNIgd++uF4K8fdu+3uy0kE0vfllNxBKHxmAmM30H/3Bw6WMag0ng7Y5dfZ
1Bqgo6X4avGFG6MT1ER20Vp3dSbveb14Fg3H+bSOCQXe4JEYl7NmYRIL3iSsWawv
UENfQel01890NalQtq+9MamSG3eTDEBmO1XPNT8iPkBIn2P+4KlZ5J8QZHy/Nl+a
uPfTpAjYtOKZ/kne3PCV6TkLic7+HM/rdOVOnUHsXDoVwm7uP4I5bYa9ArXbOuEW
UBgJfA6h+fBf3Opq3/ENlTvEFQLn/l4UM4ZgS9TU6Eao01R6jU0Uw6aUERta7fZt
rGl5ff04Gbj4T/iYwWhFnLOWQWpVgE7/zp1VsBtMJjqKSF8Bhpexua4A982ay5x+
idGMFscpXVIwrqnct4OWFE4/pH79/FNxJzSUp3ICtnp3wOmfMJPbFocG4p3e4Q7s
9jtUp/zLq+egUIU4+ZIWzsdVHFOkaveUOhUSZ4d4SA3/UWYCh51/1Ko9IIcOpku6
9RFnNerj5/LyL2h6HmVcvhO/FokbI2ydxL9j4S0ngYmrbUwarhXkN+V8kd+N+mMl
1SPhLT9RRON9EyLfKlBfpm800zmREYM+OFLGeiobqNNMLjiHmSYTXQz1I1yFTRpc
GMkRbxdHtv4lAeBe1NwjrZ5nA/NlNPeFfDvBHdahXgnAOtXYjKF7qrkijNgQ6apH
p5ign0ALgr1doJATfPMlREPzmcEb2hTwRuquOJfgIqpiG8thTfiz5y+edV+goBrh
qCl8Q2lS/XhbUf+rVdQhhPxtRX+3IUfaBHeKOFapl/TO9q9tq/GMMoTu/SXVqFGV
xz4mF548qIYLVCVUU33M2ETthJmWwat2NU4PdtvIodafSBlW8emSZevZv4ZkP7Pf
pzXgXEmqLeAfDkrpl9VZQo31wUvwdJN6TmaMzgNqYnuXULqfKf95VfCAJ9V/gXzM
EdLFjq6FLzkUfC1f6K4oSBdaEYAOq8HE0Q3V1au/2cRzsE2fEFbDvZl6skkKZZLb
RalMtNHRTfLClUMvbx/yenvMXMQu+pbiRoMFU/5Trokf2HHwlVdgbOlm5g/pds/R
mj0FqKbRjwrylyvCV2rQyxfQ9NK1EM/wFA2SEx4+LvmyzCW3hJLm0To9cw1AFDvJ
uMWRQiMaz1nVSV/dcoNFtyt9AiDGse30VeZz7r8uDf72EkoTBVKPWnYQ0Wx+AoKo
k87DKPSbkNqjyyl6cBqYSxT52skec4AScFDBrtu5PwV4ZwddFLQJ3M+Ut835VYwc
slA0qeotHn46pBqObVqJnBEg0P6ZE+YReiiRKwzL5jM7Ym5A0Lp3tbo33SyI5lAE
cAyNoTmI8KUQYZWhcW+o4fa+3oqt/ECxuKmyrLtoxtyBoyuX6Jt2l4m7623R0Q55
yiL/jlbH9bM5T9NgI1DSpuyCutSyJ+jGhHwWlNh0Lx5D9qErsVwNb2EWcyr2JKLP
pzajWXClNWOz6j4mmAT69tALMRYkfho0fBlpxNWjcq0N3MrEh49+ejSOgx+VkJ0U
dekPwcS3PfRwyIYF2yJwUuO5nKkwm6itd/5OifoDYbsy+78Er9DK1hSZ+LY3o/p1
6V257zEmG8rKt+9OlAqVuTE3ySnCckoCPY+Uk+rA1EVZioFP5SCHJ16kPF9/KhQT
FPmjV5ds+o+UsnsyantBtWCzV+QXs/B+WlRdxBrMPVbo8eePOR9U9dpB+UsycpnR
Rfv4/pYG/orhY1OkEim3/pvzOn+WhN+TD+8mTOFTIzcJvi8JIw2z/2a2FZRtexzM
bWTbH159QqW1hG6y8PyLXS2C1LdiPob0wfHBwjBUPgDseSZm+SLQEfeHVbMNFfR3
ue3DwlcIGc+5KHNktaSUMmhWs1pKiNHsAQf3EgGQAVkTqoCuEAga9W1KDsk6vyLv
Az5Th51PC9A6Bj4R6P/+ThzQGKdjYsBV5R2VM20l1mRm7gbet9HuzXI3/cHGZxQm
QPZBreXxV+jnWoHgbbDMBIoNj1NRi57dMz3BSBpERT1dAVNeKK3QH3A+0ABptnc3
JsuqXddwEu5YB4Pt+pGr/gek9lQvG07g25Lowz0SM1jCwObTIdSfcLXvQtZYcLMB
pamD0jAQiHJK7m0MOQh+6HaRgnwydN2o7uf3X50eE469XO/NHWuBnyl/nKod0UkC
sl17QLOwU6mp1Lk3gS251cfPhMFD0Qa6T0GgDN5nTBPnSKcjwu5GJqbNWQnqFyhx
6rdHiOl6thAL6FvtpDPHAeyVqa9eDnUwmF6pxviF0MOb5Ya8P+N3fu522GtYJWz3
2GuxXgnYNaTffXki9VM2jycI8OT4YfUB3+plVJtsfngV8Qeleuf8EkpbDOBSBKUW
euuoLFjPcoqVdLlBH/URFhIA83nrh/+bG4qS1vNT/xSQeUmlZorOcZ8y0YLmiqgg
7Ia0yLmfswhemBQnhdO8jzobsCkZYR9MZvHZdIMpVecUUI78G3VfiTV4BRAqn8UM
fvRnRYTBuKWsfjbi9TyITbTj2steHOpB31nzKWVFRrKqTlmuXSKhT+8EfH90bLfV
dqzbQswdIE4ISzxZ4umKXnHHP+fcnpDJ/Hyd4nNBjD0Me1hGE7agJbkuLT0O3gzo
+jAVmn7z6/Lwx+noKJUfkTCKa7pPiINb4xvxhTWKQSilWv9teFEwHlnR1m/UWWNJ
+u0hTmLe91nutErFBiVnbSPk7RT8h9C9j7K87mRWMC/fwWnOAJIGdWqDnhYvcg74
LdmUMF3mRIMDYic7ZyRvAqQFH/gmXpMdj1iHlzKbU48lTwngUnyNZHEnYeNlwOgj
8j4rTNPJ+a0fM9/Fs7hIBNe5Tf1uWl63M3MRYeG096XoRarc/RvxvY7NSwcnAqI4
7XpYeY+xiWhqyeutOCG+etOlLlcC6t7khed/XExXCX2OO6J4oTDGRwZQybssKl1u
ax8SdRVf3bF2HvrUu+iFBvcQjMHV+yV2oQHATm8CDl/kcY0mctl5ybjd4IFtRgbW
4s+OmaM3YoM30dHk4FxEYRiG2Q6levtQDZ7ibYZGNB/N1MXVQmBCern0J9bCTSAT
7przEKRo7RCtItx8NUG0fXi2WTxBEwcMxLocXCYRw98Xew+ftaB9D2rF4R4ooAcz
84k4AbZaM0YVHKVXj3jEWTVP1Y0SGPxpfr2LKvzdv7CEVdRAPNk8uHPYGe1Q/r9s
uFVtB1aG1VWDxI4dz08kN/M+JPEQznjY0yLPS4sdnCeFIE6ifseMxVvJNJ3lKiba
/TD9FefP+eTiqLVYEOcOal6P9eXC9fBKyvCwxBXm64qq4AxzIIdCB1fqozoNkznj
Uabpy4X6Z4U9+WL7V8aGn64IpWBrDhA6jBzkXqYUkTB9CYg/m8oBhxtUDuwlDUOs
LwOLx53nvMiHAUgufL5uzJMgTMGzhEjBIlV0OzBGDvJtCTV/xzI9HnuiLTGByymw
ygwHKHiDGdNoRq3T5ylGHPJo43PjYRigF/sRZ65yddWocTlEhM7sRq2TayHI1sol
j7uaIOoStkiNIS5AqvPWT0uvL2qyQ55ed95Hj1mSXCPSqiwJ3q13RSOLvzGamgLF
wit/zxnhdSTudW0ZXs+LfwPIg+KXK842JxnrtRU7pUTMzcyefCreYDgFUZci7vSP
y5BMDv02LMJFhC9ZDOWyuwwZVrajskVQyLJ8yazoBeNKQh/z8CPRqFMZlxx40g1R
Kb04XnDv7GybM+osqHnD74z+zjTqeRON/J0jiLh64MVUN/izNdOaF8RKaljFSylH
3agPc/dBw77d8IfTyYk38e28C7jVGkxfvaT4RtueZP/86I6SBYrdNZ/owO2Kla8E
yA4KR2nRSjl8fhaX6HfvG54gaYNjhUUaVlVE0UAA1v0hDnEKWBQhLvk+XhTExVrF
Lrf4rg36R16kisy9NjoTRd1BxjmAOPljSfEjCEU6uh3dT41E23wdJoWHtRS/0BNq
nkDJfUT583nbQnM1J0a/9BWFm6tJJYWK0PBmDUnAFEE4jLpAmSi8kO+61HpiP3NH
CYimMBPhE3A3x/AyL/typwTPgP0J0rPxW8ITkqvKeopa1A5tvIb+DBhxtloKoHkx
ZGcO5WFitWeDwJ+Z0aVtsftPR9lUMCuek3CsP5oftA0y2DjtYD+aW6KLY/JNDiVe
IYzoKZFKk/+DczRss02GGWb3N2fz4GOhfuD5+4XGw36pno/UU7kAKZO4Ucvmfkw0
vCwLQLbSYaZ8n7QKmlBYI6dTEzLjlIJpJ4fuLtD24iF1+W1TgHuU4L6c/F5wbkpD
z2z90xV2GvpvRWW5oVdIKJgrcz7eTwrs5ym5OuAoJLVRhBI0BCyPRnB6MBEtd35h
UJT+LwzFxAVASBNodlqcpRiIK58mtcp056X8UHC7PfPVVailvFHRbMqdQc17wMwr
5PkRbhjdpHObUSWhtq0wx63Q2E+RiB7zQtj+sSasDZt/M4xFoLCcjEnAExwZexKW
BPvX+IlV0lmNjie3ulTIgr23yDaW1TPC2eyFqLQPFO2eJGgAJABUwOy1bFVQHNJR
jvSGmUYSIKtAQuUd1oEK6JOj89SQin6kear3KkqYXNmY3dw4HnYqYC4lWRdkpbnX
0uRT6TrPcbRWFP1cJQKAyRr/08xpxXuU0va8ZgR532xiOhPfBP+EtuGnRT/TaKWP
OBIeWDBLKZQ8RK3vjTxszB4TVzFHe41PD6SNqKxV4g7ZlbJLFvXriVhP5ibATn4V
Ii1g+eyjwmHdvvum67FE7u9Njts+SMmvR/C8i8BoOsSdAR14MMpUZcvM1Ztj9FlR
NCUYwEsP0+oQ1eYinMarLouQNNxpa5JSk1wGCM6LnMqHIB0+4bXmC0RcX+O/Hzqy
tfq+oTUI5Sd3jYBP+zcEFlzbB2OjfcmH9BmljExylXgxLWctlcCSHEtT+sgQotbK
6weE8/ro3r8ljL1r+ZYB0b11mBxyFHHWGL8Hjv0NmHO6xK6WypS5WxZ2UlNN7LIH
cqVIqeMQGidtpZyLzlRJJ/azwCCer8b2L7eJzVnXJk/sD+bnh0NfDwVPHD8OAVLQ
PF0aFfcHkZaCs0muE9yvFwJ5sWGqpeKOpx1Rk7p7AZAUNSXhmAr2pysF+anlW+VA
QMwfBAaiyCAPS5nWpgVMWSEFlME0eugicDF86DImECzmGA9vKnRQUwEmdiogdh/n
MdyrYpFrqgU1klkCsveiz5ptH3YOip4+gNc7sirpeHpgrB8vIQ/yKJXXWGeghCCM
Jasz2R1IUXeNlFJT5VSmkgGsDHrSQOhxS3kQ4438ehUOJihfsSi2WTgYYBXthoWD
f0MHCI0Z5yYLlF0U9a5FWYuo5JRz5Ax5uygGtHhnttjsRLX6pGot40oniD6o6Ivk
M9xFe0A7WKPgnKy5aKhXgNLeatPJ7eeHLq6DF2xpiuVcQqtd8HpaLgiwplHwqrVZ
LGV19aqsN2a+RpULNWHx8JMNYOthErSWoOelcyI0dBcpYk/7D2yzlF4/VZdukdxr
BktJQ6DXfJeZ4xQDwNln9eAUaPf2GJ4W01HLtA0OFND+TTuIqFCehZnFDc6NdBW7
jNOMSNjI9UbsPF8A1ZjnuheLCzgDZTahXRl/nBXl+7VQQw+mli8Qf3ecdTrIVG5n
/12CA7ppYzBaWaPDW1XD88cssBXt4e7hRoZipRLAzDuRIf9PsFgI0buvO4FPeUD/
d/Hk+pzD4xWrboPQJBJ6thC0K2t8gVBrFdhAGyTDCiS+3OxxCFRyuyGu33NWyumG
zG6qxNziSIw0QOiS2om15WLYjbuNU35PCbZC5lR17KAcZaNFUbDZgSm0X5J40RU1
rwuoZJJU//8Vv+e/0m2OeI1F2QXxw8xQKwpue9YZFkcET8JNero4TUesKky5o4f+
IPY+Y2Ggua/GWFwTBwTk+XsPDEYV43RWP+ZRR95DR0D7vuzQ5dnnyoddK+VnPqtw
QLWbeffQDF3l3GlW06YqD72insjM9cZLF/ZsXEmcFZJ1Bpu3qFQ60R0045PSC+fW
IGJZP9coNS636UzVcX2bOGUBOavXwx6UAt9lMMyeisMUa2/0IqD64wAZBMkamuns
oKqJ+AO3rLoU1fefAlMf0y4s59cliB44bnSSAmZhYjkHZ2x9Ry2k9t8AexgInk9v
tBGCUOj7Z4LnoBYMKBQUgD1zKUu7LF4dTAldmsnUx473TbcGK3t8zIQVAacmDcez
c+n7mTw34HwVVFy5jIheIMIkx2zoZ5wwetZECIxXwKctElBGjbFG14WwtBx/G9FU
YsgYH2/KaHi0p+4xC7EKVSFXUbZSMHyUU5ZvdzlWp/tdZ07SA3UMk53NuE7zueuP
Cu1LEGu9GpE2j8Ys/pGxFAZiUyaAZKLAnDnqWc1aOFp0gEW5cGp9cFUdZXXHT/Fc
TAQ/noNw+UVBJn/VAzFUb8h9xpjca37UXbqxEwg7DrFhT9NttfNl9AYIqulDJvB8
zDwIiC17d19tKFqBw3GX0HMFVpOIN5CGsxfo41uXP+EUU4MeKSjIxDgEXLkMFJvJ
UTHrVUp37oqoasP43AEHH/do+tijnX9I+/wIUJnEkGhMg3EjV/YTaXpsBLFbpAuV
OHuVmPpn3cbKyk2EXyjlnRo08EZ61/qPHZlyK2ACS3AL7UjbJGppfUUe72Z/yQcv
y4yJOb+FIjsmD9t1I9AFLZ424AvRu233xg0eUd4ZpqGwknGdKjB0U4/BH1i7B5oB
wwMxY9O557ICeP1iJRcisLmvCZkBT6CZGwUbFXixYxtTKkKitrG9SnTAYAfoGG8S
eiLO5hwBFnLAFc9F97AcYH8e6t/PDle/3AA4QDuNp8CjGfaXNNr6XUIu3aLWIHk4
83aZridog3qXNtVNySxu0vppnqPjdSYPhCZu9AXhEOw6+m2qX2R2sB+0dm9w4DV8
KPXMGm/NhT+HZsYV5xNEpLZPR1M6GraRevMz+wAhK5Ew8ABCHDCpmbylg20w4Bb+
+m1C9SIk4xotbgIR+gIIbzdul2Pjvz3pg6RxTbE5mQmgdq1f1BmHXOV4kfr4C1G7
LTqLFA9jI36JWdxnI46Fl4NvIh71o9XUyhzuCNHhP0AtU3KD7+UMk/jxJpsPB/+k
ZDWvK8tTInVmdNfdDV/GdqYSzY9O8iNdYz5jRkQknd9ys62+xa2/3sEJs2HD6ShR
SbwIZ9Ht/1devfmiKyrC0iq/PsENvZH8dusRWtoujQg/I4dmRyJYCddhpOgVj9IO
M7aeb3fSBfREGFOw0OaMQbH7BwMrQtnNZ4DBgz565uAnvfZ1m7Ln7+vaV63h8WQZ
T3srK9qK9tE7YNcg/dlfXtc8ysJ7gnEnaA9kK+tUOvgAsNN3Uufyft7nwCQOOIh6
GmexVPoh7/VytoolSy+Ft60d2teJ/38hJYtzEKAvR3Uf86ujLFmOdJgbxVr8KJCL
qxzgM5FFdsTzoGIvQGCQUd8a8zO6PT8loaNXQw6YYh9qDkCwz+XkJr+SmK7CXcpJ
NOlJ4qT2tiUWNRxM/FlO0OV/YCTuTOCcmzJDdOQIQCTQ5HrVNBnXkAyxGdvESrEb
HD3UlKS4j8uq3pnvjqHAKTGcf+wm+o6vJLPYsCDmzVuZVdMV7NI+58l5MY1we7iP
KT0Y2FSwi4TARU33bdHWjZxDsHIh3JFEDGKV2XejfRsEtvdjyMHtyGjtWWXncCCH
3Piu4Kjnu9pEpKELRq+FD128Adz1EQaSTNdFiqFQYqptlm/eN3P0DUYrkkYjANCx
P0XJb8IELVf5ICBLzBHRi2+i5+6cqQXTORoh4mTP+zQuZwjyrpklEBUU1qlP+s+i
fCy0LPQgLh7BPJ1prG78kp7GJPTyMQwF+7ScV/Ww3px6vbwTz87PD/nkhM9Yg72S
oJp8JPoPn0q9ZWSFqJXSiNVdDuGPvtBn1wdjPLIMiqI5njLsDYjlp3UnEjpAiMQi
zlU+XKcJVjztnhpTZXN56KoJc2CWL/RpJm8Rvwt9/D1NlGrACynluqoBGt6febx6
k0oMgFEk+aRq7yCm/A4+8kgtRxfDTVYxc43rD3YXS+fo4SXdIHLulM5pxOup5Ars
nlMtXC0HSwdtho60zBjU/eQ70QhFvuot4lSQYtP1PxQraBg8g6ZwEaHc2Fwa3czm
YpcABvpk+7/Y/o/WDEPkPxitYeXzUyvUSqIlP6U200zqR4BHcUy/4hGnBoXxJF8G
w7Mt11LlZEMGIRcr/PBQCnPc4NG7bIhIm0wf116xpumAb8uvo+v+RYRsdEwYyUJa
WvEVBhJKD2Dts4ETswq3VtpGSfiqITFzXRyW3eoNKC4LERnRRx07KRmwy0ljf2d4
gzQ42O+/Q2jhcE3zCh117d79NHpc/lNsgQ3vxLbU0ek1gtE2zUKqSWzrm8Ku7ip/
baieDnBf4Woi9KcniK8sQf8TZmNCHiLHyHKKBoldE8zdEOQ1o2/nfmm5dC4kDXwX
B8eTPczAecWnPp4Dg977WzVc4Zs/P3HzVZ4+D/BVcd7nr9hseECfsRX+8k2dtUHC
WJZplK5zp9cWWtiV6ZxgLcpxoqqkMSPx9+J7vcrRU5cI+eKxYAYoBU8czRvyx06N
pCBOW/yxPrxLfC0tJUtAMW/Kov8T9kMMIFdCCM9h/r9/4Yo2SGe8uMzZdtDiR46J
04vqZzJcb+IxIfWOAZzI6MaerZ1FMVFEgEPmO4olLxpZrGNbhP4cunuJDX51jsfO
z9HSeS7Isc5crJ+7e1O6kSSrNmCpebPVd/LDv4upiQSjX4qymR6E+yEpuWU7/mQ9
BuJPOANOTusMpF04glqK6lrkDFMUtNLRi/yr8D48gFYsu5eumDJS7npA0MV7kTlF
PqP+yrZqblaWe5gGcG8iKNYb+jLlWPKHtn/t0vXHZ7jdopxsTssP5Onk9MjYo+pt
wqDS6GsVbXe3NSKkFcz+MORuTTTigynAoWun+K/HkmAx1gE8o4XbzqvpFlAzeGCH
olgJbuts3mUehzIKdBbNsLH12++JbMyMJ41vh8KWO2a9uzAyaZo0fXtJQgwkwfD2
JqWNUbopHrLsa/1bkeZijGSvjKDGpHwJJHCVBr7aQvag6fOdz3DrYjP3E6/iNK43
ZLDwQZNklA1X0w3wiWPo0kwhs5thsIEg/0ScMlmh0U382ILp+TTfwxV9VcvE3NtK
dSqdoy+5cnu6ODptRCouLJSNKTIXr/ShxZHGleWAuDaG/PEwuiZd8Xd13gHD9RMS
Mk720KG1NgXw6prqRFuGKy31hDjF7tsmNLVmJUxvA3HwZ1KBEJEVTgXkWb9YEvQi
bsqm8aKKtFmZHViZnyZ9DGfDVNe/iSiYoYM8J4sVhOAZWOcbdDrdQ2H6FLAPAetS
BHK0l102ux7Z/AAu1EpbA3DYNrORM/4Ma1ooNk5utukEGLJ0gAojWluqC0r4W7Fk
KWkPRlaPZKa7KEKjYMsJGSk2YUhoPy2mKobMjS+uMQ93KsIfsvufjbstoEUrjsBi
3dh6o0+yuxclMNznc2Qg7Ik1EjCNA5rxFxq+Fq2hjwv69bOT+rZDyrq1SXm+2Xo4
aW5E0Vmx37NLbdFxWni4Zz9TDxPA/P+IBPmAs8RJYcmxNtEsCFeaxCqd8QJq/+QT
xPzurKWo2opwd4PDd4+kxFkpS6M4wxuAmqMZpFCMvNwFVZQbxfm5UFZDrgC1pClO
TK/PHK72r+naMMw/4KWMquAT8LjALPCI06HecVuHXJgKor7VIyN8Rr5xHVBrMEo1
WK3yZFE4NcAcg2WyoMBaenuFKsQYlXUJpiBKXtQ9LnhdkEaUwyU4uCEoRaeblZD0
m7MeJa0pANiJwixQE6ac/562Rdo6bTVgHNki0wpPY6yP3Z8Iku3EIz3YZOgtlWGs
5pisVeSrfi9KL30m0JeHTDhpRc+zCng02Emh0T8g8sNcH1dGkIA8BUX+D/e8WAfS
zdMj2VZ3UrdXB6YYkl8Fww5s09rRCWvJ8X8/21svhbGgJuumaw0+qLEZpZUSUlUl
isPQBuiKe4LqRQXfo1wz38diPC5QgAPmIroLPNXa3RX72dKjTaMfj6UrVN5EU3+y
S+0e9HcejrNqS2PuPiUFSdCuQ4Jke1d6+qCs0Rlrh8a7NzfxmH4m6j+RDsDqPcHB
wG2O/bEoa3PhjgCD9ZXQCaRW4K7axIiIZV4YWpruJqjbAsRjIyrJJDPfY3d0FFbv
zheTrSTczdt0vJ5I8eFCIqHDlNK/f2cpInwa9HSvIogHx0WsAggr9ouQS8CrsXh7
rBLQACPN7sFk2yWPRtOH0kkz3S8JvZ0Sf9ZLEgg0IbrSfmIA+qaGfiz7ig5ZDXyJ
NkGDVkbpm6pga5+P2VdPzCwnztZC2tH5N4bjT63tsQepRNbuxXlVEME+rLQSCChn
kNkLHQZWClHP5rdl8/u6KIlPifflS4qkP8xfDa0k4UuqAyLydzJnG8+tUiW5jgG5
pitG+B4Q/FzhhAnGN6Ca4Z23uuUV97zFRGdZ7235E3YIvgFNiyfjpgPtlKYD2yPj
HN0dMS8cp72EBPv8qhPECB6M6NB6KKfzpuGtYtbpSoIF8LaSSUNcTBU4JS5uczlQ
OidhqmOEWyfOL3BMm4tp2jlFVjQYeS9pf+SBxdJv3oXaCZPAipqkLwyvjxIPG/Lj
oVeiNbLz+klFgoKist9u/x5H3wRLbNMAjB8bfNmPm8GqYY5EAFJ+GJSpLQ8kqsNQ
4pb0Ak3MNMX3geQQCb9aSbQkCXPqWeKFRFKX8CQp4yKZhi0NolCBTakXAPYpUIZN
OKxNKXfKctG59dMrb1TlVXZF+/MrXkC7JaaKY9H5BoUBZjTfCEmUzsYA4nl3TRhl
adizBwn6MZTrc4fHWtLLeQITycSSy7KQDOG/vrp0R42aHp6sZ5JWtKLD2b99ektV
KV59h2Mmzt+U3xZbmBH/yZU7X6KoJ4jcDuH1hQDX+xb7vfQ91PitWC8yDhEcF41y
rV+f+j/dKO9x3lFcBSJRRfX/C+MatBaB/bCJeQtHZhMRoxgZbJYNrofauMo2n0LZ
576xSZcDdNmB1Fl3XYoiLb4Yo99VeT8Ib94XiuIe9aZRQqAk5AmZAYNm/fbqz1Oh
kUqDdwqsfFTG8sUaIML5ekkcHWWDXqnr0GW1WgoXJdvBpHlVN+7mRG//nSRU5I1k
/yczgcioaiNpaoDMlj4NgVjf0L84Mn9Yryya8HymDCfBRjLLoHhh6gkK+fiA0iWI
I92l70rHmCWInR7q2zk1cD4/SA8SbbbfEmszIwOADgcGoX0dWYxx29Z4tBhFkTz5
EuUtm3lvfAv5V2AAepQzqyHikXjzERxbANC0qDnig+v4ke7ucxDlyhaLoAJPJjvF
/wCdv/bU9x9JwIhJywtt5iDCRaNhuusWQ5Fe55+hzNJCE8Mh12Zg2fVH/nZwB5ZE
puX72TSZfNvehNHou09glUjGzp+jIglZrzTRpFgd3eMTHrwrxqcIctIU7ib0TVx+
10JBVPC2tDCg2hiJEdUwWqI1KhJDwNyHxmYIVCSzbW0dboEPe90ScAntBrHY6Sr2
5MjpqhbuIo+Dsmdpyu2oc4RQCqvLE3M88PuSoqhDOdn15gQBblZsBU9ajTpFpk3t
U5Qe9OtShQ+hm7Zf+kQTxNYmCTISIuMwUaXmPUhYKGZoYDHOgHLeg3TRZ2wHS13P
5lEHtuPkNVSUuOX/zpg0/UQQzhl45bv+piEMOH9h9UlD6QK9kF9luLJip3SkGdF3
kRiCrkJcTL78kXt4kVvXurtV4U6ffWjvMxuZdrNfpgogvI5/vrCpX6ZUP0r8p6N0
ZGnLpMgP+GsTNCZp592u72df6Vmp7S96mEaKn5ZEJOZA0xVGSxH3Y9UCAxNxtnOF
BviEx2A/ljGdKx3kFAtfD9fjouRfe5Y448BWFgREY/Jkn8Xp411H6EpnYEONRlU3
skQqOvrRUW8xFaDN3zJcr6Q9qkYNP/cRjm3lgv2JdclEa6ku71TonVzikUqoGLmL
Bqm76JHSdKom8iDDtEvK4lxPR2QBwdFZ0b/BPdnQLTDv09zldDLEsZLLP7bAiVz+
pcU+C0MjfG2o0REalq/H+1P8ieI/zjMoW0AuQ50Tlnt/wgcVHOdVa5F5zM5wNqyj
S5orBPMT5bX1EnkKcmfy3EPLkrWt3C4n7WP0ADogJJG+iV6wWFdI6aZQW3WMP95N
FU7CkA3co9dd0ES+YzCUjV2+POySQjoSLG+RA2EwUJPwteI1FqbQ3AcKy4hQXJaD
Qr4w7fLbtUidh20mLrSLLx28SqDVBUm0yl0OzbNvMVXClnp1mIo5MXnCYyyEvFJm
IAAPMU4uczUDgQP/AWz37tLliBe8u27eSHDBFZRpQ7ThgIzhLPENsoHI25EudX8/
zTOrIAIbAjHvLJ7Mg97qj6Pv+RhDeWvFQGm8zx0jXbcqk9CkTKzCDh2dW+pcpM2F
D1CGBbSJzCG6USXdRPDJZQpbnxpR2gg5+zGghGgeqQsVVzYsPQNEv7oMpCitUX6F
o8YYiJdl5NIECXL6b7/YV9gihSp43OwSWsKtlrCPLlP9HjvJzhAI72ca3O3xdrBJ
5VSSeOsGFo3Xi/5gMLW+T7td2IsqH6l8b6017yyj2zUqjlRUZ5fQFyORGiakDQLi
EfJ41t0ZQ2PSrsw0kQw9a2bFfDQNZSqx96VLPn+FqlIQafnclvDHmbq5vAE1blNj
dPJ5At/uraBA9uVD1aVtZwq2DRuDV7I4y3SR06DDqrTNijGdTcmvrgrhDIxNUrCi
2FThcopqg3FpQDccfxNtth7dkv/cwo90ZRwi1CkzUYtjsNyNUvXGyZImcNIvnRo/
3VJBZ8gsAz/tlZ/5n464OgIANs2ctWQIFGHFpWs2nJVDIfOGzEJoYvp4kDOY+7X1
jKFhZaU2jRvsPheMZT1PKCiwhKNs2GG50jvdwUEAi2gfx9nnIsV6tBFfZsTrAfPG
kGkW43rkHEUo0WaWhp6AeBJ+C2Jshz5DMNYHpltf+4SVY+dkoDPlNURuIm7Gjtup
kQylMkTdcVsvKj7UEJrdBifM/WkFHPdwexMFCHcdP52q/LDllZJo8Jglu664eF4M
Rsfv9geVT86ruSGgSnZl/eGPlivrGseYnFWktyuiZfp3DgeweDpSwYCAdApro/24
GAwElchTQtvsmEfR2is0U9z9OOw/x0ED7YmmaYNKWXi4nFc/GVyoJ0FxUfMsFsJ8
RfnD28BBlP8trv3ha89yHJKgm/qRXV8tnLkLuG6xo4RYI5ZzSifFAOzZJMVXIS2u
oOf/rFGv63SZvpkdJGRq/yTpAMEX97p39rB4uWS4UqLTwi+5rJikukYqi6ucCxl/
vNLdHyLvhnKsKIkJ42vAO1ZKWScewEN3X73nITrI//REVxzi+p0zooYhGWzyHwd9
pc4HOF+P5oRFExilOBN8ZrWRZzNAvQYSS/kMqfNXrACNXXnh/3Tv0Flb90W8CtsW
Sk4vW2cuhulvyolfzx9SOlSgRT0c1LipQvFEQL6YBPDutqwo2aWuuaxtX4Xb0IY+
xQqCjLSS99ScuM6JxKcu91y7RlWDd6y/iV2d/saGax0ztEm4Y3yJwcFh9LRYthen
dHX2fRZnnYur/RD0t2orAFEai4xFSxU/AmAoWJFcjV7fnbDCVMnfkEFJH1vJIBnA
eHi+vN738XmhX9psOjzPi2nVXdbB8hMulmSwmpOsahvOITgBJ1JEhT1UlgdgB6BN
QO6eT3LKkp0GZfyaPJJUTfpArm8UKvwAZpInHHDHFSKeefz3rTwZiLBp2FLBRwa4
g8BssnfjQqf0OXiv5ITev+5U9bTeFzZ0xjrrb2H6cCGNEubkJX/VqlidjCQh5UEN
hS1Sp9BAUPydmHQ7z0f/WseiRKe7rrLoO8iSvnmGH4psa86C0nT5vLk/ZX1EvJp/
OU9gyzHAt0dMICgsWtw39tZJuxW8daRXhzQ1NZW0qbYekE2BrI3s02KQaSToKJBQ
a2bnG0AIi2ywIDGIIkrI08tUIb4zHUnePYf+dXO9bEsRckEVtP8AJHqstv2g6DFM
W24X3z4VM0T6Ga/CuUyE3F87c+EzMHddcgGWi3UW5llSomkq7QyJygpvlubJ7S84
gSKKpJ/qOvTc8Mcs1V1eMYlSyw8u7ZU2WFtjtcFI/48alDiveXKwEKKTDuwN6Seq
J25NKidbOBPotNebX450vur5IuQ2U2tUMHSzMzshLwjljnY2pkldHpj2PlC8lwv+
A6excU95UuM/lu0r0yREVA5s+kEtMY0pZIBQgcQHv0h9BDuuQGfXfxyV2VIKdSmA
I1IMkmJW92yEDEeCaMXNIXRRgTAEub/g80oEYG+g7L9me74ZYTLp7gXyBM5NLiRs
6kuHuuBgqIRiASjD3eeMIbPAHZaeZNx/FGIsQiHSPf80XMVM+56kFsaYoEAIcftt
Kd1H5N0I8dNbJvI2BtqbG28kpUdVHV+PBDGa28IPasbcXFZ0wpjLgsGygtC8UlZC
l9wnqtNC16tiErfBQ4mIWEmj+iWFZeAO7OO9s73zJLhI9XmORcopNmC/UnSa8z+t
RJjUBWKbnzA6i1aBA2kY7LDpyDoe5unw0Y88cAjtvNVuAd6pd8GOHPrNb3/HFIUp
sVuvfGMMnSgLTMkAZ4pZ5gPjjHobHka/g0CS9L0Lqn6U+nw08vil8AjujINB2gmI
xuRfoOMOKW3AmDpSMoRzp43aMAwibWWHddZw3qirY6qMQk82Gu3G5gdp17A5JmKS
Tc/8n5sDdeqgyF9VyuMcBg54gAaHruz/gBjgoxmyjks/HCmSyrujNWKMlEwBd61u
YGcotL5CIwbIhn8Ip6R4HMTQmx79264YMw4v1ndBtb4DGIkLAvHQQZ4SKw7s47bV
pZAmBU1sZK9I2es68Tfzr9YLOJ9YYP/OyLStdg2+jQH85i/XjvNRds17Tz1iBaN2
idtQU5zrkF1DaHR4nuta6LQGC0cTV+Aya83PIXiKrJS0p96Y5SF92POIdwvTFT28
xML1uxHKi9szap6dOEvkev7i8avtgGlRQjzPWj/zZ9v0Gv2BwJviN2PNP5QGkkYb
mo/E+lEQ9dK25LWDljrIWE3+fE84KOfihuWDoIgM+aC4g4HtXDkWxBX/u119+R1z
hXiNaBP1AdAjZT2dMQtFdFA9j4h6SQW3wzCCD1gnZ3gFPPMRd2iHP2zaN3Myxjaw
4KkhgodbywFMA5tR/nKS7asy0+PT1HzAH0cHMlA+36ImRKBawEAYrc7x6dZ/m5ba
nfI8cz/d0kXV5QhhfzH1CBY2Dp2fW5+1mEbGhDfJqSkwmXaU9ex6+2KHbHDu3I/I
otabqysAooL9Oz+MKe0wFVvgj3kuP02B5Kwp+nJoPvxUZc06g5x2kemf3W9a34b/
/sf8huWZ49V5i7W4vFugvrMC30OzRFJDepR8XW1Peh2sLfOOXVhd12TIVHuwHMEx
HOEcg/PMuTAuLJs1rO8EcnMIww/Mx9ppeKX4jsxOXOkXc7cqRKXVv6JXYKU04XAU
aZcZpmgsQQZDC49jKB1f6GtDQmmieNtnIl26MzozZ5DvXAEkdqOq02yaAvQWQDcz
Dhk4ufTrKUbHP1IAwIO0pjXZsnBZA2K+OuKfgz3HVe2ZPFFgrHNCF/beC7buBc13
Ghlj6/SA3nxWO/d+zDxrGVqVPAduewzd2Tz5cd3203ewMpin1+NT9kO0ivhvVKxt
pdusfY0eMa4vMQ/79f6X5IVGO9tmWFZtdqImGGNqKm4zPJpCp/JHdd1miVADCdSU
49diKl417ipR8RfomI5EcWE6pp6YJaNJpPUmwGEaSK7DGW0VgbBlzXwf27lmLaFe
7j+EJy2DVsevJ9l/fxAwAPao86A9xuW/Kye+UA3qAnwgSna5YnmfAfXzH3oDOwwu
3iUbiTrTND2sCx4Ib1mSVI+luwBEkfWf6Qcs+NWJl6Kpz5YVt2INplvKlHeN12KV
7uNTV5vEX/mQ0fcD3NhFFf1IAki4UgFvKsD5beLm9mmyKPklCbFYesv1haOM7Ewe
`protect END_PROTECTED
