`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kd/iwq9d0z/tMtHDoUkD7oFbA94O8J6cO53oagYGnZy9Lw0T4GGj6CkveXYN4mVk
vBlSg5hh3vVNU8TJ9DziE0fwTaqapRcSwXOl6/Yj1BIc43OCKY4MuFP2hhEWAeDU
qP0DZDiOR0uJVQEFOdMrSIRUcL7iqXDh89A+NGlU3D0BJG+qArJMwADWgdaB+kxR
WMixIJ8mcfm9ppMLQzLx4plmwB2kNVg1aFwDwlc52CJ4FrvPxYmbkIH8O84n6rmm
XSYz6frI5/1W3HFHhLwc2suShqYQXog0qLopiEHlq2uuuEiBie+derUqW8XOWYBJ
114mUclWNvoKJLzDt38m5XHJn0NiBLUhS2ZzzrSnA0DikSxBKBLlPmSVrbvFM9Bl
wRaDUBzm9Tr0Sd7gUKChZlczkoTilUUuw2oBLaq6xqJtswjNYa6LcHew/d4pPRxr
t8eoClj8I252Nk0CDljRqyz8Ue033Mhg4e/svTlIsx/U8Op/JYwEGcAYFARNMQwh
Cu9uJ7vFNoWIIHM//508toJm69SLVTb7Z0F9evRyoCXhqEx5N5imihVuWqC3lbaC
xcZcqsC/M9+AIYvxxhpbisWKs9PbTJVJTLUFzk0wPIJ2b5CvVzR2oDsyZ2wP7+Id
GOFL5/JwfoMkWtsdQRyhARLHLfpv6pmISBIu0Vz7g9j2v2DeD4VtzhZhIDMMA67D
Ma2JZgwzLbMY8MA2rakbfg8WDXjd1pcvXsGlYj2it/iGYfF+6AT2B8G36DJMgh9y
`protect END_PROTECTED
