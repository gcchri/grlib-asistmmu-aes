`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cqaa1yTVglMHH1tfUKXBsXlrsh23uxoVSA00SSRla+6phqLiS+ecGsWDb879Xpgj
pUo8hmfldFfh2K+LnAQFfLt0gwOCfadu070ZqK2JyZAbNfq192DSjPfnQc3pGwid
pc2NgsAPremIJOO73EoHIVVPCqOZIUU858RT80t6FrC1k/8tcYE4LdVHYdktvxTZ
+GQxNV+wK1djsmXpusxM9XqptQcqjHJhrKTB9X+SaeRn5QhxPSx5Jdo+V45IBcbM
egP8y+DsxGKm/TxOg+B3wYIII51WTdndKfkORN2MGOCnH+StyqZ1liDAreHJ13aJ
Swhp9h3ocvkrlh3KTEiGs2kr1Df/B2oFiOBBleV9CWLC2dKWnC82XHNnmtQytt5q
J0AkfSNrFOIn1354t930q6WkX5KHj/5EZYv/CfTFpG9SmDepWebZ74GgKcsgwb3J
eSDmpB9rGEDP6ULR4w6Zl6lvC/NjrF5QgVQoFh3ar42boyWtiu1p2/wlv4J+U/a7
`protect END_PROTECTED
