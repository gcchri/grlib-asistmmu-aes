`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hUgt6cjI1CaK9brGCr/lBE38cggsyhYX8NivzR8gkTaWjVdYFlP89z56wsmYJ5nD
9UDlyGo7rrx05XHI+2nwt0R1QazeE/XWYJIww6890Y4eJUhrMEmLvjG6B3rtK162
1nWCeYG9zLGYNCz8rHTPsAwFJwijm36yHYdZ5q9zLxOLxcU3hHJcJ9BDcv4URC9y
UbGJihe7QG5Ep64ueoZqn0wYRQatXRfDoJds2JhqPTBP0aE+Jtn3IVa2A5VRFEa3
E9sumnillS4HBLrECUrXzAdlZ+melzKVafK+40L9qwiNq2hX/7HA87FmtckIH8Xc
qOzgUrt/PUd0B1zxgtkJp6qCKLigWU/czU7os6Jy6l1QMciIHfksi12UrqpejoT0
kyr91OrwFiZ+Do2e0Lc3/hAB4WAEjqE1jQoducoZsw4uXh+C05NyszSvwhdWIkv8
vXKLHj/p2U8kDU+GtV0UqEuRThIuiECwBcsPqApUofWyamQJxPs22J1Jdlt6voEe
NwnhU7cb7mh2Ye7weEaIiVXlhkq5//WE2kkZvHeWZlE70JxkWSMEx4qHXAUd/e4J
Qt13c3ZknhVjb/XLmbCGXjFhtW2vb0jiLm6Lu8oVIr37L2C1RjwB9pbDnDAJpxvt
FAuttgX7h42soMw7uZRv9DS5aHPRa/ok0GKlvowAm15U7rZRocBXoVMGdBQoo1hb
C8sb3QqP27CmlpP/+7QMWYLrtj0jwew5KjwS3fwMNAW3Kai7QMPv6OCMUtI7Qlhy
0ANv4QlNIFtCjSPGBU2IioNqBpDObTKXWw/kLvG1AP4muWWI7I2m5UAOnzgM3kMV
G/4ou4aqIrbm6VKwtqtrfu5o61SaQtU1ym1xTk6a0rUJHjXaZGQwgrT2pIXtnNhe
4UKHaCMWa4/OCgVRerUWlNt8iVqNbUyJdiYLHHAa7+2orUmuQqUZOrLM1VDUTEE4
jz7zAtOxHRtQnS2PXT7JojJylLW7Eg0unGD7nmY0IZGv/f2OyQABrO8Vuo+8Ygxg
Kz/k8A3nMvV6xZtpI05UcT2xSxzbMa707ZIKgjeke+RypIap4AgWOiZ3eysg/kjF
roMFJFGy9nEz9DOzRBGjv2XWekOYLJDSx9RXZ2uSLfvEtLuydt/SvHMRklJ143Xg
Yti7moMNXd4kedb7yVi8g1i3zSZjA/RlbOiY8I+K6YS/tCuYPasRFUV8G6s1cXO+
ygGHofKQGL9Jv92txABDDryNZCPD5n5vwLMNTRXOkN0fFO5VplhWSZ7jXYvmKDx2
`protect END_PROTECTED
