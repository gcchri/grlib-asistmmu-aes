`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ye2zPriVXGw9xlcnqA+gg/Ai01S93r3HtjBYSecRvpX392UHJwVTa5v8AH6SalZL
7CD25j6L8atgajEyFM7rPfjTbWhp7GgKPtzVEVGRnyG3W/KteCFHZpR0Up3VAMrG
2MxzmFfxJfed6+GQg1Wy4xVDLrZgxcWsHceKK2wANrqai6Fq+gMSUzciUrQygrBB
SWuuGXrm8w+IDXPmLENWLf7MK3XoTblHRd33il6bYhr/+6vMRxtqLvWiIZMTUHf3
vhqoQc3ZITeruactQ8Dcoc9CaHpSjnRuNnv4Z4/4nUPpmbWGQxWvtFu5xtmBIHbP
ABP/J9z1N1wyIyY9hBO6dVmxrc76vp5bY1xnSeiovsqNzm/QSt5WBXqYrVlsrgAB
QQoS7OnAiak4mhQVSvcc7Q==
`protect END_PROTECTED
