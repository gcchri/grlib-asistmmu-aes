`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0OiQp5FIdKQqcjzqac3YsOC4md++Bb8Tw19Ut4GIcrF/yRrzzk9E8xg6p6qZxWh3
4+bXYBxwIjaAYoEswJm3e79DukXHtb80e43TCAeGqbCZ+7p9VS3feDxxL5t+NYPw
XNK3NFpFRYWtw24gNfr13XtNnmNPJpgp8o1AWHzR8P94MfovD6my7six73Q7WUo9
+HTOSmiW+dspxTmlxe+udVR3v9hQHV2HhVO0TnZd3rxiXcv6MAsp8qKcMZ0JBISK
h5FG+S9nYFTnH5RZpNgt/uc0w0I3dtVIooHlODDbBrQsX3mcoAaaiKnYVNFHSaSF
oEcdQFGftuB2Sk7bU0dhPuqdqyCZE+fmfsWzlLtN6p+N80jKId6hnko7XKBOLJxr
NhIB+/FIISerG/9346p+92X/k/bJ+Cvc3LUCTKZ+g7EtEBuAh7lGMF2iJRLvGefE
nfy4ABFddzu36oIxIKS4WPTqx2lYNk4UFsVP/dz4Pve9File9nIiVY224qc+iHx9
tOBYIqxDHiq1QVRfnzuqnDqqcJmfW8M340Hdh99LM0qAgx4pti12RvW7Yx1Iia5w
ZmtWu4MK3Jq96JXFtMCcTU2XrnFvGKcjpjW0XhEjkI/8yPnAfe5vNByymE7rVXpD
DDCVVzwFBsTnGgRVLp3DAO7t8xDAXrpbDZn2AZ3BQZPz+2JqgafoLA7QTouhV/wf
1r+qWgxVZNkhKAFL3X4/hUZQK3l8d7d1lEnwvfEZ4RAkC7WfZpqKQZwHpVjXkCjI
BjMCdq/+WsRCi3/qqACZa/5R1mUPiSD/RIRUOVcxW2cnW3FLHeqw8cE/qUaK5C3k
HnYervwwZ4WHigWyAaeJ85KM9RDkU8T/Z87fJPQ5T2GrkLtrfqRmkLaKCX+WBpAq
3jQYRAU/K3o76dL+NGGH/RNzT6LvZKKeBIOFGtgzkWqfxJj2+GNFfoY0UT1/2RLj
JS1iGliFy3j/BWLb7qcaYjYxpseOC70Hamnza+mLl0axPHB3c+zG9kfkyNID2Jrh
`protect END_PROTECTED
