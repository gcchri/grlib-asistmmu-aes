`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5xWTeNxfkxq3xK3KlHSNu7FWdVNAuHKg9pfBuLejOiu1jgyGX0FXNtKnLhklU70A
l58yjBLbkrtPsFpajO0NVjB9iSok65M8KdvNsjXXdeTyPT7K9JoELLtBERwGaD2m
KfYEydsjtlFTa24ed3ekmPi/Ll+QV7XyziCUplDriSmguo855bh64Xkh0ybXtM7f
ySC7Xn/R/H9JL1jOgoJGqozpukaVeNjx11KuIWCk7MuVT3PyZbwVPsOp5TDLkEfq
zhd6jQ46qL9QkE22fx3qmMTanm7CkOw1UNx1i9ZdWYEKodynJx2NX3HLGaUumwvu
Q8a+/dqX4M5UZyUH6tTr3bIE3RZ8zWtcbGsE5tzqdZbJKBEJKjYno3SzK96v4eXC
soJFJuYvk1ovAz7Z60XP86XeqeiKN1p1ZQ2xVp4CY57zCfDuzF8K7LIKWqxjwyN6
vrghdrdzrlirbzRyUjj57mQwYkGNIgtfgIy/hkGEekDPOr4QQ0oBD+jyVOKPXcWO
MP+Q8C+OZh2UeQ+plFuKG9UsyrgN74cFsRNNh4ou2alwbjreeJPx6ROi4cayWKH3
eJyCO/oGKJTh2PNR9ikfGx/dHvb1w6T9AWeXyEJ1VP4ZvmM5vpjlJtassEAB/3Bq
pT0e8I+vhPhNNav9ZJIgXQ==
`protect END_PROTECTED
