`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QAWLGpWqwiSQKN0mjt8y4+xWKuJkZP/vdLIdLnJozBa38xuyPs1OqsmaHCinfiXn
LHvMKHBbQxfhy0E0OZHDd2NDk1s3KaxGeDqdN6z9+stASO2Qk6tO6/Q31irPrkVf
ePCzCO8DIv30ZQkGJM6fGJ0vNbppKUifscu/WtVBAZ5nj0ZQk9F3LeDn7qy3zXIt
FEzpaj6hnIdVWyAp7gPyf4INkWJaVKbN01RZi3P1RRhc0IKCMU7wicbynE4ajIkN
bOFU7ij2jn6cZ2J9F3zSgpv9UV1BU8IRlG7mDusC9qrFgcTwAyRDaWTrEPgAmktY
Ski5BBa+p170B12QbHf5kVTbjrK/9miNRKKhs9oy2gLN+P0Zsy53Qb9nK5ZKSu5u
F61ZVdejDzsCHYW33PLZCdwVYYLLzQG2+tSdP8JUxjM8+9jWuCqX5xzDxmclM0vA
JmGhRJfTY1V4IMf4xuhuBEq0d19OLnURfyHb4agzq/4s3GQ70QyiHTX0HO+rsM8q
slG9lyIpGetOyTdGuIkGxvgp/BWxCCkD74Elh7gPcoV08t1uMawbIjoZXvjC3Lhx
NZbej8oJTleoke02iJdOTEiPEqriUGjzWMzvMACSH/UV4PetpxA+W+0yIl00ffN1
DZ9RBb8xx0xqaHUZvY7wE25M1Wr0Y7lI2lLeTrOkyDdWUeCLeLDy5ldaeT9xnvzX
sMhzNwlnu2zRmHRc3+lTtQ==
`protect END_PROTECTED
