`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3uF42OG/tNtjt6nkxfqviDL0HKxSEGkXUyAAMxrnuq6r0Lxi3vmcNsQ2TPZQ/fA/
/HrUKfECNM0mkooot37UVLJaJ60Di3F5MDIvIKfxamCIRT8HD9uPFBB6T9OCMaj3
0FPoOlJl/ZaOQDNPUqconwCB2/f83W1oznWbOBIJEYb8Lly8502rnJgYJ/sN558b
PWhOdMYsJjcusIquLzQRuujlDG0mSylCbLfgEXLrP+o07lLZ+5yu3r1X1T4yCuoA
fJX09Ps5aAX/0CnOLZd2GNFJ8i54wQsC4N6jCpjvY2vMDi7fWazde4I+70PyZRSN
hnUz4qDa/G7ceW0X4Da5CXQGLgYbG4ABqvHl7I6DpyPbP/I3QTbYeXtQyPpOHxa9
eg+Pua8hYiUVcmVPxqy+2wB74q4M1FJjVhtSWwdSjxT1v1MkOJxmXma3hoAwkfhl
97x1tPmRc5Hni+uqhUSQUsv+r5OgWjZ0Zf2GBY3zOhxljhp3eCl91REZ7mMPpFKN
1at9+7eFjhOMJpudPRq/aA==
`protect END_PROTECTED
