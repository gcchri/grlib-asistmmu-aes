`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mdAjlkpE8MxRLSqCU1HVORwE9ZKpEIi+USexyJ9Sbnr39oAbRVu1oE5BczNvQD+C
UlllMb9XmFPl1shXMyLbCCu5KWJ7vNT4S7UhatHWOPA5A1ntylHLTkMn4Tn6EDAr
8sb7cUdtYgg0BUxYx7ovCtaABeZ2zBMItw0qSyIbwpDWkB27KJET3TgaQgm7Lzvu
b4bn6w/mWmatvVpJFkHitYVbWD8hfhaPV4vCd4rX938z95T3lOtdUrUM3CTiDiiI
mXpSQiuCbB6/STWavc2A71LKkr+c38xGr+vmV3zHxUV/gU8i3OrZzOIjrlujDyfa
bmAtLshhMSeLk10lfGILuODUJvQ1D5tyN559acBjOKXrhLGda5fRcruJHFYmcTWg
qWe6WpMpWXy+DfDkEJAcc0r9tfvr3ojnBESMyASV3dQRrKFIVoTjBxCkY1dSeQGx
Kbff3E6tFA36Of7lxsF44yELs+kntx9aS+CZPy9JVbhmFFc2mL3EKmlENoC1t3tj
PSxNJW1oDAg0paBT5M0HR340I1SE4V+BEWtj8ovhkaeVjuP8VkWwXDvE0pVv6QtC
lAj006oRh0Z++YHA8TYjJ1zk1AW51xjCXekxLhBhnDubDxK6j7+qRd/9IZNGJmTz
G2Pz4NLeeudtWWa1UjAVIQ==
`protect END_PROTECTED
