`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4t83Xw1usXUR/G6RIH9fJj0gdE2WGN5GM9xiUcvOxsb88tnW7cUJKbJY0p4r1NoI
RZqjzWr+Bnmvu0MF/HLXapO5b5sot/GYz/S2v7jcN82bbiy5rBl4Nlx/COcxzMGo
eGR9jfb/VSd2jJ/KnP5qmyYreIZdpoeQOuEp0iFB5gAvjnNTM2dAV5+U8c+5XCqa
DFnweyy2MvbN19ntic/4+ocMupciz20Chef/0lXCjkeLdv9IRfuzQiiDZNWS9PA2
bGFoOrKsXxNK6ZErWtSOGBH6mIwX/YybaU7svvNMMvB/YoSJrrfeqoJSqHOWCHW4
qXY3HMNqrTnnmPil8JjHLrA4r0NKw5EgagfYf8iH+oxpxu7pbEBJDvQROh8Z3QwQ
O7ITs9CejDHVDI+mz/hpA6w3JyDSUm7xekPo2/SPfuq470sli4yVnkJOtx/jFBAP
cHw9Ijv12gsVrd34NbxePL9U9QJz5fKMur9aMtBhw+FPZg8MZwFcBsAozpO0kDAo
sqx9g90XmXVlW2kVvaZQ8zA3qAgrjt7R/WEsGI4QxWQRTkNtdE9JYfp9ozsP4VCI
4IeJpn7hr22LeGbt8auTwlM123U7B22da6T/6YOXjn8u+N5NFE9vGRniFA6n2g/k
yBjfbtpXteje82IX5SFelJo7wC1E8xPLsoFKDBGWd7YMjMUrNb6XZM/I81RKmnyq
oNWobtaa9JpLYZob2npcRcnVNxrwcs3b5bIWeapSidxjCtx8JqXkGawKDuGdtBnr
5dVv9s0Jx8YiZ6KktIQBnzbReF9pAwKxnSY1jDAsGXDq+sc/I0itBnCDk/GLDBIS
NP4UAMeQaoJ+5tHzMqd7rDM3+XpgTUA41UPNiOxA0sewB8JVhIB4Ydx4VwizSsds
rcBLQn0RQikRQDVdRASjPD0z/2olcZ8l7RacXeQUnMYdY7rqet1hfbsvuC5ekO/p
q+nEW9noYGg0OnVnTgC3CWrzfF71hDbyfls/Nel8BnvFITrot5MiwjVzhJ3Hr52J
N/dO7u9vP227QAa6o/2WTs6puKTRkLV/wfFsu9WCzOXGksfJzklNlqYkdIWdNc8W
VMGDXy0hOBWfJdtMG1GPikO69V3sxWYz+cQV0IsS0oO3efDYOh+TCrHglRYRWFNN
xD9FMojgw/OaH3r01uQPb7IzQNRvmwU/E3IeZcP27gnuFmZWicSX4FSj68zaRLJQ
AUjLjawuRWa2yuwVrQRQ1jB1FNFR6w0PhhI8X8VZgRy0b7V2pCLMza2dS7HNtYZy
ZDVgst8+b1tOduJKGplEaluhVavwBMsrdnew5rwFzsBHnBskIbhHwqJoS1ULiUnR
ypEjslxoWkXA5nb+qSzdsJJwoDYuKWP9g5mfgXhUvXL8dmFI7PRrpj0WotARLlNK
dDOppxZDFvyqqD41y4IoZfQo8hJknbUN4db0sIX8EKS7bXSOeJbtJ94NGiF4D4Ax
Ije32Mz74gJZv3UrhO3jnevMM9Bd+JpbHhw3dvKFPATacOL9Z5/Rp+vQO3gZt6Nn
x1BlKtKk+vj/lNkpWP/eQUOCeUtg3KuV+qmaW7g92Rwu5ZSd6AuwVRWlLNM8/Boi
wWwUymTwwe/ntxiXX5tYFz7z6Y1p6R7oAy3RPA5VqZsAGkWdaLH192i1pb9m6WyE
gWwVihqJ0673qzH0GW1aFi4sjE1SSUkq0kN64dXMs9p6VxA+kt7cf/PagQ8khHFx
BA0PUrwr3v4a7xtvSNJuvsGoOfV40k1GtEg9OhbHrFDnJA4arOrVytqqgborLZsl
0HPquHpupFR8PaBS+5cx2TwcWz0QZMnpdojFyFSC8fFeKtxpwklWz7Qcz3gk/Pan
EbOQ7Jpw9+g5ZeIFnkWwsR8zD4clAV7iEzdEEUHdez0wnHZBKyQV8u0A028eKrH3
2ew5YeVBT5Uw6xDqEYkYAjdsOnxyJoprOaHFN2p8zaIVjEWMbLHFvELDZRKyG9+b
0Ykja9rbVGKAcA18MFpjP8nKslcQ8TEW2AVeeuWmeNZlXMHyPu+HFGpA9nsqeS/J
gKjbT1o361HSE+XRC76hdEI27ToQcuTZn9ZpfPq+yJSGyO1TE778jHbha/c0ASAn
AZkh1YKaESuBKgFcBGoi7QobzNbbalXEz4smqN+2s+xT32BH/i+2lqt+6yUrGpeV
C/v7aQK3xfQeTVcOb53r9X2tgcwk0EqK7H4y3wgg/957rZFLfyDui8dO8M8GxSwd
XLKVDmBMbL/QRBl+E3VI3or6hUdsrQY2z17i/n5xAYLLnBw4EnJrECw+5Y0HLnzG
BdKyrvlwcAQ86oN/VXdfuxaH4Ky5rVRDezBM92el+kdoVrZDYza58dKIKnxBw/7Z
8hm+I0lhZmwa8Zst9LrCG8+/xX7Y+Xdnez6Idi2k3a2RKLJ29J579c77IM/gAleG
lNf6WYWblzYu9S+KfVgWeCMlyg27worRftwMtking5xHt0lVprWpfD9ZQpdbxcdZ
0/2FC/rDxzoSUcdEAxoCFVWIBi4Ikp+qKudPGHm4NKDF1b2bc99MsnweNz1UEwry
ToeFsyxBMwn8i1Hgg0NHyoIw62nk5E/LNxQIryNUmnlrUpmoYm/rYeNzSK/TzFQr
/UXqcsVsVHbZTloHcrHVX6wZF2edH7DuahOlMMiFORxWzqtdroYWIHPPONsjf/px
KN9Ml+F8EPqoK5gDHys5JbLueB95v/N7AjEPMEh4QCJjfz5jVqs2Dapo2YSA4FIe
Wusph/K+WNfUFu/kNG19UQ2VndlLoVH4r5gIsXMjbhgimvXGweFfj10ESE7jqPnF
vH9PaiOqPMl8806nEB9X5CnqNzv+yE0wPkkcLGNVP6+JwNpMjwYGv/KSkjEcx+VZ
04BX8lb/5PwoiBRYGm9fyLLXjMyNofKFk6IpBwqFYQX5jzxcQaDwuSZqbcGUyD5g
pZX9vsOqLuqEhJY4vDrVCsHAqtWDfVZ0zghCLDKyZ0/jYUUZU6aQCfqKYgS5wABi
VMWvER0F1axbGejEIjKUIHK56CBUP5+aFtnGQz1tMCWQQDzWwxHTRpq0PMeVIEhd
DkXaP7hzHBRHfkFXrVqTaviH+myw5H8H2177gjADK9yh+J4aD4K7yaPivwiAqM9u
3ovso5Ri4Hw38g37JRL/0tR/wGeGt5Ht0CQRUyj4yhrRpLllCiWeAhASRZOzBLmO
xTkn99WxkVFxSVT6RQehwdPqSKysIynq7rwDE/a20IL4dvFwopJUj6Vkuq+c9S1C
c7tTYoe2LqSLzHCC12Vic7gT3LvU+4OaG25KCAVbTnvmk1Zq8EuFMHA1ucaCT4dG
+2fdW1F8KQEKX+/Fu6E34qzsvcMwnU+QhGy5tWHGp8ZsSrq22oRfKFsPgQ4LHTfR
YTd1/PUaeQcAWxD3LsCaJzPkhBRWV8UxKffttjGhPzcwYwFe3+T+0O3AXirLaFEH
s+NPc5vMRUpnUK0ZH79j6tQtFu7sUS1YEeJ+okyj3+W2+4h64y2fP1vYP5Y+/BpN
vgIf/DUqEvvBS+7C6Koip5QxYOf6NULPsbJzJxQXYLhV8q/qXjKiZ43La3NEK9k9
WLo/vNlarhjzkzmtT0yz39Kez+ocgN7hZVUTko+uLokMtgC7QuRnXiMAxTPSj2Ik
cD/RXbOJzuMccVbDHPHQHPyzL+gBVIUeKJwydLE+jpsV3Wpm3Y9UxIswahahrvx6
XRhpQqfJaP/oRqp6ePTjUxTcCN6npT5CA2ElsUCfRhGWWkOYJm+b5xd89+czisgC
EtrH0zIBkjpfmkf0x1FuV1au4tGpjbiNch5I/xDbjl0nTPAuIMaV2b1cXr7xW/rS
GtNVNFrGUIdUEdfjBroc6yqaP+9z+E/BeDlNyvhPCu5Uf6YaDYoVSeM2BgwTchYZ
qSNOzW5/9/BpHBZRiOAxIWqJRPGMLNZ1bqxuNIusLPydCjWUl/nReemMIwahF4dT
++DuVUw4RqI5FL6mGOAAi60+Nd2FCNrlAn5k3VuNB0xifhmXS2xYF0oH8+BuvtTT
VrmSIZtQLGlSxgF9nkIrHqX/owb5ZnWOOb2hwE/x5pjaV2RP/z7cfM9iRQIMZSFB
S/dYK/Yx2EzW7B+Q2fg/6q2OYsx1F+wUpUEQjXz2AMJVutpP8usB9x7I4Yn/Ym/X
1vEzVdVKuD3NVIiHHEWBO9EBgFJ0V7+WyJ85LmShxgl2POJn/7cSZLS6aWGJarcy
hudLE5B7eVS9eG2GJ/5+BT1uqC/vLkYJeMdWn5NHvs1Hqb44mcF8cxp2kQhw0Hn3
4NflmiL1divS2DmgxrCXW1MFKB1Y5e4hg0C013OM8LDEoobUDu7P/zPQn0qroD8B
6urU/sI7wcaDDy0Y4RSWIZTPVbnDl16rPSzALONGvvANPkjzpeOVwwV0BjOeBVYC
sfhcit2FoMzuorWH93JLwtwl8JZnhLFzB+w6wNrTCwystsLReCUCSoEAZfTmm3TD
RUUr6QelEZtzF3cTtvIkdDtDiccZAbVe8F6DThC2irlLi1x7uj+22/3mq6NWObYo
jBCtceVXQiQZ1RX4SBXFzEtNKZANJrPIU1UQrbY9A2noGek9Gfvmbzod3IG65rMT
uHOLjUjORul8f5dCpxeqnRGBwXQC4sXB6szPYxRDg8e5v1SmYyWnaycs+ULbJ5Py
nKQhOpBw5zrZTvaD+LYf8IIaZmuJFQTGa+Jsuzfne4QN/pOE/gMPLfGwjt3wbz58
IszDvHT9LhlOcd7lzO62nMi5wBKeWPmOfNmnrvXjpUnnWP0Uib3Sd33bzPhmVtCN
Ki27t1oV92QqaSq09Ab7+Aba9U4zGPQ9TANTatuxshDebA3Tf/0L6B6HErHhNIxG
zxC29NJJO4Mph97l1QuR20+0o4UeG3bw8BQOexCwCMH23O8YTaT2UkgiCZ7Sdvka
rKWkRD9sIPhifAMY2Y1q5Vr+0zPsheSgKw7rXGXegL1ko4CbqIF8ETTIKCB281lu
vAvZID0i2fM/KU7f7mGV2JBFMjPAhy10TtdYVcXAIHSG2rZK5ocvqEyYmcCesNnz
SebpOjyto8F/yw70c4Du0uJuWXeTOdhjZPLbLmrfYvhGLjq7dxrt83EyApFBhL/k
etxweWYyZqT50nBNBMgSax6IfOaf3fZLOY4SSwmrd4G78lbVe7VfYtrRl3DwAPxY
oo597Lel5uxxXUejHfMG7F0M1rHQYmkwE5GU60YgrzAGuaMXuTY7VlClmz+CsZa8
RnCpbRU7R64ETezxHT2GsLyPiSpw4LVQ+0Z4zb2+HZHeoDYe8BHY91I9rQ86c4EL
JN0YqpMr2cx/eQl97Zfo6dJRjdBtsackqnFbZmzQm1mMTfn5CIIaq01a8xSq+t54
cUGwAre7VGcG1iu5oiswIl4vROjBE++rbmOOfBftfdypAi8EsT1AtidXvOGYE27q
zCuPZgKa2rpXg7Lt1gl4TC2f5dxfhnO+YSM9PYU0pIO/cMtrMxcDFe2zY4D0/VSo
Mrx+eTV1jVXoGAdRvjWIN1nsaIVfyb+7pjkFC5/nLnpQiOi3PnPKgp/U90xN3syc
FVCDakrPvWTE+2KKPo/79kQaN1YK068L/va8t+5h5+AVQ7LFS72t0bzRfhZBmRte
h01S5ewCViX4+ZhLlz6VMndiCyaranEd9SsEPSTTzBH/voCAXeZVz6NIYpmEHt+F
O6ZXDJT4S2oHVdXLZcs2caQt5x19lHiv794x4UCr02T5i37wgCqqa6b18CG3A2vx
JdyFcmOEPEO9ZOTCb2qoisPDQ4ErpC49H8irBKsHFLnsm3ZpAokX23pg7cx/pT7y
h4yjiWMtQVwRGJhs6PcAZtg5QBASK2e6YBPOZik2Y4ptrxJDAZXr2a4OgGWjU8Uc
WlkfvTBomjYBUTz5ipbQQMzvd/U5elyFHmYzGpWJ/G5qCKfpcJNTSjJUs/Hm9Jy3
uS4TrUySk4YvoiIpgU11ijnhVWe4n9z5wvHFlauMb4C+5KeSs38gJc23Dt8adBae
UCvoES2OAzKSgWpOkfrZ8HWxTroDDXJp7xOthGCFo7be8cCkADnDBg1lYpbdlWSg
95vfM2kYxeVPyCwBvbYlcVtIrUlD2w1lAVZwu2Ulj/KoOEYo7tPNC+WAiCEPQZ7Z
tnM5neD6Qwk50KiZ3WtAmLadzZWgOnXRBy8RKfAvSkzrpzkWD5MHwLCH2eueqi/f
vA52TlJqbHaMza+cjE9giIYMGB43dovzNW24IAnpuwD54+dOqaXbobycI3gO4vKp
3+Xg3sM/ixRAkNHAHCHFlMJxqT3BCHYOOSiKC6QByEU7tbXJaEoqCLlkDkOrs2a1
AodmVKStRqnTPHYdDRhBS++S2Cy2ASuIpddBotgPN6IjBkvV1xDhw9KXKN0SRE33
MJjj652n9V/Iq5XsoWSFN8hfpfsy9A7cHAhhsAGjaO+Dwv2y8e5spZY+dZE40EEy
O+AcEDK1QPbxP9M3iOM9Xb/t+eaD7QnVExmFCVV8iJiioiNXygXveFMGmukGl6Y0
/9llznTWbQ1pG0T3La/fp4y4zdUk60XXadg8clcuql44MlKsHiEuJwumOk+gU8pd
CKtE7elDj7V1JhmiLEzd1TWcXpnGhhbj0rKKpmfJLDplpkid0A0i/ui/z2Us0UCz
yCrNg70PjAO3j3w3Qi+Fh1ETa2tN7p2dgJqoCwiR/otd2eRMZlaF/QOqKYZsFPVf
PH4lJoN/AR1sozJnuU0AR2tLsIpTpowHrc41rDqu3vZOcnEt1txy00U87wEfrrkT
+NV2SwZu2H106uKz/X9M3W6N/q5BFgONHiIa3nQMRvoh4k956G/rmJZGdZuPZaV7
KyAy3R+tEMuhlwuCh1B3PweWeq9ghgz+6dMwTnHfQwKSb8d+/fgB0ucd/3LeHn+h
bTdOYqSQx2cmS6wCpgqSVkpOKit3xwgaVIPeTNkJMXkeKfj4qxMs+fj8zYSwJMcT
u+It/4NBLBoyO0rOWAA+g4OrbDyHyy065jOvzYt/yxcei87xbnpL5hSAk6cPyczb
pEwS2tYN/Tz9bn75CO3bPBkZVpXnQIQRPo5lwPxWKyGy4j7hRevvPnxQErfShXJW
1x8y7lhhSqwF7UoUbLMDj2psrlsuZvbsT834uPoNyzEU7/fUon3Ib0nx/wRUrR/i
SK5iL/8UaHVoeFMdyb1G0+xipeoFmJt7GbSzU8GOT+RtjgPUBe8SgUcvdx4x5OVf
GldGgBXj1Z5vZ2of2X7U2xuKBjXwnWQn26kxGrFbtMbjGHiuIS3rpIfQx1e5GBtr
6rWay93DqimmW/mzquVJd8oOcxbO+zDxYJzL8L2h+k4+ktEz8FJCYXVnIyH5UQs8
HlO7w3+mbUkrJbaBkLAbmBjnkafTFItQ1Fp+skC/I2IHJAW/WIZzld5rl78SOa1z
mu/D6EcKOjcFhLmLeRwTylEEC0C56KtheVaKvjesZ2h9yLgHnZQvOCnyWPKUEsfL
j8MIFcNBDGe+glI4H/oQ3T2baXWg3EBQcbdmcyZg81Nfb+ydcupv9Fk5AGYIoJWs
Aisd7BBZBKshTPe0Xtq+5noVWuWewdl1i3i5B6vGIPVK8kkTprL5zL8D53gvEO0p
i74hDGZsAk2GNFDn1radA8wlzVbmbWEgw9R+jAhdCcKHL3Vj26+C5QlZGjhVrMFG
Qvl3hAbZ0TbzO3L3dB8mV/3bAkQQ2JPwxxFu6mEFqIlALaMjycS2uqyTradLMHdY
ZCitC/h5PNMZijytDybuS3/xZjcum/B+25771+6TWv7z27SBtsFPctGUkbT3CMEK
9zeqRtiEoYkLJH6O5zggltYkCJgf3BKDIF0ytKzK8QTmfsHYwlM6e+YZog1YPKlv
df9gSaxkR7Xd3PsAWlt2KcfHlSK/L+jWIb1w6DCmyMMsg/zwkqpJVhP5HPtEMll0
nwiPBQ0OeHVdK7SS5QNWr21JHapCGrrBWZ6xjr5Qs+iEMdum0y0X1LOKhslR8Y1W
CsH9miIHcl0z1od06SPNumTf5tuwKvRhp+QxnDI7S+52y57pAJQZgRlysqwnv0qU
x1Ur/z9RJpSpvDoJ17958aTYFmuRV9ZztR67lWUoUoiizXz7ptpSe35krIB8p45a
3n4Lk9V2S4a5BnREym5XM11Z9IKE+wuuhVIcQRQPlaA5S8bsTHmuqE+dJG1nokC6
96NAs5pPXBhONC9qPxsbSmXSpc6VKLXtPasTt+pLntCPRbCq7TOxmPgdgDOodPeK
liGPieP8y6ISzBGlZ6RdIHbc7Yi9luQ9FA1eDX6q7YFi18QfBH5urwbWdIfupqyJ
Z2gu0eBIpR2DpbAdcG5iyJKXtUAIM+DcW7gzqGpFhCBELwkt0iIo1vqPqRl9VBse
rmUdt4x1cjidY4NwN2fvfeQTYWyqQ36tGsOgFQKvN+NuWGrcr/JAMB+lQ741o4VK
sz8D7RVqWcjoFDDOT0y7HuC2ttNW3ruhTnIdjcPL0QETA3GMrPMWpFtZNFLEQZHu
7EzWX3AaZGU4Xgbp+mohFqCvrEcybFJb1R+vLpaZqzonFY/AAxJhF0mmkhXN2Q1F
kH384IXngMK3NElIGQECvPTNQzjvY25g1kE1fqWSObjbwDeCwvjKkkSFTGN7zTQe
ea6Uh3Tuz59U3RCPDOaJuswWIq9TL7H+PCxs+oTPQ2I/G4L8Up5mPzNs4W71Bz6P
3oW2oqKAVIOLZtzL+GUMXUCRZdJMmtr35Sy+0347r194LvD5XculaUBz0aqRUmhl
6VpPML57TFn/9JCXg1Ne5zJbzi6MiKAP2QDA/DrjUoadPZAKFQZChLOXs++XnI3a
KCQ1cwhwzHyI1RCf8mI6eUSaf0LpZEXvKUmeT13L0qgKQ8unnFz2l+tq1REALGfN
Lj+yTupsUrbr+Q0Y+mAscmmcM7ZH5q4N3VEBkJwTCX9zXwjH82Sswli/GXckuZue
y7gDjrBAZkr9BRaxQZddF7uYM2idE2t9R7w/GLuUkyOZrU0PvCx09cpS1jNT0eZ7
gV2cdu0uafICRPHXk37NqhysOAQNjK+Bu0IJLs7hYjeWGl5gsYYfafB9KyPKb+ov
9UM8UzcjMpXdMZhsL9Xd6rEx4gsFqb3S0YXNXpTUGTh65/VClQtoWy8p9SPbTI2f
xL9/oGDHMqQt72OaBsHxi/aFeapXAmOX3duJP9L2Nhy1A5V/22Y3zeJ8Re7j/Zry
tP6q0zC6xnz5knkF2cjHlB8wLoaaG55tQOijIwQypuNs15KxUA2oTDpgawYP8LnP
6+kTHBMgtPDxymtE17njZw==
`protect END_PROTECTED
