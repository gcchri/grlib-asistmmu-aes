`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u6IUWMFG0ydly8jj9BcHmRpT9Zl5owQLmMtKWbIytmlMI1fDYhJnBtQrPfs1jnfv
SyI2Qdl6MOHnwK6R5PNg+tyyO78XGtZETIhWjk9ygTbi60LAH8iT0CAiyyUZuyUF
nnH8sbjDVRWRyDxlc4zWVPQ6moZ1UztdSJSNenZM9yAAUtzQtg5vfaKf095mfeKq
YgmxPzw6go/7r+wOWUjJ2gVpW0d8q5WsT953HTEIz6YWSbGMJoUH3v54b+Vjp+KK
q8NjjF4uYW4KMK3Vvb6vYU4H76fWgK69D36tc3gtImKudmhEi1rD4qT/CM8xPXc0
mIwxizLZqxcBPoZ0Vfljgo9o4LLwhh0Szg6/8jCBBRkwHf9Ixiz9qlm4gopH93NG
KSiiKWQlFZ10IV+FrEB4NOUTsxue4rDO6p2LSVpIrzWmCe8hEiEsnSZgqI3gzKUo
`protect END_PROTECTED
