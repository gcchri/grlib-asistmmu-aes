`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ywe1lsN2U0VnkOYLU8545ASkfbsHKObiSmaBlRvETZgbVuDj89o2SLllNNfOC3dR
4fqBXd5EO6ZmcEg2VhK5UGOGudYHeMYjMNdD31gGGZBKNhii7xiGk5j6NkOYAqzh
nKZ1aWHsxeuGt60ShiQCiWpo30T7kRJHevcFNiLt5MnuzGuFZjplcodEMbN3xhAJ
8aUuEd8JjMBuoYyUuucUXcpPibPm2OB6k5wmr8c1wc+4ez6lODo62MGZ3lCTfbym
5SsQ0Y6KaQ4bVf4OvyMNK9jqowC/yz26RspmxHNhbES1298ZkkAGIoXOY5OQrZIR
fttMJYCIvxcEgxt6NFd78MOyi9DdnIrg109P/VhHYHfBUQMnZtPqzDAfRlpkMey5
Sc74ayagwVq7SuGnq/IS5o2X7K+/ORfR882vMOgnBVdfOJ5ucK5FBEUZXLlgpTCJ
a7yb0QP3FJ7r2e2uVTp9gA==
`protect END_PROTECTED
