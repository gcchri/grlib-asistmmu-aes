`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Vlnx34QlvvjCS8WzPk49QfzZ1TUDwpHa/gggcUAe0CB6Par3zqFrsica0kTNEra
upHsKn8M5YV7+WtJSzQ6PGDxrGNkezuyZmZIpK59M6DRc09Omy3QzQchyj1RKEaR
dGi3uapwS2sH54lrhD4Rq18O4q2Goy7/P6Teh6t5GvmLhCvS7A77xkLlz221Ljxa
P3NVlC8FKO7IJByzWeFYvIBG8d/0pkj4B9ZXfbBxP+fmYtattY3ZW2qeH+Z2gwPd
6geh1wgE1t86iUlNuUtzC2TKxj8nDtNpLZaEPo9g/2HmdRsvExMywUVmiptmEzHu
w9YPYByT/Rcj4vD0hsoaCbbziKDcB30+9F+FmcePyw0Ecj6nLVJ0wo/1Rzv7YzhN
FU+0X7N50R6cNm1kYeWHxz41QwhbdMVhPLGDC74mZJkrEkEZmkwajxokZUSO5sR3
6/Xt9BCvIe6djgD/3AAlASqKRwkg3RQCrPCX3J7nYZKxH8xOHU6/yy/6/ssp8Ngw
dR+z2DAUXCTJDd/jfpGMJnDBZ4oQLfTeuDhvfC9HzDaFb81kxP9Qmb2DS9nSCO20
zk0xtMKhgZas1wrN7DNOAgDP5+V2Lob+cmmbJIT+hZU3Qo40vW+meyr7hthl9P4w
KstjcZN8LGkLdZbXtB9ujg==
`protect END_PROTECTED
