`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i6uifHZmdMxsVKz5U6eMZZe3dtVg/m3qN9JcKpCldrs5op6G4GS/QCES/tVsmyHN
hsTi+AeN+mFKg/J3CQgOedmcIo3tki5Urpud1QOPlbvYzgQ5ff1XDzMvLit6/FaU
wGZ9Y7PcLfLW4idDZNpOr5BEDL9vlDWuCkJx7YITVIDEYYaM8DMvtBpVamJYZAGs
KXfZ4poxF5NLAXmK6fHl1e5Cq/lpT4qRBw/PnB+zrtdZLqh4lMfX9uVplHFxsEf5
+C2hUBkjbbTZxHwwUIRKRwH0Kzb81ip13AnV2E0YrwGLFWdAadiIB2oxc0noTKVM
R1s8/D0QP/k1y3AaUArrrA==
`protect END_PROTECTED
