`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uWzE3QwIKuH8C9q7Zlf9K2OZXHhSluAY7/SPaM2VSJDgvarR44EIoiV/y0MWeZYj
1+9V668aCYHiMFQXFj59iqNZWNk2CxLH+EhvSUd3auP1AQ0hH61Moo98pK3HnPoO
qDP+EXGuutpp2YzMSSUAp76mrYoA3pE5BamBPtK2dQYmeFOQV88FE2Kq541nWxIO
MY4IJlfBB/tNLXcmIYqKsEhlYeygYgG2zZ3fNun1rA4QUS00+KSBCzir4JgE8iLy
7RbILNHklXk2IjwgnAymfbzqm+RjfztoJZCUTSqKcLFJalr3r8t+kZS+AgrBv7ws
JmdC7c5jPEqdr6uP5GNgPreEMTmoNm2gq9dB8hZgoJA2SAaankS+QZHXDWy0Aj3B
mb4wqv3XkblGB95KjobpnaLj7aLX+ne9rGqWZ259NNTYHdjXrlnrF94Zodi+OyvX
vr+TLy/SrHfRx9YRDZO+wA==
`protect END_PROTECTED
