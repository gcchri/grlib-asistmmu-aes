`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tU4519I5YxaBMbCls4Qfzf6T9s2Q8uXOF1H7jFcVfAnKAU8jjnp3+shsCD0WEqD9
1HyUtWkISGbvAaR6xZ7Cs5testQdObuMKKB8PJBsljMgHjcgwqxRZxS+lmPMJpuA
Zfzfus7YjaZDq/4j0S2sn+6a4QUfx8U734R+wiKCCg4InJK5hdVEGxB+Vk5lQ6eK
6y2SkGKJoUZuiJ6beNEG6dkzjDTWMyHzJ9hIdmmKjTSwYFJjBfesRa9iV80S76tj
t6oJ07NcSwme0SRDkTrC8zcy8Dcrw0jf1iUByIm+FbVb9DzzReKDeEszMwttJs08
Y5FQEqzsKhu+LGqEoDQ5Bz4Ut5ginoUp3sCDr3DY1Kp51rFciiQqp7LjVpdiX7LS
nVtkXDYJKhPlBO5KZp8hVMB9n4ePVYljIkv0gO93eJLtyUx9p2QD9UGXztDTIrIj
VmLmMuludBzTrS3AnrZsxw9Eaazri8oQoxu+PbdAe1RFEKdBfDXggLYNUiaHaAat
IEPd4eI1/hDRAZb5ccC3TcqjCv58e90AsjNE2FfUuCaX+dCJzBVfiytP+L+aBmFv
9xGfVj2VvSMGggnns/XbO1N+c7G4/UqjYp3ES16QNi86BTiSZyrEQp6HYH12um/P
IgU7pMJ+t2pUcOWBDtLv+XMHl057R+Yrb5W4ep6mTRKs+CFdtoASjtYv2D0OLCD8
NX+To+C8zdvKCUbjmrpTiSiTsmfQwJdiNaU7VkuOcW7jdgHchN+sL0hy6OXXEbeV
5W7iFK1ub5IXGdnA5keDgEK4QLXOfBKOver1V3oVwDr23PiKXptmmVOsJVsZ+mo5
KT69nAGxKkU7kzfug+sKx3rB2B/SnEeLHlqFf8aGIic326L64FL2rGbNfsAZ0ecD
slH50kFfW1IyPJAcl0fkEep1zpVxaaKmFwY07u36a11AnYJL+ZDLvlST4PDkwc7H
XCK2Va4+KoHZE6YvhftLlkupbBqs0/5avTijV19/xxdQ7bDMoQppxNV0UzFQ7cOo
7ywLaqcq6J0EXavU6x4G7uKWCkJMmH+J2t/ZVV+7bXle5RAYu/iIqHdqTEP8bcTZ
bkquuX8tu6FvM4x7xkY0hKNzEGQ2kmd0w1lTBAI+uOHtjCrRa4qdCOPdGd9g9Hz4
PraGKPStdliiKxyMs3lzXw==
`protect END_PROTECTED
