`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iiRxJFEQ3h2eRxPWCfmt2dVHqoTY4xL1luTSBASPYJyNFTX1zLdOY79tdWdP8sqo
Am5CETo6RVbAwdbmShRtKGhD6xtUjK4RPaMCVN/4+djoIiM3idWzwSxbkrQI9LLP
ngDj4zIXBYKD5YbbASfis5b4h3wTiqZWWGuOXUBkIVaWysyuRfQ2GNwqrwhQ4+hH
x5vjhc3zmci/d2Fa/BVQ4w1xrVAYFx0WhEvP92ohXqySBaNzVrXTUlGHpbbWdCHd
r/TSHtNKBg9vF70VuksXBYu3Ric/nZlFIJpiUyqCvvWhFXNg84QpgDukydg3S1zQ
sSoKRWdkitFLdOB/fUatdhCwscUm0Qs7exsRy1HZk/7cTdSiYk8r4I5xjUPbJnVL
Ge7ESudewEnUju1YGTnr3O7kKtvcGe7mWW8Q0b477UvItpPvI9zURlBhTeUUosl0
`protect END_PROTECTED
