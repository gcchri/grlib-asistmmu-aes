`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tW9hHqzA1JNK0t0FZ/d60diT+CHhfrGVcGNwWIiC0VtQTNn+ucrGjpAz+DqwpixN
0EGTWrA4QnxTgi25EU+F+OBsOe9tBlWVPekcqKoIAkqTZvd8Iq6SgRR8elnWOEKk
5008RmWjbY9JdC70UXiV17lEg9A5cbr+Mn5pIcUhdQaR6cQKN7f0GzbfmxPxFqQ0
aIWF9DU8H1oI1pcdwokiSfNpF392AR8OXFD97e2XH/YCM5HoVG6CMhD9FVLKSLCK
wd2gPOe4f+80VsojWYXgEN7N7VwRHMfP1Z9J+tC7oErsXOM1ndNGBEXW31lRFQT9
eDWcXfR/Ju7zKOL8INpytGqDXO9czrLEgPqZ9jVkioDHNGA/oI75Djg02+RRO3TC
9Chbb+JdFs2zKVKZrEe50v6qnufSN7Bi+7CTV9wnvZTRlqr8Z4AzlC/MH/jqbAoq
`protect END_PROTECTED
