`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xkYAL4jc5VkZw5kNepMHG2rf+dZynbb5/2trAHhhy8bcFvuOEuGQDTM2M3pkRj2G
jUQ2AlpC+RrWAD0yU8nTaVN0rKaqaeM+AxogdyM8QzyU6vpfIXtZHWkVjz9wI+21
J/mv1ZrOVwh5xfS7aH3Up8FOuPzsgO557R708+8GDla+AVfk3M4MINRwi5L41Ort
5h26QhNk3UwXH31u9b2rzT5H80dlnUgvTwGjkoudnJMdzax59jC843WVlDVgK4Zm
UcK0Nm/jzvSs/EtkbHc/J1VjoIR6db5+xmkt+Fmu3DAfuLtyBTQPeFTazSi3fvYg
JZIT3HRL3D2o6KVG8+On393oDF1Hcmg+AlRzwAtvMjhuHQOhJ2IRbdwWLB697Opn
nSpjKW7Ml6X3HsAs9P8tNUdnaLfPL91+q0VSGUd27ScSbAS3p0YyGBIr9M8wJuxd
MHRJIIhAiSi1L9e5dIB9xjEHcOoL+V/rtH7ZPBtdMhwxJF1+wse6qMHl/xc3HEfp
h18XWikh61IV2xssWCQbWZ8iJ73oSwYL4xkYveCMDMKcEltBVaIEo5ridcOVqsha
ORx8qroqUoQF70XhvI1wkNUfe7W3nvIPq7Jm28Mp576nUGYe3lwuPpchsd0nIRPo
qmvSuXwBmS19Hi9VztYEjJ/sIlE9XygobHO+MwerWReVfl2LCh6aooqQOHBe0s4G
sdN9kSP/qbIWT/7wAa2GxFPqbwx6su2Hd5ZNWiNYG7WqdSNbwCyNVznFuBUXX5FP
zzD2ovCv++SBybc94rzFf+/FMpl6wbtBR770e7ahlgo/JE60iwA1GhK7ETMIRnzM
+xVHMTVI5DJ9tEfKSdx3JOMJs6aJ/+xbSiZFcKsUq8JI34oLuAAA3KSgolj0OJF+
qpePFvxWv/OpSpmQlavc0xd5QSjlYzCM9aI2Pyene3YCqVFrlM5nYQvvYy9geeGU
D+hQ4KedHOVIhDanAS247hUv5ymUZvopsJynoHc/3D6i4WdDAihljjSxNulnnbSP
HDzoFoi8TEUoJag7yxSV+23XdN8G/9uvyad6uOT2aryo04GX9OjeZ/dY2xN3l3SL
mBSfoHdJ1vs9LAiR/1X/dLawFFY6PmsWGudfYdaezsrotO07E7QxBge5ASGlN2PN
qrLrneryxQ7tBuGJJ5v1mj5YIUwcOJHALD8ukyjlOjatQtpMRC6UTUZrtVDBXviS
O0DASyGT7rIjo5LDkN6Sm5ia77sLL8G7zghVTPOGurlKN1oMcNm66f5Oh9184b8c
7k3TrZTYAZ5Nc8Zf15gM9NEFkTa8km8HKX0WVchzQmf6rx6CfvuAeyBH33iDmnj3
FXx2fhsr7S8oY0pMdy9D67pSOuorZ5Xz1+Q1ftlzNvTpuWSUkPMvPYcQkjpw/qEm
MIheGTXhF+xiR+qwNJZfZJcUyiSBQpH9hmwtJ/FXDwbmrbA0jM1aLw91iuPhLK3W
OwbRvPRKSqyZqmhNKR+0mz0d/fuQHGiWo1OvWyYoBDU91R8b+gpJqRlZnA9PYZ44
QgAMR4J6+V7V8yHJKNl+sH1UOn2a7jPLVyZQtn+xKws+HjR3TafAK4Na731sl7qT
2u64q8fn+RL0Aq2BT7mC1hLzCL3h3u8h31jJrCP2xYmLBEbRxRZBeNt+t7QcyR00
fwYJRVojFf1zmeGafgWpc1T+EaIh5pDs494zBQ78gBHvtZ1K4YkA0pEZOOqa3buZ
A68AKuIaZGQXzCKYcPtLQPY1vfLJUdpz0ST2sfooU0JAzhQrGcxlU05v0SRkFGKC
0xX/nelUO6+FYy6KXtfKv+oTenSFITRBrZtPsIeCC9mPhSwMxQcMM6OkdmOqmCfg
IUdUfVYmxtBy+NkNGzIytoqV9vwAlG+F7F6Qo7KZ2HuiH1PZI7pc8xUgvtYNqPXk
7lQDtjCFAHzjLhQrPK8umlB2wTA6q69MB9kCkaJINvOn9DquAzQ/Vg63kw1nezDN
v4Lcggzyq+x+ZBALF++0OraklXxmKX9HrorDRRx/Zu+66qsUQtXfqSxrpHP4F4YF
x9W88Y3gMw9tSl6e5WUFtY3QYsSno7SowUyKrSrtaD06KBztahx0P8d0jTsTzGj4
vh0cXwWSw7O5vlZWfMffIAgVzhzID2KKCU7fop60Lal/BAwlAIhkdB4eYdCZICfp
`protect END_PROTECTED
