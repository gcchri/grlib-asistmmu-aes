`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wuz3UDFc+A/tPL0AcD5I/o0+AiMHdBcrZNKappjGCOftlEQcdjcbI90RzH8dO2fp
Szvcnw1Y/ovz3bJFvwJKLALDL6+DJJBOcDueh2SlNJCebF8gwxFPV5nFUjBEvCVy
lBIiDgTdMRJKSsXvwV2U4YrpzaI+uQZz5wfx94NZzuzPVyqOQArrZHPSRLCGRAPi
sSg9tbHtyUXSvs76xw5H7hZqYfO95Z1fWUi310FTXtbp45ikguoI0zwHgXCkSB5/
p/HqChXoEVArMLhgam5yK/kIMfopMjo5uQiRgqupM1S988s/w8NT+e3+migvYMkG
RYPa6avuUANJssexa3JDVf2A5gNslhRqf+D5ceptMHYoXsc0wjVCgpX//bDyrdcb
`protect END_PROTECTED
