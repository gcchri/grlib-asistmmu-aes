`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wg/MY09WSRzi0Bh2YFEw0c67d4Kzczx+/2ahnkTDheISyIkVuF/0Dt3hWssplF+v
qxWDDOWr87nXVwgC8l0sKC2lf1hEom/xNPEi9N7/DVS5Cnnc9MHM6PIQGkS9LC7K
aXxIEKkzFt7q4w+PXps60pALBAI6xc3u3iPnjR6bZpFYNnlN6Ju0/rWPhLSKNY3W
XiqIz8HLGalHGGvpRvksMQ2fJX4udVrjV0U6YRi1nad0DbKWW4FNkyREmR0+F9Ba
Mo3QM/6S69nlvFoSjyizuDDERvTzRdMKGOpupsIlB715mrn8QFhsWtUxF87CIksX
Exol49rw12dI8HzuZ5q+D61dHd1M9Mn8fNBsyo2RFd1T5hhwLgtcwutUa9KCAsNJ
pBBWOAphdIB3D8n7wLR1uHlCHcGcrYIS+xOgLVke2ccNKjEIHUdtsS4FIbwPxGNo
fzfVwYBua3nnRjuzYbkKARfJeSjq7TGa110tYwtij9jxNismNIv/JC/kJ+QSDptl
H0htvwUmbcsI5DEMm7E3KpesnJiLrDyJKgVZAJfKkPrnqfm0dqJtqmSE+m40PpUX
`protect END_PROTECTED
