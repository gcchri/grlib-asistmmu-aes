`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5q6W4Rcu7wVKrh0DaKzMFoKVDKqZKNth4+5w9mxB7FDBsNaAa0LcN7Yurgl6v+Mi
Qt86/ouw1kGiekhDVvcj98e5gCUf0vQ3RFroPn+Mt9lUIjx92XNPOMQr/u4spCDK
snUcq4KogJoDdTgkhHTj1fJy2ZgdEp1Gk6PUzZfQSyPzqUi/v8D89laZ0re7CeeI
K/kQzZTJwMJ6U7gLWmiNpB/gfEZAJAJIgAfvorEGSACNmlwymY63/HoZfFulzIYK
apUPO2ULvMhB1+TQx0G2xn8Mbk/Ah+N8dvUjqKkYp7BtMiPH+BHcMSALqY7l+7ek
AnQz9yPmBepGks+jInBAP3FOmgYq8KCjr2KAGHK4UdH6k0lkcfGIC2PI4izGZBNh
QkBvubu+6x97p7fNe+DVSxPCXA2G1rMUXsW2p5HYEY2YDzFKTvolIuMz0y2Jz+5g
DfdypyYZj/IIJVdZ0BgeZCC/0WoV1N5/u1fdSw6zMZa/N8E2c0QNUdOmzntGQtNN
sAzshYvm4WABbt0SFZbZRkum/vvCqNcn/u6kk9TZL/p/ABRd2DntKb5voUI6GUbj
x/XdqXEg2a4QRJ/oyLFpYTDkEguLDn69yP9IuHgcHfHhvF0BVaLQCUQ+sC9u9Vqf
0rDsehIX0Y2bEVkPTVkukxYx8VyX/uFdojKNpK7+CXvl1C1e2VCsJYF4DMSzMh07
4BY4FBmjTSGWnLAnslwUmu5E5Mi2Bees23gFvy1DZUC+tcbj+KdrIXg6tfITVyKt
RgTsh8Zf9BXY3QpFOrgWJN0DBoTZ41lJEBrjgRCnmCTl06aAuWsNL+N87oeEQxjH
He/AG//bWLc9om+7j0OmAWtPnztooSH54Deo6T8je4DSwXJUqduVTbsmJBu92OGo
5dLb6TCmldt+U5t0JvitnFtnGkbgfwbnvW+cJamwCeJPmXVXx58KI5bK1rHB/2t+
ZB4FdO5KEkPq2N2K9PTroRbF6zFoQJeg1y6ZglrD/ThFdVWorCqxw6Y27DOzOS+8
oFLfsRVu8MOQqTzw9/NZP5trpvXojhHRVcamU/wQndDhZTNJTZR1Q6vPnQTXndLt
yuoc/+YuNaIgsIageeHZ5dzdycG68vrCmaZBdexTwqRPEPW8hYWFaDBztWZ0Q/Ba
b4dbxnv6o5wFZAHPdmu/+a+YYBGEZqVRDa0WvVUewN1jTxpC9kZS7emYDbHKNGRk
opKD9zqw0aNaYGf1z5Tyfj+DyyPrU4irGsopllnX1M6tZNo9Mkp0KtTPaJplPlNB
90qcyWykjsD+nr+xJ2wsBKzIGtO5DDIZjFtlhYH1UD/Weu6zl71YoObXaoBfvTzR
ozevERv/XH1unqPWAWj+58yF+SrmVhxf4mz7e4swH6sI6sAOb1teuhxDBHEw0TQA
Xyix2a8u3oFI8fwUS1MLqd3u4nFqfPazT1Wl+RQiZ1FNcluYb24ezYbDgFcfUf07
CXCP9UJyr2d3d5OudI57MLQcXoVnGTX+mh/oB42Hs57PamluFh5SgFJ3iGgNIsAU
HLoPzTjs/72qiE2LUg7qRHa9tBZoS4XDLtFI5obc7f+da4K9HpdeIFRsvxSzt9+k
y1Z+Tiw+5i9bXn3qdvS6sj+8YOlu6k2GQn0vPyRpoVG0jD6Ox/88pK+R5Jlwv5Dv
UVPyUr3Y5GFK3lBcOVXwMIPtP6w1OBPaInhAWMW2L8BoiCQn5Enz+a/Fi+FJYZcq
`protect END_PROTECTED
