`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wk24Lf44r2WQNxen2QS/e2Kjh0f0GZb7wnQX+/S4FZ+anb19wMIvdXYwtHqiKHzK
rn6mCvtO2aUMpVa9OUzo+SWi5aIGgSlHTR/CSMORJ2ESVho8B+EvpBo4RSmzg1zL
20b1YWQGSN/ovbE01H2wtAAAvV67cQeNiPqwToy4jEzBaQLIgRjcAyx72/w1pTJN
LtVXeKIyEZn60NT6SuZd+7k6/8IjJA9iQtkIVL4Q4Fz2lXteVe6ePYNrmafxhCu8
H+1xnKcoKAHZCO8ZeSeJsYTwq/UvV5WwLPDLZE52VKVZEa+J/WIWOmACYwdwwTDd
h30XpBR5/olySO5gToFW2fmnI/LyLNXP0xTMA5IIZLNZqDRtwtoEDtc6hb1aA+VM
QUz0T5iqAecj3iWx5QuyqwaK8/cGmOos5aWxz3hIfrU=
`protect END_PROTECTED
