`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N5svICRetrjBzfs4vD4NeWAkTJwdo4mpsU7x01vfv94rST/gTaafkJ22/Sc+fZKO
+61jzwMVbWDhCwHhMpXu0rwscGPK7FmkF5k3LfZx1c7qN2J0am/TfNIg1AdLTsWo
Kqrtre0gKjozZSkocKdTOaSx4gRJK5Wm+zlTtKdppiM5pzbTins/JO+0qWlbkkf7
3QWKgIh4v/Q8lorEOZ8dyeVrWoN3wfRG3musomGWeeydpv6pfGkIdMgJXObgakeP
QyRsrL9DezobNhValTrZ1T0HhyNuusPo/JuD8/gmRAjzCdUljhPj5D0118GP/GzC
XvHJsM1pjxvNMkYpmludcz7ioBzb4319WdCZ7r+Ws0ExjjiEADYCMXQt1t712BW8
Xp629E8Xky9PWfL9LOJSmIkBbotgt+edNo62hQNchM2Asf9+rq52ePQ8ZrYoJPZz
u4aPGmM2eeEByA/VoHIJQ1s2Hh/WSIX5V/8t2Le1Png=
`protect END_PROTECTED
