`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WiaL0FgHY0L9AKN6c7Bm7rmH8gN0R7oxdRwOpxI5xqwwfcD7w2PX6tdWy7bUs9Om
wG5J09QxvsibSEN7JwelpY8Tz0pfefz7yV9iuwLHYkrhJoJ/ERGZpjvrHjY66mmq
YDWS80czwKstLprmhFGqPqgrxHFT3UgwXVXRS3fOcI0vyyVcO8R58vmLrrfO42Ib
YKu2QHr6K24KRy1/f7GZUZHl+y52pZbcU3NNpDNMvbY4TR0ZdJ2srzQgj3eEIq75
ee0eRUvWQ5yTxdrxlG76CzoSzgmQ1DynNEap4cpnqdcjWryIRMloqLx/OHft8+SS
dtOYHicoQZYn5x/of+8wUcq2Qo09sx1AbTiygcN2gHGT3IU2z7Hr8KX2jkuYgbZ9
fuf4mZ6vig3ok5/uZ/01O76WKEk2zmkIVchlsYBtWQGesRGraSlupj3Dm9MrZx7Z
Lh1u3d2oOfVgK4wL+l5tkq2zJ+h3CMtPUTVTL5j/m8iq1wmpsUljDmIgU9XHnJvM
UVAukhhz1MNIOIjZy/MP9z6vbfNgbgghE6/A4Jra4I2IdmdI+cXgdOk4o/GizaLl
`protect END_PROTECTED
