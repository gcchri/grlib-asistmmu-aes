`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D+6ga8a1k7ZBvIg4GvSGWqO1MHmgaVjiE6qgWobe/XbMzU69sR5bP0xlMwLHGeNv
v8yu4qkMc8+st5IjLRuAUnRKK9e5DT36JmPhJAd3k0NwH/ld9/poqajDLZ0mye8W
ga3USXwhYIcZqGj9p+P6mIR2tAqD6mHJy9xpPgP3attbj5zRGR2g4griagUaEyT/
ghqHSl+DNpOeFlqUVXNWNN+bCckJ4H8/DkCHS5tvdd/BhGdCZoOnvZ5Zsl3lJcWO
UUUZA/HEpFLS4TB02aeyhTSJJphOK0OdRhnhhtiwQLtOrcK1V+MyA8NTurEO8e5+
lSLqQ/Xa8m2azRBVJbtiYFvsmCGUdQmwZNwMHeJNGdvlUeKJq5SVDA/PM/bv7OrL
Me4fpi6z03iY9Hz5YM1ziMaGGzMJfbS4vOT7GdDAv2jhVAbZeJED3pJuChgGGUaB
lMLzsS1FgDndQBqxthJjlbGYR/o3z+wDbOKppab5K31J7DgBVnt2lvoVVxq26kMu
lVZoB1oztV8rd6o/WbQN1W8NWK+8bmuJDtEXUffOJwBFI5/micZo/+tinMkYUA0c
hLf9RuzTs6EBTJRkf0ou0YYQOgU03jbAHQkHy/XC+IGqsIjAxLs3yJ1YqPhxAti5
yUs16EtbXMJUzHwSzzRknpEnd5Vn6Rb+Z4rCkN8NE+SQQsGyIlWCOD0CvKszOkHL
8yn7hQNVyJdQgrcDYVr5qAaY+n1aH7gTg+iYIb34wSYjr7q2VjzIil+vIKI/aa9S
4vSNrYa0RwPOz1bwYtSs5nKFpQaCh+A/+TzTIecqla4ewAWX5F+XicKE9c8MWIdA
aJ32R/iDeurlK5mMgbZfspNtvNQ8bwaXFIUQSfk5qEClhjrxz3RveVBR1Fqpfl6Z
DrmxTg5UUH4MmQ3TqcNjRXcoVgNC6nkZh3cDifbQnFGY/JSJfthUH9YRXLFgqStV
1qGE/uh3MlVdPw65aTqfGTApav/tq0ycNW8uPqVnpELTtEIInMvmmFB+sqZVT5On
bDiKufted8iVaJgHwupv0A==
`protect END_PROTECTED
