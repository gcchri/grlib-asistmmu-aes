`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T6y3FDXkf5adhypQfQjWnVgfYTQjQ9Punqfd4mVjSOGbZ52VPZN+pnGJkJS1ZUaX
V4WJHcK1VX/8zk8mT48gGd17x/JmnDIbdcXRAmfFK1lTzmuVBBsCrz8Ptqz7G+tr
BgLzHgPHjg56/rsVS8pUBbbss9aWd7peGD39aE5g/zZRtCcvd7GjTmqsLCGyJ6co
cexoLKiCBOV3ttCJiZcJKqGd1NxW35bEf4AKOGKjpiM07NxGG4yzkuHKSmRln53V
5eeVccemXPiJKiGzk6Kohm5u8BnqFCEubZkJhOge/QHuEmo9DcmJB6ruC2/VXqrq
gkfKLbQ6JeJ71AxGEZBhmJS5VrBqnGwTFgxJkh9Ysv7qP28RWJ5LQdkv1xFIIycs
BCpZJJCzI11Wlfr+fJYFZrOYSk0gtsZ2xhosqpBuS/EImDLNRarrVnpWPt5SfF1E
Ci82udT2SlrgpnUwnviK0Bo+o1Yl9CaQJDnivTXyle7Q+h1iBCfSjVbmrOLpLcfW
jAdh+gK9D3Rz5aVxS9wE6jt+FKJYgmSPMWanGSAn82zVxI1Ok9mhUiBAdSGczj03
i9UyvWCWYauEU3pIum44Vr/lKrCxFQDpfEfQSQdARQ28FWGrOy2a9uHeugxubWu9
5LDIYfRSmY8WMqhMXuCkEIfa8PLUmmE+mu4jXy4vFZWMwm3dSwTJhW6C8Bs7l29C
8ZYGAZSoMHVwctZgCoESgytYANRSdghHGFBShZjwZUydWhzD5YY+2W9Rrwh4aPu4
jK3o/JzigIbvw6KKTwYYihX4eDBRqkFsEt9FtuS3T2i4BbVyeFS2z9k756Bpjp0y
MsgS8dbRkMmJifoQk+j784uTc+wdimgmvcLlvA7JENnR/mKA8AvawXlVtGRQUImR
CcLG0c/xIz/6BBLIII+rUi5H45sS1DIKsLKf9nvCUAmqbHxfV8eW4+xe6RpR41C9
`protect END_PROTECTED
