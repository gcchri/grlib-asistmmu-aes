`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YjhdhueCLprxz0qnl9KVvnmhcucZx+KM4fZRBB2wRi8M8LG/twmBEHEkU4FXXviv
AZSTnWXoD67o1IOx09dn0ttxohdWRqNVIsmmxMl73nxDnv+4cQQm0zLc3X/3homc
LbQ1agQzyeMS1eZt9APdMa290crnBe6A56EK+wh3BizfJ8Cg+DLSwFnFXhPy6UYR
w8r4zBLdT1oHza+lxgItrA5/rDdwHP4bv2F3nHiHImj9ANeZeWzmJAZHD/lfPfRf
w/eXxx3LHZfrKSwtk2sd/rpq/16C8+FDSmp99ra37KiItBzhW9EPQM6I5QzUsct8
CemfPNOBk2tDYAKdlFkXnkSKJ8IrIg6mnItGFXoubxyHvj+5WJ319/PMdsG0rq/F
`protect END_PROTECTED
