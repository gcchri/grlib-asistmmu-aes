`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+AFzK0QxaOMdWl6TMh/jyrrJysTl7pdCGJqmkOgbcRMOHcq+pwm0tMburIMJH71E
wNNRWnQ934xbRbrTQd4GIawM7XcyxgCTcdC820yvE4gLVWV1SFIYUY41Z/jNYSw2
ilrRcbbBD48kT9DwDC7wxLR5ALav1q4GtU2BOfqfPueS00fObFxNDFoCq98d/Sp2
H7CbIaUR2o28VeRQjCtGLnNbV86w/ZbT3hyAh19jB96hM/NS+t/HcZcScdWkNI5c
ImXcVwN43QsUASmPqVITaNwbzQjtcIeEBhgHQlCvUyA9stRyCB1va14yHhurKIhl
tOYYxt9RJsZQ0oSMyu7jZA==
`protect END_PROTECTED
