`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HrZO88+wYIoeqFHiC/FyzzKTi3cH2jC/N+LdaBDPHZ9dWnoC5cFBYByyBADnFmpl
68WJOXYUyLLH6K8PqTHKcEKpO92ZgfbBJO2zf76f0DsSz3ie/UdvMozOwhMyBxA/
KavRSHvcQOmW5/UlrQyYBBiw0NfsD6E3kDM7Bvo3DwQCr8p6eKb/bGZVRQ5QlmYA
h5wMKpiJQRF9LWwxjClcb4T0LWYDNJvWvQhAj7fLFYfl2F7n4MxvNoPPVuMKOBxe
2JWNV9o6+af7ESAaJ56sUTiM/yp52TKeLrlu/WZB1PShtX11P9yIu5BGm+5Abyjb
eDHtGoasOtgXk44y4jzqpBJTbv7o5ZLeMFmPvWFTGL9tyev9WzaKRv6GdHJsnpaq
5VYcoR3ECVQtX+A9zVNlGaAa9F5X+4BsY/NCPfRviEvCXjReGFvdIAqFj5y0TYvK
OzqUOJR7T79/zQjXYXpKGA==
`protect END_PROTECTED
