`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Hj1RVyGDnPxEls782Axb/DNM4x7oitO0CSs2Q+d8hJdeblx5jFqEWqYv4/5PU5R
j3hBcnUPRdTE6r/X73Z4N8mPs/xhE+byfmDrNut4nFCnQECaUCGVZEYZlhgEbNUg
paqLT7Lgtv8Y7RzEsLZatyYsXBf4BaCGr3q7AGwORIN88FamAd7RY6glWMCRgYKn
SUzdc0WivTy9QcFQObD6BiOUV2hhdYsXUENoFi455RxpoDFUPMaVbbiguW36GZW5
yT9NQAxmLsxXlz1Oa56GVht5jjrcDTBrz2GESJ6jwZncifZgTwDs9G/oA/gg5H5w
`protect END_PROTECTED
