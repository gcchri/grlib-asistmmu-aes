`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RssjsZzovkO3oAhyDHIpeIAdOVxxiVvIv+mDmr2+fcfqy/nGscHmceZDQhJ7h2DG
pqNg6/iDQNBG6wMLF8zvQkSYwcULluX9KDis3XSccUeTZVhIuCgLbXDd/e4CR3UG
mSdpfHfLJqDXZlYeDieHOKlfmz7DGHgUP4xC5MJjqIVE9UFdQWOrooCeIKf0b7VG
zmZtCjz1uFTBWOgaAtUj3JrFMYY8y4VgkOvcBX5jVXmrIq4qcs53bv+62+9rZqgZ
o4gS8z+7P8G+iO4jFtLaOlLcO/8Gfhnwpc01Rs9LCt3TkASHibJEb5iiu0IrMN8J
7ZlF+V7x12GUYouabJpdNeh4jcPBHw2qRRrmO4nLSlGR3RprOKCJtNsrcLmCoUk8
in0dFf3/XzYJuYSd3k33+RS4oc5NoJhP1FbFYxSybW9NiUfxhzrSlG5ZR8JtjKfo
s8H/75pBKwE+m0oKoaBs+LcujP5ABKLcfpf6hAsA89R83/F5aDIzseWzml1PE7ZS
7DS10+tvdiJzN/o7rFgEL4BcXSLU2wW2EuTIfX32TzC44DXjVA7sEJ+2C2yY/00R
f4rRffDWaVsSbxsQXJVBmPY1VvHY6Qfd87Kk073hQXzqgCMgb3Kdeqg0JuXI7POz
P/p+S0fiZB69rSB0nXRnroRJuedjQgCQvmbY7/TiICPE3GTxj4lkkGcxU5TnQK6s
bQ+gpWqd/znEbj0V+I0uQmGkxqS7cFTyLnYj/OuMfCVX2Qql0QeLb8yUxvxP7Sph
+teMpB5/gL9lUGKZIHchawJOA55Jda2JuS0HUB6HUKRh86dsaC8Xaj82Q1ZMkWS6
bF1BYRdPMdABVcySWzcfGEdVs+htytr07gsPuCaHaX4qk9texFrD9UUAYq46KMpg
52XKZN1dFcYBDVLc9cp07Iqva/v7rhy8n05u3dhDQxfWy2cxCeJVJFyxh1h7aELT
pekIvcI7ITMl1tXDbl6U0fpRxgneTrCZrTnNuna7+Fb9f9LnTRf622oiwfC8Rq8L
O2gyFEl0CojtIBQy80Rzs4PHX2qa94RuVgD09CYj2nCC7syDkRPAhMBXNDL69a82
85m0h0t1sWaYDFFqgX6tyqs8+xj3kpMi9rlTvSto4tAOwen/kn8B4McHYaA+CV64
CRzFeIAwQULBSc6qakaoSkH8WY0JRqM+orBoW5SDQdjiV1E6evhGRool98gP75Sg
MvwcwDrxtV+uLtnQmcir3MXeEAyksg6to9kRrLmEIt/pooLKiXwY0vPh8Yz2dyww
`protect END_PROTECTED
