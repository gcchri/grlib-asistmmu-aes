`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zCIlNvn/oixP1ZbRGkM7VV6eAP3MTIyKvSPpDdLME0U4dE1Dl5TrlF7M7RAxkJrN
DtgMaj9xfccLA08h1IM0cuM9tQKN8Vi1AZDu3Z1lhs8BKQrZvFIeKccQRtY458SD
Cp0VLARlcLh3MJCL92nqmupfumhqDEkdn4v6kokcEMYzanDkhc36FurULjglWQdx
EWYCvPmRzyFLiKeo84kxCjv6eDbE3BMJdiy9lxloGQ+tHaq003hbZ9WeuPk3Ok6e
AY1duxTL6TUcoaIbJ9QB9U7JMoxZBifPG5lpP2AfBgcUd5ORf2zh3gDUVMk2aaBi
B7+qNK/6wAn+ztQ8fH6zrZqo1CxDI3kqZeBsXjCwK+70HUJfSb7zzmAfzgLvQJGy
VW0ECplk2InqL9TnXLAs7pM/WP2/GDSuEpdvFour8AsSJvyRz0H1Zd7pcXXB8J3b
`protect END_PROTECTED
