`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
behsdGYlUwOkrJTn/WSH0T2M4fXKuH3cIg4iyqEtw/VonUxVZGuGuX00H4dya2P6
TxVmBh63+/XqP2ojGCstRQv1lsKzUX83glAbt/HrLQYiEFoI+I34X9fTT8xnqoyE
7jlUzuBdcdDph6+PmFrhHFF0GFj/u3QF+pTvGHYDCHJCY0TAnvAXNPtAGX1Ytl2t
MlBruC+VtllKZhH98jswlWQ9WukwUi1G+QXWmXOb1XYY4sVGrqa+va8VtTeb7oOC
veRJZaZraxfjhZLERBsQkDUM/oKkDZgqlh/xfM2V+USiK/8TIQSciQHPkrTRHoP9
4mIws9hn68VVR0XfiHewaWeuOYlj/XcUtxljzXrIN8L5/IqHIbn8HM9XM93YQLlc
t+zFojnGxgjSJBAKS7VVYJfgktu5KpNEGfFGU0bHcQyJi0a0D9XVBKdR3ORBchT6
nGaKWtERTn/UsbtRyx5lWut8n/JXl5m70Ysps20MjDvPs6l2R9Y9EMQJmGcrmqjE
snpCYoo+FfPuFiNTyvu4PRtrhWB50jV7EEL+Acpr8ksfEz6DyaaAARf7WY7+MP1f
fR6E7Z9zkL46CVWjMur+W4wgKhqj1GskKMdczSkX0CnnAZkhzeqBqjbfBCYI3wr5
AlMqTG+TL0ENsi4LEYXOJZvc+7kTooPtXGhNx4UtwRexzQCCMzUgr2Qs2rHbScTC
uy71j8UDJenk9h01CLeU5eSU4IUJE8mWxjHO9r5momqzpK/DZ/UgOkOoVn9AUTEk
li/0QjJM+S9xjC9viqRzJ+un17IJhcRHPZh5DhKws2smNjxllhny590++MsA4IZm
PB7sgz52q1hyxxjWV267vIW9S8CEb76HCLzdU25lD4lDwTE8uodqem66+dRvWcN8
+pOxaOXCYiFfSfK3snzJsheyP2f6mGfca5/yqZ/V9aHk7/Ou70QcU3yku7DuXLXU
4Hag4tvKTFGCwKZQpyDFpnVEoYG/TDzzEzf5nLRlHTyPYJ0fkwUfYlQBiegg/P1X
edicPI+TgnjPjhyv2y4mI0QDA6SBX5iRlfgYpzsaZ7cyTClkiptMIBExHyMnMmNi
JWtDnmrxVKx/j1FRoKVWWfyVsJiP8EiZVZyjTiAZJP4QlZKD0++lwKBVis52HwGh
PO312xcpaCR8vMMC7Tw7jMOZs2HVOHNNGTSsHseXpI0Jj9IJ9hxe+P4zgypsoDE9
OpqhG+dNzOaOBBq+kHm6lrDZbCVes++Jz3rPSGunRmMQvMnxCMxR0zrjORPEP2IT
bLMiMy7BmAJs+e3mGlj+YJJxNMFdS9IZoeZ3YswXIxgdW5OmzFCg1ftGSb6Wv4Mq
0mydgCIJ7rgizGYZ9PD8TyvnZRYvQufQ2N99FRCtF8XCzg4XyTHJtsCcVoYp0I4G
HJByDITThg1EK13h5fvk9DOe+L7tIqO28k/xbeLJUFoR4FCyGXJqutdcD6dHolYx
cPFQR8O91J2qv+OMVbj0+69JFDrKrsj0yA7Xjyq/nN5Wylogp+p2Yw5RZaVsTdnV
fpyuerjGzNsDk46w9/TtgW7kSAbFzGjFk5+hP+C8MQLmLVNskcIEGRf7buXw42G0
AQ5XSyveJxOgxDJyWukr6sJBMrP9ZP2FqWHF3np/ojUyrIBjGw2FOLTNmNe6XTM5
oQRQBKUSNn0TrWMxHyog/a7wUAx+HCaaDi893dRzeoZwjDwqhN7Wmnq2W8WDjWpq
wsyiI6/0GXgttxzf3Yq+73Afb0kACVQbwQE5a4iMHdNIuaGgssiYgFsmt9AnVKPi
J13e88++dYQCQLi/RUuBDs9aVQ3EARQdVhWzM5OmAr5pXoHGi/tF3dF6bk0FJEHO
LDz04jxNJ8QYli3BbQvgrMHxKB0Ey9bG2pW1M9ELVZtC5FfTUExsm4TM6Pwc34v0
TCV/pcfby6NL9Lo15EzpGYkqXfNvFNc8WUvooZIQtjY8yS98awKQGIx6eC/uKG18
CkDCTqIJVtPbhgvlJQat02k69iNwFjJT/QvCpGKCGjYzlk40JNoXFSose31zwgwG
U0cW96a5i9XWTXRezpM7lG66G+VYxUTcXYtayFyQyx6Dd7E34XxxnzABDibnaplR
tsGjGc+k5vuuu7K72vh402YqG4qmLuSf8vk6+hafh8KGxfVD5rBELzOEU1Uwmdif
avxYIP6QHySw6a7bRk1KgB6k6GIodpP/5ztXuTftSVmLM8kUv26yijPgFZv9XnjK
EaixA3PE3a2Apiwfdu42vdqt0p48wFd+1AcwgcKLQlNn6ZDDpsnTTk4i6nwGeSZ/
0mvGP7Iy+NIe7hRE0qsQlOQFlNQLCnJgaCehe034uD8rjsQtbDBTvreu4+CDQhdG
rtuBwQoMrxh1KsW5bUszr0o0wN5ixuweV1wwTK8mEdV6QStFfKF4n2Q/HCh9gZkh
bS2lmmyyqKSMaGH/1SVW2lBh2BUtX8bcz3F8z6sIQ62zJn/vVlLFsna/0YP61O6M
rxylYHKhLGmL7UUc5DLzKcRiIlhLAkc3uJg0ObmHq/YOoTsciL4laulV0nuA9iRt
UItRbvFejR9Ik6qKQgWoJGlmq5ac9CzPCmydqaPXxzBSgTW6fMt4idwbn8xy515N
vdYKK5HsiZBuZVgk9m91qMs5o8+otve5iL4AkUGVD2fR9Zy4/VvjVPV0mg2qvrLR
qLMx0U3GBhUgYH7bQN7GwaE2qMC6+s9Zo3P94hanyJ14hdWHACMU4UfePgbn+Lwm
fAcgrYW1DoHXOzKoT2wIQP7/tlyhJpDj4aNNmLmmDn2Pi6B7Z70HTEDJzkbMX5W+
lNr+JpIPzBmN8bXKS/Gt8/yr9ClvMN16jRQKICBmx5M22MLdNm1tKfqYs2XvfEMF
iKvf+cbvK4zHTbfiG0N6zGkMZXiBGwnhc5HpW0YizEZz7CO0L3e6aSnKJ+R4Iegf
+vaWgKPbBEHcXEa+TWl4HHxVWLpnF9IUGM3ceELAKSsr/x33ozeU4+eQ/nP1BhYM
RZb6zGy2B2HS2O9tObYZzQm9Q79jUWouEgz+kx4yubSbKDYZqnoF6ru1l4G5kP+d
35CcdKMfJZpjIfvzzqz95xzZ/UNT086rwH4qy2PJtsQ4MWnoIsBOCPuuhvjnS/nh
WQ/hAg50amdGuSlCh4dRErK/3/knne0qIrD5P0kFYIR+OOsx0OAGoO1P0vxdo8Sl
mdwew8nEsJaY64XdoTIeHcXaa+Vzi3j6zx4w5rKh5peGbcZIjTKobJDY7D3BPJud
2tRErxaUSyd9VlETky/W2M09VPDwOhmSOu22dxUVVo2gkz8gNONbRbZ2vvMebSMu
XQj49fSE3Jdk77BoATGJwq8MVJFL0eb790ftXGnMX5xrXYUsdecOnQ82sMjJrG6E
qmF2Y7Als0PxQ5PpJbgBTua5BGT8TSasGNmMRVFYoqvZ03DDhj7MsIh87Xz/n5Kp
tInrGmFmdMvPYw++BUFD3POYRAcobQ4psUpnkNE914uJQkmvONRuAQCdQ41L5OHA
C/oiWCEVA55SkDswQmqYrWIfCf5LMnEGvb1bU0bO4TJWU55hIv5xdXym6vU839jS
BM4/UOMBlYs3SIyQSeljuV+0PsSLkdOglBPq8Z94lwxDdH2LB83Vq8ELdCpWwB2R
vRFTArNgBr96dq1dRVe0s+yZb3/iOjPenqolCEswT9Hv+hbvBQXves26gVXDAZtL
+vApvODb0C4eCHZN3bLRpT1CtFDRE1F+3mml1G/zSZmQJm7Yej0/DhgTiN4WPxBc
oWJ118zfS7w6rx3bCoRFADw7HGKdapHUvZlBO3KuJo1eyqn8L7zaw1Lg5J+oMlEI
MwjNFb/sqWJ6yCX+1sNBGaigzPaLNx7Cc8qtNmhw2O6ZgdurfpKCFWfZm0Ip72nA
mEWtB8w7iU3ieyg0k+P//riBW8uq2UJQFR0MiCIP61DI3MXYfA35juRYawwF6+eu
dKskspGYd6kSEykqu5Y40BubazZThb2la+pMPxF6VZBZcVuFrHAz4PZj5dopNn5v
4VlFMOrbVhkZ34lQvGiNrhK4ffzrTKHHaSXLNcQtW7Db+HL7FYl6zAcgS7ThroEK
KpdjI7j9YPyLqkQdcZEkEQ2FDQBbmbiGH8gj3ioJBTz1oBaBO0zvDfsiqPJJO7W6
noLSrJlSdDV7nBFJl+/QCBNBDT4VjyS4SpH2/5p2syAWGBJwAGWlbqNC2gDpZMMO
Fjvm9dYRZ9FOGr7MDssLK4bmtjrMnDvXdPdvnVzePdi/7v95/sft7gVFlQcyiZp9
eTpW4rijMAzLVorAUF4bYKmI3Lhi7T0b7WBQaKUxKx/tvejNutTE3NacJTFlgNac
SXYv2nXlpxMvcrK8oIEaJDnt6N2zB9N6kND9u0dpRAcp1B86PS8Lceo9voqArFDT
+SMv5855tOOXwMv4yQ+3S30R6V7AUILP3QokcwbXh+XLWEG99UlZSne5+WxoObFs
hjzI0aFhJtII/iWqHNbXvFLwe1VwgV401WiwqsiPEGRBVSK/1CilOhJMiHMXvULM
q8sUIFIgf86W1YefDIAcS7TW3sPy9Wah1+rC520l8EF+WI3vW1RXdUjBos2La9eD
TETmA0M79mROcHmypuTplwmkyYPBqw4ML4ahh8whU3UYo7QLuC3pzPKfsKwCY5Cd
EBeGHhRmeKLUJhQtY3GokIrp7FZZ5pxFg8ftqw6MaUj/blxUviDDiffNC1XBbGTG
KHVOTgCyi7wpVvHVGgnm3cxliPZqemVDl8qfZEjDRrPBx/fe1zvtY7CSn9ZmZfQB
CbyzStwKMjfTDG5I+D3ap8x/t9LoI37Yqke8JbCJ7EHmKKgiWKE26WlrkdVzGQ4X
MTJRENcKXgAcKJ/XQqzzrPE2lwTFKniSlk2vPIdK+TL6oY5s48blwP/8LgLJzUtP
J6AN/nnFMuIn+YqixkE47UEypGaP9WJ1GUpr+hJQr5VNSNGfIB9pJohkJKZTz3D4
siir5huBetR5n4mO5smBWOZkp2UUh5/eDG00ojbkWz8/cdtgRbl94vYGFRvII2TN
AAYSHGukYKUsB9rVhEak2qSpuTw9hcSS5Aq3iMp3WSVvbpUUoHiMAZS2IsQrxD+f
JT7SXMnzpl9xoLjUSDYPYSbH01PI4Xzpa+bwByJ0PnwHMhGMXABpQMnOWDrG1zw2
tPd6VdKA6MI11JTTWjMuAXWwyQtLusJCSMUSK25ZXk+vFA48iKUE50Eo0jTlleJV
Byjk9YJy7MXi9DKLxHu1K3L9OzbtQ7jnj36e8HM768Yqd+9wNJ5FH/Gb89RJD7TE
oi9CtTrp3PdU5G0fcPElrxCJotnns+5laWd+3/1XxuPrF+VhC2IzFth/yqkk7itK
hZ5u7RzFL4brbTxKopzzmdZQ2DAMikqXykxsyj1wL8rNws11CVnFF4zaq+ms5UJa
qp5GBjrXBiOEXAtKhX6dhHmw6JMg/MCXvcyvd5VrKUYZYP2a75uXKcQSuNyva3CI
9gOBKvptgEiW1oRdR7BCZ669GDFMcSQqvdEBd8G6Ut3DyAGNGqoo7L68su1+9s+g
ruSn3DL+EmBzHxr+pf2Aq/vsaQlflUavgzHYYtmZFrsyrjdpyubK4+yKsu6Yp9gO
Fr4X9PiVNP7zM8kBrjBEELG9oxoz/imtqYIonTBix3Y8dJQoxlt9uuXY1SGvKZ+O
6KNDvZni2gEaDecnlyD7a1CXda9aO66Zrwk1wgqnsaKSXavTQMjKLsELfwx9nvUw
IVskHAP4RGe1xFLeivtJxESxyOm45+80neyJ7HVlfwqe0xeIrdOil1JtK1+h4PTG
BgTKMjMXpsCDpxvSxd2fYZMak7l+vNBlL5TdW2KBPkrSV6rkes9YzRdgd5KySX3g
R4VBEqwTO0B00ezlWW9szuvm8JmSFf68OLKSS9ZN20WZ1TJncSwPX8SP5mudR795
bV5ZSteaWZot/BtGOxs25gxF1S/FF81jZ3jHTJisAz9/ULpo+nq5/32Vd5tLxMiy
Stg9UVzsBY9Je/Hx76Qi/PkAj0jcNq5R5E5xJhDU82/Bn6GtTUNTdQG1c102HyDs
bANvmNtTYC8PMjZBkm4p/5x6PgNlaBimCGEZermFrx9gzrp2snfpm+c14gH8JimK
Nn2qqMQ/zCpdypUqXNJlJekOKWwEzBHJ2t960boAIBCnORZxJStzhHiLUhPSLbP4
Pre/XBDAYO3oYC+Gwia/7tZS5TcKu2ka5jWX7JK2kSlY2A+NHVOreGKZpWR0yzfY
NcJz0+BtSmp8fFGJ4S8FYxJvIXcI/GYOfGjS2VbOF5Pi34L0Lc0GBjjiNKiusnlu
zMPpCsWpej1THxRM8vpMSVRq+y0+vGNCMKlnyaLKbWL1L0TJr9Iqle3YP1g3SxQw
T+XKXsm6yOqZjMzzylGgtqEPfHtIsRSwy9m9ux9ItldiB2Vu3GUGrvhxd3TdlkLr
dj507yFrxsyB+11U4HxSJp6IRa6muOZGPmDfrYjqLlcSILbjTfOiZVI5b/5bwji2
botaLrpmjLARrZk2oxd7hC0zIVT9rnSyxcGpbznmF9DwF3kW4FAKj5v5FOwY5IPc
MZY4rLybjvwUcfw6BfnHn1EiS+FgZDnehFhkJr2b9DjBHtS3xq1oWz6audGXv9Kw
wLB9t8M8/znpW3+8PwJ67xYHVxpIyBpoQsomGzjf6Ns/r9sKxKr40DEIA3WkJokK
g+8me8LWIxTooF9/93xqT6dOpqfLmSkb7D4KNnnT2Kt23R2j0JJrk6oEL1ppzfGb
diI4Od6X19B593OBWguFeLHjjXefeSAYydx7aqC1qJLZfCACKIYmW8GpulN8uhoP
vACDp2Pe2A7n+H7RFb4tFt4L6x5ZJZaKZOJ/UTya8jWsnBLinitMU6Iaqa664x+X
d50GQEyQGmG24euK1CGDhW6Mk/UQagq3k1AdXjeYjdh0EL03lDg4uG98PdTxoxfM
FwW0T3L6LBIrkYy5cy4OkntZJfswlR5b+z+8PX1YkidU7rIMGVKKdbqcFYFcI3w8
a6Onl5mri+/d2uond8F0r4srI/Grb7TEdNpiiskYbRIu8oNTUUfUpSkqbK+5DhB0
d3WHGZnVT1+dDOPJJV+zUk6pL3K2ixi5h97gbYMvy88LoN6Oqh2aZ86MOltzot3Z
2sEmJSpVt1llXTvUis+M9dBOqBd5h51Q0EjxUOr52bjPh+hyLKfYW6Y69oNRgItK
ccmf9jHzR0LrCRlzFS8p+3Jib3xZLbCe9rFp7P3FJ1T8XQlWvz1Ya9/YcRgD4QTx
zRsPBxtloRbDDmvBIsl+YYjAAWaz9iBU4KCLLPwnLC5XHdYT5WrIvtAL80WnzTzq
rZosWpe/IfQewKY9pnfX5ACygX684d3LohTPT6ffTJLgtv6xyQVtQNUWxb3lpkaM
j1Y+khhKKr5cXa1gHaACYXIsOXdanZ5XAZq09+HEexlWuMNbyKA/LpJuspLcaPGE
DAGZfG3CBVUClNJqtCykNAne6WXFKDFRvd6+8Bt5B8QJjnuxNhOZ5fzUgciXqEka
1SYs9/TE5rpLn5/JbEpkv/nPbZXv8U5XXsX79WndhsCICWJ2Rko03Xjh1860ne5Z
gDgD11c4WaJKuCxm4Zsvvpk7Ea45AoInj4wY2jDcVMYnwy1ZRnk6VMyZf/b++KYw
IEI9LMfoSHPjOdxWRz5+8KziuYS7DiwCj0K1tlczWdRY1/Iy5yejpltOihzSZPkJ
faLnTPnabmQrnyHdk2I9YgohTXFbzyFota6rGkfL3G4xDeWJ2T4RYYj4r2k77Odu
66u+NLE5cHe4/WPVNJvsAsgtbKsvjSvA1sVpOCSjLEs3sYBGZaaTXxwBIXg4D4aa
8KFBTJF2eXag6bki7Yc0xWEul/KwCZdpzee9aiBF58SeFPig+xAlRuXsfKN/Hu5+
wDGnZHTvOxz7pRYjRZd8F1xkeK9mhDpgbIW975rOJqEckpzYSZCFWuWO2x2OcH4R
h55s45t9ubS99XO86XX5QsfTy9nrDiJnBt77r962M4kplAmnoLv7DPy2a9hTSU+c
m45b1klbPyOmSt4DRUirqV9yRW9TfDAhbaTU8LziD4JQhkFzrTEqDw+uh1YnyXaX
qWp4Dwy5nF/qNLzG0VBNa+DxaZIJeD2JQwoPYmmy3FoLka+tvZZSI0jLoFEcMvuy
fw4BYr2gr9aB7fH5huEJYdme3Bep7MCF5kSwDHcLl40WS6Lh7qK0B1EV3cWX9hP8
B3IL6kvVN+wTWj2cDEPX5U9HpPrMvDQrF3RM5cOIY+4+4ggMFPcqmT7w6KVVIuNS
XXnlInQhzPSmbMN5Pt9h5C9qPDeXw+iC6RvVBd68Ju7Vu3QPsFMdBscpRJRnMI7/
d/AplWQdyVlztc+JmzaQQe9qay0v7mRaAp5uzOWSKDIHJF+TIXf3n3QVAMdgK6Kk
bpoJRbpna/9FunQTlT+5y7d92xIUXtk7DfZuH8dpemJUdSzqdrt6KVDVvFOkzjXN
3wmzMmV9VOhQpyMjJtObJ/ICc5zTviaNkY1SOtV6sEZYyMhiSi/CCZVVMWYJmCXk
ZF5gU+Hom5i2JpjCLgvH/TelX60JNLnEsf/N4E0Lb5F2binAowdWSZZAupwHtEa5
4LqVDG/q1f3P8yEGDR3QhB3JnNsw7A+3sTqwABN9Jx7dX68Z5FGKC0Jr6YkXf+aC
BunlHM4xI+XHQvCJE2H1QD59Er40pa4NAKavFKNtDMf/sy0liASDTHvzeGUveE0/
xymFDKNewNj6Q4RHSPBszWWTegnhS+IccN2iY3aji2/i7tC2wH1EhXQy04gq4zxp
KradaBtN7lgaVrl+Tm4HDBAh7tBoE0D13REqMisVhlVvslPtcbxvKMeF0Ink0iZh
kuezY2jqSTAPYsaSz1PAi7nvSy1ZnQdBZUvwmRFIULNQieMHH0kbQ7nK79sCtXpN
0lF/OBCmwrYPw9B3rMwiH6cukTpPiBb8z3KcGi4LAp3E1PHWS6plncpKS/koEBvR
l6lr8zBxwQhjhgoC7fCcRUN2jeprFu3xommFCzWZrCq6h+bOS2ddkDD2FnPAWVrL
NQWR36lO7Ja7/Ht/o3mLFrYgMPdQ4c4MeIwCDnc4CPwRgGW6v3dhydVy28iU0I3B
cpDroK5RxY8ih4F7UItU76y3vHZERNjq+9+74Laq/eIrXuUXL6ln2Zxq7eM+9Byb
qFMIkmkIc3OeW7lqoUbtlJoHMXEtz9PlS1Rh4aMj3B6Ue3TlnzsSt5NEmrWF5VGG
9XVTlsGad6ZsmKBMYSCZLYs7qS0jeb4I0zGIIdWTsnajMf/r4sriPWVZuODS9/Wz
UdAvLEh16CL/+MjUb5NHMUBwlrtZnhjSrDVJzhJmBXZm4E58r9tplXcceNpEAxzZ
v5TVSeGo2oJaYfevhuIci/Pi9boCh8j2j02EBhLWOFmI1w2urhQIPw1xLk6Dp5Q0
p03Z6PrfYmfcObtyA8mWXHqecRsDiDEZE4pgk7KzluW5UtZuDu6L0LfdzbFJF0wK
pABsduJdByStroHg8QL3UbqWt/i9H6akNFoWfInFL3TaGRrOg0nBxZfk/YrSIYob
JH1AzT08E1OVogJmewGEWWBTjPWhn/Ic5UycTwlUbGxfyULmRPwDLcV6ZS/DRnhD
ZfwH2oFYLCYpqhoEaHJKZGqgFrX3vG2445GehJBNWw1Qa7PvQ5WKm7F74KoMcFZs
16S9ENo+bOSDoK5EPLqtRn/AHQbyVctUMo+GvRE5or0ZUlL7+RQhtIJxweRoZFiG
Ua94ekm4YLQRr4S+mz7JvDhAd7ILjwho0gYMCaWyk2mkY85d/qiY17wlXIYxowRC
O+9Bo0cd/q+sxX5qZEW8vH95LnLzNWRS3GOrdondhdx1LDQWk18FBli/lQuxnkR8
tbHA9Rvtm1SpXkYJfnFj86rsM49D4USgp79gGUQJmSDa0U/+LEY34XyCv0j5LI2S
9xJWHf3UYgft46xwawacqSpVRPsi4+Y6rr89h6AkTnLSTb8DhiZeYqthTalTjEjF
tPRVZO/Ng3ac+HTUbrva93dqsoah7dDEb522JwFEHgn/nqr+4vwU7e64ssPv2jzq
XOYkBakLgMjWQwypvy+S8kYAM2xINgsCXG4Ym71JmO9L8N8dv7SXxSOXZ42XoOFA
brAvXNBrQNus5dLp0gC9+LS+oAJlnOEHpGhSB6JMuqlytlUjiPCZKm6SyErw4QCl
qx33eS+lsMnv0/E31KeJHgVyvsvBpWClDYKzje/ijNsXDgHTpl85Myd1B/SWFYx1
QjRoA9T61K5du57+j9A3Ho5by08u3WMKjidjrRs0M66eZfgNKkALeRWN4QTWQR5A
Wb7fIqirbUE5/JrZLVQH+9jI3qzR9BxTHVbwUWJLxg2esv8UBD2F6Wnm7DB2vlUJ
lMcY7xcint72E38JdYTc5zQ8VxGoefIFRUJKFJgoFYqmMfsxDMKwaXMgxJmW6noP
E4Hhg4XYCQivZRBIfjoSCgVb1ZyWCaA6wxZft4JZ1IzVsk4GiBWoKnOX5BowDIvX
590hmvcG5DJZAH1z8J28jTqnzIBMPH8IQDUAOTIbqoU63ohhnt7yYAMN4e8uGk/W
cC67Q3C7j52pn/oks7j2aa6gMO3m5YySBbImMPL/gxUECt5QUGdrrTILrY8YU4gg
WI/+0BO8moOpXCbgaeYljDGIYWZ2ZV7aea1y86vsr8+2yNbOzdd9uoqX3g+Oac2g
eFXUU0D+LekXUTF/3GvWR8NcO5FXlOkPWI6OFuLWiQ8q0W7xp9R1A5VanMrTvcMi
k0i2Gy0WO+zSr6iRlFNkz9J5Pcrmu2M//5MJ6110TDba1A5YYbj9ltf6IDheAfJV
TnwKfl/Xsl3ykx6uEz7yTb96i0ot6PHnH7T0ygtVKILwwx4n/0ED9dKM79JUhX2P
4WlkWcM8a06x66DEN/4jvVTJ8wnnkOJTx1GgmFNEt+S0+y+x1CindUqkaPQxJDKW
zXITpALQOWpvuEY+r8LyP8Pr5Rs2aqwvQysZOxB68LwiTt/3BXvZZoMneg8VxCJw
XA4XryeDVhrlnM1MDGJRFGWIFpoiwRDa2iJ/awsMjbkqDrdVY7eQPgGplpnjjFc4
uICYPMHX/QrLMFZWN2iV7ZNl4f70JWLhMOfKo12sKvHZmnHR4nN3M6tkkQKU+C8g
D/IaMs29IweRIPJoSN4fiSJa8kzv3QCD0eDaKxJZhzVboEhXG9EFAW9IBgvtDgdj
bAQpvoGZagkG6FZFoG0RdnfYJAd7XDxtUy9Zq5yT2gxhdh3mZ2UTGkkJahB/Hk+Q
m2rC+gbVvVrO8xO7cEe2SMa+Ow6MR21YXOxNhwJTYSz6sDi4xpSz9WOwrxoP33C7
iEYTCxPJQh+IDvD4NpbJwDP/uI/f9ysQ5HkUHCO41Uly6oQnnoeR38jmU1wkhN9F
83tYO0uCAiIEkTR0P2UYExMuKskq3SGLch4q+wDBpxK4ATPqcc+1BMztk4pSP6sP
L4MASorrlAVaTRfrD9vpJUFVUKR9SEKccJs/u+OQkTp2ruRo3+i/NwOMYgvXl76M
acM4vQ2iPks3CTAQv2qwmnENqxWOyIu8z0Udpdi5U+H4IfRhXbwrbWR2HhrNKxvV
viFfp99k+DW8AdGdsblJaMeDOsPwYLwncCFGPMXV4iJKxumIYx+zTvE2COiXT4Rr
81qZU6M2jOb9oEmsW1OU5KD9Ssh8ueQ8XQPoORQsVeoZmqWV2fyC/rue0veAkRzt
f3GYI0Rqnzvos1IFosiJwKDjjtMxaAFHS941QAAbve7N7309kCR4Va+BUMmgYHfl
BSCkuUPK7lGF1HK3csXOHnKJdSQT1TvJ09E9FgTpP7QP/Z5+xckETgHzZyXFfInF
1WrmzEigDq/8Z514JKwzNoh9ONRXpS4qcVs+rciOnzPzvRXww30mE0wAk6LjyRwb
TX7A79NLsIlrp3lBJQ9gE9bBI56eME6+rYinTTZ4Wea0s5GjEDWVI9pnf8VwxV0y
pI5j0QvjDKaAlsd2s7XdUj9ymvbCxFI9OTwdxi1HwYQP/vKhHmaVxlhABOqVQT8+
JVfp+egidvely2V9OFoZy+lYNy1hA2jjtBOy0vwF1ipfpA++ZaR5ES0oX/HJnxxt
d/kYgGVi6rtiy4CsHFw5RjizEJDuV9X9rU8HXyRqkTb7UkxeTYfBvV87kEQqBm8g
B7DBMhsjA/UmgzP25l7Kp+R2P10/L+PLMDOc8zH5/OUsStOo4CkeXSMrAzhrLDU9
bZ3i7av0nERL4a7Rr75xM0c5skAYKJIHneZ3cOVkredpfSUm/159buAPDoRerDhy
FYTcpP+qwUSjEjmxMzsxVcUWduCCi2aqikNylkqxWcxoFcmqIrP4lP7VP8tlNZ28
GwUfliztLNoEzd3lWOBW7lWeCYbgRgHHDyvTmtACZ03sdaHLyKstfv/+XIPFFpkO
785utya3iJeuzrBw8u1NmFEn8teKRrFhGqw96Dtq0p3gATbEAHMVhmBmxlmodTOL
qrvFvEGZTWJEQqhWknw5Cvg1QwflRQnUyc/Ui0JG9r+WlrwEXT9SgSX3vxvDpT8K
NcSccHhqoa/zZ2inMM7T1lXqC80+JNT2TXRFw7JWDzpwxZdco8ZIhnTsesZqavY9
c0s64OOy1d+3NAihqRdllaHzebGD6zxU5rByEix1kOStX/SMr0Tr5Xw/Ei7X9LvT
9/7p0PPM/3brkg5Fj+R2OHculhraaEGYodktG8ZFMMrE8uVPcOUyme7Udbdotb4R
6y20THQG5NA06Z63SzJZ63ZZnM4VHZsapXPEuyUBIEih5TKTVWyp0cTdNsD6BBOy
C1SuRNVmbqTuEwDKZ/OsNfERZWh1SK0ChM1veTofwC7OH1dT8P2kRTiMGS+eGXxl
Od336tUyYSUL3SV4dGngkq0/7ig7/OSqeQx/bDfagFLL40gPXXWtUzrMt9xRDQj+
9ltwrMmwaUC9hgHVfJRexsLi/msgxUkq6exFiqJCK+OAsrzKKYmd1DemCIa9IOr3
MWT8lfTr8yKa4gJT+EDhfXwdSKKYnDyXVx9RkxKSNrmATCLbRjiqZsaWx2BSmJd8
wk0coI4FcGDOwb9xFKweuICI8hBxCIVV+4/9Mp0ist9rxTErsT9CpJX15Y8Oe3DF
NwxhOlvQ0t+mf90JJQYkn4cOxSl9dXdAwl6oeqZFlz1XtI8NUpWyl84dXvEvyVpI
SAUmlqRe3xTIe7igstWVaH+JTKoKgdPWuSUy2Ue/HtJvL7ZIGocURAdHktEhXpXL
1ixA7efBfuJ5Sqj+rtEotMDMzNYYx66/s5Y8B8cUJcBf0R24/aMCBCyXPnRSvrQr
fnmBwkrjj8M1I7wOKBAgwXXNsTA52OB7IQycgVEc6Sn1WiFWXJXMR0vJ5Ix+uiUm
dgJeDWc/5lKK8uhYa4tQDPpX6RkOuMXHavseRhU+3F6LlW3eahyo7bXT7EZRM2JM
bd/BNxIU2r7LDlpAnc7V4nvNQmRzR7xWmSrcZFlbLxhtIc295YGXKDuahd6ndQ9A
XrxsX94AWkPiwG9qVMbHkdfLwsNd7zXOqIbJSm5I6KjRp+3xcXBJ9Tyv6TxaGjzd
qLkoP9CItsv5eVV/osibBaJjubpI0FUuZ3k5Iatp1cxV/Unx9/8FKOKdy//QOM7u
tN+Vw6cQw4Fl5p9X6EWb6II7Cu+5r8qHB7w2CMkuGNCTt3Y8gJmGVYbk4X7EsKdP
h5jM6Cdfp1QzApaiZxCqHVDISHQ+uB6ZTsSch+b9X6h13SyGWegXHsY861piwDgJ
kifD2STCrpCQIuna2z5fHg1FslhoDYr709RONXLGI+T3D+IT77t07sZPvUtadqb5
trBQHhFZZKxjHzrhixOTicRaPGDn3ivtt9usncj0HY2SaFX+hADZBnrIYregNmsN
GNZiQyawt1ynP4ECmCU3Ct8xM/8I/ix/8W6WGa67t3d7Sml5nGqXeWmds5VnmqHn
y/423PoKLjUBsenrhBqsa3655NFJ2t1OMF5d7IEST5+uiXlJW8KgokGAMlQvmYAm
G4tx1JC/w6ELmSNXj/+3jiEVROKlwRmASn6v7r3sutRxDdDGI8SSHRo7E54ADvFR
2xDs64yVkd8E9RdnNmgam8HoRcsnomwVcSTPvRA60alsCd+9175gCebArXktW/AG
zSU1TcTjRFBCEp1cMyLJFKzsRCz7R0Qgq1jX0RXvGznGMCsfkCDaMe7otoGjsSVK
cwBliUHQhnOKYXF+IwUvEUg/ubD/Kr43CKYZT14tV+gWZA41JkzgkZndEwsL59Sl
C7sIR9S5WCnTLUJGIwODm7+Z+QpRpA8S0dxA+rp2l9Ag9fB7IUNqqVxjJsrT9uvJ
UcKGeQ2iYu/5SjDPwrR1fJXfiQTwcBrJh36hxX3bREVVikCq8z1/yuUQZiJzmRII
ysdiu9ij1YSdBhkdQoyBGcW9RmIoBFeMErNofFU6V49pxB9xY8yd1SlL4eMnYWhq
taBA1zTxe6xYMp7VQyCVK5kfCWJrf0fWMmbn7uklyVrH+KdU5ywpAaFvBlTSGfCr
zFxtx84txX1Fa2FqFTXZtv4gd322AZ2EPIs2KWG57WWBr0BafAsrDb0KoQeWh80Z
cW2bThQl4pc13A24p6YjNgBd1fc1nr8PWd2Q+3KW7wWBS2aaWySBnsK8WOqoQi8G
GrpKq+b1y/rM/ata03xn55mWOUQRu5xwdDe1lwNyMwv90kRiBYVKTLGAsLmNWWYw
ktohEqboo7qLvb1JL9q0gdahpWr/aZEadWQzxk/3L+lCsEbrRIqYVr30zeWfzeAd
fJVMzFmt+j+yQR3WfT3lg74F6+h38u2pZi9WJeOSlMVTzOiJhKRC+8LRyhmJQZcF
F5zM7GLTxGa8B7Gzz1p23VYn6cwQgFZSud0pBoV90oOC5zzE+o8RAO00EdizwtGA
zRrv5djZQoy8yecUKmdyUAwaXxGkz+/ql1JplN7UAfx/5yOxDR7q8SK8nj/xowHf
AKM0kfNnhmO1d9mXUNlG6e6OwbTOHO4DNb8JDKXFEhnGs6wOtaLTMTlG1nivMqd+
uxSGWo9V80qBFirLm+O4AgIP+oKsoG2F3apmuXGTjqp4I6BsB6/kH6ThXLsHEn0q
pyhDLzZCQsicKjlSrqhChqvGCJBnbqlzn629Ey69fwD8aQdRN8kxSzBn0LjNriQn
2wlMeQ65dcm4++TCa1T41RMsIk6XunbdBs3OaxCeMCHn2cthkprWmCUQPT0q2JBY
z9M4PXXcLe0QeUODqA6ZqUCA8PkLgDk/UOxlsaeMOrn+6HtYkn7HjZ8YmInNbzbc
kTxDNvKjYwNlxa82Qq0BCMVz2+RxuynVa4wrhNbbXG5JetqSNRog7zcl3Ki5Dxne
DKg67rZTh7OghQyjv7V2n3qoFmhhfMOY3bglXxV85SjzZUlIRTVoX23YDJkXugKh
bwUM3wdr2AKBFI22UNNkHvOBb83eGB3qWqa5cCHHw71GMMMBdUUr0NPsO83OWvgu
SEDXlhQe7VPZWKoF8tV0UyWZFm4tibgE9CDgz04QlarOwR7zZezdeAfhRrV4Ov73
JfXlOtQgc5utPCUavn36ePR5naSaeqT1pJm57CDs4Q1QfpxWk89l3YP7/M7Mn759
67J7C1Hxg46ErBxY5LcqLd7ZEVyqr/X48juYMeXp3OwQw+wuYodi/FDksxISOSWS
EG9drtRx2ij9LrtdUecfQHWxRxA7J57VLHicOhVV+bUZ5NyJnereeawb56LWbJWk
q9bg+LEwPg58c/m0vgvBuw+PYhVcZx65SUPkPBoEn636PLVenH4n9t9VWro1rsUo
M4NNVSfK2Y3XX3uu589PcJPQtGd6K5yb69EzAaIqcR2lJhKkxvT0jEIYFWjWNAfY
x8ZPCUFa0ApkZgzpRUKUh/tQKtCJ1l+JZiqEf6skX12wdE25OXroyUJVDEjaxtKz
oqbCJ6nLZSW3M4f7iQlv9nGiYHSKzre29Velix6p9LlaSn3PFNaKsPT7ZtlHtUuW
TbBHkF59pvA9xxeC2uUEfMuArK3q2JEWvRTR9a4j4FafFL+HOwEYH5S4RPBbBlTM
Ric8Y6zxfGZXaDnQbRfEQohdtZkphU0foBAGBYlaQ/b+w29KeU++50K45+bU2ftg
wYnMBnSGgd/EmixqWy2f28YRNVOqMHjMV6cVR+eQAlc/ZJzEi11bbMWn3RS3V7yb
YEFMoWc5mVFGrogujyvfUaN7gj1D5lHq8f6FWmTDTOcoGt8oFRl2Cg7YEI04Jr1e
pwDf0jj81N9gcp8/Y0RfmTSynKIY9pagvSp1ZF6keM11hEPzqsENX7T4T+RPA2zj
6A1TqGcDsXWg8W1Hav8lAHnWETNX55TzujAoj5bA0V7ufTdrm3yj7N/QKbIcyc1Y
UIbaXzIY6nUKaatIRyzi/rjSk+/gKqnOKl6qefOxoT09z5BF1kmD4RG22+ilnrl5
ugLEhVdpLYt1lXebiajnr01xCDY/zP6kpN3XeLLeZajkhfwGcOvQU5f98VeKL+H4
FoPYMphjlBBRNywUnuVGiwf/+pZYaQY46YNwcF2K8G22ZomRxFZAFFjFgwtjE1po
uabY+v2N6WefI1Xd6NIawxYeGm4uklNB1xP9CIW33m2SimSnKxGkx7gOQYD5dnEX
OlueMxhe6PyFCelYGrA1UMIwmPVHosrnESaW1HKnEjZmvwUT/i7c9bpzF+0tZjfr
q0+nLJnEcwYE87z4aU8t1KC3pFoHMvrwxEDNl/GB8H55OWNzBvGPlZ0rWB9Pjcaj
1HwIk/egndMDewukd8b24ZMkSLrZJhyCm4SO+HAY7lVsDUvnL8Nq1DlxiMuXISkM
Usddi0c9w5y2qDP2YPPCNeUSGDDPw6lTJovXA3LDNXOPdY6uGsKPMT7XqIqlmEax
4YkIkuAxFiIUL3F1DzQatcsnjYrdd+MUochOiKfryuA3NB4v86MxJRlxnPXwrKpp
EC4kVSy+Me8FMrc6/Hzm11ZXdBtrYIcohbGBP96am3KuSFnP5nDgtgmRb4DCAEp2
I8EjS3G1+1XFH8wsu60126qBVaYzpAaKh8vHRviLcSLTmrESzKmmdLCJAXJbsfKv
5Wel9g00ZUn8s5lyK9lek9D1trCqLKPo/MAym3N2WYIdbrYTTZ8a83p70TTJH/wH
iMEhrEaj6Lm79JHE97c/5AwpR1IFRQVSO1/uAbHcsKdNPoqM+958Afvk6c5n39vs
7yHwkw0/9XtMFkP4k/L93frKAcHlqbRPSV0Bzqg3wZrKi9W3i2ejEKUHIwKFrMvy
Yh3VjRgyBv82nslPfOJsqiWKRWCxWjVg4+Kmd631SJlf4lSh4Rtjt4kVn0sN4dGf
FPXrrQcbzEQRAC1q0Nco/yQvxeOlIsmr/X48zrjJZUTDtwIlkunVoIyZkii/QsxA
HKLB3Ehe6tOyjXmey6uXz1f1zOHbjSGyxDi2k4sUa88AFx8ggm8lpW2wbVpqPbHw
NFDE797nBKq5fA1DFew01WeEYwHYLPG7JYFulyr13AtSaC16+wY9EV2QnNRXl2vG
ChptngFRXm+mQlWjZCXXgtldTote0c5SHl9FtC2iNy8LdltvTkohFctVtjLKxoXl
KFveQNz8Mj/cjmHK8CcOQxORwky4dO1HbxO42wwk+gR9NgiB+icrmdQPK8T2MhBX
6VMS/svGnBS6sLnTvIj+Mwfk1F2P5klHDiMUETMJJCxy0nv7yiWGNeHB1qi/phNu
i2qdaDod0+Sig2qQX/yyI8meNXVvnzqBkLZ3vJzQXkzW2RxL/PMPASnwfVcx50dP
hSDw54/sLlGSVYbGlXERFaKK210y5Dk1cYALSM9n1uZQVAKplx4GDcOLShztYZFB
64+8opmNWaIDc2/6hH03ZO/SOu+VDe6xwgXLdJHYzIAWUxCB8yxvbc3QY5o1GIL4
Fn2GE9fr491OyfLBoMbM3Gt1g4lqeXEmzJOcve0EufrTF1llH+44mFY8xJ6DCRvc
X6JQh8p7gpleNkQQ5IpNBGv6NB6e+qFsgGEQlVMk8InsD89CCFKY22GQ2nKY4n55
L86TYDv1UZK0hY8wPj+Q4LPy6Sa4nu9CdpyVejZ4vw2S205fgiHKqEdoKj65YNuJ
Tv8P7zUhLBr91UwkRM2I0VHVRkMJ5WrZNywkAJIcrUSiSORn5+2EBnUTDvebtKDH
5jBbMoBatQNodA7HA+B5V93KtJ4yVmI2481NfBO/dkhvWNF6wY3W7FtjYNXVw/TZ
dcrKUhZ2yMpXgKf7AcMyEJCpl1HqO6LwrnZ2w9uLKUqtqdHL3sYpjzVSn2NfPYz/
AotJFF88mm4NTMqFePoPjOh7u4ybgsPGjsR4hj2eKrW0UbW7xX80hklW+E/WJIrB
NLBlYIdMCEft1N61tJ3Y+anqMeTzCgmeNVjHzCIxHvbhshd2f4sneKim64/fxCKb
UDKOWBtoLXJZYu5npXyVNnDZc8ZTnAosnSy8SBVscMDSkBFa8U7SqUq+xpw2oXSW
IcPw3cKw2oaTNcIfAv0wexDEHdfd6MfHoJcYYr2EYSmhZ2grJvQ4HdkbLItt9Ju4
A7fUK4Klj+4hPVaGMSJbT5Ov5J0nE/8A7GRUB7zKt3dlupVeNVQTOt72AixjZLZi
U9g/i6JwE1q8tLxE7Yn4PSWLCgZvfFmr44Ud4bOLuhC3PxZK3eg39UMLdyHyEBDT
W6sAawyrppbCBOeYm+7MHy5euevLUhEudgL3iMPuQ64WMchhE/rHChLyoF5fxLJK
EQFdjHXaq9O+V3hT8wlothx26AvJwjNbpOGV150z7sp9M3z3G7XhuM2SXbG8/jvH
eCveENt0qWh0TE4zSHDHgHTKUCQkCcB0spmqKnG/XHtg131nFKCJ2ARBwvrIZl7y
bOXIUP+5vSlWWmroVV8sl2R9/hjVVALPrI8dX1SiWIot9at68T47p6y1JKxa5k2b
yu1sqvBEkK8LaQfdspZEFsb1MjV66DvpJUIQnAQfWt4qwUUlcPluticXKjuxXOH9
llYHxlys+4ZwIj0JotZvDi2vi2+eLbyFIGcRkZ7NFWgR/H1obhAqxXAa+2p+KpVu
pLYNfr0vREeYLH7hymlqx/H0jLQLzy8yEw6JgS+haY6ZGky/q/zJ+hz1yy66D5I9
PRbzflkM9QcbZu1aIjTd+VzYckDy/r3MmZ9E7K5Q0oa7gY5yPLhadNgFJ2siG6Lv
p4ozd1g/BOFDNkqbbW5Ji5tucFLHCogCUmyAPANoQwPtP/g3f2Wc3/0PpiIPohYf
o//6/mNYBTXMSTmem3r3mhv2aDOoLuhpJpGj0IeEXm7VqdhcXkdLn4k4+Zrcfoyd
gScraAEbNM3jJIoi/NkFogFdMCtbt9Gg82u9MFiGm5sP81hflb/lp5gurajMB//E
RijRu8pFazYNHeUI06XaAHtehEPsd2UrDCVEWXDufDtRQzjhabVgoQxmS8PaUcWg
E4TuuQXFf5nPHxNAZl7z+nwKnqZVtJ+ljs0RaL56Uw23DYbtfoB4f88G/YfnKlea
FjfY7JcIEH0qmIn0Vw6FqGIhExuSN2cBbnPV0yGd3loBbDe+5aHYX+dws4yV/ReW
t1oLJ3p2kOGy2otY3vRN3x99DDeqBsxOHCNJH0wNQElxG8QWy+pRUKYC+fuEZmLa
D74La51XzyS8NedkSSOkzglCeB2UHSo3dRNzurv97G1ILfHUZC29NJZKgvO3BJwW
hhI5Xc8ygvlki4exP/HXem6TjUXT0ApttMsxmA4cYmB67CTmc5TVgn8L+66CPRou
yccmLniJ+QrHYBEgDcwf6eTtpBo/6xqapK4foiXfE1+NCuBGgZPFHfYQwOJZmp1w
88O2iyW7uhFueubUhT1kLawXgPCLSMqYzftr8qAPE3GB4Nvk+ycVLud+ybiqrKcK
FFGZuWqvOa95ZHrcNghux9fEDgj5BYvOTLFmmR9SrSbWbf3mJBpnde8HJuEStm4Z
YOluU6L/GTdquwkguOwE16XTX0bFqTQyRpDJW+WFMwm/XPT3algdlSAagauU1XdQ
5t1NuSu99WNFTQ1vmfzZ/VwzmTylo1Pp9JVM7oI6paXgFFoALl9kCneDD6PDFqTi
KTlPnbNX1S5AkXYzxqYRxY/HZd4bspWJfcWTHwpkVBpr/111POZvcpHrb5Hc9B7W
LxAn5HdkvmCmKXTbuyLjdEy7hW72lZVhO+rQEkfkCkHV9xbCbs5I81Wcw/vK33GF
kD6HKUOI74FyhW8QxDN++BT9hv4BZyz7gHsB6cEMe89zhOWc9kFlOLVJ5rvSmW5n
Is0fBsd0ITlWixsiUnd1o49exrB6rxNPjxXouq2tvPzJoE3vcqnizUl3yDkvkPAU
GNNXvEXt2wLbNrlTGyOn8vuWOAGUIPkw1aSXFn9Pums0sn+8mTaVcCXd+mTTCD2S
OI0f5JtKmgfhnWaxH09+Zj3RVCFzLFj79XE3DuLOesgR3SMxliNCSLicp+2QSx1E
gNMWh0u02RfcuieaSRVoQH/k+zJeGo7qkfOBOCaVeuNOzSX2chOtWH70hCqLFKVK
vMIaK2sVcUTJSu21+afbFXvmlT/gdrhZOl6NiWaVHZKDou9ghX6YL5mG6JcKqPT3
12K4VHV9mz/aAYZ9Do6TzfUNthF0AidCx4sdC5TJVYHDoGUuE0u0q+GZD/o7pVH+
pWxikqvxPt50wgXsucVN/tejlsRdpX6e1Uq3ocfkIvM0c3t+LLY9TsJeD1nc3FBc
hRzjDNkgStZnDUScP0R5e2cgzrGlMKPRj0+rGzZsefIin7wjJEv4lnBrZXStbzPe
QiJp5Xg9yyl6+gr0aUc1f2QhVYN2kvZyh2yvIaDdW8nLuHbpm+5Rr/Q7rsz6DAdz
8O2Jo0LQZG2byFud2AYk3+OrztrU9vEF7UAgEFcRvopKVyMNk3oMqnc1aZM+Zxc8
QBqpE/J4BwQmlLYuLYMY7yoK1S20riCpmW/DX7uiyXBW1qV6OUGQPZSFoCbG2uKQ
xfqmQAR3WKb8Yk8f5cAD9LFriPQcdL2EvM8nokfdGsiJx1SJyNYHqIVjyteHHdhs
96r+wRJvYOULnIiin57Kng7cPO7duyq8g7juPnciI4Y5gXqSDbRWBSJNRzooBZ2z
X8a7bnI29fnCIQBAXw3ue4W6jvdP1LWmHlPMebkHE53w2rLWYg1lI6lhbEsHr31v
c3btSdm5nUGQTv+K+C2NagZpV+buFqfd3UWFEc58ozDZO28aj1YuBqsXMAAe8ZZk
QhY0d9jRbUQkmug19bB3haUavC3uMMyuonXrmkJelc4PN/q/U5kMkZp1SjwhhBF1
pw9P034UPfhAyCElrFx2rz8/fsVBRno7xYhVT6SuCPw1Fy9kJgJkCQymAFhWMzVU
6FRZJV4TOBUO1mILjqRbvjD6gQN6xyZnvpuMpXgeOoLL32VpD9/dr5UPvzB/aHAn
C0hSzsZMovolcuLCDUKj1GvpAiD4Lx99NKL0zAlIaaHycWdMLctWuNpX/GBRympu
wwV3DvrcYjXGezMvSIfkDd664S7OrApM/N18NEFeVVOFEIdHYLxv6Ya1ggBSDLy/
P0bVDwMuVc+Tl4EGAMulkqyGvxuty2j4xVI9sYzS9u0Dib4eyN0HWi+tJ63+tVIj
3WRKCy2XoIyHzmfsRTpR25CYwG9rExkfGEgr20w7xJbu2LkavqgxJhRF/3dcDwLV
HGDlXZYVJg+BlG0dQNYki1o8ub09R8DYG4vgfsSkzO8muJIHykXxzX5VerSHAP6s
eb7IlVxr9gR7lnVofGRh0rstbeBeGT2PyZJm0pxzcpx2Ir6ihGcb97pGZ82cbfXM
cBiTP1FJlSsXtl3e9RKwj62wLWyUBZge9zfmF7YKsjEo6Co9nsn/2twc/n/Gj1ff
gPFbdDbP26g4axsfuSCbLcckotGJhK1uE/x+vVOtSaPO752McANVhxRaYEQVBYOg
OG1cu4r8wwz3oWeGa4Hi/w5oAOLSV3Wv8N7JEsqw93GvoV9knZXwpYBInda2sxfo
CreRLBE7hQGPxB2lEobOWuyKw0u4Oz8aObVhLGhJeCq4qQs38iqKrR2uUSvAm3KQ
XDTS2Fa1gOXhBN0rzbyxp3gXZDBkWFb2H+rYf5hhSa2HEsUY8usAjWcwO2m4roZp
/84+MxZpwGJC1W5pX06HA1iroeS+u6nQH8+5CWM0YNKBjsDVG+HLLDavlhtj7XQu
iwcN3AaCIqrzAuyZp+OAr/tWRkwmSXPRItNl/eKdC/lxMvzw9Nz0kr9Ci39ZkWMd
LowgBv3HNhgo04/ZyOZj0Sf7Xnd0KabnI3pmO5tRaSvuXT8eY+iB838NxHAXBzx/
R0xPbC6Zfrl26MrXdwFxIDNKGQTT993bHgosIFTUMtcSZ/0osGR4ilPooII0vqiD
OpwDcw2Xu5wRUGnijtH4Y8gvsgEw6f/VAmzfrj1+fdxF4S38HaaAUVVHltDhBksd
J3wsMgZNWqavTIyN0M01CQfBBecbYyEs4XcFr8MQmUbi9xA1J7eGM3T7XM7FiJl/
D2zeMWDgUE9kXIFYTxkbpKCRLG8fpFGuGXtZ11kEpNNxSOQBkSQ9euB7uR5/wVcS
ATVtzrrHFe0FyETUrQ8kG2l6TjQTzrMdyEHyqTeTD92TMSFxN8cLwqtLxXdd0oAW
0Q7PG8I0mUJ76PR505tlEL6doEIOPzpeW/B1eJwN1y2t2G/1+fQhLqyrJrhlEp/j
BLzKkmaaKIG0Xh3qMo2NatKRov2Nk9Xi+DBOu1aN28FGm3X33JN6y+Hcl3AwI0Qb
twHvxjU3jctUr2WsNLKzGoKKmc48BVzktFPAWw9BAYiu2h7v87NWbCQ1cWt7ki6g
lY++3m2qSiu5yIy/Njff7hvhoAsIJXDF5wa/+CIDsTtS4IYPqp7T8v65cL0VoHmH
GzVdq8JkV/oe2OSFB5lqDzExLgII84fKsRdc3NeQw+bRkMvls5QEkmOtEge/sImQ
4XdtWNUF5X/xRXYHdx9Of0gFvqn9z3sbYLIu+i00i4llGsSVItIqF3amPsG3Km68
H7plXIvfoXvNnR7j2bV0ffj99bBDCG+RnIF1vgMUHO40Y8+RWdjXti/vkQi9Nr9D
DERCEMFfc7qmQjP07y4Moi6URhC7W7J5JsXWvgYxiNibXcB/4dwY30e/5++Mde+t
5X76aOAg8hadbymBi9bc6xCVg5W3tba/qY2JR7ADRo7B3s/mpchZWsfjIKg361pa
PHRavDfPIwkfmW5h1doG0Rl3vGEclRfOt9doFpOa8nBJF2rJJ4bfgEbyiPfVUPJ2
lA9uRBfBBjDayh1UQfzNBxkKkq4ARzkQpznAY9JJCZDENvWMiTX7tkDfeQ0axxAu
gUo4AdHs7deYq/qLH8AVfBKEuiF+fXM0TXJPLtTkbhM0YxQovwtMDAGaxHBBQ0wV
CTMksFGtrJz40EczH0eg4RqkcFw5Ys+m+bVOOreX8q9sY6MmIxcFwvyAFBJH4LWH
q5INPsZIsvyK5L+JP2GGUWIYmx2h1w1a+4u+CVKQjLTq8w711ZlhI5BvbuEPQ3qq
gEwuFimObKwNBJQwSJ7LU9RjzeNC/83KqjrACOW5a5qlJgJnnWhOXfVEM1yHd0m+
1q0bWJd1xw0E9hImrUlnRXn5XfFNt+PDKS6qeVex4aY2WbrPZ9XWXl+d549aB3Qq
dgMZJPEbHkDnVWz/sH9+LSDLVolhJobrSmsBrrYa2H/M6pTZRm2do+dp7CqhmjU9
gJ4brxN6GJ+lZ5dG7feN3oy16XkK6uYYK9uBBZXXMdfPpJkhIA6vs38KLPTwhzr/
Bsh6LZaX2cwrfyJ5bCrB51FiLo6CPR6Pl1AxOUfRkKjjawhbIY0MiENzMizcyBGQ
IKTyx+UrpCEFEkf2Wm+agwYczS32Yis8lNRhVXRtjKQoYJuCY4DEClBkP5mvgh3A
JV4NzIp2eTOwQMzQj/rOoeq8vSzulpTBOAt1pkgJS/Tv6988KnXBT34otiGg0JN4
KvlhSyprgCnFRDmpvZBt7smdh16MIDpu0YUHG0NK3nwosSNwc+8gyLNAF0+EMCQE
70imjQyR0iHNdMHbsC2h/1wKOeryTXDayEdzdyaiN8QnGfyekvnG/SIiTYq1Xuyy
iBYWqtoUjAeBb0FfbFnNpDJ67abSt6OqoP8R2fWQbapuf3ywCtTY0/AExh+31Ur6
IIfSCHphGSCQnozyOKPw5OXdHL0r4HtEJ754X99v59Sz5gviK4WCcBF/psFQYmNP
hf9txBwcrTaWy7yg4JcLoXIJH2F6xGCD6iZW34/W6Q7j3uuKSXV+Cg8S+y+6WqoU
dRSPC+wzHyrM/fIgOraZKOxoLaS9p3FU4yUhmvin3o51/ezBjsBsYCr5sQRwGaEz
k1zdWiuQqfaJ77yab4RkD+7cDVn+o0zegY2T6M9zzH7JODDYeJCTQrGrbil1oChe
W2Opae4gt7tlM5z144LR3ikzzMclLgXmsYtyeCvPTO+C9OjPrZztoo0g8+HRB/vV
OpYJ7kziRUvEIBdJK4AuptoBbftJ7hpCk1oP1oSWTCKgu9Ff/PlsM9Lo37j29bXw
WlC8j1ZOkCL5EWh8Vubvy87pg8J8GgBuLnpORQzc5tHqelAT45524lN0R+k4TR1s
7Vjz+q6PqlKE0rgodb0atRYgxFQRElj4Q3VARwzRUOzroYAQyAD4kNzWXmAtCtb9
VgOkhsN5i5p0WwhLBmA9icPSRKomAgTvdhKEOSF8mMlEw0SU9sqzmiDn8V+SX0En
3eUZ3NKVeVwmXIDtHG7nQ//IIqNyK9DrVAHUYp1Dlcma3SNOhc3GIZvtVU9TUkWj
yOggMhgYq3MArbWC5KHz1MDL0sBqLMn2jGVqchTxFoBiO0p8zBsYkK8VHA8PCZDU
UfKFIqBiszYBY54lWVPjgX7YZVeGs+jzR1jyzDLdyhnVIuZdx+AWHqgQR0lTQ5Ql
bMdXvS7FWa0Hm+69BZdfqK8ARmBwyVp6QXSANHvJ0CGGlnLXIhZDaP/m87avK/eu
E2akeu0XHZ+Witr24CsPtXfTpL5gCER/OtC5zNoyeM1+YfuFaxA898wbTfJcld93
85gluHY0qGSqMPWau/41h0iVgetrc2Ukvk8zgOqlYNkeQf1VZMORadQd49l1G5GF
Y/PoiehrlZ0p6s8U1fOhVyxUPxkXI/8dkGAsKf9NcnlkIniisu4dAUQxYa3PM4uV
YTt9y6VseIMfUJlj/NBApARN1GdBYY0oJxS2rqGFzi89dfxaY6LbuJGFZxhhaEKh
2/ynHWwBaP8rO9Yq84Om428scAESI4NPxQjcHDVI9KwLue9x7ZXf9HHXY5Wth3Xo
UqJkJ8BI9dfkAHNa3oStHSuTnaq2ReLa6k+eVBTFoAMVYJzzEnI+kbuCeaMSO96V
62AK7wv4yU3b/md2LHN387li9Z66Ufgy5slX4u6de7qE09EmnVc8H7AnvAh8tYb6
SRMHPK9NmSyUWwKFbk4Bt0WnDf4zDO+Jmf3UuQeG6xrNZCpfVE7v+5PXzyvjbouI
qnu/ouWlicl39h27cJsAVyYY7QYC2vsvObyBW7XV1FG68R/nRlrL/b/W7FBROd9+
diEHm6S516ectXvYFVbBSy0mSC/BdNOjPy9zbaKcAGHh0ajxcki5hdmWHtrM721E
BdStBttIkOkgTHX2yoN5S7e8mwJ5yh1e8l9Bv1LLmS8melnavrpaPBDkey+MEh16
KPxX1Fc3ggXZuCwumGc+T3oQT1oIi5Q2uFkMOlGo/IkZF+z4ta3doSDso5SJRI5/
qX18e/i50uJ/ugDK11VlpoqStYADoM10xalFi7ALhqX5+/nGTLNFbF8mb+sEbrPg
mpFtMyH5U/3tF0cswoSrmGb8Dxfmp68AvSeeJUOY/QwXzLR8N17lryhqRN4NRp/4
i55vwS35F58m2fLb4zVIWv6JTbR/xU5pe0nZMZu4yOO41LxjmAWagRTlcFhIaKo3
Aya8QEcYSFhr7M/aXaQVWoBsdDKN8Yp86e9SoR8KeSWXB8F86ftDQloIvGVCULzH
SE5sAg0sxN3/Ju/39oSZTYUtwzrLNFw/bBqr+yi3lAeFF0I4/qsPBQqH0Q5nlUQz
JPtZ3YUO2axDihsXjJOZOdBPsjdf2DMKHDAzOMZIQWpto57VKgHyBS03p9e6yZZy
epOR1Rm5CVIXbpm+DcfX8Ymn+wAkKyQOTx6fUBWfqCzeigcrDb4k2cusQCn43cN3
fHLL0q3XuhK732ob6kvtdJTMaU6uXyKOgB8MusnRRJ62AuZQhygxOr2UVURvpyD4
l6GtQfou7u1tT5So048eJHvTG2MdRfjxFCsTqQKJHoxFOA24MSKjOAZzcHxzjGZD
o2k8QThjPiLQ+kfExadJGJ3ro33eg+B37HBBc9rdSRwhNv2nPT35uXweQTPZ2biq
OQA8GK5R5nk9qaYkuo404j8H0ZAqQwdQek1ZCE4QXbsV7e0bAJuS/mNIaenfVHfX
+9A70x8t8IxrmAbU1yHli2LXZXE46HUs7Cj5wgMkC1sqge86nThYBccVeeeWarIT
NnTtMCudXfHazPiMMXBLoSS+ZJ0wfGZM6r2crtJfzlTUtFMIq57PFEtMtH25dleL
sAiQdsvpnQd7zr/dncs++XXDeciYRcMgBShsvBS4QgANJW0DFbl11SQaOJMr6ahF
sCG5u2EoWaCky2TD2MnDZMuEZ4gNSvBwtRmE5SX1Dt1zvqAXY4iDuSMXksuC4/1D
am0wQt11X69zXSudvipymXJvLeAob7hnmzk1/lDG1Uvvz3YmlJlqAm6BoA0tUdqG
B23erLXcKEvpznKx7jKRrUv0CWI1Tz3Ioijs8DeUdenFZKP+sw+HhPI7xB8bIWUM
xTHnnQI5MXhjAI4fjO8+S74mgjnoFPzOl+G2Eju6JUzpGuUEFyw7hSu14iL2ge63
CGuCjMxc+OoZGQRh24idplEtHq/PW/TcncbrDOV+8kYqMqHvbQBAzBOBf/ZwSkVj
xGBfdwBtKbyHwh1tSipR8vtcvHPmSy1PArddTUM3gSo/7g87HwEz75o2Sba8covV
Ncv4CCSVlvES//udGyxFAQmFO/pe2HIHJzb47gIqPzXPyIvReBuyliZ0hCbfHx7E
wByvL24H2Te5lX/jX6R8OD5aMRCGS+p27TbR2kBe9WBbLB/xZNfoei5HABJFh0ad
yWcf2xibJ1qVmcBqvJrfEAISFTpeB8Oa87cvtWSQl4LD3cQEJC50gKefxS6BAg6X
K6XxODT6eFx4Wq7YUgqnDxDAIVhtNL0hLHC5zsHsky5fnNjDd2WaQTGyARuo0zTa
eH8Y9FoqI8nMYS0Q58dMAqySBY3y/nHI+CpnFytK/Jcb3kXAAo6yVGXDyyOXokqP
rJweCNe/wBoDfbCsi2PrW/GnWZNhi7SDFcmuMxfI7UU8GIVZ2zRLb4Ym/pDJKFDN
NlYnZj7Rx8FvY2IY5ZkZi5ux+O6pnzuG8gzORgR93mGeUTd9gQTwyCWkCLBeJZdO
RmgKEq3xjTgqGj2GaOpA74eF83Gc6+HT/rf2C1V5UzcHCZZ+lsnuZfqpEdQwNo/W
PLEk/EBucsZTROhSkpl9LK4tW5YUtqirMeehWOjc/6sEDx48G0wQP+boDWryRMIH
DjpBoZFSN7iIfOWeDzckZ7xwYnxem1OVHIE8tk6GovcNI6dp6o4FzirXOi6GhHBB
f1GeUY/GIa3zK1JvSS8oSsTJjvfasfIWyNzJbw5ufJrxD6YEqfXfOLQg2Hs6GiTX
atDUfCRToD+A1ojeLuNO0l8PzDV0aM7+GUjY4nw17H9wJFplcAIENxMh6eD/dsgb
HDnc9lR68g1BHX++DHqGxiieDvUbIy78MGcvXB8TAlX1hrJMtzA/kjEvswdo6jRF
52A+I+LboMVJcQ6S5T5+b6dNRvsnW7JkfG+gp9Yc8YSkaY8XF5W2dDJrgD/v635h
dIFBKcLGU3Hji9b8UPFom4UJzM9FdITt+ZmljtjRGv4/gUn/E150C1tsZa3mXfmU
Hk09krzMnHkXD5iq0m5FXxIfygtPww8N+WN2mrKmLYtDByJplgXQQXr/HtumusVq
Mkgs6vmxv3NxmNXuaPKklL/yw7BAocMDizEnKedRnpbol47kA5wp3UCOqoQBpT89
LkEzRPpjJeXunSaiL09xpXlf6qBSXoYOz6KR2hENAf2QhWK5a6NLvCGcieQAnLyG
OOIrA+K8wjGOyVNXHBN6j475VezTHCMa07eRTE5/xoiVpSfWE5tzqOICk5Huz2fj
SviV0H/oV7PoU/gWIvv+jon81Fr6edYsVjLCmArK94hCCV2lDSdr5TSRVrx8QtJw
vDNqT/TIdOPd/N7n0WhAhvfyYBzx/idg6s1VRr4fY7j/8rpKZpZ9967ax12YjwPg
algNnV529ZdeNcrdynqhwg5+58icgw9ibXE4teMkFiDvmPiZbKuxo9YAfoS4287U
VN88GaC+JggL30+A5EOBVNk4Bi7M72RoeGz0qza5dA0a8EVCi2wgCNcj+29fDfIY
W5LPRnqRc55DvBecFijDwrxNn0UnHKciv3/JbiVpD7CzFs8UvMJkWvmQrU5iRarX
NSoN/UGNCrv6VMgC92vfIJ+76BF5z8ALnsQYY0W+PNMwoQSdF0cJ8SpERqDKiPsV
8KI8+kcC5erltdm6frHG+hoZO4ps2tfx2j/d85JCjjV1jxBCEA+gfgoNrDueGD+P
MJwWbyHzRuR4EE5TmrPoZnDIcr2icfXf67mr3daAwPL1SYW4UWdnpUG4YkUgXTkK
fn9b/aclYxf1WSNSV3c5QKZ1RAU4/b0zhX8NU7sNk7/n37nzfZRrIqxtreLWos9Q
aHuEzH4WXj0eegDYor23M5h/x0lPOFkvO/ThcNMUu6J+W8YFlxARJUWzEYKtiWVD
97J902yjJ6juFf2yY/d6nFzyQm8zFnEkJayDmv38f3WYCL1yAhuqwbAYT++pD6qX
5O56Xa4wQ2xx43fKulR03GV/38VDBA/gp+jf38krO5Ilrgnj/wFwvjUaUXdMjzea
bhoPKDKIFPYlqd8XqE2niWDGkyk95qjXWxxjk0WVPDfYC7ugoEFgbUdWnswebWvN
2UVoWYXGS30BiYcs8TApEVgFsLtEdaIw8oWnKW4hnkf06gTSU/T6LrZNYf2uZ4JU
yJZUu+2Fbhjsj28k1dkG+TE+Zg4PBrt9Ck8G/5YnGe53JtG+7YxTleQPc9k3Jirz
4gI9sbDBSKalsz3EujuczIdr7tw1WYWptO0sZKELHP69Gj3BsCG6HzhZPzs29osa
slGEGS2gd2+5mTSfc7CbpDKgCq1kRnTiuM+so68l3WJodrTNKXDLa0+jhD7SK6pf
SocDgZM38oyFMGg2CGPhCHDxYvfJxonsmYQ6AAVLudhm71T6gD1YjyB6kcWcU1V+
uXQhqsY1AybhWfaVKCrctSNKKny8c/HvysuvXXsE34X48cu93ip/KTUvEm8sPdSC
BXHRN9RoXcbJF5+bd1wz0GPbvuiWwh0KGeQ2X67YOTOiOJ1WZ7zvpRLuGiCK4XSz
n9ClW7G0olZPqLvEPnsVOZLAZch7qs/dqgvEJ9xXmCEY+e2wMKmRVDKZYjw8rY9M
aGGokj7ufBpxteYVeKaJBZTC8Ab1k54NOkZuXG8gidYQ6pPopzIrUXn0waDwP/yp
ZNlMkfiyb9MmM4BuaEEJFAYc6CTk1f+EAyfta83degYPmJAjQd/nJRungV8I+l5K
uw7oLG8t0Dh0LJjoCQ/HmqUGT652d1FB4J7A4Mq+Ad1GIu/u/ceiyb9dHpsqlMZr
YcChOXk/tVS0zJOQ1AQfl+gt8tCgl3jtuDsOPeNsmPBuxrcD+iFIAmh16flAxWrW
r0j6tDqd3EuiCxBzvKNmmjVvRWiYzY4L9CtGci/CIG6VkAYoCdh0FUXMawQLD5fy
ssh3tJ5y1SieW9bnNPk3V2HnGlztsXOJaPEKhVqJVfpgyiekX2Y8sDGLKVB/FTSz
NuEuDqOlmvTsQxPIv+Q2VaTFa1kjRsupmAvv6NMfDyh9XUinwlk600/x45BwCFaS
oTEhLkGy5hUOrPEufPOUgUL218DgLaC25BO65b/hvBu6CRUcjQRGEuPfoCmJRXqF
BM+T+KRSrsgs+Afg6F+KG5685LULK23DiASr4+bFnLkyfLdi8mTBO1Xm9woRpaxA
E/rwcEOLRukLdmRNoq2AKFJ7yeCGol0fOWgCf2FJhUi0QmMcqDkZpSSzpxKenWba
jL4L7mhPBFuzosCUK0W+GdLOxPUUlg+P/HnW8TxbEy2pkQWiNq1/H0PK/FI2jvRN
wywlqgzU0gUZF9f9zwmZdHaVDLZuoTNH+QeeoDjDyFyfgCiHgUPnqI2YaBYY9nTe
xl/q5oA9jcYuysNoi7GzPN/11UXB8zdzGRBO08I7NzmXaG2ZFJSCfTnZVfJ/zEUx
6XIV2lrsyHf695Uh+5hiYkiB+ousp5Z20WnWhfzMYdtZsSPDV4tout0yQlfYxV4b
TslzFN8OO6GVdKyXgt+pwcYskb498I+qqVEGuxj3IZK4PstfdoCLhagRnofstb6e
9npoy3y3RWHQhuKxmFWeIBGxtRvGTQ+1yM8mOm9jL6kDYQQ6T6tQGbbBOO3MTe6e
vGH36NzRkbjBrR7+7JBIC1PN+AEbmgjw3SPEpHELCYwyxWVqAJNFdcLFTEMn08ux
t2CT2KsndRmjLu7gVygg/A5K52+QcXWOuxobsr9i5oJYNfkSueAKvAdUMSNhqMcX
UsNbaymzHMA/TR5z59YI8BTe3AVs6WtRg4uPWd56Mf944mEvznG8b5LuqTD81BGK
A52YORmxVMAWbyA2HV2PX0AciSLKFiL0NICgvtf1pu0=
`protect END_PROTECTED
