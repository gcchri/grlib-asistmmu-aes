`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ig/NxiZgxwRfMqEASCFxre2dLv+mugeoPrTGSchbJGjRZuPNX333fF5SWziyfOSp
BHxj+VoN+OnrmDaWytz8IToeHoVBpmhHoLssBLaY5Nxm6cC9zpk4DQAX9n7VPIUM
jtid37O1xkVaUg55l7260avHF4D2LN8VMMPHvRGWAuBQmbnI+UrI02UR6XDCtDhB
dVf3ZAj/SPwZikVeATYQP5LEruWlhwaHOdAxfUZP1bB6Y3cOqi9xwUQcAJpRV5RF
NV2fZSeH+x6m6qvRsFcuB+uw4I4etEUN/LIO+AJ2xqlcXobS483+1UwR501dZ7C/
6JW8z5Ue4mTxb4Lx+6pvJ8vW7Idnn5iGgcD5Oopsuzmr4brZsr1WqAA2+WczpK1q
W5gV7iDckDfolfwMaVDk0q7YfBRoVhYMxDGmKFb8+eYeYqgDw/YKWlpMX/LS0IMx
jmtBno+RZslyrtXh6t8X+DaoBMmVSeuFyA9ionh8mlfCLqa9h2IZpaI4ABcGTLbE
Qf6BXqWorGdsi/vVwriAZj5EPiVODrjzNnGT/e4vruqtvDOoEJSvCCg7ANb24/Js
KelRs/f+8yAJRftjxZlfjDH95M3R5JZjdALTQM27VZsP7ZRRGw2+9WlbHdCXHqH+
lL7i47taRkJQV7IjUysTv39KO1s4KNyznLNyVsnTh7xbxN1dutExYiikd9mB+DMz
UZ82WZv4uxf+ZbY/YyrOnvWEh48ZamGg4u/n7W4N9MllkaSK/8/HMNLC/n9TJfRl
vhOg/XxcF1S4qhMkECoIUg==
`protect END_PROTECTED
