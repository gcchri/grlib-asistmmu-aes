`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ex00DejS0pPe1A5Cpu2JBnP69Ex1kd9GJHbgwXNGTQUn6hBl62iJAyFBDQM2YhjM
EtV8sZmrr8vtNWY4E4BE3vaPOkzySY0nBKrIM9g8ioz3iypwbtZY7hdaMD0Mdrg/
/ooho+IOI+Jr9SuUR/DEPGVC4zrZ1LEG0EVZFQixor+1Msn+lk8i6tWBcOeDdHfb
BTO0hVGYdNUydKTOTmlXmqtg9z67h7Pn3gpoYdA5g8Ssg2BYvEy4DQVvNJqki5Hw
d/cC+d+H10j+5cwZ/kYTrRAil9HjCXuimnBjsTCedVJdtoBH1fBAfd9JtMnWd0bx
t0nc6Mz8z4Arj3cLV6R3das5HOqHKar9YLLjlTarM39zAtODWvytW25Rt7OMHRLp
Bqg7xPNbD8WwBEenJMfWVzfgkDd/lB3Z4yiDotgpUagsTmoqvzNAY7FX+hqb/w8p
CAbPeesrHtdgA9c3TFPow56qKiCv9dc4pLz32Q7uMHnym/DqTsyLa+hCsxY1uSb9
WJtAe+3CwQCb+i5onINs31gG5KNFnSz/Hb2o1T8BpXlJ2ot1iqV6fygOObFy5Jpu
Y/5FYi0Wbx1jW336p6hZvw7/mgzBIorOdwgNBiKcJ1BqBgzUqTJhPvhl4iHDo6yb
+eZfAMzz9MCO2zWb71OQXP5BU5R9WTr1HED9qBetJydhEgNR+HPod8S59ZRAc6kD
fXZHakdgqBh+D9q9xhmD7+rYnKJ/dma4XNErfvC3uhq2pWxp3bq7dCbZqYmc/SHw
kLCOdlRn74u4atoD7WjNydpBvZbaBRd+820APVvZ/LIzqos/jmXQ2ot+VMJibFW9
ec0lywagl9WUsi1GF7Jx2XcR1zJqzFPEstE5sVjVCjNkw1pxxvPbELX53WbFsFbQ
L6LCtJiGvsMzbm7jJnGxHZswX+0dEKCyKtXceeDnwVrhUAYFzYc+S7jrlPgiDrJj
gAtDr2z6DBvpp0Ew2MohhV8XHQ7K8vX6nbBLUJaDkIVf7dNEncBerXCwUahMU1FJ
yT7CC6ACDY+B+u4PrbNlsT+dFQ1yclblFdlmehYLlsA30+DXI6KnxAV8/gyNqK3Y
CFmWdLoKHyPKGRmN01DfqpwgbmwOJm7jQgf/6fQsPAUEW5Jkyr/PtnsUnI4oI7VM
XAclVRMLyEYgrFmEj0DuC4Il01cY6ie1ZXAqe9qKnXGy2xAueeqLGDwEGU+OqFUq
wYy5Hi/ri+gg5KA0eq2wbAhh7iMvjdNI2r+wDS4nVUfpsqV+3nG3bLDEmyPDAz+h
vUczmEEvn8hOMOVeGicZKnhFAXH9jkc2BY0opQZmFnGhV7hvKF8hmJxYhWicT1ES
Nhr4QlUomGNaIuriHxaLfKg46aOCpxIEe7HlCbptZcUaZWfL6E2pyZjX2OJsw45x
9F/oDRICshNuzkB1+C71b1s6PxZgaPWeAoPpyrLIfXS3UJqoLNEqq5tERgAo+hb/
bzN9PJwr4rqAkcFjbzZb9muj+JvaYIS51HVB0TfuZxUDGkBBODF3fhIEJ0tki8b8
gGbXutCbG3lkwh7BptbBeMXU8Lmw9WiEXViHUFGzzG/kiv9GvtVrWOEx9rFfn01u
861eHYuAgf7RVI62TikgCS8bYaFb0i/Cy8aUmk7uo5ly/fBQwwqPkp/wKMUUU/aH
`protect END_PROTECTED
