`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2KUhWrK8VhbI8aOhodJBsyHSD+BXFayNmlrzTxt9J0fC6f6ep3IunbgjtxCsgKLD
x+tQK15LD/WnYxZH+izUAnq2zVeQNG+Wvx1BdTDHLaw52msoyv2+aexj+4WCBt2x
gOxnMdP4kAzLNgjG/rsPQlrFkCA5zRiZp7sRJ2kjIRpK3lEtLosyfiWdF9vDXvks
Kb15g1g1dvM/A3u1k94UFIeL0WLlnDNjkSR4hqu2z2atWg62miI2GTIF+oZiot+d
zpxrwhnqwwWK4y/b8Aa3dwz3fo4unv4Q2aRT0pxZfPRbOXuYmq9Y8nXHkPUiDQOj
DqBIe/72p3G54K011TrzbMRjEt9hM4lKUIZjug3A++d/aqObqOWp7Xd774D5FPUh
5HhnzFlPKPU+MssJokokWTQufchM2Dn3vzdwEScARjQe562pmsHf/zDlSDwRRKhk
EEpW8hGqIJ+wU+pmAWfuyueMjq0vhb5FNMq8Hlpb1Nmpynzh7amFBj/DEn8ByZXD
ezr64RJn5OYk5pmDCU7CXwrs9pD8TbTj7zZbQuevncpddNFOyGIq5FsL0kFHMxS/
C8wMTBuohlC47f9Of5f7dm0T29dr6di5KABjZZMZkbxUdFRX5p+9p6uBcXeE2o/M
l8aYPODiMm3pVw4Ze6+acX5rl6i477Ohrf33CS5s+WSba1m+htJQuu1uO+nOb6yn
ybHr4/N4U/oBcWP1lonyYDH/lPSKQooP1oPfV5Cd9IHT9CsRkuvptM1lzthN3j//
qNy+3Qk1FgzjVU9iL5l+JHKxEl7oalMIP9NElGRujeyVidyPs5hIvA9dSIOSbXg2
zzpewadD30nugId0Xnain6yVFqaaJ4gBaa82QRKho3GpBswr9mk1JQKOa5yx2M6A
y4HKWjvl3T0Su3jfAS0qmJw4PAVYnP3jzKi1QyNF4y5zN7PT6L3CPujB1KDb8Ibw
/OTufENz+2E7Me21Yq4GjaAc/MepBOpxz7pWwy+npiRL91rIgWQjlmWAqHvxyPF0
oSUaxvoCslIOGTlAV4P5iCQozBfkld/Dn9DLIWotBC2SkPj2vG0kmGR24KRBZBNU
bH4AFHsBrAXCWFvCurNGaosqRY5YrrO48m6/TmjbjdTq8xKP9JTChuSCxRSJ6JFN
2DVC4GeRFgs7g4qkqZMpW17u5x6K5B8H6sawMDa7X1S2yrSYBCqCo9KPLNFp11lm
50ePeATWBSc1M3KafH+hE3vi2H6Oj8qU/8tRP5dCo/ZyVfiupqunOGjkLZxam1Ce
GMFVYb+EL9uYB5Vsqx2S11ILJ8ZVhCNXtL1peGa9n+li0f+VAnqwnZhJ7rXoEUcf
eN1TC8xYcy2k+8ibgLBUdXnIij6er5pmDSpxx1ZnDtL7pvGBkVDxdsxIexLAi0Kh
gsvMzDYsz49Exvdr8m+dBCkkub3/+AJ331RWSbPTcmo=
`protect END_PROTECTED
