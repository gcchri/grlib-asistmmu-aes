`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xHueor8Zb4nF8QHIIrl1QmH5pJmPBdt48hKr2ajpF1rWQJtMDZqIPG//Zs5rSgJn
g8HKKtdN2Q1C+tDLeuXpSLRmkMaEIOKQjY4uBHCM7dX0coTm+ZAr9wiaDxk5ppEN
iKjD6GPx+L9E7wVPqU2uAfr+OkLQWFxhu2qjBqZnFqACQZqR3e8vEM0xGwFyrzml
Bh622GBoe++HHpxWj9TSi4/LVCHmCBKDH14sHf8v+HpHjMWhqdP0kX6ROjHIFs7A
UQfVrK9tOavRhT5MYChTek6SMPKXE/IndhMoySg7ymOQR/RooGxm8H0di++giU1+
ZvpBBom9QmHsb/GtjOeCupb6AldQuA8Rwa49C7j1xUKgTmoVnzpeHVX3HpnHD/K1
qDZJCJbwnOLKlkF7FUaoBEg4u3FREEpziAu8pMeKHEHYfxwhMFUBmvdKhjgnv0Gw
H5jlFkh0oclkzububRa5w+nU/tL2d6tsUXYZneEEW/qBEpsPOXZUEW1pVbdpvVFy
A70h/+iTilVh24u1lMncrLu2L2szeGL65vMOVFsEHG/9C74vKlVsP4ZZDr5iNjR1
s71IYDGOQXvLDvqLDYwfnpWsD8fN9EHXGGHCZ77ZrEw=
`protect END_PROTECTED
