`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l+v9wT3c33yn/yVxOzH7n/IPtAQ5dMa+jiRKNkiF2WNygnFOmZ2R1VHZxGWXSxzA
A0GlzfsslEO7X//rwDc9+u7/uXjLXD5o7tN+Zfe7Sn5M95DpnFr5tpa3oB3TVDd6
PT80MM6+J8wK1IIHWqufWu8j83wtBkU+Ruq2cZPOSI0oG085WvZCkC9CPx6mvVzr
EEtXT0A/DM8BllMNxolffr9wyjPsgzzFlshv0qDA652wmygs6HNgcsMF61lR+fqJ
VLB/qFIHwORQjaCxUWC8LpGD/KawzAEcsGaR72ZLaqQOrvu202MUFCxaUANaDZmy
5cMlDOHvs+YQSQUTPOqA5oxYh1RF4sTdyqnMPOgFWIqqjGzBw5dnbhTFPxxuG3FJ
I4nuBRhycw0wdU/B0Dja4UsTrsKbLaIrSdCeMcPH8wJEBZkbGUKCgw0ON/sHfll9
KduVDdVlu0y0/yPtaIQh6RohVxn44KHCvC9dovsvRBXpn1vQCY2Ug8PACe3FhBwU
ZFCMr4viNNyIB+Xgp9/L75OcPgVgIQXASp98Vz8icViyKmQZ1q2Sx6MJZl9FcYXv
MxGmHIWuvcFXRyvMbkxPMTZpW6QRFTgEf0A9GIpPtHZaoi6ioZF4fRaZEMgP1N1d
j3ZPScbuxYD+ex2WbbD/ebdMmh8HTs9WSB+YnzN53qGhQNlW0Ghb+OdKVnzXE3Pa
rhW6j/0K9gj5ouGMVJPPo73SSMQoV8ToaZYTRe5wpkuEbTUp6tKr6FmeSNz5xnI8
PuEqdz7X2atQkSTAvHqHuFz6/48S/gE3alyrCZSTxyorcqWzh5wykzA/QJG20nQo
GovUjXJMySKRebm46n3mGy0esXP0LtV/f/irxt0HYN2ikZ70B63fbnNS4BEHalfv
hhAOcDKqxxa4aiYm0T0z7RSreIo+CE6CIg9Rzli1vZp5YOd3ABzZ/Qiz1mHZeUM6
`protect END_PROTECTED
