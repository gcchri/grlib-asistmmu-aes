`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b2MajmZVgqMJfwZV5nlfNm+/Kdq2ffF9tqjvI6UqQYOR5mowLXJUhqHnUOqxd1WX
4XhEb2GgfoSMZm36/m4CDELJad3nJeqVrb74XruYY2HWZ6y3mnDUde2L0nJvzE9e
03YmkDd4ChpD0mZ53gUnvfc9Wf6pGtMfNbvWymjUkp6ogNdDsBlRcGriKxzOZqt6
3e1ns9NKHjXDnbUvlQfctMvv4Y5gZtCrY8xU+EOZut4zI2wJ4KhkOM/p3c52ykyN
uk++tu2k8c3fInPnCmf3iPbifY5T2xYf6GknV7La1hh+1MRpU8SkT3oJH05OkWrN
A8Wu2xmfAyoTduHxG/I45HbGG3ALp5dYtSBXiFZamditnUPfhSFuR5cp3nUWzZz4
yuIp/8734+U8g0KpLRnFZrfYpU4FSzgNpL6LQias4p6lFJ2tzRMtOooIq5vk37Hf
4uC58ZPhjnzv1cD0hdYpAyd140ZORAWueUWS/KB6411Act0ItY2wNKGZg5Iv6NxB
YiwIH1m2USdb5bjO4nVdhB6v6KJ8hKQBoSJtjXdOaradfRm7tVNglmyEDiso197+
0qfpu+iUw2yjKulrVswXv4Y1Q4vHrF4IRU8qKs226D2gPVHXOQFvP/jkjoIEWwLR
WWONikNkrgf4c3GTOb4Kh1hXl86yeqzua4/Q7H5VdEdz9JzmMGg1JMQMJfHYFkk6
7+V08utKabZjl1PZBWzPyD0lEi7mVNNmRx1dlfqmM24=
`protect END_PROTECTED
