`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QpCoy/Klcfq97+62ijiU/R2PDcpv5+sGAd4wXxQB9r+DmXZbxJK6GDDlL2bBiclu
CM4aUJziQSa3TI+cswTAZ/6l+XHYvJ7zYNRjYG77icAWVsqQGPDfsIwFvhULAqG0
WlmJFK8T4fGurD6Li8ZOXt6HluBkQ9F8IULMXeczVUXx+a4PFJ2E8Y3xo3XfETDK
I4S8Lngaprd9AY1FdRcIDlAp+17adSve19LLA8DPtz6itM4t7nYgSt8EvMcCpt4e
DydOgfvqcmn/rMzpEk5dYfQmPdzWoiM5GHaQVd3RWwiPICwk3wmqs1ThSN9uSkyX
Ahi0jgwrbCeVeqYPl0xt5NDObAF5opPoyodv7xWvIJyLGq5xWxJRJ9q75PBjFqxR
eRfHB1Yo0R878Jld8K2CGg==
`protect END_PROTECTED
