`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hFRHe3c1Hq7IxjBi230tPx5ObvOvHCVUSw0U52wSamDQorlSJI6+vZAZGgfAciA9
6MQU+zR4+fpr8j76+KJvNNlCf8jYJlp7AfVVDXQW2+j2+NI55XE5WG3aR2dXBddy
IzIaNbomyWXRDUY36g6v2Mj0dNe+AiwOI90S9Ryumg+L6ZO9BPOSoiSWPPpsTO9k
7adoXaSpGhtgpaULs+BBLft9WqcH1n3591qteiqkiiug3yHi4ttkK3FHKEAk+q2W
4XGT85tYkOe/tPKrGShzGUYZRfKToAcO3qY2yj0BWieaR5VF9uxtYGTpc+oWwKdd
MTiEk8rw+z0JW7HsowTDpm4Ld7+GTBo8NQDQNFW3O2ZRpK5+jLvV5IDooFOadQhs
yPrEaznUfA+iKkM1c5+FKQQoWEu4aItozmTnIMyHGPi6OjslVt406dC1aNFFQ3N2
yEuRAtzO/1zNPvWP9PjkM8XfZYPyvcKEvfNPb/ik/laS17ca+Q4z93TjAJIrggCW
`protect END_PROTECTED
