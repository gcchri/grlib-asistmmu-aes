`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TwsZ5P7bj4/Ou0GeOgbP3TUP+f6XCraMWVypAvyby6xYuXDQMEhBrzuUgqIUtytA
orMpXr02WdL8sDOH7DYU+ybfExj5+fOUJcEuFp+EVPcgt74v7JHNywEkhO2OCIgC
FUgC9ivalXUh3N/kZW4fcPa+lLdczQiEBMlWcQ+8242dlH90aR3rpG3JEOvK+mL0
1A+Y1IAN5IUxSfZzCiVAC5FHAseQOQYQGC71z69VLzorFoViFHSl3GwhgorVcXvU
oQ0YgjegMBgws3BKZV5kXppWRbH4eFaPOGx4cr6NHPU=
`protect END_PROTECTED
