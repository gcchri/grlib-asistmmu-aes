`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pU+FyuAHWOGMqC3CODU2Qg30ghmXTDDOR8sPTtTIMGnBByc6YFXMKVUcyn1Aqbqs
bDuxMFE3SPLHfPuw98Jooexr1UIqNrXbrgAcPpJwsQCUiHlz/+x7fyg6pB3r1Wwt
7ZXCT6KFhOM8fHjHh1MsWMTa+v8ahWkVOg1jvJqqRBVj0e/1KHD9wIQEekxTjeUp
ueSlUMDCn+fsY75RgisVO9sYolgfveuOhZJaPTPSbbW3VMX8ciHUMRtEUeMdzpzG
9xf5HozqvnZcgGjBIS0Wcun/tj7rdZT7cOtnKw9J1DHCtBXbV2S9Z2pp6PpXafNL
HoiSCYC/yNuYquV2xuI8W+GHuNw1PC6crXMErLm6IiBZIvvRrSc+Q1ZzON0OWYEb
Aaja5u3XLyI7wEnIgGEFlraBzBHcasXZWDbck+/R1bqhIE8SVtESkRW0mt9nI5rx
7paaUQ5Z5u81f3wyXeJP9OSdy2p8Svd+U+PtZRpMh4a2pOgm3AZVA1mB3BTe2qu6
KDZ3e+I7aAvIL70sX0zEqbvyNsqYnTJeEfrDry3MWLqZRdIHHI0GuQH9gRu6AS37
3Mg+W7i04kLLSjcPmyF70cuQ77MP+wS68Uemv/pbcPlMKBp7vAmFaqDxtSk+0vyi
hW1FC5vy4i/K5KT1/2O60ChzzT7rej7TMYNdvrDrwyYr4GLnqwO+N1fTXBiXgB9R
D487oHlTLrnKShFteonfzN8Ur5NbJVFrib9FoO5c7v/9E4nEIWYzD2Pb++lCeUWE
muC3iRdL0/w9nzveQcgzvcslT3wL13lYQPUo0hC6aRVwXld2z/eX0vPjGCwrsebO
qu3+0ptHxY8AAsX8TpVbitskCIEsuyVsIsKSWdweBbnuK+nc1MUsX/sM5CTV5v7m
DEI3RdalkEPE0pDjhREbNXX/m3hIji7jPzmeuALzCpQd3XGKF5brG18+Rw4kd6rB
IR0AxCWaqphs97Ep0TRc0VaC4lTXSkzZafp7naPz6DyWAX5cd9RAkLhixhQikOga
bWAXLpPRiu83y7Av5KfPjxqX9SedKIJ7aaPC8SzCGvNmWGN42myspBtgVgZSEA/s
v7BjOJeC6jfA19q9UNSyNnwafvm8SndpVo4/CpkrnCJ2kFVxja+cbpb+lY+c1MKO
Pb4bBDpoMrJr9IePEMcOkC0yFo+Sg/7Xy6Pw4CS38SzoiFlnOxZSaShIRVH8mSkN
lYtVc2/L1/E8jZmgXOJzVt1QO2Xn63CaVEmleaX6wbx8v/RIpFM7pI8XigSlnl/D
3dZjgs7zRZKr2YCEeGKO57zhJEdII30+zfWDVpJuCt3zDNfSwakRGtsL6ek0FtI3
nbhxsm0L5hDrHPonri23Y3tBSZbYCaQXaTp9SMIxg7xYf+vRGRhoXg+f4zAJx3vg
AbQLFF4YgAfRJkV40PaD8tnfAZCBW8rAgqnqzfD64+tKadvokITEh1wqEY30F7O7
Rn9n8ljQVOTxaAlhM/b9g+kl1De75v5Pmz2+aBiALsKOT11zNn4j7UH3zGeHmFHD
BSJr2yPjVwFyvY4LeyjDVlA7WWkcXDTrpHKknO8HxuRu9VpyGPOCsE80KizE2RSw
afykxhR7nKGF0Ky8Lxp1F0jNTj/Q6VmC/vqz7u4cPbVW7+j1VKFZd1zWpm2rowcH
H8pi/YtKflXQTx6quj8LIKK2ONNBbpCYvfF1oX8yT3o9uaXsvl7RjrUq3laTT7y9
ndMuScqdp2O6/eTPi7+hugw7AEz5cOmDYBe0Fz1KKPsDam8QuNVloFnH1j/bfRQU
jeNgzaurkR/6JTNaIV72NMYjLW2W0MHN580S864EQaSzpZmGCUJy3atI3BFY3GMz
y8rvetFTsEjQltN6wqqVeFH6UkmbCLKdWoZSUBCTxHuHokiVjgvVqyVCdhyBYsD+
p7UCDh+WeNmXqlqOuXcSnqBoADxd+lHXDelvCIVHm+WYaGi0r5rKBKSAhJx7mYaP
G8eycFQlsMNLw0wkU6/BhTseN8GVebY3Z1xWlAcTyzLNhRZ+ahDpWSeHTzTByXQx
buYbddB84CA8qV1T39oZ1cQPF3kNjQ/CchCKmjSwM1eRuVEfd0pj8WERN3j4w8EW
Lit7Mt2afdaVcltDfOJjOYgDFj2D+BCUDyceKLqXPg1haeiKjHrqof3PL+ABDHCg
Rr63KErPNI7tHi7O+FxYaPx6Yx7wJDWT3qC7eQUWTnqeWk72aE2jBuOqqbCZ4eiT
4BEQGpPejTR4u2T0efYbfP4l5gleWHOp1aZn8bP5zBb4iIBMMJ8IR0Z7LpaSbuH4
IR61UrP6Tp2PbmWDxz4g3jBpZJFY5ylUrUDJk/4pLbFNdxN8TUoAxY/t4kmPWHhc
P3+5JCNh+2RsWQNFSfcCDAXwp/GP6kYKuDyZ5+d2rZ1txAHdG5jb4KP03GUUADUZ
vXR7L4/QNMXGRc1+U7DxLQ4qREUuyhr1Zm4S6GLj0SA0iP3YtW9toyo7RCYkZMr3
5V3VJC3mzp5X0Cd2AK8XuswJmcAFPzXtSmDD5oTrJcWtiO1PHI5lNuOFDQwtp2SK
TvbNqCQdi+Xjs8H6Pq4/RAEzlMHWZLYsg/nT12xK9yvmS1TQn+MB1IQABcGSV3TC
lhJweQHWkOp6Prr+jc1gdhNncsRMMPSVa3PbosOUgUYPZBx0VylMl7QSac10o0tz
wyIq8zf94sIEr8kuk055foeT+YfUIN9VENiR0ZSi94zqGx8r9uHKVAHY7H7bqdCm
dndfO3jtq3qb2U1+/DPvwOVl2eIv8AhoYvEOS0l4hQ+es/gIeaF4o8bM7Pu7W+Uc
eHND9E7Pc8arajF3ChadhSLWMjmnYtED0Y7E0zQTSIqOOTtD941McTBqf0vAY+7M
xvQnNNxkAamPtSMZnHVjx4uD37wgQbi5YZX1DxN3pHferN3zsR/DBgJgXUdZbKKv
PyEUoNgwfCxSGrhJZyyUG5LkHrJYUp2TVi3DwjZloyxmZShA8f9LkKB+U6hrFWi4
MDyGUiqbAUoaSzyZMab43lRQ4EMhAewxho0Mu9Qfk6Owj/APe11nNVySkCVSwJFd
MFGlE2VCBz/E+NbelupgNhNL1JN7+Yo5vlk2h7x+rmIEBmKv+uNrMeFqLUCTqtHE
colHqO1CEThQ7Vn0lFi8mSewOIYKq3ofBCGq2bqgMej3mFzeOW0KKm5uzzHvN11v
z3FFbf1yjjmR0413WR59YdZXTzqBH9uiygtkNJxLQq7mksSZLBHO25e2zQIVtQFE
HWd2sksKTujmLk9/TgbPEu4mHFSH1gRIgddj6ijCzFF/Aun1zotTvSpGecio6ElA
g8C7n6fq8b3UQGaFJK44fQQxg+Wmnwg08oGbwrgGB4YKAXrm7W/UbUXwk4ajT0hD
kNI/nQ2G/auo2lyf95nuhaJAeijISPjmAigt8qVvjz9/aZ5PZxWke7uu8spQVf5v
u6KPDS/+TMvkk/hb6RK5cH+PkoSzHl46FpkAUmiv6Ly/xk5jN/UkkQtWHXbT58f5
dG4cDhMhRSlI57HsyYUiaQiJ+0yijY7F7oNaodt9aokDPixEkIxIVIyTtFMDBJMH
OtzV44OTL7w8KugHCe3pEqeoIW0gtoZzDw4csewTzoqcWDWaJuedOT/EFrNzr86F
D2UeXcQS8QBScGfmquiB+lRptsqk2k/WfU1jZkFhNok3CMRpCWKXRtp0JTXTm0eX
l4j9DQCezl5eNvJ8U8DgqAIefnFPigHZAZR7EOcTQyw0t28BBHEgsOWPX0Fhjdjs
0ow9hWUFqRd1buB6e90JL/xTvtrGaUpwh+idw78F+278h1CgwBZE0egDu04aKdz/
FtScnP4P5HySGetiKPQE+2BTZxqHFCA8Y5nHSldHc96o36e/bDnYsqye9BeyvVaE
xm89JmNTdiVk44p9AHzeoagc260VUsMNYNjSNHQIoqeMuhnM1mMcaMjGFoh1vqaa
MG7D8Qf/7AxJoHbCUEkA0Qju+cEkJgsqPv9FPr+JHc2wn5AdWI6qw+AZDupWyaTO
uAs1XmyQW9R3OUBitsqUDZDUR1Qa3jgPslqKWs0H95V5C0u6z5dz6uIzF1r9B8Qc
bZ12/BC5WVEKa5+mKoiawbIdDKfWnkk6gLPxgFfAY9UbNGLiwZXsAYjCK35fMxn9
tVECg65EcmC1C8ejP2kaNbFTlKfbw/+SIsg8XSnuLr0=
`protect END_PROTECTED
