`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c4ii54tBIrwOKJxfjO1oOB+0Emnv77o5nUqFHnpAGWdHg9J46BzIaYm+iS2bJlzp
55csLEx2L0J9xFXdKLVo1ymrevy7rtOxvnHgNhHoJMbrn0YRPlqeg/kB7qmaw9fJ
97BsfbVPU9vIVsEoIdGCgV8KYV77Era6UHixZ1YY4PNnrh/h+UWH9IiFPwiWqcQo
CwlzajlCPBMIdZdGT5cnj6zGi3NWrXeGGfZzp2ky7t3Nt7ey3HUltdOsVUtc0t+Z
tH0IYxgCbPQkYKPjE+kF66WiGnmJn1B60hHlrtBiEd9+R/kgnPRkkEJg/QinNaIf
dazWjU14MWPoduK1xFHve8NRrboyfbYjxGMvXvOFuLg=
`protect END_PROTECTED
