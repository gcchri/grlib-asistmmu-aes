`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EHd14SIHgjkiQd3FSg14d07ItIBj0/Y/Qe2crtXKdCRldeh4ecNnza9AQ/Kw6ZFo
2H1EaO6pjGZr4BxLvYSGpnOEZwbHEPmDHRKKpUcDMymu4wk3QFD9YG+qHd00AaqL
M39IIneXBjrx2i6wdCS3cGJPBovDxFnP3zhxRMCo05ZGM9MS8WXqnpoFIX+pmlId
9LZ53v9bhLMwF5y/Oq1OIKZq9gYwvkE4w4P2f1w+gc+SqLCeY3AdXXgrWnwfuuEt
I05LSu24oghr5ghYD7djt3bnBHAhdg/1MKcCPhiv9mfvAnmMnuhV7GAtKT1/y8mA
/R2NLuKNzuSDIaZzeQwc6ak+NqlN2Ess5apHEuJe24YyRWyz+cyI7ifyzPOLM9v8
1Rre4AswlR1hzvRPYEk8JpSXezZ7imqI2T4SM44c2vmsOVCMiNQYO+jJkpTIH20D
`protect END_PROTECTED
