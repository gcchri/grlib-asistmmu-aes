`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dpyd/97ShT/4nu/h0ayi2gWckm94CGollwwkKXDSjvCGDy18BQYI2zNahkVrgQP8
AE7XcRTCyBO1e9klqIMkfyMQgthnyvPs9OuqFF/nFcYkE9apf4aIJ2e8rgqYY10G
vFK1K4AfTBlfY9GcVdIhSEmRxnoc5QDNFT5rmSg7r5rudy+55DjeFF91LulIXbox
KqGgY16+kK0o94zJweO4nogPvjN2mW1pKiHTUR5G5MBHsTP2hUrfnjrdno/85CKi
J99U8mXfiM5UmvNcakEw9PBBoJ6XyMviqyQIt764urcKC/rBg/vLYRfdhZjpJ8vG
Kf/MRFfnb5rSoCBFIqwizoS3XMbJl1N2tlRZsU4+net59qB47BGYzzF6K9NeNSQb
dXXOHkXJrj/01xr/pldO6X3cu7bClNccihoTOcqlhV9nzwNqviCqO3Xi+6kgGe+k
rpNcmwrpy5qDX9YKWuSHI079Ue2qPhj4iw29ulqRiPMT8msqW0ip2PEc5a6pT8Pj
SEbcXmO1iGE8GM8sbNsx1rbFd8h3A31e8Z/sOepW2fNv13THNGwUDUtDcsQMOYVo
IqKobFHfW7bHkt4ILAViUPy262mAyvamnMZPbeKOEiS7NoIk4KAnVREyRQo/oeL2
rudpowPDdyrvjLC30cSroITRsF3g4jphEp8gMe9KfLBf4rgbzryj/sm7757WRgVO
wDFaLJuXe1BDLlRvaznZJ3WBqpvXCjgd6slfisHfPBzkmZ3Rcn5X3nxaqXyODPGY
PIGIBTz31tFbMugXlOp4yFkzrhVucY+4/6NGZ5p52fMcwHIPSCKCS7NYKBw/P66r
WgcLxw8iLErfSdwuI3XK6pmUUJIHGTh5QoG+Miiae2lC8OlyWqbt0q3Pt/R85sGS
cgReMVLHWSEfujClLWSmtRhBxGxW5kEitkisXp2FrkYZr1J+wZEJgR2xmxfiDUSN
02EiptGoPcsqVY1SB0P7HXNyMwsu5qnh3kTTiMfdhP/IIFeBH5yZV4FW0oTw7Vva
Z53xx/CgHp+EQKi/g86POhF5TRf+ImSfvSxsxN3uuAxjN4C350wY1eZrx7KdZ9YC
8uj9D90TuhDB1A2OA2tDCouGYjTPNeSCSEAyk6KsUsVmVk7fI61cR0oOEWrdu+8J
fjL4o8eOXGLa7FJRiqNT2CTd70/CSQhB7v9/sExeh24pF5A+18u1Iy7AsZFdsGIx
uPssDPMnOYRp32guSlBQF4Z9UO2OaK5WQyj8EOHoiuLRqQ8UX26cfCeT7wOH5nJR
dgYDivqEhGXNUzvXkvik45VVLZKAyrCPufj6eQoSqpDeGQS+RJIHASxIPG7/7whu
ePzaWGwaTR7x016Q59GDBkuEtPvi4Z4b+oX0jpi7RSKxWhlwWm4mN32b01MqBvKe
1jolPMK0+pq5j7sh1oU1MoeYojIUPvL0OQx2EFQa6nDrb3DdAHgma4u6XVG42yry
m8k+QLYchrp7ILkPjATPA7a9wok1c16S4KqNUz+XaS4QVjivkbXP2aVKlSLN6+QO
I7oNm2qIKABkwMfCxqTZrFIt67DgnTmcEgT5ZfxWhn/x0tU7RL5yY9tu5q35yAcs
Cp/gzn6dMtsQjkaFwkFQbIW7/EE9p/7ZOY3wu+VMVK5qG1Zw1mEuhvzf3u0Afw8I
on1uaKyQKtYUQgM9YkuQ5VzdXdY26sNwt1t9+LDbLbE8OMBXmn86twnDwH8tCNoC
XwFs65mgfMKjw1d0SiH/XS0zEyNa0J2rdoZgwh1IKRsQ0zRxHcI+f96UnJ1bEC6z
aPOlaq1uyVH76zEky/Y88gjHNvxesnudQHgkZOlnlu8RjebEYrxbJykLPXnOrJCY
hIrgn8InGJQQQbprZdcE3RP/6CKXTB9oraypCprAnpFtqObT3Hoq/YV4l1k2JVU0
zs+EGCbLxL23pixP6Qj1JC2Sniey6oxEPCFRBu2V1cSI7x87q46EKgfwBlhUuZoM
kqAzqrwj0xNhXJ6kiZ4YW/jA6fp8Nnmg975sjUZeUa1LThouuMdzyNnYBuSD5QjS
XOGGOJfKdvJ1U5Ro+rCQucuy+M3zuJ6J1bSeneu0ASECmu/BR+m1Z+9pBX4Xt65t
64253zmzoyMh3O/TolGNu9a/Ov433ezjwLYv2kLVLzlVMq8FMa5gckzObqeQl1qe
jTdHgvr2GgXT3DDC4MN0109qGtDtrqU0FyXkdUouzBkw+s/WwFcDo0MUTr2vqH9K
auw8dx4o9e/1ZODXVEWSzw5yp6lAfs044/dtUGlqf37K8e3ahqotfsN1FKMIVExk
aebshPp5sDwYNc7xcLQ4GApACGsJ4Kq1CCIFnHcdP/G8KfGWohe3huu2TOnYtahZ
wjWjDe3CfkdM9kHSzsVhN9fSg5gV/0SgUo4Or1CFOC+44jwLRK1hWiQX6SbfMyWa
y6m1cRQG2tTRyyseW/F6bEUjXZdwN/dB4ZXRCoVNzU33plqTEAckxu4esYXWDuBv
9CXW7Y/SE695QQdEE7VzjYcchB++RQ+Nlj7/mj86hOflCyZMo9R5dm09ApwSyAX+
hd6OSPhYosn4x1dc4F8ka99FwwnkM655CASHNDJKJouIQ4NQDzV/yOo4Ob8V4Hf5
euuPI/Rz7SUm+CmAt6FvvQQbK9jn4L6CyTRo6woL5IA2lRc3ATdPy5hxHjg2OTT1
eYrpniaJQ3wv0mbwdIHnnOoujtF8gRaYNsdf7zLtHVVMyeUH822TLGrc4AIyQ3CN
SQMP+hLkaUNvegUjwWo34oYVMkKwcYERMxWIx+ftrAfR8O4QPvAWHLyPODLcAWdq
I+SkcTiLL3Q67tXaw3JH+6KKEklnGF+kw147k1nLxKnKkIfP7MN91cSPn9zJw+BQ
BauvqLXLFGtZteN9/E8GtT6UVlwb60hNHJHyIso9fW30EFNLTjuiyLW9drcMRylG
bSMHywSx/BXzNUDI11riVODoBbZGX2Zu0kEUatC4PGBL03mnZZi7QtAZ+a6tOngO
E8OfaeiN/29W7+x0E7GefrPJVUXiLgNFjx6soepkNwprcZBhM5+1KMiErAA22TIE
AJrAG3E15APLoGYS8P6Tf3AlLrnXiGj8ldZtHMdYw73t43IfNmwzjKnXO+RVm3Wx
P3S8QoNKGa2/kqMdPyA/F+6ZjJjqsmGqVezg9XUbHuWLs3uRJpMEI/XS99LZyYZw
dRZfO/mN2kox62XFsBJG5HbeKT6d8C026CFLMwN6VstsN7+TwKFeW1Xz4SI1W/mA
hGFYspPNdbaRbU5aJR2l8p+LuTCJVPyRElaX3ZCmwFwYKBDtPl11vH9IYo4gEv+c
d7jLVEUgEW01K9+w/ArTjcvfqW0EOUPEZxWo45EuqIf8mfM1CjDSsJibn1A5vH5h
dWHPT0qDpQDNNut466dX4MUqh/AvpSs55hZoQX+bnqEHoYt4PeRimXfro7+Dw4HA
+n7Yg48iqGULRZbeU3ATOq/0ym8RiCGA05Q4sXLLqdqQ3dQKn4MOWd6sRDadZo8t
UMThbMKBGyX1SprIQfsxco6R4O9abjw+NaBDUUBXld/JbJby8qMk60n/RP1MumPv
KlDvakpBHY772/tkXWinxmPY4hw5X+B5UFx+XnSVc+cjUS3djasVDno0uDFOAw4O
`protect END_PROTECTED
