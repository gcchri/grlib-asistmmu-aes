`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
axwx6jyTiUnaKzfiYcRMbbeYe4XEh8TqCEzqYoPyA8tfYDrLcevGr2mTeFF8gDp6
0R7zFCyyG+qvFAc9TjAE003gaQ6jaQ+LsntCzAdkuGkLJUOfE/EV2GFl6onqd/6r
S1RitxDsRQQUbQ9zfh5WAbNa4DJjm/bExPqZhXX0LJyxlm+BB5PiXkYFuvmnkRrq
zH7YZtL1wkdE5NKsUEmMO5WDV0O1AUDjW9MeGrRpJpDVaAOuwP4g57t+ijh/HsEI
cD3kYri9HQP9Ojd4mxamyETKulsyw4REplbMJG+mwHtoVwLwtfzkUW/Qk+WyYctt
I2j7Ic8qIL6lobnWtRZFIadhaRrxRKFBmKUQRlbRXZQfZFDz/wYYdQfKT4pKYvuZ
jxpMCCfGjtMl2lhn2YVjRQHs954LL9VN2em7NyFQzpHiFHYejnT5cRNFrlaNh5kt
/jnlnWAb2YoPYIJtJ0ShZmdhZYdquo9tebmYOgGuqanEY5ExJo8PCpdc8WKbcOIj
`protect END_PROTECTED
