`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
87cAJDAUNGhr9l+n0GpFtzd2kz2rdOqtnAbvoyeq1LrOtY6jHc2F7ggAbThOW2w9
dd/4jWpW4BTTFCbf08cCSYNeCKxY1x7dhQ9Ig791qYAzbJxjRvSPVokr/MSTqzZC
/wLcyc2aXAYJOs8tqP8+1UiLLISSYgBs85Bx0Au+uIbav7syNjtBtf8OcO8QirWl
fJRbXLWsmZiAJrr2/7wSdd4UnxviYSRX6aWTOv9Ee3PzcWKSOzB3R/qQF0GmsYYh
TtwU7hjw5rRIUyl/m38XXVVh+FhkLEJ/BBSwnElK0Qxn8AwhTKlbM8zanIYd2wzj
zoFXxV6NAle4uYI7VXFBrcIIadfGNeIFejGUUsr4vZtxE6syQMjsQGORqC+K8HlO
naBKjtXWhH5qjWw2obK+pRq77utLDNIz5lCKn8uZycG2XXvhLn7p51BDBwNu+U/B
`protect END_PROTECTED
