`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Wf3mqGH6P0FfE5LA+ufwWGFaTLHrWW4WVSodDHGARYbYQHJV23PgJVbtTZ8KkN4
y+VJZHR1DK7L8Cwu36qYaNYJKY98iok1RCJAK07ciWVW5CbRfE+Uu3dopVKEdWO2
80wf04U7ZLSHGiPGZmyUdeU8zmYWuar+8NmPJizVDpwxBC1ft9NtxX6FN6erc85E
t6J4ldnj2j4ZS+uEDN6b2u60xNWuBEf7eu7rgO0wWUN0qudWzTcj+BmT0mW9rPqM
eqRQ4ACqnnRTjmoSxJQu4RPqV7CQLyfXKNPrnR3m9TPTdhFvqOfjMLmRiA1rkpb/
sNhxa+Sz8EsJKW1Vwqxvbg==
`protect END_PROTECTED
