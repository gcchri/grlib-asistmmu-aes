`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mFEPSfiWQh96NdHEgSOTNL0vY2zsvL8cl73w0qARGvW1cOeey85/e0oJAQa24vb/
/ymgxysPScIl1OAd22E21IMpCwd9oTsPUiyqXj2N4V+QmJAxt5YnUiXKWRafgSZ0
VVenk7WYtetiEAIHB2joBQ==
`protect END_PROTECTED
