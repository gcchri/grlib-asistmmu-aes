`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3YQARzYJUVh30WvGbCILpb2LZqeI0k6FCsj7SGeLuDGqmaK6xvDOAkDIwEUYDWh4
FPAoKek30WoCaJiC+10GXN2ZPeHvBWJp4swMBPUsZog6P1HzU50YbVWQfYR4/8b/
dDmTueeWRFWQmQDgHa3TCL9cxwITJpKZ+pLnC/y8eK6WLCvFBY4FB31+jye9RAIv
5/e8nX9RzyZb5/xSTjfMzHMv0BfWJ7R8tiKILpzE2IkLXGdvRkC8jTr0RGY5PZoi
Y1iTKC0oi0QupKCIqoo2snGy2hg7v3WxxKAELfFCaJV2Jx1dczvXNoAQVBZZQKLD
nsMAVRVnZPIG7dxtP8lqL9DaZO2RpLW5WwiZKF37rLxkaRu6JE71YPRRG0Y1lbmr
035s87sREkKpicG6znyYxSIsj0N1uxRa/IJJCJoxnip/Uur/ZX+hFfUr1bGicfVp
RD3KzpbzoY84hWkI6fxZVVOEWSbI8GM4iZRO8K9LE9g=
`protect END_PROTECTED
