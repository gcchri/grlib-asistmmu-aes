`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2O0xNz70WpPRgQLVEfqq9/nv4ykLUIAnl6FLXIwrJbtbc6tEwxXRgJKojRQSVU4o
3COd42IzhiebLaXNR995kmwu65t/h2s+Oe+GMzIYnOOAvrCF6zW6guZGEycNd+7r
VuXFTzTnGMI6iJzPYI5YWBAar2Tbkd0M7ut9A1ED6Zy1I9kAaV3N2J96ZStNOwvg
WUCFBHCooB04SIpFZXVjxTFGZeeN/nWnfBHgds8QzbLnbnQsMAQZZQsvmiLF+T1Z
THh8/JfgYvTLVg3iEYiCdb4/kwOm7YCaTx79l/s0p6eDQycInciWoxvnOMqA8Y14
a9E6KJ9BVRrkGHbCL4ox+bYkWJA4WJ8pFfmp49MSIOaRkWchVmM7ekQKomSYWCEv
D7WxCVXvKoC0NlQngHUapKc9m0S/i2DcDCfrnIsXdiLRDH7xzJQ99lNh79BzXfLF
8Dvpm1pmjlQI0+I3VVRschLMl7kdSFzcfeGVCjqlmluTlo6zx/PLX8s/+kTy0S2k
pWA18D1uQJk+jHMK57xrviDOTTh9LpqmWqgc0IQXNKrwazS//+S1Lrqu7iu20z1f
yIyu8HJScDCf7t7wo5ZHnkZHA6N1pjpTba8aCqKAQ6rV7MPoM7hmhzBETiJp199d
BfCfvNKjnzS+9FcKHAse92ec+jJqztT36g0WfrHSnn1e98JgvEuYrh5V2aaHR9jm
3RAdawR8/cEPzW6UY256a0NzJTOpR9tgeQwRdfMz5GbulV8DCoPa3dliwKvgLl6x
Wvkc51JneEGvfyHUGtD9bA==
`protect END_PROTECTED
