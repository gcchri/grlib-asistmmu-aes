`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IGMcKrVQW/Fnz4MbTmNbKoBieAmOlJ0VaTjJbIvuuvutAsVaBRMIYzIoYIOwE9LQ
UZXocWFzcmAh5iPFEMJxE0c29Q9XtkpU0IYNTNMc4Zz/jSWuSa0UmqYBT8WH94F2
NiNYEQ5gPt82UwjqrO1L5Zqh3Gz9swELcLJN7fJjEtWR4tNMkXwBcRdoRta5h6vv
Jw4JohqwV+/PyBFN6uC/1Jez0OVLEhdUVlmzlZ6hqal/krUFq/zbJxDyLj/f0fS4
b3SKegl/SfSu4gRO807buQSFlqBZbri6ttZiZ7MEYuQrah6CXhkOiS0iJPRP6upd
fr7Jvpe1PRDUPflTwMrsp3aQucy9j/9EEzF9+NhjhVakL3xu4JylY92159r7IGXI
IRbxVxQe4cbXea2IvGpv9qmoQIAWzVLxjqgEOBVZ4mlacNHkbOOsr3hFz34IepbH
hhuJMT38yKu3MNPQC1nmWIkmDyES0zsED2suZbb25aLuN6jljq6QbQHoQbEtGw3v
orgYIcu0uRyo73x/SdlSGOKs/BnIZOnRAhL4C+rEaavSTDmMUFX5kVXLXXcc82iz
6FNtt8uL+Agq911/WOwsbrhl18JbMjc8WAlkq6Zf4P9WIz4tyRsRPWkr+dU2/sYS
hlL5dn/7kkjNvwK/BHSOVXDKLosCxd6zCH+gjuYyC8/5qRwuMvaivLFFmtGGXl2X
fy/Jk+5FIW6ws28pi9UKTBmdCBRDUhEOeHdrua07is/W6wQ5Lg108k92UUUlFe2Z
XVAcF5bCrXpmBE0y15Lk9Rm9CW/e34rPEc/fx3aUu13bndpcvyWSLMhQSj2tsVEb
OcOcZbpmWzQBOkAE1pHZiCFpM/fzNHdsKRnPz92HeXmMT+kwHjU/rUzkZGcEmnj2
hAzOThX5W/e/0oiqUVXuZ0h1ccHzQSysfzwDjgR280hnC/KGRM/iAVvDVV/V/pIL
IxHeEDNTlimxvlVPSsVzT1yDz4W56c5qpxQu7I5wLerCjHkImS+Gpa1M/aXADkuq
a3Rz81kjydqphr7ikDu89uRzcAiqE5uuFtaceuz7HlAoLRVLK/gd20Vm3HnTn3o9
LpjyBHSWJ01M+46FFUI3yEYIEpnZbIG/oPhny5ia6AfaE2hpZVX7F1FsYtEPZAP9
bW+VzTHD+Vs55J4AmvMhTjjdeGGKhcbtfLFQRz/uzhceCvHvHxw9KcOQFGxtcd/k
zyWCpZpXmlCRIIx0uvHb2+Z/pZzUWpuTobVl5IG1PJAoCiLZ2TAqP6sfQwMaBIDW
`protect END_PROTECTED
