`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pn3iGu59hYTW/fuIRs1qsPH8JzEMP3/C35SBIloPmMmN1cV4r0EyZ5AF3l863wpk
v6PRDZ6vl+eyovfM2755A3HKW+/U2JfCBFGKR7lgbaMPbpGQmlw+enX0zWnvK6Eg
+q1PRWnSEZwrTO2nI6y4wBed9pFGWFCT6ehZxBWDwMzBeEDGwjp61xpajtqtubDj
u/emgI4/FvGajLPlvxiwLP7kqesrxSI1jda6+mT2/9VfM4RtnkFSOgRk9jVtErmb
msIeRlNKpz8sk4G4Z5KbDY0FKS1k+eRfNzcYekDJmHLY9eIgESxk2axP4e37d6Kz
kqF92pzT3wUyJJclnPv5m0uRAXntvnBLzrJqO9w+xfijvKUAtnDxJgzR9kjpBG90
URuVDLpDtImASp1AJ2NZ8FtwCVg5e9hy2GieWwaAdVOpwi+L7fy5amtR3Z04stHl
dBi+f86rE0tDMK3F6Uk2Xl9fGqb0bdDN4yu8xTD5h6pPEQaw5qgWTXoE8Wr0SZoG
6wUCIzwClffqTA7TvI/OCyXhmCEFc14UM4orTasYp4Gosx9AH0EhQymolIh83CCB
ogm22V1BSDA2Tzq+LcBO/4fCBkk1KtB0xJnqb6c/P9eOqDTkry9G/Ox8EL/P4sFl
uK+hySs3UuJrRcthSUuphSAIcEQxIDk1E699j3PdAsXq5Ktl803dIFbFQynWlGcT
eL5CFjui5GmSQf90yK4Ai2GyVaYN9HGeva3jLBhvJb7jYVM6t5ETsd7VWzLRiYBX
UrHfuMhyBu6yj21WE02R+KRk9JCgMEiwwbvdX4cQ3PW8nK+eaunAGVtY82CBOIxv
l3fMklF5quLzdRPe6nSsvsUGc6B0YJ8U9Fv6/g+wVc92Y6yg2uDIqqZhDMwh/1WZ
3ANbJ9H6e9HU6xo7CRIDqwUVyO1o/GI1g9S7vCaiy0X/hBiMiDxmFluDnM5zuEzO
xd3MMzkA1+f5626SGD7lfcWMWbNRl+uEyOaB+EAwOhHWxWA7xnzB1pCAdxSqZ5u0
OfQnT8heoNRv3Wny3SUJ+p06cUhcphVXmhud2G4pxGZUp/uPjAVj0sDqUAsSfia7
4ZqE5eLRJKSTkd2XoEdwK9l82P+2hTyV19emNY0zGInraAnG8RZpy+wfaV8WLD8I
if8rYx0M3zBZmAgFBpFNgn5ZlwKr4if70l5co0UyiH1VmMrRr2kd8jYxMax58DSx
NO7O2mjuGXu4C8wTGw3WwQ/e39BB3VJtT0gZsIaKZk3PtbIC/BYoIphEsASi6/4H
Cd/66Doaf7a0AihR5XEhFonYx4IB46Tw+L8jZO3NaeLfvFBvUV5nNg8wGh1jNNhY
NvCA2uyltmT04AM1gK1ogi0RuLPnJ8uGHVxzUefHRd+qQWrFpiKDvAGNF96GLJ9e
HMCERdPujNep/taREKf9/J9lw4Bg7IBkzZ1/UxyZeHEc4Hwci3fxTXt8xS5OusLG
/0etziP//aJLhGtZzIoGIOID5p62y2h3KMkArg8HEYmYt8Hb9Jx/Loah2OctwTTB
67PF7i1Ec3DQ3TjY2xN5K7U/PA2PisLdGnSwqCLfh8FLNd7lh3PJ+RoPlfTq8qV+
MPsz9uMGLCVOQsYOcirSL2pg9mmtQOxi2PsT7V1ACXKOTBtmQuuOLBHMUt+TbTLq
a2WXN086Lc4TQFTFku5xodbUtcOkbP7geKrvqL2MhbzeYPyp4TNM5V59AvJuHPXI
3ErG9/UliMpxck/p14GDhDsLKd+Yw7e8ljXg0hxjMPvAQnLM6fsPtWf7Sk2j8SD8
VhZks6t/dZEKKukm18rl7Uc5nVNIkTNdyrGYsJOeePkFDkW/Xar+RQxZXNzPHTsN
/LpYOVmvNZPe+Uw9J5Jddg==
`protect END_PROTECTED
