`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oV5/KS7X5FRKW18nZVv5QTrI5mdHx0MUnrxnVYwSe6xipdoMwfhKP1m11Xhftadx
Cc9DBRDm97KBN2IBuaCejkLtcAmuzxhfRwLZvNgdaWvsUXgnqqNmDZUVcWZlCyiH
D+dfF1UDrYLJRiASK9s42r+Ic7KE2yGYLspaxqGFqveXiwpI0DvSLs+z42EwISE9
RfU/PTuyyCQdNvy/ZjKmJVrGqJ8MaOg8dQBPUzs4eIsepm/lk+Z3D+jv9ASVpGOb
iCftj6ZtZj3tGJ3L5iFKQPXtsuxLG+NxKLh5bzk0JMJWXlRflwjWs5w9S0KbbRgY
ylLc11O/s+OuFwkOLLnq+uW6KZiBOAoTiCjF3uEg+9k=
`protect END_PROTECTED
