`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kgihv7lK9ZTz0rLz9QTWidBdlXRwjopRE163DQGicqeHM4VK+BVx8fZ+otISSyKa
rfpJD/vspV+zcvZz3vu9vf2X2SXRfTqyuCavbOdCbxkfGP5YBz8zZj3zbphTMuKR
S9fAhIaRo904LIz0TnRzxsspi02Ikfpfkz4mqEi9t4xNEII9l4z2L7X4YJfkz63C
92LhKhCjcZ/2FybymSFnTgALhNUM4p/qER3E1/ArajGjqvzIUPsQq4p5A6U9f5Uz
E28gZ5tV/bxWj4qiAQN8odwmX1xduJDlNLaTRQS90czY326pAqKMv3AsnkwO9qch
Asq/ZjE6CfA0eYN2rj3GthWZ7dLpVzrunHpOxpdPyEJPI5Z0wWOSd8DUZBrjVpYT
0/snsAOyNgPsiXi7spPfd1xHJ0VuCQsybZ1+iXdGX9A8UTU1EBfvLYAKHpotJiK8
hGWyIZ9gOsRpNXP6LIxmVw==
`protect END_PROTECTED
