`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KYowr3xFH1rzt002zgZSET/XuV/dFzpJZ83oDwCpCvb2axDu4ijkjatzqT6mZ+Or
o3kVNF39yoAymCIu7BYK9AhqR6MAGR3gnhYhZxk5HfVOwvz+BaGxtN7/adIQn3wF
cYZ5K1FveIbcH5h6VuoF6oO41YfyNgTSEo3h/Y27iaZfWZyvgMPGWWSWVhEWddRh
0DjPtalvS/q3wMeFFYYYBNMS+r0ozUuN1/RdlNPqKCBoT1uJvkgxNOl/XId6VK2k
R+HlkO4/n0W3KbDUS4kzf4ehHg/dsKdBTDVHDnuHTBCElVXtB6CPzU9QxVstqsLz
`protect END_PROTECTED
