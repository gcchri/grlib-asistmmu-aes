`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sFrvS2bCRp5qGoffyI/e1UTE9HlW9fH7T+nv2pUQ7Rih+KP3IiCH0jLwWX393dZb
GZyHH85yNdKt/ZJ4j3YZndhROksSPBHi3vGC5eZ04Oonb6xauBB19jJrYtH2gPUs
HAyf8PciBkAitYjbod5WOPb/vPk4QI4/nxBxsbyHpHN2mMbW9k0vqPnzh+GlCsoA
2ncT7jU080GVTf2Q2lUVNI5c66Gj0f3eESFVLRILJSUBT+gOOBo7vB4vjmw4epBj
I7/lsWZQg6DsM5VsruNYYCF8kY8mp8ZI4j1/4bpTQdUxuEBUFVJfPCCUGqk9OtoW
2RpOXct7SzU+xToOhJakzeJMNZx8JPjnGQR9AU5t7L5VRiDjCV5u8zdem9ttkOe+
dKJUp8mVs7F2wOUyxLKDJDty5c9bX9+zmtb9EbP4cX+UfmY1k+r98beOnpZBAJKO
bmXlcH82o9phpMLsz3t+l4aHNcEenHlyIUgVc6hOmyNLgl6i/7w9WgQ7YjJGc9th
G14kXv7cs0o5wdKGr4Lkh7JAJSUOgr5W8ZbxgyZA248Gfn+wIAet7+sDIInlyxZ7
8Jtf6AaEbHy8B4XQ+bzUWIgyDwb8LjfpMsDLZ3sW3Bg=
`protect END_PROTECTED
