`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bewLAikS/RlmfrojCE9onsFi1XsAY2MHWurLMJ+hUZGP2x9h9uy1xVnjAfxqmHax
LhHdqGrAOWF+RDn47Ecl7lB4EffQf0HPSG/tLcj1Tkwj3uZQT5Cs9lqAxgLzqRhk
TQtNLPOwYdkQGUAOawgzxkSNfvXEk7szB4vxYHhtphpVQ5X9mtM09h3HQFOVXXyr
IkTh19h8ber0Otkb6sEvO+4cbRie9tOJJGX7XtPQtBd0le47Vd+XX3xaUPEs7RPg
Q8SoKgaFnM+QjXItyYKdxRYsvlrM/BeXh5yEZIo9HeF4V3eLVADMKWTisFNv4Frx
2IPcxLUUbUPnfF0eFYdPxSYs5m5ZkLEm8VumjJDSRb7FKWePRBb+8Unc0tWEIXSx
JUcH0Mx9QxykWzNiW6RiL3fP+L93Uk0GAODYchRJyhs=
`protect END_PROTECTED
