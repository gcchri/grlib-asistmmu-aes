`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HK8OclsK6zzWmqVlf9xkhgiehSpoAadtkjUFMRMRYfQieFyCmP53w4eD7kT8Zhgd
An7wXx1VjV7WQ+yJwtRNR1uBL9D0NsJjQraGZH8n+wEflN8n2o+PvLeA5bGLdKnS
0LI7geWs9v8Cf0H37zEQ8g2XgOfE8I7pkkXfJXfk2JWT0nbt/7Dd/E9tRB3NlZWd
GbkFQaJ6avAyxLZzm+pW5NcHExdK6pVBDwZb/8bu3o2c/8qiAUcPmcpSn+toanEm
GvD418qZE+Dj6hoLqyteqHAYyQcfFtdh/FYfJzopWcTXrC1QMSG+BePJp0OabJvP
vz3qrgeLVJugagkMTAbnBW4nDV6AK3gPzOgoCy/f5PCrSE7MtSl4cuHEZqc36AYB
iO0oMmHI4VnPIOFLUggLZZLKyI1eYSPMdiFAD6iWMnIqTVkFMn/QrSLqdR/IhgZR
fPOhqHFzD9vcMSEcMA5MS+1wA3ZAVaE9t5xujJQMQzE=
`protect END_PROTECTED
