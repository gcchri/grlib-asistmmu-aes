`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2mUz/gHN7rgVnTCMr+ysh065bzXKIKnla2SaNeA/DZQSepipkphLR6SvNvdHtNKJ
BRM08H559oFrnPPPTOQBxxe5N+CdgTE5v/Eg3UqwUb/mjOSxcb7kjwsMnwam+pWs
JP8x7CkUAfU1hsWABDuA3RadgEwXZKzeS4bsupBc+2ndZDcguHfvIMxIGL1467r8
oDmixWccXcQMVO21NXPfGsOSkhovtUkNytjwXSFCJyg8inbNiNXxr5InrFOrgO0H
epHw7KHI9m7CfAYsaLxUrfEFCnrcK+nktEGDJrGghTV/cAj8Ur7eT2ZIzohvkH2l
UgqIc8w0RpFx31Zfze+nwLDSPz6YqaWadGrEY/rvx2MCu1f58rKtrwRi+Ks78hU1
uQOVpwd/SySVWoz0wOlIdmRp9Y10BaJxoViE9NAzy3Qit++nd4hS3b5FfDvzFeff
wqm9NhP0ONnXjTlHK6+X14Z4BrHmqvgCzKbBC856AwWeoBWpsqPJv26wfJqg1/gL
FnamE03QOaK83YNj00b84SzUoae7xhJEDPBgq9IzO3rsLU+wdzhkscuaw0iM/8gp
L9023fS4Vr59QPco5PulnOorXjrq1Gqt0VxwIzgKMKZITikFMTJto1Cn1Vt6pCud
EVXIh8Q4NeaQ+zKrgNb//Z+JsbubteX4sliHp3MgL5+uF6DBgJo+7s5Mr6rf3f0o
LrVTBzS0+jpuJxCahPIiQPBASqYkdWkAi5wDFcwg8l/cVRNLchE5pnKiFyiB8T4x
mfkHyHUUQ1fph4M3vm5iWm4cyRDpP4lgfPs2digU/uHVGVnQXPkOnNonHuDwJFtF
`protect END_PROTECTED
