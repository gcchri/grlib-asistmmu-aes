`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p9hO/m+QNT4aav/vwEyG5KLOmZJRdnpHFfsHdsCfy2IPb32bZnhijxa1h53Iy+Nm
BBS9nOfXuYD0PYTDObRdT0Afo5N7vlx260A3NT2yhHkkKWjUg9lEOZWDMqhW3nyF
9zNa5PAJakwmCCpxlwWuRLgjs9Y4GEUfUT6sHzSOIK9ySJEPFMv5gVzGFCLc5MIN
fRKs/j8iQOyvDkfGl4tAJ665Vf3uSsAkomYlyCMfP6Xgi40+0Hq+Jc2U6KYr4Z3c
kBbOGVjdd5kRm83556UNFIyJymScefEqoE0gPJXgYxIvIkLWj9gkttRMWc/kcRsV
CEhBRjrLEL9t/hZ7A5Ig/ZbS82p2owl0A092netxgKOsMM9oVaEhAlAvD7VDJRgd
`protect END_PROTECTED
