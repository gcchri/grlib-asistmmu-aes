`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2yQvMLScQc7pMqA5ughHXL969cv/dx8ru7Vsg3WMxYTfXdoqAFVZ22p5mKLdVvoA
sCWiSWx8p/09XlAYsUGK7llm3tXFQYNwuYBCx3f5WK+5LuYSkf+ITSEtwUzIyGm3
oqJOUl/UXF63Cdsj+QHGitxNIHIlc4fqDLGEHIRC/eIeb+Y2P3cDLaC/HyMzip/a
wgVDp1zEAygDYupUG5nBk/csdes/vjgWdZkTTZasU1WKAjDF32Nh2ou6E7KCOoKs
A6XHwbEtws2Umeec6VhqCNdrvpldGnUy4asR3UxUfpmAyv/Ns3nvZrsPw4Rc635d
+qekliUImzTprKT7PTUc6S+QcLX2qrbYRGa0VopgZhkiL1KiPnTpep18efWEm7UG
gEWU2i8EKFMA0/WzcLDR53piQJc/B9EwMGhlpnFHiX6hXff0HK9k0hN81M0qPqKA
Mjcvq7zwvR7+u+gck39eJOoPeckQfE6hqvhmupPJ/rO8+bYGPpGSwjhaLCi4eUOB
j9se6lKgEqwARuEC95IhTB9QeHTyMCW3f1nv8vMWSIOXbsNV2NlGsL35oDU1w6No
i31AXvqtyXOtUosES38jAaPEFccXG4j5AL3QkTvg9BWCfdYjof045HrxPhcKaGEL
oCrtcm/5WR+bBzF+oZboLYSGOiqdGEYcKCKkfAjY3lM6awMJMnaSH1wfMfUmQ7ye
`protect END_PROTECTED
