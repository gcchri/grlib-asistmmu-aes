`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T3IQo/a0f10bE3vpY4e3sinIKjVIYoPdevimZEhVP8W95pRrWoG69J9aV4O50tLB
hMlgudKSVPssjgWT4N7VrRTMNHpGlc5i7RfEgeslM+ILp84kP9MM4qdinZzN73Vn
YUbKpjZOAYCnkuDCekWGGQWdb2DN5Iuh/N4n6+2k5nCEmYQ1DzPtseIhNoPlDTGz
kA2gULWjfWcNgqEAAkdwzrQM19HbLBvPJwDON/GxYH9ewRAC9Y6jML5E4ZvZbCcp
w0fUv92ifbDsFc9KxsMfiVrEcmje46lZQg6puDn8ve+NMWSUa9q+EeVvREqsOOCK
N4X+NdgQdrEp0T37W6ALemUInB7rbjRCl0wT4/qDWNvQ6FmBb4F1hctiQjrkvzcc
lCM+UYjV+edBt1s48VxR+g9F1T2fw+ua7gMxGue+lkwIk1YVLxoy59mY9Ev6O/bl
ldSGBYPU6UEJGks6SK/6At5sk+sLv49TjIrMQeQ8GBhB2K+EGwROwfsGwA5iR5SQ
`protect END_PROTECTED
