`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LxrldtQPMOf0dN6+ARytLkUmkI7pkb19bnz0n75iwU5qoOqo4rJxWYxOF24de+GV
0+76XzBxLs7HV087pGOtoAQ4kvrmSNA8SQXHcPjQGgPSZSNXxyQLwa1lsCE+UkKl
zu5c1j/y/ZXPTLGryVev2ck3Boluct7g8MlpkrX+sjGnfBRAszt1kkxRQaSNzhwe
idHOHXKqYYeIcE/ezOCmDTuR52Tr0aJI0gZTObY9jEAZPsO7Gupu6nu+5+B59a+e
Z/xmloMSeyLrUOcPuQnpp5GkmAOMnjNZ9fVWfL0Nkdcb+nsPf3fAvp+iP8CTzyeE
0AuqDHe+cFzqlaiU5qLWjgbxfn9uPu/LgV40xRiumVSH+44HMjYp88ndevMF2sz8
ywuA9qrqM0yh+ALJfhOZOVqosGCQgZNoWMmwvbs0imNTNVdtcHn3nxI7xoyZLJsm
GvYo057Ovyni1F19JP0nlwmuvr7zGOX7xWJfOBOmrp9BFa/V6JCUPtK0t9nnrU8o
mKcQTL5WVa69L5rgpcaVv6Q2i8QXKG6gZR6KxX3IUJkx2ccdsTc4mmdZ81gZ9cXN
XWBXa6gusTU3jGJgm8sirn3RQz2GDvBAViiGlmWwdQY=
`protect END_PROTECTED
