`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o8mLupsdwDi3Yf+QWAvu4cQNArkKeOiiFKjyKUj1sT/pKM8hRQLgTretbyjt9oMI
iaIIEbPej//luMRaxjs6iIBaXvynOQd/DdiUFsyLaGvxO6ue0i8LV4z4O/acXXPw
Q1ow5ZgjSs3dDEh70W0KZPytB06AT/tC7U8GpOC0dZmHimaq077ctNIAmZ4HhNuv
xQQxdwDXW6C7sPSUwlXQkxW4DPiqCqNMursgo7hVUjnAl8wL1TM45zRtn2wGm1cL
f6iYdSzv1rxnsKTiivDt9hokcgiSPqD/COdyIQ6NjjORzsOoUClkCGcSsn50GbKo
D7Q55fl13xl4cQQsOSs7eH8QLhXfj4C/cdeT6Hs5ZO6yBZIFv3EYZuKi36B4DjmT
GPD4Pgla5isOdXqTSDa6Liii1OwolLQ7d+D1bBd/xCn+u4qnluqFiUlXOO/lsyW1
v0dah3SVpqZT8nnOrARgv5gQuwsYFBGlYt0WG6ANQBli5MonzoGxPXFfv+BaygF0
3IXuGOxBKtBG+gPp02ZVsKMOFcE9zbF4fpRaBnBsXhrRtssdXqlQNIe4F68jWtYE
VPSKAaM0Clk6bKDXW/wDVF7W1A4efTCu1HOKGqvwO953t7q8/pxq7SK2kxoUJs27
RWpK53W0BbiTGrPadpWpcApJ9lBg3Bu6EQEbftdQHRM2eEI96jJFxr7CQ5YESiTX
qnJFwQ/NwR6W8ktcxVxmwVCTB5ARRrtOkQrJI2lqzubEyeII3+lmjec3Vuz7CJBV
BJco2Oi9nOFrWctFhJgf/g==
`protect END_PROTECTED
