`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3rbXevt73vrCQ+dPMGDediJWdT7jCOK7RaR8Qdx5Z59M9Rime2/ErWMhX/QWgWCE
0vmdI4dBUmXGlU/xqmc3TGJog1gfJwmkpOy4ZhPhANX1x4NeNGtIHWjeeM8F/lOU
TU+A2Kv+6Rnv1PAu1T8eKAdHhq2/TP3w98wStFcyae6rCueqoBL9P1TzSig4Kyy6
RZlcdvltdrprtSq61pxne6QnaCXvz1oIw+qVzeAykRZ9+ZgJ+/eOvr0Gul4LGGOa
7INjuVOujJsx6S85/5Sgj09yzkWO0+o/6bZBrsypppxZ9GXInCk0qIJOFORilXFv
NBcoJoWjkprdgOnwhqUD1w==
`protect END_PROTECTED
