`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cOKt+Gnx1y4Wu16DiTE/Xp6faKsWWcwF/+w+ExZxd2cA6AJsPm51lp9rJG8qXQtu
bydiDsEukn949d2oLMdP5FCgZhf5S6S71m7G3lCZ23OZlSk4o3rfj42Y0flxda8C
19+sOLlGPyxyBvHrhE5MGI1ivTJrE3icBcAiwAwgnMs6VBnf0FbufUBpz/5V/YQ2
wHmzTerK+o10BPsMPOSyhcx/3yBIRLc1Okvh1dHcnei20RcfNAkzlLeuMyLMe6zu
5DIljnqMGfS/usjPo4O/h33aOpqw6mMMckkXSzimQyo7lbeGLJHYNn9ugnjvM1yZ
AMu2TYxbwm3fHxZxGdqnanED654vCdAf/qIkF2ek9c2LNsIELjHI1qOcD4NivKej
dKQP0pI8JzxO/dtyAbVoUyLxwayyGx7Ui1knzdgw+SYLXfUQSY9afwRBaIqNQFzu
A7qAXI74VcTc6uBK2vVnJw==
`protect END_PROTECTED
