`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BMqKhQO7W523Qcs7BrjRSZVzBwI13513aGqWyXyFQjc8No5kGpbdMVn1/98jUoF8
hbL4kNSc3dvAfPN50mijqmkHO1N/W6C02hvW+4QATGhfPieu71a70ufvzkaYA7Rv
zWFJ+b7JS3xf8ghP59o7VoRHSrVmUayf4eZxLWtSW9T0JrKxvM0aplHt/dSjACCP
rYsBkp72XTqwZqBoI8fckoOA+GuWW3MYFgCz1dKP7/xr4Yy1yIQ/l335+VoHqUCd
`protect END_PROTECTED
