`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iXWnpAlVmA66/x+24Z3BpB6xIak3y/ZPE2IubhlSlWbFdsLN64hzdumk/PrktBBx
in2YR7WCS8Ix6y59hOCZy7DNGZQKf9e/rOPxwyEFRrXrP3VizdsdORYp3XY17jLn
YIYoADrA9LR+QGYwhN3whk0cVXvhzjfJDM2X/axf7Ac9g5fNmhU9Mfm2b9r7LP+f
0Vjp5Sb4ClQ5ILzh6mo02V0xVNQJ0w91NV0uZjrVotyT6Z8U9/twamZwR9U3Iufe
vch+S7vp0Beg8/uBUdZ4z4t26sQ9F7GeFceHs2PwjKzAI8OxkYZIDzfyqPqvcnHP
OuY5rKYtbeU+L4v2v3hX76Hcxbtajf1QnuVwsu0dXjCVkaXNREY92Nu7gUkz3eTx
UjJ7Im0SuMSFk1MGPKpgmkVs8GacYV926fGN/H6tH568scbjFHNIkoH80fAqul8x
8Jr9cPG1rjSGRDaOQsV8YaBIO0aVBJp1oBvvoziKXX57qNImlrygxapBe3ixCi29
`protect END_PROTECTED
