`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D6b9adOsRxwdMsAqUqrL5GkTAKVzuwUzPzRvbBCG1U8I13GwyWRHVN76dCCitOvn
FFMzehFpfTPcV5zw8shPqOrUBGC/x8PEodIWp7qjWZZNTvQo85I8aHGUp2p7zQfA
8XSUfj1uW38vqdHVq8F26ZyaMYKpXqqdUNTXR9q7CpheAi2ChbYnKBvVwGRe0YDW
9dASjQ+XG4/j7Ohsz+Y+drg0wgGE25COXViToK0DCd1bB/x4cHk+lQ5lEIYrd04F
UZBALKtUTIzhzG3Nkrmz7l18Z5bmvUHa4Z2AJirgufv+Qq0c4HS8S6CXWEFkcrpB
1LVWi7rNhAtdSNnDZoaImkPUCqDn3O9q+eNXcuZNehPuWks3f9mjXSewnINnbT0f
sMSAQUOnj+ssn+Wqfq1ICSfRZQJRpX3/LSbFQDgCquUhxAkgUt84f7qNK0iGXKcB
tcNlqQVqhaGHxcCL3UP/lO8UM611DlGEVb5KBxRy4KPQj5jbJpfttyhrN96KUEyu
QmVX47sT0lhulAnbZ6xWclMLyzlhIgPQ+CK4am06Xc97Rn/z8REQ4+t10G291tUO
`protect END_PROTECTED
