`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+3yMDWPzjaNalnT08A7ACdmwitK8Nas+PO5jyma7l1gyyqNv9aiv9yFf4nagLIGV
9tWIP5Po7YDkrIJgj1gHlV6QZecrcHH+DAZTsHFHMa/2n74s9X4Yxs9k5jEmXZF8
ipuv0dmoZ3sMhkebptyYyFynqO42oxC8ZcC75m0P11WjaGUkeJpnEXhYn2z89ctw
Yo+xMGknsdcieR0AaiP0kN7RihySDv0+4HLPtnpFxrsWYOemjKrpcjLmaXd7Mw2+
TGadOAkD5OKT9AueSBOzJFqhIg4lwvHptH8F7hZgWfBAEoQlvvAyyGUV/4x2K03N
2soA6l7xfHE8Rdvp3kwkpa9Q0lVAzpt1H3DhzNJFUpAKPBaDABSaz7ldLDzj4bAB
7Tq2XEoG7Eru/d6Se0fDUwEHl+96W/Ntq7lMBFtCgKXPf2ewiGcps0dZHRb7c+rL
hPclx6AmaFkNez4Ljq5qWovxNsVU1xzoAFzlFV1io+lsRCViByLQlsKfho4gul2R
`protect END_PROTECTED
