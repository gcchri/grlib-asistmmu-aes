`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vkj5y+c9lr3qLOhom+qBwNf2/VXkI0SzPPvNBr/QKZeJHdtJxA9q8Luu5MoPtDs1
n+5XDk/OwOiVBQZ15XTHNBTgvx/FuT4282pzRd74cfHfuOq6Qr0KELa5mbM37qEB
H8c9t4IwCDHY2gPB2/z3cjlDivPE2KlS0KTeXIOZsvZRaNuqhitmqmHewLB8ZYLq
+39Ll6lNgzhJuDQUcGY9lsKhr68PP5v+Th4BOlORybSNTjyIpCkYNNXHlEC5yfN7
X88tdVflTDiv7fNwW6BrlSCV0tKHfwfu1R0PYNUhpHcAq4Xz/fxHKc4MeI8dQNgD
O5Ojz+iK7i8MVNygIn5fGevf4THn+d8x3mcJ6PsUVomh8jPnzltsOn9U6yWzMKQf
4zyOqksxiCRkxRIA60PNIR7NJSInxLiBMK7XI6SDCaGB8yIlrdYJ2fAQK/crJfNV
D6XLz4GFyJZ6Am/PvSP8kfv5wr2X6HF6G1mJAPnA2kgEvhcySfBU9VnWS8mKqD45
qOWKSXGCfbndtXf5/x7baL/LGpSLOsi8AH44qUWW1wuyLL+yL4ppoalGGXmeuSbZ
NdI/g7h146h7fXEaEp+PoT1i7P1gw5CxtW2sv/ROqdgndLYLvkCDs46d52k72O+A
NiJy6v0YbYfOu0u1KZwP7HU8shnacPHvwuIL1Mhmqu4INd2xaJybr/tIhO3ojJHb
9b30Yxt5a9ULB2OeW7lyJRX8yhSNkDXJvfpRnSWpDF3vD3jbqSE2DS/GXhZpXJfu
L5UnJUpvX8WR/60E30hmO3F/oTZ+rNJYA21wjyiaiO/IQCalErp7esAZPCFpnX3f
q1jWGDJfDqI/QAkk2aJEM2d5wNtnKUc/F/R7ZJJwBzwADE7oZ+pxoC/kzglACDPr
e6/aP6aOj5eVgtBJ25dpCBstitywOBJeY5ENmqauKfb9mZFgbuOC5fZR8ceVJqaW
znFFNAB8yW3JqLTBDX9ZEw+zNFmVu8zcgnErxeFJsIxTJLiSqo4o/KzQ6sKIW5ab
0C01x5vGaCkB3Zab5bpwnMjGIJ4KNWRSUWZihtolLjyVImHaUOYm0lHwuqiTXrSg
ZoUSQQotPxsIv9roqqeh13qYYP4htN6vu097WuYKxkyYZjMHCRPkFxtZR/wkF/9r
x0A0OFlHlUEyUjfJB7i319n3osfI3QYi/4LPtlTCkYr9+uPdhe1p2onMa7wuhpuP
UBiqnFLbBywMyVWH5uGe3E1ghBaD1wmxgXT46C2j+1mtLG8pXQ1sRLcICYrXh2Ks
VkrVPuVPUHerrYVrmIAV/DMvOXKeWsBwhnH0xyaup4S84fj4odWs4CZjvOgm8vdT
A/rVRdMlXvWwKURXB156bv1+w1kMaAMZMHMPXU1LYbhyLJSZRqmKCwe+qVwJ3H9O
7yvvjK58pkpk0dQvZ0EYpPpkzT3V7JZP1+CCJ5DWc7+sR6wiQPj3oDgf5edr+k5T
GNXp2qs6t9ZymtvjB8Mum2+6UCkqMV37AOHvY/xRC0CuYWRi/f9mqweu/E1QMyrM
tUJV6ui4a0ZVgUjeIewiekAO2PKZczX7TIxzdyLbchSzCJd7Z1539pkVhGcBxAhL
5eilrX985GfFeD9QAKrkh9MpD9FCsVYVQvnUZlmz5ma4hPhSQOC7zGgjJ4A4ahEf
tn8T9J4Dftlo9IN4tZItzO4VSRadS0hABquZjxGGban74rJE16Diw/cZajEk+Xs3
O1PRx1+0sMy1QQ0dy7ATAYn09cIM5PeOX68sulaDSO3lJa2TtI8D61gCs8En/leW
aVOt4Nmwg9AsLg1/KZ/ZPPzlxFN4J3S4MzPFRQjwnjV9fBHS+EjCvx03dcWEfKFj
UXPwYbwEusvYPzieuRhl8QzSLwZWoucdz8wblQkm6w3Pm7ej+inRZ39L9sLP9Efq
WNWVo7PpAcOBOy1ldtGp7VuUPEqQLv5nVN3Qq1SvJplS0b12EJ95kZCc2KonYhSX
CY4Nv1mQ9xettj3+NgLJHBRpAwqgHAc+/weHwJpC2L4+yrwbgG4VEHkcDbo2/IE+
DFeoaMBDZ+fPC8m2LzMhrI9PM6uSr0/VveFGP2opwXHvZQzKSp4PFbo7WG2ttGHw
EbzKNx/2GlJ7gb6Oj/2FpEBepDIdYcnBbN44wYzaHewr2HGaGcL3QJ7QHBHMbZbs
WBpTmIqlIySthid+m3Jy9hCV7jX7qfAsIfWjl92eu0mK+m83MpRtxgz05V/mj/DZ
PjfDZ6LsCSld5t4Hbfb/1I3iacT+LKR2bPIZ6TcotUNQY9CdLpAT6yoomy+T7JdU
cu3+WAmPmbp+Y495ciQBG4EELfffWM+bXNTLuPO86Rm7lBqjVi+CFbx1JqM6qvJ2
dm5Hzf0QepxnnMsIfFBX/f0JqPwYhc3znfQb8xy2cAqg9qRt+8bFLvJM9GaVtTYV
AiQ48FyJ5+DQZ2n/E1c4w/w6wCXXX+n/TQ+nSDTrU5hnIudTuOJmJYcuL32JSSh3
ZoeqQuYDHyFjVFUU+8FSqwnavh0+OXt2+zwqfmAv2KJl9i1eIvzqB00GKCsGGDyF
YJTAYpGe8+yDMbbhtJi1ywN8XmgEl3cv7LVgT/vaMRr9ZWgMNcjY2DcnczVyP3zW
aWYSZ78gTno84k5fxY9GqfaYbaD1VL0dW+QYM58sY87lqAyFIawD2lBkjm+73R3a
35PFesEE2RRB2SEb/s8kzucgIeY/Ypu/INWtn1rwIuHHtcbcPoJn7Uqn5rrCzDgT
E2y+L2/gVUGCe16Kbr82czySkj3qQh/SKpDlbVU/rBGkog8OsyqDjT8ip6OcI+EA
Sn/oWxonD0d1K3GDzzl0be4tQ4ntnDE8QsMSzsjVbMrkGmyNNlsl4cnq2nVxSFfM
kITEGYAjc+3O8mQZAzGKGOO3hlBwDIvOxjV6c/qORfDHXeTSp4qN4Nz2cWoVoEDe
7uliJMIoDi/8sabzmRMiuwSmiW/K9mMLwFV7/PWfp0c9N54mS/6lTmPTFfFU+Dxu
4inRAtRkvWXACYgOpvxfdOs056m0vHcUqZKAo1JB1eXqpvC2zhn6I7bIK2MOCA4j
zF73Xi+M65q3XFiWh24xhx17TaDhhuFtlH52PjgRCZUEPRzARis1nkecQBgTSCAu
W3Z2uyA2eSFL2/0boYIBw3Woo+FhF9V2P+Ie5oLM5ucydYR3NRbvt4eoxw4XMPXv
F9Xz0mf82XrAsk7Y8q0AGeKXzgLTR9pXx5XkfhhiLFxN0Z186alnTF7D0M7OmLHG
xvEXbrwkCC+Kh1o8hvxTWqQ8fpSdlYRymHJzMB9PV5RHvsXA8ynFUYb2DjdgKIiR
Ov5Zp0lNfl6vqLxE55UBGF8m8FT90Ya6w8DkcILjUM01qWesZfSENJ8mL/3j279y
bWUNyZuUuTbs1LPV4WH+oGM6szWGx8KMMfyMpyNw+1M/5HLuVMCX5XM1UiiX0/MS
9aNdpb3RwwQlIS7HeFlH8VxkA2iWMRxYzRajd3xg4wEB22HLHEBSxwBoU66KnnPJ
R+mLJ22fBa4Lvz6FJBBj6Q3YwHcoP6+bOas2CqlIDYl59KQYGY0u3GozXe36fXsj
ayPBbeyGGpg7WansvdV3cqaVdgnsRX3m1P1p0mMoF1V94jG1kwOGs+fqQMAyDyqh
abqJkYy3ag/J1g/nBKJZHOLbDIPfiDRxT7Z86hSlfDjofoSl6v/hlZ/77nTnyMse
vDsivHf5CsRcnbPa8Ahh2AC/SURz7vUIfvLSH7/QR/nlTKo7xettgy2I0NnIPwwQ
JkuyzjVmxnfzOzN5s73pBaT4RzlfXAZKDuRnbMyWD8O4LTcuqo9wVFS+0R/fq6ON
Sjpo95DzTCFvsmWHPf+WGWRn0GkIbvNCV/44TWyvw8n4FeEuTFoI8sclQD2ywus6
Kht7RVjD6BiPnhBuDBizB2NuG+fTPjFNyqIupYgMUVa/fQPaM9jkMz8jufCLCsWm
/7dfNdmyZnYG9GndpQJPGXoDkKaxGlRYBbVet6lcktUQM2Lixn569Uyn3NoG1ZeF
vRlaln5ND9eLq6ugiN/BCXz6yYwt3hUziZUr0jzmEbTq7BMatLbaJU87hrSl9B0H
UBubr+p5V3noim0wBvqS9WXD0iNrmPM4qLPz/paVwicx5owknO8qHbdtFlwi4PU/
w6Yt0l8q0y46ZxhAwC1ReywZJeNBZM1xw/1jLoIzdYFFQkATDdEfHbTMB2kQjW7X
cE7glJ9nxwSHVghPGtx2nMwwYcBmwJKk2lA5pWI2d3d5uH0hyStna+tYhi4O+HQF
s5xUwpf27B5s2WaO+HneQwDtU2sLmYQ+JpODG81z1DmFscGTaY48iM68N1u19efB
HTbC52zjeFdunQZlv8M9wdfSLY/qnlXBt5Hl9QUpXUAW5gQP9eo5zyNJMcjH9C39
bOTiMxcI+uK32nB4STU4E7UDfECbNvE/BCy1PWAbVxdU8UHdw/YiUG3KUIp7T11Q
hAH7zBMzOjmHT1YoROz3FeUfasa8fFAQC3g7dY5kwCsoqjaiqFTmYa6wBvrL6b++
Otdw8DxmZVwLngCfydIEfb3GCdVT4q4xaD7uw4ZkLAqCH47AiZX8DvCbd52MPq9K
SNSMm9P7qayc9+1xiRFoLZA+WqVeICTREKbyuNPQwRcH+NsHlpRpdt8QiLAQ523j
+rOPhuKo+U4Vrc97Veoa3fMkyk8J1LxKnn8EaQk1JmpnIhwfYUGSH1WglxWhj74j
sxH/rOo0qt/qCyuNRoel0+RlkmO02S8aODAZwALn8EcVwZpdUeOdsIsI1QA4mR7A
Y1sxjADH6SKEMzWRoY92V+XZzxDbdRmxEahMSeUx7tqI3yOMOU2PO8JNtbgfRUOF
+0CslGEzHzrQ0Hv9q9wjSIfu825uOpxN8es4mgLk6oBy2vSBKbzTNOx678CMgYCY
VZFHfBCuM6VPp9EXm6KQ8BrcZqCGmhvgeQ+cIBelWGI1tQAYDPl6fqcpTRL62C7l
A3F0W9WtHO5REJHoFRVzrR7ok4X+6q435MtEZ678J2w9QlC3rVwIrHG7DfX7PVIM
O6YLwil3niqtVBPKYYBzClHLYSFF7ES+xbLiT3wzxTe8/JZQTPSI+O95nPCvWYMG
oqdNkDElgkjAwehtamEopqvijKLVekLbn24laKc0wESaOU7miE/okCCrLZd146Vw
uM1Fa7FQxijt2VtIovCTMt4fo3nISVGwZGkqykVMj5pvucPqN0BM6lJAb9VGOlLH
wSwPAXTPnpXjJwq8jwiCGwuVU7UcrTeoXO0URlwpoodUOkXUpSigvQTGLPY3xW4r
70Dw8w1bIyfDXfwvu1LrXHRVxkYPj+o4pN68zUWhphK99tuyUvn2xrCoo0+Jxsx6
3y4IoURhP2DPtZMCJDaNgGHC9BvX9NdJzoiFmaLynWMRMVCKp1qR3uGivMyEi5Dc
9GJ90vAdmVzsHx1bX3QVHltw3ImKoS0aOUJSQzkuBAqw9QpVP+dhpCayjqbBg/mx
ASBixG0a8GCuEqI/gGZnSN+kEOxL66A7tx4zgvd54iqgmHOzP3ZGX6JhFHQD9CCT
BryYGw6XG4c/tE02slJ1bU3QU1uGDjc/aT2zlBs7oQz8RYD7qv5JxX9tDVlLqvxs
Y3596p6HLwsDT2IFBRw/Sd95Y8hfL3ozS4rC+3OUm2TbMFdJqCBDoHz61jRI4Psg
F7E8y06Y6PyxBx4OBWB4WdoNGMborqOE4imliSvN4E4R7qJ7C4q9TbtnM3tUZdKz
Y0K2Ka4nEOh4gA7STziamZMTwlGZhAw04myQH0Wk/6sK8i2LwkHMwcQ4fi7Yctaj
ZBvx6jP8UxNZzrU8fvVeudhh0FPM1PuscP0QXL6///sB/hcPp4qwd1qZNwQnMlqS
F0rTGcYsRgEDpHzR1kCeo60x6hRJuN6tfINQeDAwT5BFPXlN6Z7QdnIXHuMq1m5A
p9D+btbeOns+GQa4ykvBtyrNZK+j8P8HtEIJkKGIL1Yxs9vBlNuCHh/6Ki34GPSX
/rMfMOp0fj4Lmq+WU0o8BOsaiQy/nalOO0s2+XKNzvNq+QAJalxCmNLj+j4JV1ZT
lTMaEw2j3MrbC9mIuBAJuuqkoUj1uO9TKIUrXcu5Qy4dYX3cosXNcqdMSWQgWWon
ZBvcRW9e1f7VcP/fNqngwoUjK0seBbgFVYJLhdTRf/m/LWzCtpglf+MfNNY3LfOm
7/gN/7m+CQ02DeJS691dWZiq7x8V4Edk0289aAoVQ4E8DkdcC/I4WKOGopUsqn6k
3sbTua6Oh/LtCUtSPukQz92K1PbxMVtTpBvifijyT3yzcJdOZPu1+aytlZgc7w8Y
IK+pwh8OuSpcCF1Un2x3H4UuEFxyT7tCQAqdOb9/WLtF2I3tdYWwSx2VQZj/e/we
/QpPK0mePPugsuB3lkITd1o00inzQu9o/KUDvQd3l+yWSG5WbzyRyK+4JbtUxcMK
9YWNCmJ/QLQWP25D7p8eBeWC6em939aE2UARb5MZwLQ5QuKBlLL4wKG4hn6VsR3l
VgTDWk+RhUq+zf7KKXH4YCkg9eha37vuvdu1b/Ui88PU8BNnCihRxD79SS9/bBdJ
LxL9CcScp7pDDU2DUTHDYeqm3X5/hmQSJiEhzXdsbNc3zKKUVU4gUYdILahklHpW
+dTLJyPwSHQGLOuLxywgog82RDvFRYTm69DRIPnFbwJ+0o3+i3wQeZRpIGiuBjWE
PPf9J3TX88rYS1FccfxJC9hCJNDEGG78bH6oMxIsT6s2mFD2sOyd7Uu4eh353qu4
Hgf898L/j8E9pdtgegsatEG0zqZYqrvrLCTCsFozVjWuG5G8qQpb+00awd9ZMOuN
8ubFVnSRXXJZ/KOfJM54SmSLxDTDu7ze4Nz0u1jW3EHgES8OTcjjOz2OKJIlJBrm
Ec4wTt0JaCT8Y83jP3Ud2KFOnUHDAJA2XSBvAdCPqCc/UYJfz+3EJRzRlq2fCJC1
3Gv+Tks1cifQ3392rTYPHzRKXCi8WjWBHdUFCMyn1GMlqXzO5LVn+nVGE+rZZtoZ
Wml5ryb/5II1pmGPMaHv51S/L/mwXJjyedHleX2J2OtdBP1D7tffktJv3dEubLKZ
t58G81x6CuOcOTZLs0e88a1FAEnX8eEIP8wpf1jYSp+oU6OoOffGMvEhg8o0w99W
JyJRyi9mQYfSdiT8AqpUALkvq6YYsm9HrJWgDRoePfz6KJ+pM/aeWSZMkFBmRGWE
swJxagRT19bNBXJDYhZXDMpnzscRqdjOICzNSNCEqSrK5iYSZR2+OG1AAVx01BQa
MDOgMmOp3368X6y1+OLEKGRvAAdaJegowRxGceDGlKqg9TqjaqDy75UlB5mjgwLG
bimk5Hzz5R+gxoDdB9BbitQgN1n1V5WU8ouvnqmGeZXzOXc5sIh0EkjbD+X2yVlo
jnvFN6fcCbhNjZOaPtLtWJwoOi7eTcsuu5UlLOKlumA5hsCeU/bg6wvYeybn4czo
MFXBnk5MbmxpcUYKtXkkR7wR0ZfjBsFbkMJwQdeJCMHKuuIzy63wcfxCmM7zMH7i
XJ9mg2oh5sfav6jckVGBd4cyKL+tjEwF8JbXlqZ7qpaINReOKdmK9wm7Xn9SzzI0
PoSyEusaVbv8fTaPrMM/MN7oLCnW1Dz3DGIMEaNZ99BvCxMMJRgJbLlBlvr1my1r
K18MBl5xIitkCLP9+5rHNle8Rs3C8XYPEkoTbV3nUGy4/bqhFvnsuXfmerp86QSM
ccHaPxtNnbciTphc+4277VEcMA+IUPdPESSYAnZgubFt3+NRjNXkQMqCQBfxitU+
wscbwQF7xbOpFJSQMAvbz0Wl5teGViR1hbRs7jqU2TjY6xA7fHgjIjZruA0KZtgf
5LbaHTrLLTkbx++iHyOBJllHNJisiJrl6wXPY0wFMTKwTcGwTBpEU+XJxJxmCJcM
cCcfUTitUhTgFtGFGd5DrBe1IOstyubnHG8wAMyvEvjlIqabmalwM4EmI2K0rvYY
EG4E1RfK9ZFu41Mdbj+J6P0z3ncjc/AWC5ONTjqi5OHsN/872Tbt5d1vgpy6P1vR
wXIyk8VqF4h7XusuUxLeh2a6LWE4fAqMUTYBxHJP/Hg4Bt4a8E+XlRE9tlhiz1PH
NQkYKrKNQko1ittlO+tXycYzAjRcjW+6TomOVAGswr5yO0fRcwbV7enTRsIKoz3i
sPVPOXZWN2CsSDXXbgKXFhIxj36pwDHUpGFZs1282PscBQV3bEYg+cFMr+ddVTk+
XDUeq8fj8sDm1W/2ROyu6/LYcY0s2ReMhTS/PHMRl3JNe1WvZxaadYb3KpW+aO86
zSJGaJ5uUlGLsCok3JnSe4Qg/aojjIHaMreMeLuimKmRQzqPQT+AvqI5FOklyGa9
Y/8Sd3QjFEXoC30NHQucBlH0wbnUWIRmUtuFCZnGMP10yu4dixp41X8eLwcQWUiD
SKDvoe803ff+AmyZM8TRn78Vi1b/tyAJrrQXkBkLfjgPVLP7We6bqQFOXpRcddko
8WyT7h5Mg1n/G/jJJVamT7OpNJk+IxGG9Fb0nXndh2aNYcE/lXMFF+a3Lf98gRyj
AOUd04jJXfvzS2DRS1bH3LBC97JZvyxYeWBam4rybcccQEAR2x7PSN46fks/LMrc
EgjaBO878fGp6R9OTdG0zpF218X5gmKFAWYdcLQl+V3EWApcvmlssztzeKVBV0un
+3fyh898gya9d7PRkvNvaNrTN9jlQcUft21I48N8Bt7pt7WkEkSVdmCqdWn2wgQP
JNHXLsewGBfwz+9sVLnridF6d1qWcm6UhRHpU4CyQuUW2/5hHe2ZvHRHGnS9dIkB
riIXpCCbigCSBe6wzd8P7/bjkMJZyYUsTPZT99ayQb7B/GwHki/lHtoepUNXXWz8
EAJeHzR3NkgBp5WQyyq1NfZjJHm7yGoQJqX3HHtnpcPi92Ry7BqB8IhuBkE2+BIF
Pl2WgqjLq0I2ICOOrhXVKzGm94xKbZ05ZJULLekLRQeCkA8hIOwPDwLCXYBephWo
y1Cp2PWCZzhMazxBFtN/jf/tQTHHoG+MzHDmQ9rX48ymjhNH3J4vtPDtRqq6a1E/
b1HlFSUkDdb8Z7/Ja5W44RCHrjDplilxZETUmsPDTeNRn+oMdCN+wIRwWiu/TRoy
OD2NbOluhYeM1UNiSCEP/aVQMruJLbUzYJeF01JrpUFWwGxOa/9v2XRzWEQlpTpV
cI1d0WB999+nxCyyRPdrpei+snXDLAjjkKwyPQ6qmemYRXBl9aUDDGzWkzV0swGh
hf4xCJBuL0mmgyD/XT/FGyC1nJf66MR06LletbtU3pUai3eEAUydTvBtKo7+lwqt
+SwBaDIYCDho4Es+k/El6RHDzRKKbRiFWpJLdKbZW5/OGox9So7QHxlZPwO3uCGD
Dp0a6yNY1CkITbW5F0dbQ1NIP5RGd0UnGEUtHLvZYmkqS/RIPcIuSAMJy1qoZH68
QE1rU4//RWr+AjZkpJY3A18SSZmeILPAOoms1m1kT1uJ3oQWcEwx4EOzAJ4hFlX/
3ksHS/5lfWwKWRwHHVjc1zCRVXPg5iI95wGIK8kXS+r3hc6v6QFwLQFoKbCKrFsI
wUnpZfoDP4c70rZAifGdfO18eRPp+dakdujdbQOB7uh1F51UQjgnWLkAI/6xmI4T
y3iEv+PBw6/b94d/hLZooLn7zWYytUF1Outgp1bLlzgQkRXVfJMHUtmtdV9VriXi
OlwtaE/0Z9zWBHQtP1NloJhixOQN4qomD9ZDufZeoom5fwycEBpDAJfcLvKUIreV
A06Yd+rW28UhxzltTgQRLYbGL08FXBlpXR85Sb62JJMRLkS8oYpKKJ9NA0ixvXFS
c9pmQcly49VAf/TCqpUhgaOzeyUOdrc9dT57Egu9GtLUxoDERgpypjI4IRhozQ2P
YRjSs+fp84g5m9yJFq1vZNk214VYqWF834fX/NfipyWv8tDfTdKE/diaEID2koHV
iXRp/nA/v3dwtFFWb8wLn/h1j/YEWzqUm8pBvPY7lK0Tm//GKyG2r9I72GWHFPM8
IlqXM/gqkEKRQ9MoAt2NyXbJbvS58gqRaqXzZbNOpIxfKBPLceFSQ5dzx7esdK9E
SCNgx4R4YgJDpWS0n5PF0ZSgTxXRarl9eKFLkb0NzN2lZyh7H7FZFMyBLoqxug4t
u+5VQ91COXFhn7Mb7BMwdLQiJ0N1qw74JuiIMWMNLjLGihS94PBerRFX0JF1KhnV
31ZnWf8m2VznlbdTvnyJv6vQZl/WZ9iuGIRcPAfaMroJYzNmkUN8G90T4a0eep46
z0hcwV7doyv9bvdks2aq4xsXikIBdcWVwKebKbB3tBMcBrm8IZ1a90ACLMjLBLYV
Y8icuJXvwaaKNGZ4GYSnlsZhH1CLbP75Dd7Gq3o3fuFsGsmUoA8PYM8ZXNMennCx
ckC1bUYNTxO6O1F0ig35Gb+Gim7IruDPdIa9JUE7i9CebccKYrgVhvt1Zn/3oUxC
tOTr6WkPnSIrgnHyFZXbf10Cz2owN0nnm8TnTEBHCOm6/wJ/TxwHw6LFnCleqvjU
Eqoqg5s4dW0Ha+9SxpTrIdMpBzWVlfrqZAkviPsD9WHzyAUWcwK9Kl7O8NGE6Ei+
aH4i5Oj+to951fEBMnVdfkOOmPi/JL4pD592hV9Z6gQDpn5z/xe2rcPrzrPvMjzI
OP75FLbuWNaTs8OjFrsgSGlm8+QFmidiTRQ8jkEEpShoFQQtc0okmkDBqemCL2xx
q+v+7WSe+mdwg8YsvffzOFZBQzyfuVFOHWydV2dUItudfCLyKOX3WKVUhRDHci6f
2q8leVxqUZNCZXYXQv2mJqASSzvZkVHAtYh4cOce8kkKLlObLjDbeeUUOTMO8O13
gbSAblbBEeNjHs9Bf9VF+sIXO4zfFbGJpdntvL4LRTIpj9vAegQ9x2FTyk8LLDZt
0GUKJRZF3oOgczHRHcuEFaUeCIVqkxhxO/QPuWaCPGJOWjGQb1MK1iLWwNKoPPAI
WK+fCe00aehfrV6mMfpjD59S0cq2n+hH0xZlkViiXOSHaOIqK0zvAEU9leysQxV3
v4OuoFLetvke5Fbal3gBs18xrJSbIiWsDnUYpO44i2H5unzoYLfQD/mCQtebI9Dn
OlerA34RodH91/Pqiu4bhAZ+YrNE/kri2dCmAZJxk87M7kKBcL7z7vUThCmZ0hIj
p50VUkwnncGj6xFLdDfW6HjbxvIQl65znStm7EyxBdZWMlqtEcYVlnRdxxKpEDXt
/iejsPsTr/xm0BDM3OPO7AxSYosdzS5NhNPMc61ZGmOcjHqht3rObLv0O/h7oraA
AGhr1kvobKBwgLMsfPwkdPwdU8Lq3Q7PYZA26CezQR5BMo9sRliSiBEqKanWcLZx
bBhbXrXMRohQFVtSs5sKimcjxhf4wFidT7mh0QxuZSbmb68RkX35R4JATRkL83m0
TEkBfzZNpCEVFW6mtO/g3+j6bj6prVb/L7JmcrVTo9dRjpQgyYlsJ7c78RCnwz4k
K1A5fAkO6bf48PJOQYTuLaGyrn3ZtVWXOKevObhMSA3Gbbn8Zduxfjqzqgh447Q2
5S6zaAzbqTCAy1FPjm3BJWtM8bkVxMR5kaN8xfqjnJFx3nQXMxKeCDr5MbDT9p6t
QVIRjqdTA5tB4tVoUSp5jpxaty5Hl4pjgzksrnBj0IhGZ3XqCkoqniJbWEB8YVgU
6Nct7I9y8INNJxyY3iwK5mhQ5w8WzAtpSdxiAGNzDuIEufeWb+HiTB5bhLs/2hX6
9y9Mp+vJZGP0cKh3r0jxQbitCiB8nq2pbR3xQWYkYGXY+IKj1MH+ImJhKNEE7fdW
2IQgrIVWC8bfjk7ojyiFC8bLWL9DX4S0aaS7B0oeQLetS1gKBll18nOjbBmDY9ME
8N0XDQDAc6sVhVvfyu0hTkfsEQ3AVywNK11MYZgOlzZHS+sX+MvEGGsZvc+y304K
8qgD1u5ec8mVolfrnV8XH7mfd3Qd8Pe64/O+BcwTydfZg48PXgBjgfsW3kezMH2m
w5deqcoef5SnP2xVKjluyGeBE1d6fupUMULfUF1ApQJNhH2zNxecWgREAD4VPjcW
bWjlboDz5yZDqdjmhWWIum6izcZPawzDM3aR0SuTJ4jXUWQAWHWpTA8k5NgRRBbT
8n6tiIaPBInzxTV2kI4xJ4Gxe/njRr4JQZVAc1+9o8ajclnp4egp8StNLLqxFD04
TsiyquB8RuWYl3JvjwXJ04WFhpNGJt4sE2ASc+Yg8bUy7cqZw/rKMMeYNBl6mutp
HYsHyEF7GVfOf+V8xoPiwwpcq3EgPxVkPqmqCS3c5tLr4WlIP004QfajOokqr8nV
mp8lYAq4J1JduV+IA7cXR9IUz80bEme8/2UOQ6QGVK7e1NXs79veTUgjoLfQi5cO
kPfJXsOhA3yl6cREbP5eRNQ6TdplNQyKj+IYdI5sO7B/9iZ/j0KRs8JGLSp47fdq
DGrtwRnxh8Cb/VOid5B2uz2D/5UrlSxxOut6BQayo14lVO2xEwSQZJNmxjjbONzZ
YHzHouHniakyDgrM5nGepzTYszd13x+v5K256FV4of/sF4DCHsu/ea0Gus2aUY70
zERTRkBKLzsskQVtv81IJRpLPKtIJ6sXEGMBmXxF6uGQ8QPgHp03RmepB8gqEtqO
SDSJ4Buj9gNS+t+EhNQLZ6NcCAXodY66WCtIfb6WMi/jPWZNoaJCJgr+tJnTnFET
dPd4DloER90u4ejFeSY4PK3nzeyctSScrTGzYOVlTFNCzc0XHcMW5C5HnbK/fq6F
FwQAuFfa2pWOSuvOJbaIG79yqTVVxqXvSxHPRrMB4zW72SPfQFAkjwp4G5kEo7RN
uQ3pVAZ4DbmHVUhZM3TGa0afhooSqKIzJ9hgLqQx+dfyZo2sE2g0TnlvRyg7n3lD
nEx8iGIr4blqLoq3RNTseM9ycKZbio1Vri8LzRmwIJIbN2H1wdtytSXxkZzbZ+jo
rEVUVTN5+XAONpuTXPy1GvP3WUf6r/Rw+vg5ArBWTnJUP+XygoLqKsnWtHZRAUtP
S0vWy1gy3zn5dR/xvadOiJCwjCGE9xvsORmY8wJBeaHfhAyQ0zDnOK3dypOdibUQ
x8AeMxrhALwJmZX7WxF05V8FxnuBljaxrjUNk8+wpVdlx5ureNaHTdG0t7wrcLd0
AbNcezKBFqknXYbOQJcjvDvrdp0WbmWTyIlhAyTzRuIBUsohKXS9EJ+TY5jUke5O
yY2dzLO/W95xmUckvIK5XYk1VtDFiDYU0dlZ0ojg584PjNBYza06RP11G8jV1Cug
cpH2fd0gQOBoxFrn6vyZHs/PiLAhYn+yCKTcpZH357NaVT6LWLl6UQ7+T6ZYRves
0W5VLu5xpGDxhzLlvuF5UQ1vHicWbh13n9ztOZsnWsjQi+fFt/Ivm8Y34rbZRsFX
wF1GmAseldVLsGjdq//YLUt7O8DbYp15NX9s5yAmzrOHryB6VWzzT+iGW3H8pefH
fSjJurpo+QiwlWB81RAfDlSN5FQTZO7CIaxiYMvljAnu40InBM1SLa54Rm7S6G0Y
aRzV7pD6XNswR2BpOK6nIVTLjd3Mzp8qF6cJ3J/n8QScM54DkoaV8d5RLEtTnpLQ
xdolvxvyRC0dnfRkqASfyTz2/Vsr7HHiOlauiOWAn4OLeLAXh5LZR9CtWEVuSrkv
rmCfzHbw+fISeIWIODlZB0unVUGV386oYQ9APuS9N/OSLtZTPUtN0IBn1J7PKCU9
TL8TIt6frI1rrsko8cycTIKfMX3RW0R1rn8R4uZ36V1LQRY6tSbgXidfUUFuoDMD
SFlBFOx12WIk4QjU8/BZ8Ej5AKWy1DMU14CR/VVyn5xpc0r41R968+a5Y4cpn7C2
5Qc5a3EBsWHlFX+xKV2wj07wjnMtnqqQBZiSHp4BpC2SgchFAednbAr+QVC7ODHf
zELO8DMtfDmIObeCcC9rfY8UGyI2+6Am9LLswi5kytHnrUwc2LH9MTrLo153wAx4
ov0FRJ/PcL8W4Gulbn77fRA0cwiEKnXMDTl6Nb5JO+SrJ+8BsGGlX4lFXOxlzqMF
MUtKD3gAhFzcP9K6G6oH5lHwVM7hiUef2nS9NIPYEgzAlPooicf1kYV7IvUc44iT
vIy85BBTojscKxQvzK2fTMXYNSBtUiFuD6EDiQp60Nr34wwEkz87wtPXqJeOmOj8
4yh4XAcfqf9XM0l0sD7UOpB1ygJhIHkBIUYgu3ybwdK92XnMKHVBzpNiPAC+c7r8
PYD/sQ+tqno92tWTlUCh6/QYFud71hGwiVXI8RXZtWW0T1GJ+FyNqKnrovvgHImw
KEctBmPyBDrzhBKUm821MCeaOkmppqBXsodmOo1qYuPFKgWEW7lx0QeWh8z5LvaG
qIlkWzFNiOmANh9DjIg1JxSSKAo0PEEq1xb0bakagl7vuzqxc3N2g7HfLNZGLG8C
l34rQWFFUKfIMel/MjWnCL69bMxivH6P6jmnSaWAbuDChMWUGkKkIGqbebyUHFW9
5CRR6ojLt1+oOnnqYIT/s4YIF+18QUBJ7iAA5/QJ41IoHcQwriWvZjeviz3LhQV0
Y69vXZgjFcIVpU5SBpz1u21kxfJSFYMw/ddxcoWwXWBTsftL2Ylbg3pY6osm30m0
SPma6V6v5oWFOtlZYK7bb1ZEc+pdWQ5jcpqVIpVnOmOaxJMSnH2rbJIyg7Chcy07
Q2H2p6mK7S8HuHmrd90LjdRhRqz7ty+u4Q7QPG5GvGWmZZ2byDDju+mBDcR7Cnvj
QhjyktRAL1dusjHG0kGIS79rkLZHLQMC5GbZNYavPf5bX0qPKkYdqDqI/iUng1B4
HQazSy2R0IO7DWzuTYatyH2iJO375njVgHIDtxr7Z0j+Kff0g16T9WTRbmACl2R0
ituV5eQ6GQuwdSTuPEWSvhoRx2TZ0f5viu8Envj4JyzBW62bvd6Na/lCKex+lQYe
smAnowMxG3zgXP0MLDOJPBmJAulmYDPOeijpPi4N7B0PcyrJr/FB3qi1ZzubnRR+
ITNZhHfiScIAOrktZSsrFCaG4QlO2ePsgJ96AkQ3Sf5l5HQD3euAuWPNtXvufhaZ
vf2Pp8/HbPCz/Sj02B3pp1Rk6EUq8a1GhcQ7baLo4WB82QnGplfAQmbmo6+6yMIt
O7NYgsonpdlitJ7zEisC4g1MRNims6kMJuoC59lmo79JagYNINo/OVFq/DUezAye
FvSMKB5976D9BO21bHdRkQXW81OwbzrzwQarZOOk6/bXCA3A/09OgrJdzATzDxUc
2GI0CZY+hRzU7rLBNFIs508CR36BSz0FZEDERCsWLZJwmzHJM+aanIaatLmSmc3c
MSbetrq8GZTsKG/+Q7XQqY39B+RpEuQ6HvvhfHP7KeJTpd2FKj5xi3+1YUe/MTFc
Z1zMrLTBDyrbB+LjjwHaKNbvaMuGBuVuDqbNb4/57ZBBR/X3PsNNmEq6sAweki66
9oxXLSy0UlMAtBRDdl0J87IR6HhZvSwi8aVQeton+JFOze28+KKyq2uR+zaZSzGI
kQrIbkG6mbidA5r8QjMFnb7v5d2PH/WXvwXgDCMHz00HFy6mQnwh4T1ALpxFjzpt
YKmCif8lU1Lk/OKtxsUYxrOTZmpMFW4/ct/medTkeUnDP/+cUfTjRNqr84WJPLGQ
2BK2BxpnG3myxANDMKJq6C5XsZxuL+JBb5wd3hGMI59cqkgFOYU3Ec9ypcAqBwpV
zKyfwMDBL8dzRXzjYps10psPkw0fa6m5Brx7kxiR4DQwro0X5HXdy6gxT7L1yXK7
A287ezitDZ5hOA5/FHNOBiaAdM0N1Ld3wpX5Ws+6Jm4201xB4/umDt8MjV967PZS
sYS4U+XdJM0kl/WATMfa+EHMe32CjMRwGyJ6UB3VTx5HDIzJjED90wOtvAfH11Eb
I20YieItpKeLB2SB5bfXRfhhWji0Daqvq+OHGQ482Gfzi4XK7fX5trNQ4faxv9LF
b5F6shK9ve2PgggnrtnnO3gVB4/poyjG1mZMPNmpJrLQhzdKO5TTeO8T3nrKTB/P
OVz+9IvkAGBhIieBlyNpS8npUmCpGzL7NXN1XmUQwlzctLe72kGWw0xTg14qywcI
dETXiLfS0wIm1gBT83dq7/0/Nn27ELap571MrzTnelnMnCa/Ilut7IT0HOqTyfXQ
MTcKztbhWjqS4d98D/FcH5/tjmyRfrEhaLilUeC7z9E2T0cytFuZHuWLX4ZmRZpJ
HZjN/vbQ/8PnL7QBE+/mdhlNI7/0cS7ehdHAml7rz9kOybtl0I1GrAnNl0OKlgze
hrPZLY2r3YxZAzy1GqlpCCRDYThkavnGUHRRqJoPAZ8Ia9WAiS1WT2mMjV8TcxNY
3xm3HQ/75ASuuehpNGixYf6jJOAYI+ByxxAuQQ/iWE4nyzCLpRLfXxb7Mqf/PIah
VFBGeHGdrAXDa8s4wbqmfovG6qkZ2mpsK9KY7jmZrOOqN9ZlEFsH1sqHM5+Kwjls
NYn4xbgfU2BBx011sMQ9QZrUzUcpqdB6ABjbLgM5BnnVEu9ZkPVchAFS1VE3WtWt
aMnESW0yA8lL9onJtA1i4zmbh03F/++ERIHpw1ov8ZWiqxMgpqW2YjWYJqwm5qOV
ukEBv8Du6bceSyPeAauvIvEvyOUIHTJlG3WoOhGoOVL5NE7T/oYOqStx98XwG2vE
GS6hYgqCrKqJSoAmXvpnaKC7Ld7SGOeAoWK6+TYQLinI8cgyypYkGkVcoCU20IVM
gFVhA5zQ6eChnwtnNBGRV3s1y7QIacwjcQrbFDAk/jAaWuLR49Xz8bip9tJH1CRw
6H9KDUMY0pDaGyw1WeK+8KzZ9//JkTx0p9Dvwt0CpnaZkaI31ZQKelhXSFKzicNP
bRJ/PjfscsTzKFFBs5SD/h0GLnzaRywDJ683nJ7P8NiyVNTkVBio+oPXhWFhLn3M
++Jxk1jWmv+a7ILWo+3m0J4eSG4CIFmCFtaSUulywzDyX4qnGKuhI4JQqk/ab/No
KN2YMg8keCLSD9gKngccwh3XlJi3/UY5gFFh0Vl+2q7BjDjZ70wjYTL/Bk0FB6N7
i6fAJW8mUqB5q67LEDHR8jMwxmFC0/xZgfNijyBgeYyBcLRa1tVdZdo7ZFILE90h
tnVzrRl5CuTNVjl93FMAjCN/FE8fy28sVBVtMEeSuZ0tg2RS3uXV3RuypNQlQbB+
QOfut/M0Ci70WiBsaOx0dEfJUDHFrQ6+/taj/yoT2kueguCLw9ld/adSlFtzlB17
1phl0+14LHFAwvUHFLQ4ZnacsmsWnaoL16g0Drsos6hxHdX0d0jLVkM0mC1DTN6T
b9IbkFUGldHM29mEmNOPHn6sjVXJJcfoM9xKe+0/R9YS7rSmyFX2WX1OHpS7at7Z
k6oryAig+nKCdnJYfjje74pj2Flw4rcaQj75lDYxiTrIjfqdjvxK2G1XTHPLxN93
PWTwbXp6/lMU7J/IZrrc4cF3LCNsh0CyN5OGhDCAz/XBG8ySyITX677MhFQjmfec
COITxzBm+xY6oAC3MocAaZ7FxE8U2N2pLIguTtYiF2wWLgA7idtbc6EvzhI8fpDI
T5u5Y7f9i4NVlIS2pg5IDfZuV13mczh+sLcvkbnJRanw1+B+7sGc5WGDcgDFzDNs
O4mIZDjOOzEU5gua7QPbjtKE+9dGbkRdBtNjoshN+IuqBSJunSPFq0OZCi3uBCW8
56DatD8YkV6v6YEud+gyr6ItgLKCaRs0Jep6N+CwH/shs8DcrC9r/VPVbWf1lqtS
T8jvK2FuFvfCVDggwOcm+xk5OI0Px0ahZBeHJ1tzU/cnJ7GkuNHLbz4qNyL3pcgG
LXp0mbmriZuDoT3Y9gVObq9lhXB9HbIYC096hxPKMfH6W7ix9J6Pp856Vl/M9zNr
DMc7UCS+Rkxv8At72vJv/A3cSN2GX3ycgdkBjovwWty0sfDC0VApWlkSzMvpkO6E
fWWD32YJd0X+QrIPWRTxwQUvbLdRLfdUIUkNLtOBd5XB65w9hITxW7CKGVdTSOtJ
51a2Zmrm+LqAplQ47EMhL2FgOdbTMtmJtuWAse4VQHTDQ5I9c9akwRNffvxK/6u+
a62zpx62AF+Z5CdFpZfHFl2SFrny9cPeZtwKi3YQbxzpLXKmNAQW02MF1LMEYd2/
hWFdrxI9JQEp1iOnKi704GaDshHivS2TwKwUVQEfPx4x/pbMpgDLBfcc+HYY1SoV
+JQ5nJdkXhJaK01JaO88QVRPwl4lOg84cNTpTbLGdJB+lPSEPTzutejse9w8bk7H
jIFyrcRJ+8Y7md5HUYcDyb8cg3+jHHEpqoD5yTxMFuBmxaURnFClHu5LsxrzdIZ3
XgrCVAowFHsWC1KPJLlHEPbI3U5DU26oYB6UE9cCgnlPeE7Ucwa/gc+MxEH6C09X
3bc8yj/elgDw8ouZgtMzUaXZxt98krW8Jn/yiDQK35Qc7baRmLbJrC3KjhMK3Wgt
yE4mZcG26WVrgVUSNR4xWG4MX8U1RsWYfeXELHrKsTriyJKzS3gccMgTVtrTzIrc
TwmzOYC6CybL0wuYxfsFVjV0IJczIDVJbrQAkSPTSM+L9B4b1BO/hcuKTuLpdvqr
tM2vT62W0ghlPVuLyc9qRkFqelb27gmbDI/cJupEsYxMZLJBRPMCiR0UMp0ppRfR
lGeUryRbChl6ZtLdNPzUi8++TJuB9ZRGLbIWY8jSNs5z8YRRFuMtbgk3i61zGbCK
62o6YOsiWdWIApejVafsZfzoonecWKTbxTMuQ5pvSUZxQsYbH2burPdYrxSoKPPY
kKtTHuAZw027iG1fmVM0kkDP3wqklYMY74NncBxfmPf+nYouV4SPofBTmA+ArdGI
C/9OK4xzjzyHXJsk/qsP25IRSeMRQ4d2Ndi9eQ9PX2pT4wLbZVm37APBTRcok/wi
nKxITK9CmnI1XwIKsGSSMwzvb2svu5333eSX+rJFMefrV/og5898Q20GPk4cmChe
+kkosqQfsFjKEVv8gXgBK3OAAn0PuuXUS0OoAmTELxY2NLaFG69vDmuWFix8d9Vr
S+2rA+HpTsvv6ZFqg7vjVXLQrfKIObQ6aqWkKZoHcjj415dgrJl6+4Icf93NGQ3j
fKajGLcgdRKhOymgHincEos2EHU/8H5lDdCB+u7c/3QeNXC4Op3qAUxuO117ffZq
cU9hT8Lq/KDs18ZZ2qW5jKMCGGYLweFIXYEBpufIAKGPzGoFaNfHhQTcDXT6yJ29
0Re6SBZTHJ9CSOSXqyIe6eEOcmtqpx18tVrVZOZLggUGH1tivBFLS4OCy3cicQV+
ly5P4QJnKSxrgNOxDTLPQCISOhZy4kmhIHMHPFKZbX0iv08rDVBwlBGXBa0WGXTk
aWgJFCjzFY3ODsN/ZaE+IrUWm6fY2XZtjgHyoFiLtXZbrk2Ocb1BKpWUKX03ZByC
Ru41kySjn/Foqkd33iOVlrYTwNMf9UtW/W6YC6ou+akEvtLPgOPom/LwqGesgYTz
FtScMJYSFqENuJu1g9VJT+d+I7ZQwgkIalwGT1lfYqD6GMyieus38Kjg3MQ0eDkJ
axDbt7Bus5sd1yISws/9mupL8vxFtVVvLT01wAKQP5JNINWstOWl/giEl9XQr2mG
vODADcxOjHWSs7DGAw30RARlB98GLbyAYq7eobCHiSMdQi6tj2jp+LwBxdIJy437
gmt8HizK92i031NNgbsoB1/QwxuS4nvLDM+zMcenVmyY9Ox0clpUVbrvYq59IU1c
fNIWGEMXnKhvw8aWQqvqD2QW/rRCyQG5Xb1qM5HVhS868MVAd7Df8Nn8Dn37bV1h
sljN17SmWhgVcLb0JgbeGBXpCNSv418mXdwcxIEq6xSNnqZLk01fOKQl3zNNmAMZ
tPr7eJk1+5y1Ob49/jip4Z7XsFqrLpBlaZgDkPotTJ2Pz8FS6zAIfpwWHGWcFAlf
5FexpCBCkGlVibsafodiGj1WHPMiuXbEyRHtz3OI9Cu2+X/oWmdHBYlTjyI34OC5
Zz1DVLaxpXqqUuFz+8MHNRWKc4QhPbOhjgdVGav5AoMw8QnyL9yf+wng9d2oxkJ3
BIYDyPPTS+LbwNHVsNs/vnExOiyWxruDT7lqp8LCnmeEvxZwxutyDN5HN0Jfrodv
gXKlu/rBDm0oWtRL4FtQwOTxpgv9Hd30lRE5HJTYkBVo2dHTt4XRgkVdk12UyreI
klRVW/24akqtJoMPxqOUYX++3Nfub4NT2GzvMffHJb3pQ9K+U3tnYSCpIf9Vsuqk
sSp+RXuUtu4IcHVQFZZBM2uMl3c0KFas0X1ij+8zjO/+03gmFtQcuDWnD6eJ1r5C
8Cyrl4OPo6n7ToQmlyGa9tkWTTx8AiwQCXw6/2n6jWxZyt3Z0KGLS69LdtfGqLIt
fVrl6QoDUF7n3dEa5w2/WtVQ9rp5XO6+bsQ7f5N/N5B2G+UvICGgML/BEXHRazCv
WIxRsSkZM8dirlZ20AM1IjPXi7b5BSNY58F/8d26nxdrtXT8vDY2qAg6kZ4tmqq9
zbqZA2voSaQvjJ04XmnPu0aLz82WcIrgQHniYsoCseqh8Q57Pf3+mx942VD/bgoF
2sxI5YJV496eU03dkYZeSIiVMe3JY6r2cEWHej1NFSfHVXRngy4l0bUlneLR1XWB
hZQGGnT3CHO6l5BfIMqmBUX99xCh8+MizlTz9SrY3AzGpC/9vUJQCJe6cDw6MoMx
GXHeiTQpkq1CB1kPBG0N+XrLj+swkP8fExI//FkX4J+RNWvmzCauUs3n96pSNAKg
eh2WFASjWb0C4Auh5O1jvW3hYudt/RSziT02DT6OtjhE7eVaoAhsjBFTecyYXNsn
WpTUXULdfWHD6HJmcgnyiVdYCwVoFrcNtL+Id1pmDoqtb/2N7bJlECL5hZbrVmDb
bKKzXm6D5ntG1+oQqO15VC5AYkYCUyiyK+/S1yWHG4DIrTOibnvZBToveaz9xf6y
yjkyeh9Rr9JcKuGSbfG4m6CHP1XEe75QTiwB7z+9suav529Z/+l1WtG2tJv+cdcg
cOzA22SpvRybp1JsPYczRA94xtUgFu44geupYXPD4bI/6SfNxoVeAFphGkCVmmnL
hL7ddimklQsNZVFUQryLkgmbzrHmh0jl5ADEcGBhO27Kd36CtjpYE5+SX5YrIMaf
dW8WOkNf+Zh0RHWldZu4BYnzq+j4joGAvDlHL9DNFgFk1cSE18VV4Y0/ZvxxhrCb
+ZM9DgMJmCzPshG8Bt5qXLoztijMrjzDKd4AOGo2PjRN4ISqu/hLyJNOu4Q4oRPD
2+uXoI9a3ejldn20al9vgEsy1e8xTdhStY6YDq2YRClxhfQEL1YBCL5C56wgXqGU
LjArjIRWRJpESN/8sPnzdeC5sPvnZSBtVENQxabB1G6aooH8Ba5lKYcHHx7jNqtc
1soFFm+VtBzq6dSZBL+kgdilgheTPmFzE26sWNYyyk7KSw1FH9hGLXLnWl8UCKtL
AifsRonGaeKeywpIP+9DbjFW5D/Ls4k0kJdtMk2liED+i1LR4Lnz1WPVxGppVvSF
89SZ2xIXU/ygAOgkptAFJa4ypLrSWbPrEhv2jIp7L8GMdxrfl+u4XnM6ZSvVgJbs
MzkmSwNP54zh5DdZbFBwIl4kb7K9gdAFrF8W0DuT67ZFm6uFmaBvt93+FWyoZr8B
6ePjtDDTEH5qH1uef4/aItJiGcDHjIeDCkdornspKLW6pTIid7uTH/dvRpWM3sgz
sAeRv4SspeuuKYYPe6hrR9Sfj6yUwYDMosUA7Kul1eR110ys48OWOWKdNUtOaWsI
KPqVLIlbUpiYEofw+MeqvuloIQUxpC84x+Fc/cU7Of3JPszZUMW2snAlkrnuomRS
zGEwIJ7lzSuXd+TG/iDUDQQQxttyAEec4wMSBVXWvVdu8fikvBoCezCjqDdvvcNn
XUWWXBFLyDUpoXqD6GRLTEL3syMQjbqQRqrrXIYdb/3cn+3DmkfI/dcNCLGcUtbY
mAfS//8c+YSLtktyd+zPOkuR4vONHx6wrYND4x5I9aVxU+Jf3LhgWlvIfvS5R4PZ
/BzLUOGOSz75jH95pwO2KA3x2mJm2U0/s2xO88K13ABmYn+3HfeJUB0DhWEVAIWd
J6o0L0oqt+cYnLc2Op7ECWL8CxJFb5NxSyWaudztL0BomN0yEqweK+oMqOrK/aLK
LcL5zGmKw/mE3HwQhBhw619VsejUH0+Qol2CJrPLD5jjFbAGrEgLpfsGKRQxG4+O
/akBh2wiLmemhynPjyLfjxoHpdD/wisfWXuw6yecNHCdA+sJhIo+Jp7nDGW6dpxG
GbvONy8bR4pLhruVFJlN3W9UXyUmSRCneTJphwVs5iZC2Jutb2E75usBf8lFnoZr
/KWkFe4wQl3bAOi9UXTHNYjh4VhxjsZmKqsKqY53HB4iymMT9oced7nTvAC4kFHW
C8wlcAwZ1B1h/Y44IQgKCBXJLat+YJiUh3wZ/6nTCkSTuGLLA7zhZ5nv4mTr709K
N14//VIh639T2B0NOmSlUlwOxxHEsA3NhjtQcg7uu5wEdR2VBL1PwG9B8eQ72P1E
MWH8jMVR/dt3j3Pd4d2Im8zf51+wH56gdUdRcpcB3Zrj3BkF5KGKlDGuLm1mZOMG
9S58Z24QF3HAUlCeOxQ5zw8POoF1CMvSb5GjiqUKSggrFmvn6CYcWonF3fDl/ceY
tt8NM1ZDSBAVJLUoo89f/VCmixzqy314I81Ecz+Ot5re/MUoz1dESr6vfJGx1Rtl
dgtjxpuqn2t22r/OnMrum2gk5s70OuFEL1saQylXz2fhdUGKHZQ209LKbyVDTyYU
SYuVg9EfIZbW7uKeFUH4DJJ/GtUJFlideRoMp+AnUtJVOYANSVOeczYAS1Iv2w/T
ST2V9+AKiu+rHSI6nTNE1fFEa060qEe2eOWoPMAcWuxyX/Rnauq5GvNwaUY5cCLb
54Hmw6tLwT0t15ccbPXTFRIzKqv289OKboi747UNmOM3r7BFtSHFjXmnG5DgkFfU
hhGp+C9Cdpe4X7ycCBFYjo1nQPIiEsumXLPWpL98OZDQx+wQYqiEKZjnNk990o62
w/wqZrBMRAq3Wo0S7cgd+RgCtxzxeVLeJIk11SMILYrmjOd7KtoHw+Zy4LzZ7Dhv
zLF8owAuJlc7kzlLv/v5J4YFFIQR5HNqyqFBkOapceKwX3s+2LalvEXwZUjVSrjy
6mFBxUtTe3j+v5JVxa1ENm/+3psZeMgJ8eGSE1kfIgPe3GM23x0n4BBQPsSdstzj
bVkpDzRP6TMjdpnasPL1niCwYkxBgNfVfp4ZvmHgbEO6pL8OjtE6fJ3GKa+QY2Dd
6Hwlc4z3n5I/St92geB9jvbz63CDIJmWOpa/WqR4+AVsgIu3uXUNKrDNi9dMWhAo
1KVQWNB2nbzuwCHCgmvntaQlLcIDt3jTrVAjiPmb22UWpBBrUnGB+jgZ9bO2Lc9s
dWAMf9FDeW0e5rka6eeQfkpSF3P7QplprEgzHctLGb69VMMPNn0Fq0Wps5JvJ59T
PJh4F2WwE+RpF/bwOZvVAbEKf20MxY/EE2gbKHA/nOg5FVw3ICzwn1CITyeNdFU8
wz8uiwWz1t6YmcM9xLSWMZwiPbaqxnUUjli/2UwazKIa90ybJQmaMUjCu63VsYT2
Z5eUHAfBvSwn3vtaUu9tG5n6AP7YF/FyKf2DWsfD2mnAufxjb29DPyp6K1nd2cBA
W10Iq1x5qSciTkMegKUu1Yn9pk7O0pKDMMEq3fkeMPMk9ScbUFhT6vYgrFMIl/zP
zxkEUg3j1IGOmijOXnPZ/ql42+OxKDbDsJgnVKwifxN3oMCbhb2+ygpily+Q+Dvn
Vn8OSs1eAAY+nlYtrSw2HMFzDifpZKORnSCeOlpXffpKoCGKyA3m6/4sLl4Wks+l
LeLoUkAkZTjYMkEoM8NpkKb8CcIzIlpWszXy/D8WblXvoArHVjTUOmxIRAIxWqaw
fA2EQewspbrscVMssegcRWbOkr4waGgubVXhjt/5V+DuFfXOJzS9fCOUamfAWU8x
70nDlPPOPG8oll0MANO2k3xh3V57+WdZodhp6bUGIA2gqvlFqBYqNyIG+nslnoLP
3FQOhIw6o+DWQAhRnjTbaaAsurZwo+Oc9CcEmKflwQHcq9a0z0azeCVH/PBbgell
uJHXx6ZUUmp+FAGV7ZItDwdqmZVh0UeGVp/3VEFNB4fSnd9TULfcJ6FL+0x3hSS7
xVi7ziJHMR0aAhqewCJ9STYe6EzV0Gdcb9ogXROF5yw2do1NNsZjdrmKX3RxLFvs
yKc0c563QD3TVcRkpgVQMP+TD9WPwnUE3wT25ZjYM30xD/FY27ocRjZMYvEB8Uri
QD0QYoVIX6avFp34JAV27rqz9vjMkjWxnSl0djwWyfi8bTmjSkA0jSrzfjit7WlX
JbYryfWx5h83bAYqImgibpUhyIMTsrw0TmDTH61xgGLSkvEhlY4lniZSa0ekoHfw
wq92LKffdAoqh1Bv0yK4HTPqqxxr2LA81+MSgnIWk18HBcjvw3hGxiYchuNVLXEk
u6ibkIiwIsZVL9/iKseVluK9Na7vGCMXEbA0QRzLqpYi84wvvrSGLpGcqkqnGyJt
X4REcmKYs+NMgQKXNSxxsAAGRpCMn6lq9Hq5BY7ap6tWQuoEiwOnZ6O2v+Hvds8p
HPid72wkMg2DLVFLDaYyStKRFProDi95zFYsf5kJHO4TL5dGuPqKhr79eC8JT3Wd
4KitiNVTNFonZXzpDAmpddHvcj4fFdrF/qwVQFWYyg4F3m7Qzo9XgrLcSepZL7C1
hunnuURMi/HTsthb2XmCnS4CgCDQ2RkN1QFFhf6T40hXjlGLnXqKZ7EKIoDsIM9U
3rMfc4iEz52uazkqb52KQUXBlT/W1tMQStetVKqu/mc/FaA/8QrsvY8KNJsruO5z
qvVAN/mmA4q5yeQvlH7k82beB7KuI/bJv8gSPYW8dgY0w126HQTyfF/8fSI7SbFz
Jr11yBGTucGTqiGoAiHzCJKRqOBKS8nrWTQAuxKbdyalpbCWKzg42u7QSJ4XZcgp
QhUwoa3QE/XqCliPqjpsCcvmhxCDomaOlGZZ6bDR7fDQcb0FnBSbfgdOrF4oXomD
Gnlfba33CceiFkD/Ec3u+/Dz9K4XNHHvizYfbNlibBkZAECRLtZgizNxSyg9KQSf
RpCppHI3onfAFz9jDTCiikKJEiwmIgpxnqIPchs+0p7bIjqgAnxQIUMLP9OBdVKk
dFxzdNjZAIF6498kl4mEryjAMIESoqzrY8wmVWczPl9WmErVhMU1k9mHeCGe2B0b
F61fyv87usQKWRsRdK3+pWTzzvZg2s5sQ25cWF81+5K0NN02c8Y3+u6Cr+9B8oie
NdpYff0rgvGwPfb7IdWKKk7cG5poiIoFJgTknCTn/7e9h48InvZmDSqM+xyEvh3F
ET2YCEA6vBbpBctA2kO4Xo7NkTSoPb1MvDAIuL30pV7y8iq2hPGUSuGbIJlFYyNT
gzcZnnX74A1Nq0hny6WtCzm/Ut13XA7W+GVyTO9GyVbhcET4TD02xJk5JnuZ1Apa
vSiVDNgjAFnjaktpFYZUKmS4GmqBuPXFVTA8Go6iuvMfXMPe+roUpA3P3iTiJ4ms
um9YaXt1C2rpV6+XIfZSZOf0WCUDR+RhcB8tqBn0k9uGP+KCSjkPoO+CIk2BuYXg
c4TZMBMRTi5ckVcvzqlTVG9bdkcYYR1sXpXpi7piWyrizLIkvwsBtwFE8JcbRSHR
bICIK7V7BqmZSVfp/EtYiKFY8diua/dRw2AQU1klniXf9+tl7DiCX4Mau7Duo5s5
QSIfif16We1mFT/yqwwn2sdayMLcjoaBIElKVbPHXGNhuByAVOhESbw5Kfg2sn1w
4xCX/FEuewM0+jkukm96CtZqNm4fJyW74pZ8n0gCdeB5Mo8VDcuaYQq7kNQsjzBc
cVHcSYP4kQEG048Q04euMuLGiSBtr1b2HImqFVmReLBERPWVD/Q4Qa7SpwoqpkgO
AejGybcZ8wDPdQr+x8y8a6109tlToTdE7U/C14s3intpOl8JMSmQM48aOsFvCEcN
ow0+JhOXANtxAef9HiMZ7RpkLYX3qrmllJK+FLml4bnnyk2rW5Y7rOgtaaRQED9j
f0EHogc/rUCnRbYQIn8fTtqPnQCeRkOge6Xh1jUx/sRMLOuofaAJJGTyWNvM71sL
w0DUix09ABH7bqsAx7K9GjVUQCGZhohWjaeFQM6CYIRTEGBgv427Dwy9w5tdhF7a
A6RZwb8hZWPIiC7K6XYLXeox/Oe1tBKs7FlG/z+tVg+X59xOgzGUnkSro6DGYoD0
1Na0fYqRZrIGM4O9n43z7hlld0Kuomcod74h4ZWj2vaFYlrSpR85Nm6T1FbCPMBX
aHm1N9nwfH0uLHCylPuI85VLyZ0Ey2M7bVjwWeGVamIhMExk9MeL1FtNRgsY4dNl
FiLveB7aKEPpvXyEBUxXfiA0QdQXKtBIwe3q32PmbnlbpVmVXVdyYJC1enrsW2Ea
L9e1fMvEIF4J10r8T5slCjHgXSm3G8vkTLMhDYOhCR+HJwx5dxxRrgacLZLh9WKu
bi6u1STCRisaKw6zT/ihV36Lt+TpKJHt9Ievc/UY18SBIFhqVawdhJDHosbn6oJ5
eoH8l/E5DLiKeLBxNJS2mmzsU9CO/DLOIvOSD9s0Ah8YMBbtmAuX5SBbACgjDQPe
WTBB1/aRa9C08/wXgomRNNmcHtqOnH3/xsEuIfO2D7RwUomkeokqNxtKbQlujh09
0pCcTWJjg+O9ye2zJaD2D8goZMNcVTlkOZsB+SDLcEl4weF5lJuCQxWXzCQ36SdG
BSsUne5A0GITZA9ZH4EQE0Rx2PdWWwMMXvm19qeHP9/Iztz+Vm84qWRBw0OfO4Xx
u402XNYn8pfzYxC6H++3uSEhdy2TJQfr6UaKu0M5KgD5ZOWNnmpeZ/hbFCum7yGI
wyyvn8L5narc7Qw02uNkWHpHWZkdy3LdVPLCOAHdyb0tKJACHm9n2fBsEhqYonm9
iDKwQvFLNFAC2PKpfRmiDjsYI0+b2OxrLwMoQQYvdqkViGB/Yk2KGYnCQSmBNWXv
XF8R34kYNJx67PCJ15BijZwgu1llXCYSu+vbYe9GKmQTlOQSpvOyTZ7yTEEXiD3N
4oqY9/mhRbZQIP2L+UmfPJsdsxuTSRUm2Bb1cCNdyfQjSNT8eNd/ZfpUHL+LkGKs
E7UtLVJ+Fg+kdN6bcIUgL8nY4pAWydVg7k/6/wI0BW1vfKpf5L3Q1DfNkw3rd27G
kWwoUgfk/7/eVsopHp/lCpfo48iCkRvMzS+exqx7D+bRZCa81RPuoxhlrtNpaEfN
w2krciJ1afAteKJ1/k5Z9P4JXfVd59pO1w21vh79aX5BraQ0LslfVn+oTI/ZhjUB
/yc3HDUp4lJG3I5lF5k9s4pGJUrACO/djkMJDpj3eG38jMk0DbszGK88JDjRkRw3
bPv4AD0ajpkExJOfu0/iP1/uKuQTVEXcwej4kZzBhoguXYoQXW35FHr4BJ3lj9s7
csaqMacDOAp8Au4N8xn2Hf3BXOdw0auXT9TpwciG6ineHR+UA83lzj0WEZ4pTemS
6syfEJtfcalYtW9A9TDnvSlji1omI+/8hXbg6M6N6V4IsqzOfy0u6Ztk8LRHHsvL
qZ5WRp2t87Z0QzDQvi0GikyPl/kFSl6tocj6WD2XK4pa+ZQ6DgQQWqQhZOnq3XUN
ZQHkHIIvjrptH3X9HE1xuz2GNTuxG4V0gBMZF3guAuw1lIyGq2T68YCXBMu2KKIu
3eueNZwnc1W6+oVPXr/m6LLh4h6KPaomvbgazeLPehDoUYyL9I33mjqlvug0cMAy
AlPNkKn1LMJAqR/eVomtPOz89OjMyp4xUkQpwIHVSvdWvr1hVzgwtD75VyRF2mn0
vFRXBroRq9WGE5tQYRQDeeEggwPGesYjtKtbIiyVqpw2NF+MkfjvKsVbtIC+y+l7
mgUCZhu5lBWom4/foYDoRwF3OvwzzUb0hZY/cXe2wibgToVFP3qhuwjvZ7fhQ4WH
ce+5c+RJQi7QPAiwZpNpyVg5hFlaWv+A9XvFhH8aEw9f4QfoCumqOov0YjkMoNTp
ZJZIuSKe+og1FHvTpKOmUR5dvTKkqLK5VUiCo2OmYdWp7nEB0NY85xpX1Siz5iqg
0oAMFIruKDECD2Fq41S09qvhznVnkcDKPcBQ+Y9gqMnPXxqV4D7bJQWuFFdDLlCH
PxHsQhKmnjKhd2AN39nxxN/QMxgtC+MxEHPh+z4rJ9V4X0yDoBQ9XfGnIlTVKkw5
X+rHa5GJiAhGRb62COtKlXE8jMGxik4JAhkoxT0aLLyiVjPwhf8u7XwcOqSqTaz1
BZaA3HcxnIdcAJCLsuUdcDReuYw32jRbjmw2aHIAjhC9oFkwZ2vb39O8N10mPaMz
fLGfp6cN+XIA07y5dL5H9+hDMqQbWr2Gws1HEjGI/erH4JOG5l6F56JCR17ek2gc
dKZOmlKnARodPvx/yCR3Flh4c1zSZgJ6miiVBhHhXly8xdAFWcXLoRDmSoVL7jNG
wT20J4eaYgHaeBpaUy8ihOt0Gz2G3WHBPt2M2DXqJXKgNlS5szJQTUiHIw1+ZsxS
+5tk4fdg9+m8bIeY22dXD+Jb47Pi2Qub4UBeNXkCTqhr4prJWs5pwLwEO4rw5oAy
uFOiWBOMrADQfNpYfHRG0kl9v/3JkwEtaS7RVmY8APJKWke+L2MEhQzauUsfvSL+
VfyaJ+r8LblqPKzy1fQFTWnljrfl+h3RlGa0euT+IKNVMdeki3FMZ6kF8tmLpo6c
Cp9VFURqAXABT066/TxEBZHF+tHw4gQXM/+yhQrFykg9ZsuDwK6fUgy6nPmsA8qu
01lw3vYJerIVPr3PZcaiGvUf4gBLr8dEFw7+XoVjIOzs3Cw1En1tqKP4CqohUTk9
lYsGiLHNsDr5Nn27EcZ0+Ldkj0oQaCrX4hFXjSteoxz/57oixgY+Pc9McdwBuAgt
UCMfCqYDbJMSdNydm/M1OsMOMT3ovYBIZBw0QaF+xxABL7x1OX+YsHMmldmciYX7
6ZaRrJbaui5+jzNT4kruDjzahh5oE6uhu2ikDtOSGOk8h+PlMGsOdZs7oKL7J9O/
583VVj0hHihxveRn7oDnnV6tHmC0cBa1ijN5fI5r3xDQKEsmomm9MMkGK2gUzMS6
5rIxTxDaZD2CHI4o/IKNUxs1InOIcMxINSvqndpe4OsVhvru8WQeRFECGl2NXv7g
7j9qPs553teWmoQYg84GtV+c+GBXaHipnZcXQSK2kze06ZiTwG8CXNTC3fNiMaV/
tsS7jRnNbFJAGZKNuYN4WH2NE58emxapYjqRJttiZEP+VBnzSkw4va34CDN5dY8c
ysuFu5tsF5X499V+Jwpmol2c7Ur72Rl8oRym42AcBa01d8FAvBfy/001yAkIaydh
VuDhL4jJvSo5pnz6dTys0L7dJWDVkmKao4rPwC5K29/k3EUXijsQjKaE4ljr+8p/
eBRPcq+v8PWuEo5HeyFGK1L77fskRAT9sa7q8QkDmcfKL7Onu2/z/3mBVJ0tcqjw
eZrXk/xc8OBfLGdO2Qvhy1my3qa2uNJmIzyV0D9TslEtafHGkqB8tJFVwrhIFjz0
upCXJO2h/IZo7uMog1tzV3AKr7c9BE6so2tFGv7x/ZZU856ZJCPwJNEsfcDkRCsF
vxfjmue4u18vdnVVc5BuXZzbQDUl+6W42lTmkMhNVkwHvzdY9dP11ZakQkDR4nCR
dYL4C7SkOYOb4RG5uResCelUY32xOfr+L7+iWHA8Jmk0LLENLuHpQsEsznuAOKtL
ByRWb06uWKA5LQyVEu8NzS83teKfbBm/JryE9GPB8sZtGfMS3Zvjdfi5dOfLjsoU
k/dQjzuSCoi4NrWPdPwOsBXGMPpxTvzrE5xM4aIQ54hPA3QNb06RRrc6bUOm2x1k
K+p1MdW/yq5zPxve1TcJvtZlGVsgU8WkfVp5VNeb7wRJAHYCATBKRLe/em/7uopb
8YYx3YcCeMHH2MII2GIWSNOEYVsWHlGAbho31GogeKyQ7C5qT79l4e4YgKgspR/5
2GRaQcCoKNtM0Z0jo7YkJ0aS2Pi1fbpQiDZm+ftJiopY24i0qfC4uWsJaRN1vCyq
NwVv8y7M4BB0qQcLEpWAnfcBJqDamQeNqaVRDPbMCljCj1hSHzngOwkNPKXSYQlE
vw4MGMsfSJBX//0W4LSrELpFzjmvLiH2BiFJ6NgQj9WcnmIAKu5F4JrRaVSmsSh3
bTebd8meweWME7+PLnqnUTve/4mqyAsCgUVEnO8xS3xU0cMLD+7m+zVaQcseY29B
YL1jwVn3mv1CeYvxPvLGcYpVRj88P/wymRjRQ6Kf9L0a9BtX01bIgRqb59c51ndc
1qte1DRIO61fWZUXqxDsJgxUcHUTsLpRBhCsRD2ceka7PT7qIMLol0B3tQRQGt3O
rsCjVKkeJtumNipeRG3xqPh/JERSLzVnhzF410FiOEaGcM8MEpIalQlSs/ZMeTFT
BiLF03Qy9C65cgaZbYAdi0pyLgLC6zQ2w0tq1KbhlEHWqYKJg97Lul4ICIne/Zw8
UH5t90za9HwRS6URhdldlkfr/jOY53KdvHED4tp2PQ04zSYivu593EJrOtAObre5
iRqnqG94f0u7fdA5EyubVn1UyM6mVO6w/AHVDpRqusjCCd5UFmZUndMxaNw7axaa
YNp06ou9EyJcwRJlppVKGN7coPmvx5JMTvDVq0R0FN4mpMWC5D4ATuYK4Ef5Q//r
nfiq+TzqA9UWH9oHKt58EmEL+iPHmDbwqK8VErdH+kspnIOX1M04sc82kFZvRD9+
dn1ftB0SiughNLg5mRrxGvEqe3znIwaPJ1ogh87BMkNOB6x2oiX1CR5gfu0X3hzq
cMDfvvI1MYNQf7TM2KITCG34hWslByrAD3Peyyn0Oysj9m7hnPyQx5vTfgMrxmyP
M8qgpOhVkCgAtwWnF+KmcuMiI6TPVquNOQ7m+geXJ81+aUOtLS7PTl1Uz62UDPp4
+zxKYcFDa5oz53NqEsG3C3igzkyGoFnZByieBcL4PsJg3fh8Sa3jPQt73Ap4cwqX
OoKU+QEB9wVIj/kR0BlAYguftJEuIAlwkYty8pRWzzMnDvVIJXf+Kp9S0xHolPbz
rUKkF+xPnD9zpDZe7eoNcciKtq8f1cQAi4oAV3/jMQWG/KqRcj+VajG9KV6u9Wy7
dP4f2yhyi7LqlUEsNlUSmXBgRhsl09iITxImGER77MRaq8e1Hfj834R6FwSHYoY0
cdZydWWD+BlHsQOQYcztWdZa5Fpkzqj2GDVQrkt9AVJW0sCJExSlzxVCqjGxUMgB
Br1DgtCitMCtMVORPNbzjwi6of+OiIljO7HWrIMYE5P+jaQUHX03/suDr+qVmnTm
/LXVNS0WR6fHN0Hp0wPIZgEDVwrl9/jHMr8rOHNns7ZjxWNHNBgg3Ufut3d7sg17
bJuh3U0RKrPdYuI9NNwPaJVoO/v6VUDXds3ROhAbevWbB8HSEylvOsVypchr9e/k
xb1+uw/RzSR2unXcSBhMtaKjaGZZfAww2fiwZvpwkhOM9byQICpu38YV52cNbs11
bM5pIdgZUsGXKSyTzQJBQdpk6UzLRo3hz8PBRLQb0Al9tU7ML9enWI54k7JW8ORB
0Ycm6FtWIh/hq/OOj/HU7jriljCkRH82SujcikK4RHTk9mMPWhNJ7rhyBFJYUQ+t
JhX/OHgI7xQn8dUZX4t88RJZh6s7bWDyGDSjzKYuQ7wDpJ3wxYN2oYMvvARkjOtu
lJkUfDgVf+dUyHey8f4yNczSWhZuydD0VZV7IcwXaHuG1fkYibaGlKzdA2ZP3t0N
Qs/bMGDmNXqKs9VzNJKg9vWJ5HDUH79t32WNqeMNfLIQB2QtH77K0g44LiJ7CUWr
oitgeaYgXiS/MtszP+MSzo8Nfiiun2wh007dizVRmbGbieMYR3pJhZ7YnBXq0wXO
4yTQV3GytJiMyWPLwJML2yteBEN870RGHzlY4/mvMKTW9uKWhuRX2lzgYMWHg1LJ
+Vq0U6yAXrwPQ1WhD8abFL2ldp0hbgWDPJzcdwcLIRQpB8CnlJ8mTkeSOJXaXI8j
GzntVYLWjSf99QbabLkPzpyNZE5djHcTUS+XrKZzsgjDFWeIyGRtySdgNImZrEiZ
lby5V+Cm8Ta+dsOhmD19L76zkFrSbL9rJ2NpsCoyUE6+f2izP2P2i/uAxtGvvwXT
PETEGYheA2HfNMVpNJgCg3Pp/p/uMzvKB9h+lXH3nicTRlWZ8vwwKhKXSF2g3czS
eZoG1gmw/xgwq3MJcK/qAT6tSHf+w7tsOmPJM91nGOilFqTHSc21zxYhvuFA98s2
kpvL7j0OmbbEH2RLQcFzWramtzfHNgqsU9t12ri/ta6Y4BppABux6zkLKKc2zzhb
X3NmEa3F4W9zQ90qlSbekd8eLtidMUJR6BOhRwYDHfOeBIdYoaU9o/RuiurhH9yO
bq+NSryV0lfHsUnxWs3ZUg1129kzFahtdQ6y3lXaAe/uMPGMsl6x0bvP9HMXOO8/
F+KFePt8jzZb8Y7fuSrkqmePKUyhE2kqIjrIntKUUOgMHtDCjtVYdLHaRhIIkrVY
5Uo4+PQ3TmiEB+6pkpCDhyv1KvxWDG0JxC2FcWux/RCV7+yEmWBQtRwaMW95ZTi7
dl4sQVVIx+BPzMEdpZ/nfO/zkKPCJ9QPLsJE5AEvu645plvyZBjoEOVkBaRZxDg8
UUVF4h6ik3zzt7yirETAt3Su/YoSvCzHzafyytAmf5BFCut7TGGTHhHkVJE2NlzO
kedNoDvm1LruAxl5hqg1scBOGCzWgTTZb6bLkK+kcfTDtJXGUQAj9vFfxEqJMemW
D4natZyN+B6iA++9fQQP2i0gOfLbJTSMIj18b28WTVaW/YQOJwGpiDJtsjQ4c6xV
MUi2ErfetfLzKbR/LfD4s2ewijLUeV3wcH65ukxRmpETIij13M8gQ8Uid5GGVkxi
peWM8HtCe2wBnsObtOYUmZe9VBPc/DCGqPVs2gaE+9t85CU9VJk/hYYrMYf1FnM7
6iXhHInz/zpzJom8EOjqLfG5WDGIQG22Fuhf/MrNW9mbBRCFdf10QT9Ig/ut0s+6
PHWm/t6DgsQZlxfn+IrmDANG3g7IRsyQuchs5sLnhcp8xIXhkpSP+b1Dw62/sVzQ
1BJUSyLfM64o5v8itbJHJ/VjLHwNYhNcVZv8P01XxHnkJe+hRpWspcjf6HnB0ELi
qDl79PoXis0y8uYnE/gZ0Sfhb90nVO1s4fu9nJCJ5tLgwnc4Samb3rOYC5cvBTHr
KQX82yQ5QFt3Sj1UxGwusg3HJuV/e3/6QxoX2uTybqh/sRaLqq4+j0fgaj4DnyHA
dz37GguCQtNJVhtRKqE77img8ymIS5ptSYdaLCK/yQBkuKgpGDAmXTyXTTUQ4HG+
e9m4m1oSURL3kwub3xcPlUEGGHYmoGO0p/RIutgiolVDKE7jGVRf0MV2b2CjinLq
jnZrhlvATUjF2F5IF6kJo3gH3FbS0BvVXy1Cki0hGnX1+fqUujy0a4oql+gE3ldm
FOO351N6AVv63q2PWUPdbkn9tjML1DCGG4ioHM7dDr8x56NEJ+pf5UqBJfpZ9r99
SUxeq0BF1BIUflsV54t8cbPvlVQWeZgvN35eA4QeY/HZeXuO8UKEEhyr5alwwben
mZE1OfEp+V5bVqqKM5WB6Is34XKoOqcBCdWySo2MIbthfHOvHyp6o7mhEcoHc6y9
167wmb/F2Bpfjb6c2mlQ7BtSicGzXW7f1RQwNInpEa5a0tBIOw7jV+jd1XYi0RSA
Fq0+jZ5+8sQ/X078KTP5i3euHsnmAB1iG1y8Onb2iXnGFDjRRxVH0xevnanFLyhR
IvmudgPMoD8jNRlvsHB4ZwQHOS7bBBr7QGBQLKC7fbemLrYnvALaaLnzCIMfa884
Dt0b7kB/Q9L+1UZ795ADoJR0bdPWGpqWMnausLv261v4ORQ7m5fcHoLpbK/uwU8C
2eylUBwwzAzR0c0OH4pk8eNukjcV1AnoebGPJy7slTz1oCLEz2OkLcRILFuYJjap
NQ2tJyK0bJCZULXhUW3ZIps/+2/SyAzW9MzWvKs84SbHSm3c3ESzhWn/LmknngXa
hEW00ABbJbafwbpmGeqHutsAYfGvLVXxZl0Zj5ARCYTkZX8ijmk+h4Mj0d6XdE4L
SozmxkDpvNVQGSe8YliIMcpK2WnSRW+qSV47vbVT/w5PN2pM59wC6L44oUX39Gs6
zYCjPkfHWJJIWvpQrc/Y0gee/CF8q0my38pl4hR1dQ7MMCwJUqtJoi6B2OoeyMUL
jb7IQvluHc60inqz+Jbc1FKufO35GIY0O7x+gnbVThApyeMe5l6cZAAzpDwHkIFn
+v1ZmSs7YTI6jIW7u0NzdUaiUUGQP4t4xpInwXIrqICl7ObK9l3BuYIxKnbVcmJY
9KePnx/ziASykPxWtvcaaTuLvbca2t64pqdjTnGzjqIcQYD4Kgn2pZX0UIzb/SBz
6I9Glv+vO3FVApzXi1YiC9QXm1v8oIy1N9Ofo+5bToX8lblXPms+Ab8116R28Uhl
kHBW5IHk/DUut67HCpCXh/B+jN+aeUkTtKDeaPSCwJTyef/jIvk3XGjDNwLrwA1a
Nas3rpC8/r089N0gTVfSQLDkoaeh0aPPOlhqzQGFfpkgXLN95z+OWUE9ORR2zwOy
L964PfH3+umn+rbM0AeB4pQ6j6bEb/V1F5bq66cSb5aN7p3N5fJRL7frOVuLR2b9
sYrCQ1kdVA4WHLbyn3+kdxiBEqevQ0Ff8Nz556jqZsW/FhwRpxuvVNcEZxK9+H1h
me3rJ5pdz0eeB32ga3BVpbtVJDhnagaqf0WV39Nyh69kQNp6IDQzkXHOQpRg82BC
lTGZb2USTHv51Mj/bKa+sp3ADs2yQZweeH2fcDoUi1+yJZqRUXgb1IocD8wZUF5U
qDJq96WB4o+H0uTQ+E00Nqpaico0etXZu3fJSA6POXExzP7LGhnhcroUqu8cbYFu
Sm29X+W7/KcUYnyRc4ZvB9SBUDyt/SpuK9Aw6pGOAqzWMcyl0e0k+nsWgkHIZpVL
1tBl5TeE2Aglo+pXy7Rmk4Y/0lUJW4XnpHFRIe8J88I6S1LSIftsVWF8/0Wsiqf7
cxalyWT3FbNgWFX7udk965Rtwi7z+0D1Yks7KHDUp4Q0GJvf9AjIChYWqeB9mJSL
thaFtP5u0xRBbyV3+P55iIxGq8WhBuF51if+LUMginQdw6fd0JaLrrbgr7/qQYge
Qges1zS5o5VrtL2tukFk48XKIMrnJ5v9umFPZS1E+9t7olrfQzNsNVeU7AsUXJYJ
z+9Yp+STwdFh4/HEniNOsaIkRMLSe7cU6ft4WH8klxix1IrVZimdZ/Af6rqEReyF
ptqoHEdn2Npjg2mPNuWSDCV4aj1ctBZqrQdh98tj22pggvgFzq7mKjSjox0lLy61
9n3kocuz3w9EylF1uzq8r2YBWO1pI3X+AwRlCrYti4wu4mo8GoyqRZpAtLYJzFor
dv8osvDNdWmn6YD51G7ko90/KA7FRG3RZwtzo7ycsXsqERcl9qPBDlkM+23iQMXZ
I8RAFYqQoAYWaCWcJjQ1pdlXjSgMWgVJgYRq6iClZ2ZumRioMSF+VllNGxVMlbI9
Pw1BffoqTmHvBhdoY0AIGZlI+Q5nmHJGvGuzKAqzTRZTJPrzBo6r3wJRaS7+VIdB
PWsNhP1ahJ4OVN1TbcrbEgDjqvZZHwP81XsYkpl8jHa2gTMl5quWHvIwK3vA8pNN
uyGGWs1ifX8SuLauxTI0xersXYhz5+bGs3RMaXpzml9MAoqYMkdChuQYA+CboaPf
9XFRiXxuhTmdWzZ6+j5SpFPL3NQ6jH+BVFn5SdK2RDXZ/VPO9c1zinMU17N4xEL6
yItY2hSbdBUiDc6pEqoq/Iib1xQNk8nDHu7kcNESuYVRoFNo1jLAD+seZwEZqO/U
z9H2BDDIlTfMWEqxVBPOjDMvNCdupWFNQerbbYn0Gm+hZNRCRFRTDQStnHTbmzmK
zVexvplVr3s8GSrSI5gdxseffZSCHa3ZwtT9uBg0nn5uJaE8OEi/aNKVZhaSJ3Q8
FWnWJdtJn+2ZuD7vMsjJzsvJ8keBPVQ4DX3DHqLAYp1MKsheHxIZtceNz2DFD2zi
Iz8icq3IFVwpZXKynCi52Hei2c8VqAqPifgNKDULp3nFLOfNyrY8hzNbIWtZMlf5
rR51I2NEYLsOvdqLyy73oLQ+iUmEM1EJgOedFF2R2l3ssDsMP2Xo2sT0dG4iWw2d
wsSgZSgKU9i2E3QncEDXTYvgMIftXCacWpyNKSHpKTQUkAZy2cAAIft4JcyC4nzN
omsFbLpZp2wbW9dOwvMzZEANLkL6wiQkbBVKwYZKqODm6SNM7GLoKTkEe1MDKAES
2k/7lNqnwwbzKFz7c1qYQjnPwA5M7aaLtg1M70Q4rotDjbYTloMMv523QQmeTNZr
8nivFqwXf5Huj+h3qYwMBQB66yt+AMgCiSHnvO9Z2xFUN4MpeW+PuR5mG4A+u9ft
tLs2eiaqDygVSCSiaX6mAPAcUDZ7lGw2/E2W01yMDSYyAyeqoeMz/AnlRQBn7dx/
iuz0WssRD8rDD9gQYKJNZ/6g0s7K/IcLW6el87BS18AJSDVH/+xC+WVR+sTEB81q
LqpCBQy8YrN0FEROTXrTyxhYVVmabejfgA9zRvnR3rxz52BpWZBiTekzcOhp1CIQ
NsV0lK0xLwozzKSdNvys2GnkCzYoENhK/3Pbx+SdyVvmyYyT6tiPXUbADv0M53gQ
OLRbmy3gcs2h4CvRJgX5cclumnBICXJb4Yeo210YY7E0L7yGYgtqPMc4xLEwbezf
IvQJCVwUX482rwUxVm9nZycesRB/5duawmrmUGGnv+PHP4Slah4Y083xpXhevKgR
l/3EpQPIcigdyBQxph/5ZtG8G489obx4W+WGDb0pDzgsBgalGuSFqV5LfcY01gzn
rCdH1NXD+TYQ1LmE6wxtobUNYbFSW1an/OBni+0wZJXxyoYefhiQJQZ9/Jp+NTd7
vyWBkI+W2URe6cXdZuhvWgXg0xlWU4ezP/VKCu9aG2ir8K7+KBlCsxiGrTqUxuHb
QUsQRsfwqIdp2OZnJIJurTKO9fMcIvGui2Qht+c0GNGs3oR5Y/757Zzkl24xyw7H
93xwau4Q0CcQj4ALu42n6qB8SAqW2nsbZxFbe3L8cTr1sDLnIp/YX9en0yrLuUWK
Tih5ZeWBDJt2nyv8ss4As1jSH/F6krOavUjc96F8zMWEDb2o97uNf2ZzUtavV1ok
zs+OGySEEAigvDbAaIniDfUk6s3AqgTRXCEO2X82AHC13GdZWfwjzB8GIlFxnYgk
pav2Y+t6Vr42YFYcGE0fhPXZZ3AzG1bAOxOb5dn+ZUaNMbJgZdGcYjyDLrr72mGR
ilIoQYNe2pfDV43ppbaPINGoC9ZcfZ7UG61XzUXdDQ7VFyIM0Fbl+3u4RFjrrOHm
RhCM/yeZtO2VY/6DfvOUo4ckXgmsXU/2ThlAyAq8GCgUaozMEiIv9Y+sDynMC5D3
eUFUNvhd/r1inY9I7NFvhU0hlC/KPJ5xkIgob0/0ZbCn73MmqUZraoTAQOX+/Z0H
QCefdrkqxAqo9JFDVn8dDicNqMaOOXu99Lh4SJc/sbhCeRRIEXkuFE2993DqiW9I
ZI2qHrjTFT1LVQOlB9faPT2yB6tKlRDjQoo641F/4N+VlpLnbCmQGsZNLnG9kXUG
ErcRjthc6N4aTTRke263RG9yv/toD2IqoEVdkKN0vz/0Gu/CzXwzm2MG3T7bYsMb
OLDglxAGojYi701U5IRuf4JAa+uTw9SmkTBvajqvkJRPkFLdPU1qsrgqq+b34QMR
tra4o6Z9TjmtGilPtd7wkqlrlmrcl1kJY7oVd74xng6iCKvr32UlFPBjqt0RaYJe
TSPeL7zc9FOlNeyEaNkhYyJ5yhAeQSNeCuge97L3APjkNOh04eM9kaN3V2ugWwWH
4PcAgeiGDwQ0bjbUeKw67xMMod6JvqRtxmEiv334VWP1pFkYfytdwUsD+h3a3uFJ
LXDMx88+z/rs12YbgQNvAKjCr4TSd0A6OHPCk8s5hY3VC+pgy9/YRl8aigaYNUAy
V+DGpAUkuURuTZv1cGlMuRQPsirLyjHaR3tTT0BwDvGt7RzUHK/9bRpZeqNwF7PH
N3ElOxn7dORxCy7UFub+t+Pt3l7KoTTCLjjIz/dKolS2tM6FDqH9HZZtMNp1on+U
qzhmlxp/BSUhEVewKyNUEAoKoul0kQRUqRnarPz0kaCph30nXJOYIsAN6Lscwq2L
OxwjDYEmTRgd4EkF4q7oT1qMTWMJeudEJShE+NEKnFH6MNOUnrF7ScTJvYD6AGwK
hcvsZev+jgcg2OITDmkFyW3aSW0y05IpQk/cHB2bHfPy/Fgqk4z0VwuTI6BvNw42
zbSh0iSPgiLnjHsrra/TwhKc14mSQget0a4ORD+is8CqTsjmOkr/whxIufbCoWHq
12xYLqN4+qhVWRMOVGu3YlHaG3K1qOX0swkGzP/6xqdHlFnG/v9tD4+dUAwHl7+j
vq8mMEb1jZo4PzY+/YYOaYJhZdAxIkhyArImxYffT3oQdi/4GouJthDZfwVLO2YW
xaznKrrDgU2kpgP2fTA+J38b9N7Vr41Vbb8voWcISPSjfw1SfmdUTGiYvOeWV0VB
3ZmZzGRXkGFLX9Ks171dipFQ6wNARE+cqp6l8b9awag7pfPqeA2fe5ZwnKlAJ2aN
YOR435Qz0XVv1Hz51iCcGhdkZe1U7KWWZnXA5SpSnmfJF+4kqJuRix4idBAhb74k
OEs+iv2yZn8ceqbjwRnOGPLBm4ANwOAxLbjP/8gvxgOqq5H10pXUrjHgzuK2Nnli
XPDlpsyjxg8aHXv03EZLfY0j3vGWOoYrEzSdAuEz1wMlueXyu8f0nblvH73C6uBp
AcfvtZ3Fv0mrfzJqE/hRQRuLFoTOIV353fB1gjvPEx1/REvjprlpSr/VAdvqi/hg
C3OrsLUv06/i0sLyEUhWc30vszbGDOjIpQ8+7UJN0VJEwmZuptNIdfNcnafnDpf/
MefrsKycIEcEi+pT7TelVW3q+IK99JzneZ/KWV/IZZrP9wSfvQlwtrSoUguV5Wm1
Wa3/CLqJ4F1hJZ/wpTIkKI119492G9Mol/qzpo9fLAMhqToLtwq2weHX3XPFT8LU
fI56qswhIHx1q9xuzvh0qS58qRnmMPQT7fycW0DSduR/YdCR0ut79Sujs1aSNssb
iYhRrjI+xbJmsDU9S8RYgP9oQMQblN6srKuR8Nkv7FPgDGpZTZyeWyj/XT/dzYOF
WQmx8pbx6zBr+W78ErVORm/ECw8HUaiNVPvZAMJ2Lr7rXY2WEfwJ/KSFsTVsaxLo
zCeiLazlyPsl3f47g8Dw50xvfBW1Wl/X/nTYezKaoAoMCxbICJLdpzP7k7IR1sVE
sG4IWVUFEK7fsHVT+l2v/rUMfP35o0+JxrCvOtMrBcQ52atpggSndzv0VxYSZ1Qp
pcCO/UtcnqWyrpJtakyNIM5D5ddA5+uoRklAovJ5W3DNjt+M8/O8s5ubooEc1yA+
esnTxVnBG46FFjFKlp0AW25OrSHqgvyJT7YFkYzD6Jj1qM1LZcmYAO6+OPWlnYcH
KAJUlSoeObANKcpFMN+s9ssK5rDekMQQRz0mqMJlX/m0s+rgDl7Xi/JNpWE306tV
5CaV6hw0XzMrKZBYZIoPIcBMpNhr5rUq7DLUvVqwdls1h3q08aK48qw13ULso7Bi
RjWf+B0UwHetqu7A45LGgEjruKgBsFPl7J3FTC9/oIoz+zCx4V1NC7+ogUrZjLfc
hcVWnk2yAT2ct0nKsmGcViq8fJD3CCFAy9zDPn16ecQoW6FcfkL3gLyx2qjl9aRq
5DHD8GLDGK05w5xV+wv1ItxdUPGnQisNP51eB4IhxzxSFirkZCqokNKEwhpxlvxs
IjznhBBkTcWAqRLqeUudHv/8P+vecrH1QPcAvF2Fs2KJwTlRp8G9D+wVk2waLxsN
i84RDkYJke1v9lKEqWSwtu20GyIPZhl4F3/WMm2AA6zP+pfjp6V+JCJElLxvAREF
wuNoZp99iJD+z90kTmyyQDZdQFGpFvX1V78Zd9IBtVh6u4xckONZWzYz4g2vnx/3
zjvPxX1ZYpgYyw4iV5czl97/HYB2sRWbGn/6vIQlG6bIJIWUi7QxnFVsbcugHCeV
NHfU76rXjKCQzpn7fNr/qUdCcZ9wUn6uWd6axt3+/+xzXW5S7YLVqW8zDbyS1wo+
tPKtQOYmc84qBUFOxRIFvngX4YJyAjt14ACqpm0vWKGe6b5Mt9R9ZgHjBIdou1Np
l99NdpqZOjQbiDv85noxUmG6GvzAyDmp8nc70xYvZSTNs+CPgD+o6T1wOSzTjRQN
dhDrB3Rc+VZjc8PPNKtp3YuNJ0nAlksc6xJux/J5Uf8uWX3PwLN41dPk3RCrwdhK
bpRO2VbBh1ElA4XuuJMtOLDRX9TSFUsoktYXbjEreAdxlrT1tqtNYz1gvPPXXpRo
215W0hYD6r1s12CNo/ze2nI2lfG9Z8NXUY3WFFrLu1fevyn7uMkLRjdw0X/X9G16
7lR3cD+GEOBwV8ShXvZSsgzvseZaWn3aztE9Cvi5JEiWTQ5pkuBnBIh2lbJV5KMu
IKxTuAmUQZD6YnptAbj11h87INsLFjNutsFgrEgRFZQLghkXzMEp8tU8ZpHRPN9V
tjMs35KoyacykfWXR0N6MEzYgYlzTMFUJTz1xG41mpGvJ3wynjYQGPYhlH85GC3h
NyKbLbuOUY+9nzQbG/XQB5nPTfYpF8dMrlr4JT5iL14JGIdgspqcc/L6WdeVNT36
Hukuh6tkj/YjCf7hRo52CaFa2Y7fWc84tSDWN+w13Yu4G6Z3d/wPJFFSXmgZl3aP
Uz1VkJZ8/N6MZRuWGNpM3v/c9Sy4JYpjDH1BDQTc1qSil57k9Yjp8BB4jK/XP33E
M4Bwgpidi8jWf8lmxNUpf+ZOYiM2Gz+0Wj5ipdrFMRA1J4fexN5/pFl4K1VkrUqd
m+Yrb0A9Vcj3f6px/q5TWT9BhKqzaUR964pCZL9u9i3iFGTb1cwbnqj4fKHfv5Wn
nTt2JUA75TM39Y1S21g39U1GGkp0zZDaBIjBcp5Ivss4Q+bpVw9SD+e0XDsuC8hy
UzqggKNEbfM4NcPPVt26XqKPDzV3YCe5IaptFtilF9Bb9ZxrK8NJIM7o9XdDbMoW
TI/nMk+PdyXYZRHatkNjynMNeL4pBm0lndl2A5UbGE4y+R26lXJQRGsuLz2PE5w3
N4Nr8VkHMX8mcBnF+lpVe8fpj/0fJuvK0PdeE1JXf2p57AevGhO/2YRh4/udxWNa
yos5WOJw9vmP6A30vEOQsxYMQ/mSj/GxN7K3NaTYeMaW0/e01aaDSp++iI6ABAyd
FnYx2kKMWSsL7K/uUpC917gpwCgyyERbbBiw0TBZRRvpN5juZPElpgB2JM91HJBP
G++3PpkWUK/MBoJ/0+HYyBH3nCUUtj7wKDHkK0+CdjrE4ixacdWBgcUc23KHluAw
iX1XnzDNacmpIxP+w9sIgsjdKIbVVfFVfWuzPVeW6iuEIS85ym6YfW3hk53JnH2L
5AjLhoWXJoCTzrkje+1YJzkGpRdRzWfqsocsCCF93zUVdCkCg/t4FkIqyfw0PEH/
ItxKF2MDt/rROLWODqe9G3HbJpdGdSk2byy0N/ON9HlvNDplV2BPHI8T1EG/QMTa
o4ieu0NFOb5dPbgKS/UgbSO4HEgcoIlXp0gKrv8l8lsedyxgN7sZkmls6A7lAD8k
VnV3C16VnGrzYDQ6w8R1UCmLlZ0bEJgfsI10+IBAD2erAe03Y8npJKgJOaeSpS7I
SB7hhPyeB9xyisosCjPT3TssX2f2ljW1MzHlSXHweaGtX/jKE9bIr/YpTlIikW9K
cr4SYLQDzO1T1YDNl+Ns+phjx/DwiFF+QlUngXafrBixV+tq6UDU6yuOtbpXBNrm
dDZPZ1CxjczhssOv7lqmsu5P2f2J4Gc9AoO++bZ5CeVTHpCL5xAC8Xwy4vyfnWf2
sn02o2sVdaNHMNyVjwv4iLE481KZkYCgcWeM7SzmIYKkjpXf01+SmEsPUjxhComr
yGayj6qFlVR9NJYGgzRjquEQsNodeogp0B3x43LcnSU6XnnSH55rVDqTueZt9+2h
lRPVVCGZ2xC+mAxiIh9Ojn2mAchHYEATEcoL8o7mPqFn98RjTCZE7g6bCPGGENV0
4yfHlyzj8EDe/0h5SZ7iZp9OtzMVfiMt5BcRWMJZIHf+gGj8T89/0C9A8RNZZvLu
7Hk9LIgnIPr3ZGgzMCJLjOhqqGI/xokFLAvKbu5HbACzaERYnRRY7wPQApba6ZRW
Am1O9Xb8wVNI/ZHov+BmDrr91p8zrpRFqKrBFp5gTxsQ0hOM0TKF6x0KBMpWe+Te
HjkxuD3B3GYJFxIMBlPGSRUbNZ9vTxRr14oUsE9JG+Y5RcCSUUowtZLzWGh8Sg1a
klVvH8hM6VorQeWHB7A9GgNAzKCA5kpBhvhE6BwYoriQvFm/dU43BN+4YBDZxNJk
cp1/h6IXiz4qOMRFFGpizz92+U4zYITemE6a3CV/NeY19ocT7oDL8fY27DacbEW8
Xcd/XR2KglrbnUVG/PSya4W44oYlSVYA5M5HuEMR/1MlKmXjAujrocavOzVDYyIB
RdpI4Fo2oUXf1Ee+31z+RA1fQpzs4elAEEVZK0JoMJdr0EPs1Px6yT8CN0DsulHe
HQ0NWjPAHUU3LAOXdrHCeBuyg0XCYEUiS+x4g0lgtRWsFa+fLvwLAws8YQr9H+9E
fDDcvpTssH+76RpSWP54xZHTI/WVpJsEzVkKEx7EId7SwGFgRtGzxIED43jLebV0
qqIUvv1KEZLCMbG4A4NaE++sZjBbXEtQ5YpkHHMyagYmsTNU8H0dNzMaWMEAnYQ9
aN0/na36FimBRNCt4ifHgxEENHiryDlwtOCViLuiR2osn0IiZ9xYugzSKbcAO8Jq
5FQqZ9vX5grkEfMHLaRQMSErWsD7wbhdy5vmh5PcOLuCLfJHZkfmd8dnClU6GaDW
4YZ9R8y7VoYLw6CW+l929tO+BqfS/Br1CAxR9lDy+4kx8KOB8B6SZ5GkpfSR240U
zHinOGM/zGzzP0ESxfGgKaIK7nBJVI2E0XLiP/X5ZrXC09h1U5iKKICE3CrMhXL3
D1c5Ynmw68pJee02e8dYYHUsLR1jOkblSWZxj0gJl+lY7F6ZoLd+PRstsQmsoaXg
mx0X4IEmiKVZmVRuj0bXwLt25d7ckk4bRD9FBOAiA2VcDMCaCpSPAt1S7v84jQM8
HhJSyL1y2WUROv/yaRNwQoTO0yexarZCuLoUPNL6sXEvjOyyjgMr0jxuUrk2aNj8
vHANuUj5inHlC9Zm6oAjpESAp2OOrYHYZjOpt7FK2Cvx/zTQPv2s4vIO/L7js2DG
HeYivo3x4xYxlTyb1HS6cSkyjJge0thTurqff/pd0K4cJxdXnbe7xx07CUX8BxDH
uawOPpwKfKEn4kJ9hDE8K2uU0Kfu0MLp4bStJetdy+ixScEmGOA51/uBPtaSkn8W
hlyGMedrZdcx+fzV9PLU7pW9Moct1YEpYmKqb1m2I41FtBWvYjGIMxaegfjP6Z/w
iGKw+x3mFu0K7CEPveQuD4Jj8eMEDoPOlDp3rSJWLbDMzPysB1QR+l4/nxMXDzNs
yfYe7lv7AelthEy0fI6P7/+4kgj9DgHrLmumbpPEDv+prPOM7tEcMIhU69W2T8Ei
3f9zJlZLt501Sqo64V4QRyiPPs4ULBa9wHl/i3XKbI0lRIJOJf9dVS2A3fErvgYO
WBd8wV8YygPqmzOJGbfnOYFqPJGvstTSoo6vkO8mbieMurEptYcVb+YEvb6Su11d
87iGKQiqSQEGHvH1u9HYbCPVGSoJamp11qaOkrS1ICpPnlJek4i4M7lOrIrrIH9/
Q3nleBoN1VUDFvCazdpBY9gPAcW5MXtYeJFFOwnyMS4OK8ueq5PErXk6EBPDRSuK
tmqzKjneN8t++QatNHcosz6mLnUOhmQMFsufrro83oSEyUt0oM26ZsYM7OYz+o98
rBSPwi0T5jvFRvsOJkbZTBj6xFx9O3C7KIQ6Xgqujd1RWpMvkK7E49jnPW03/oI+
6EcpNMi2o0CUKiQzHJ15u1+gaI2yACn87jyzAF2dZRAGVt1kSIyWwFWZvieo5aE0
dcMn7+sLx3btuDuQY6jijVHDZqV6LQdKdIK3Fn89TmHn+BfhsJaVuCba69vYtGji
piDx0WQUnbjL+Ku3vXu9ZofEgFn4ie3vMkuB13hfiNdPjewIg3vTAdOBqpTh06+p
NRQ634h/7RJbpgkHxb/sOUdAMf91RMtoRk00xY06/EdlKFRdMrAXKchPueVHHJcT
Yh32u5Pimi9i+zYhtFPc6HaHea/VRSt5oNeNLZdbD9niL4TG2PoG4RHJ8xpSdPSm
TbnHMYtRWc1M8UjkEMhys1/dxqoQ1W3rO/sFWE5yvssj49SjXNKdTgm8Ynj2Gfiu
Vx6wfHg+5qopS8xUQyHzCInJR2myeo2FXrmSXYL40khMbr/vSgIQMSSR/yNPPjIo
O6En8hPTe8Jy8rohaSpB2hKIpTAjfEvtLV2kTXvoOuIr6BHcAe4+82GV82vTvcuP
Z6ufihrFTn0Rj6ShHLYhbpAztlFaMB0WqsB5Ua8lVnt5K0zy9dk2UJgaxn1bEA+1
fmk9wbpr7N3A33mjZOVYYlQ+d/NhV6z9uHh1FjcZ8PjCJbX9jkSPZgtKHOgW7Efa
kvtUwPESCnebiGqYKu/sa/ZfVK/5ZXgu1PFFsZFPu9ycOmpTCSPjHjJa6WtGmPX6
DExlmIEif651/XiriYhIQOJieCOio+mnd8guRYahpDaodTpD6bB+rFvGziJAbWfI
4smsO52AsUllnQxB3m8sdS4/ezXXrgvOqb7+IkgulQKGrRHBNN7I6TNDX0cUFAt0
rUffPtBOCJHTPqWG/gBrqxAJpiukOgOULMYoeeB2B7g5dOoMiQlg+6xnuFoza2qR
b9u0qZwT4b+NFCOt3A7ZkvX+hDFUS26ths9Av1tWgViYXF9r4Nn6V2sWJglzmqzA
dn7kzEwicTn+xr8kIskLGZDasqAOnJdal7TBOGnh0CmHeEX7tUfO3AEQZTQXHH+g
HtpxjdCZZV0+QaiVEYrJGa5lN7pff8Mspui7ZVtk8+hE6HWkemdAKjJeDpX1RNVd
q5rdze/pX1t4BDFBjYcVJOiSSa+HekArJRsgsHwSPawCTEo4HJJBlzCo5hwYXnfC
Q9uJGFK3Dey0/XGFDEmq2J/V6Qfp9SXLHY1QEPfwBIBRdiqOQPHjs6jx6i6hJU3n
Nx6AxkBPHZXWI3s7FNwNNySi2k6X2Xl2nlNmWUvD9SR7TZzAW6H8YubhUxfEoquQ
BSESQDZ5dyyiDhVoKyBw3eYgdP66fJIwjLLQKF7iBbw2i3T+iWGbw69MF7jJy1B1
tVsvDOETYmoSLyBZBDGOEvzMB9h4IA/QpqQsaFaZY1w=
`protect END_PROTECTED
