`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
60L6CKO+WurK3ks7VVoyIlaLcvuAjgV2LALySx9IWG7BRq5j7vEpoQpnsixzyl4U
nko551zGHrgAlKDMaS0b9PcswABwdoZgAU1c+5rPpjRlfU8cG5+5TwF07Qb60jYX
HLRy7wG6tBECGI0KKFoAUHnpjtpNqOoPdhdYmvnPyRaZ1KJboteGYQhgAIZSLSsT
iDmU08if8Sli1DDyNqOqWWRLMFHj+tXEwJrzGNVgftR2+fQ/GV6t4dHIZvTbn6Vj
hrsegsRCzxKniXfhFPzPJu03Pw1qtLA3+DxTyi7rQxPof6mnp6XEIEOnVQOIegsb
pyuTZKrgyjgJ5nwMJfGDsJCn92dh5fXHDqYbM/k0r/ye6J/rF3i+kuS/yIuPLdNP
lsIEoAbtqW+v/cB6IluYqDPY74cv/3IzL/fgN2TOoTEU5GZgFZhC2aG3vW47EY9H
HriaGYmAhG+dUzcQjqh5N8f/xp65EL1zsBldBR3xUKiHsH0rbrA+w+cuAr5B3VyD
TgyOElJcta+ipOOdBSDpte/6asxy9zoG9JAJoBGfi0IKzNcX0U+gl/wI5WteSKwS
KZT/RNSi9RFUbCPOWajEhQ==
`protect END_PROTECTED
