`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3FFVzBYdAjuFSeMwhZ/NxVqjYowfehe7TwqZBiRWZ4dORzqOsLmtqm+y7fm+PvXd
3PpD1ZgWa3dd9ZgkBDu1k1hHdiy1e2it8uOLZ2yYZsSBkocbJ097X4o3K/jNWKTr
YVjdjd4o8O/ROL+b1aHvcU3DlvGKDvstgVzoPnqA8D9gb71Blyj1CLu5v6ou6aei
wRGA931Qe5+SrrO72PcsanOlJVBtZkMuCAlnceP0Cgdk3/sg4i0NPZt0VKLceSBB
4JhNFzmW10pgJtBFHjaJRZDmOecOEaTR47jhuUGlJFwf4ZGdJ96/pBwqphDaa2VN
XyvQoOOOA+cF+3h5iepSwjd+//nqp2DWdHlNLxOv1roHP2ttrTfVMDXU4vTtBpBD
oo+L4NDeVFgsjiGdDFwF3cBqJLUATbrr9wXEeeBQAfC6RknsTf5X1UK2LR57noMr
uZGAOSPgkKkDK3CULvyOONn3N/PF10SghVE5/wwyoFEt3AnTuRMn7MS0JX54wtrX
ohi6Kg+bFvGPsoPzLzvqsXK+OjMMSHYxSpY0jlZgeId4fa0G3TTs100ice8eFkfM
steKUyBx8Tffm7KN5TfHxovafq0uWfJTjyYjmeoUkyA2SQgeeUovjFypgdMxrs42
OUzHxcfzny34mKEhxwPyp60tCmVvqIqoOCJp32HPXc0PBvIyD9wg1ziK0HQFewNB
HKX67ck6xhf2hl7xZLQbJQpHTKwt9qdZ9JdbBbcC1LgOuDSitkRbQoxSd35+8pvW
e+2G61RSSWHBDWFVrQdmRei9qUKZ9L4DbKnjwN3JaZRkBvszsldpHFE7icOhHO7Z
ljp08LOxxpmiSFmMIEV/se7Ad4UZb5LcCmea8mGkxO+ukXBZ+kJeO5+cG9g72GjI
DuEA50fFBMrDPsYQ2a+v2cUn3dFl+cTmaNd/udB/gJzvu17ncRpQJr3fXlZY8CA5
gURMIHh0nPPYSxRroW0efjG8j0Konmesoy4sJ+AitvNcuRKht/6CGlVIoSp5WTlk
KJf3pr7xCE+dMH8H8rSlwi2v5+dK/5f7FyrhWCdQdsFKBXaU9j251S2vA5+M9TeJ
gWokWH7uZ3xV2wZh91mxyLTPsVEkW2Y7r5v3CZwPk27inmWrqXJdmLhAdyS9FOLo
w/PHusPel6Yuk7wdhWPGgqqDLG8yPgYs815JaRH26YAlzjcyELZmDncgjjWwgoPV
I/3LID2M5AiiaSjwtt/fpGAVnjJWL207XetC9J89WzJ1xg2ZCeqhBvuHGxp/Uwk8
EQRWnkOBM2VPMYEfr8CqVaBOaT574hLWwTEokHa81CNQvoS9L/J0evl7EnQLT2bj
K0qZyUKUgL1gaDsiAVpfV3vK6BYPK8MXe9uJd8m/YhdFSMdib0/cZOxifnoWySHh
PUgI5c2e3LlOhOykkYdaG+Uq/ECI4LH5nN73Q5TCEcgp1U1fWk2zV/fYdfv8yZU2
KugEUgJ1xlvZD8FOpowUhrfBR6dC5RYl6RK9z+f01l2Haad2Tcx88VgjazZoILxe
hbz0l0SEHf1b4Trgr7DG5csqq6k3WsCwubNZ9nehjhoiADaxtGKgW8LQoKdPnZiA
De6XkOfSGPM1cU2IX0O0HW0WGd+gMO92MNCmbyCey/OUUW7dswxcAEzzU7TmEblg
uM0yM+a18jVMUVb5TLJPisT3lNNkURG1uxIFsJStC/+sFKMY2Xvmj4undFEt4+9u
A4I6Nd54bOnNA8kjsu+G6QBM9X6a2WJUguIAMY2SpMC2CAvFuOabZVyV7M6LXl4A
t1VZ1J6MHWCW8g8LBwhy5TAFddhGb3IewOQX5o6wW0RJMDUAxEKhQG7JHM2yZRDe
ijv/8aiYVXUY4Nk7G70pZ4gflJhUdkBItrJTOh0qMF2KZjxjPa5JXxIT8w0rzkho
XF0aF9JEf44TLtJmh5ofmk+PeDTtMlRvTNx6BQqKE2WP9NL7Mv8Gqd8uMfEL1coA
eE5VVVoHdN6q+cO6CkXOFDYOO3PkjNDE8TEcSlCjM0aZBqhb5absrDS06ACbZ8JE
DKWtoFH/eU/vxwIb1MHmwCBlDZY5tQK2THYkTQE1ztZDfVHWZjIxWm8qHXi5egJC
FSCBSsYY7e+TB2Oa07ECo3sjPZjH193mp1VHeg9kGlB+lMxT0yiftWSfTzPhv2br
PW7x8FMr5MIPnIhA0d3PsOuOTV/d3UE+Yr9aogwExqeRY6aGZ0EPf/6mC8PzbYuW
H9WDCGgpv/Q5AIcJvJl2ic95tbXroIr3CRbKg/bix9FctNHNcZ9VBkgLm4SSfMIV
lWit2e2gtDMq1mGF7QT7NsVXnHlWJl6lF+LLqtX9BdGHrToZSciv3WXb3V1YT0pD
1dO4CeCt3+T7eqThPmTZQJ7voUwVVFOUs+g+2JXgbjxnKAkyFX0Va8UmMcfiz74d
fVWeJdOJHV1V6QzCVLoGOmnhSa+RQiYdCZ2VCFX0jvTUg0FtxJ0roi6LeAk4y5Gr
NUoSmHtFW4qJmVu8A8DCl1+yJE2nqLZ+xFMYDRF55VGgfzJ5X2QRrjSNm/Up4vvj
r5IcoHecGV4PlJCFjAdd+o2Ii3wt3uBWOptkiprgMCLegfTrMNZcd30RwnuBHfjz
ruHAYRfbfCpBLZy0yB7xJShtsl3XvbPuWnEt7+HzMHnucmwbU4QrKxKm2dCQvuQg
m3LZTxCw23e2k3o70G/5f6DsBTPTPcXjky7ejwKngok=
`protect END_PROTECTED
