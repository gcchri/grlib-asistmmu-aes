`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OKDQ+R38aTqjKem989XLt6RMQQ/f64RLvVD8ibgC4KjpLLGRvbXrr+GGSXl3WzqZ
cKixOLG3w3s5FZ1iavV8I3jSS0D49qRJA7OdbXXHoJ9TGsr/UTtm1CJXOHIqXTAf
Y2W27GYin9UUpPhRfDBwSmK9H02wbTbMrqnjQa6qJXZk1aCwtLqyms5AlNvN/Qwd
YrAy15Pppq364WKSzgN/w4mQctOICfiPfIra8iTPxvdcPr1fnKiTbM4RX/xjaZWH
zLRutaSuwTDRfzucm6cgzxQgPnX/M0OPwmU6suceUuk/EIg/G2o+DdDHgxxVJvo5
gyr6VttZ3Moh+StcOO3bdcZIbGUK1bE+7zw2OeLOprqAgUVEPemmyT3PpdxBVcC4
GFQ1FiQT8WfN4au+1MMxZpMxdPlKdDuAjY0mkG5yO/rjU3me0O1et0V/58mpMTyt
ItkJrsV4IZ7MgjaoHPsmBMEkVKbWlz6YQVn6u7+B4NF6vxNGJ6kNpIXepSQMc8KK
NXkmWHdLOz215a9q3sOhRMVGcT9tN5ju5VycBv0k3lB+LZ4HhJj8tKetjOE/H8iI
wai/5yRw9+HMrIjTd/bfSYdg3UsKf/D4SxUmin27MX8=
`protect END_PROTECTED
