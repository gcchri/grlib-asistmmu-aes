`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MNPHaWR2mBAGBiVGYfaTohqioJDwr4DdvOY39+KkIe0B3WSol5GHJmfG8oxcdIqT
PEQe2Bd8AGXrvg+gZ5AI5125jeyiQUhEcIjpABYmi7qJ7vBW9OxLLhdAWJaJSklI
djl7pxPHwVuv9mdD8qtckeDKTBmIQRcU9H2XIPrE0YDsH8JTocn7ZSo6p50PnlAf
31AEgIjMZxlBBdXi/3uGW6KeUM+Ma0Akdcry6kxM1NR+RvndshsHGiBfBhg9BSO6
qJjnGpdqXwvtyn+Lh/5MiM96MVYVglTMBh1wUCDSUw0h+m2DrXPk97OlU/n8+JgD
8hs3c1LcMZEbZqdgFHCC+LpcarY3BqXgE3ua+X1ycA6yfQSbED+H1ME2esavbCAI
4bieut28qZTQdohjrHPHTcYm3URgrwa+K/0ZAKIk3EXI9/mpkQ0RF2HNIVJTYoA/
QZTHw8xOz0lvf2hSj9HCBnqo0QzL55tZYWLD3472/yhlqcKcgVjHL3guC23HLyc1
39Vv6JppdwA/S0lINSnW5HI/4689RtN75hPczi+egz0=
`protect END_PROTECTED
