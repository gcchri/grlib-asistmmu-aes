`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/PFNYoCZOOnXwwrgdVdYjaUpZKIkvVax71QT/99DqwWB4XxT//8P5ITjuK0FLMR+
+UKVv0bxrGvDVfgTx7B5UrswXm2DGNx0IT7qI3cbVuqlc+sInGy+uG5x79k1C/js
9qqgxJUsm0eTGVcYDLbkD6Kn+vbyHkxToU3gR9/9cxrYPqZXBlakx783NEwy31oq
qA0uZUv6Jefcytb49hWnWYXA3na/l2FlqlZe9mDaMm5S/By5vNGWWFhxIdUqCSQ9
bD6moX2rn6GeT6e99vZssAx6tQ0g5tSRT7VlnsIdcTUW3izc7Qnpd74KmrFIwtL6
OS9E34mqj/TNVOADjGSnsx6CTRv2uWanGFojAubQvqZ1sMDFsZfniJis6SFe/n5+
FiMQcv8yazSooIsg+ixK1LLQWNtcjoSQhCzSc0bSGcY=
`protect END_PROTECTED
