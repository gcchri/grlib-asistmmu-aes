`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GQOQ+b7PYNJ9fP0SMVVGX3sLHIzwKUPG+7FSPO+KZoOzfwda/Di/AdqY+7e7f8Fk
uD0qTQa4B39zAdZrm9KNRleuTP69OvVsoj0BgUpJpvUocA7YHDGz7i5a6whEi1jB
eVXwX5SfHvpfv+o4YPXy6xz1vT6VDU+TMRIt8Nveag8z2DxZqjyEO2LiukOAo19O
BiccI4hUQEJNart22u5sY0TvZeQ5ur5nUJ2TSyvGwKW+Cp4UQMH+BsT/zKN/dgtM
srVuDh5VaU1hThBelg5Wh99PJLbve+gvitMv6yORjtrwwN8daXedTbeQSbTrjN4H
J+xIJ4dPxcPSQMoVjoOg3Z/Of1uwN1WI1JVGP9AKZJ4OKrWkTnNXcUA4yKABqiTp
WdvRboyrKLsjh/XCBVSx++2QZy9ZMrvP1Pv4555lv8v0MYSSAt0MnVuR6nKYodWC
zdp4lHmaYAJ2LJFw19pFFT9JTY0ItBpkpoUicdTKwfYokGMDfJN19F+eIHFUAafv
d5ucCH7PA19CvEogdoSmXOf4nvgrhSRiVXwK/0bAmRO+MCDD5DgpChm3vlc15K5e
3Z3/X7AFsmc2Yv3d3EEX2uCAP3C1ECAOGHSLTa3THQEQw1ZcYTkvOorYnsgm7TOS
ZHl7bZvxVEHDrdxtAPiXM/Og1dywp9pFxE6RqbpW6YW11o9l8b8/T7M0sypHrHX1
Bf9nXZIsycVnM7fvTSXxgZ4USoUpHkcrKjO3auuk//eCTyJ77LgIa9MTrU+s8wIL
w3lryuuL3/6XcllTb4ooMg==
`protect END_PROTECTED
