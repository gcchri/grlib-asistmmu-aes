`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P7tzgiE5HsjnE8dDdj+Y2PJgQQmLLRJy+jkmi8gmyyYTVNfXJ5vT4UAfaVakfRUL
vtX951ZfeCiK2gCtiVBFBK2y4mZxydn07Q80O7tAw6dgzyraDIz3T43dJQaRgOZK
M1wuIKfYE9Mx6YUTFxr/WXe13bPtB+a0VTwQTNxjGMjrdj9T9/+vHJl9WzSVBApv
rSgpKpZLFVxiPU5TdHRgSGhC63+rql0FCTtU5wdZ1vykHtaU1gl7biVbSwq1LDBP
dFZrVFwNpqcjq0Kj68BUtNQSE2bVHnRM+vWh1n64u/vUZDggoubv3Lqwxh84Fx7I
29PROxqB4KJPohrx0m3mpNE4xgAkaNbvHLK5SIEDR+18DmW/RjBdwopAoDcsPAZ2
jxwqZoHJf2WhGD4qKuO/FKbSKgMASQiBzY9DDsDk5WKC39/axWcf6jc+/KBoyh+p
wTuKQDsKRfgLXHsUNQo1EHlSdEXhL+5LSbUs9/ndSP1aJijN5vxVuyKZ779ovB5s
lOsfVMicLjq93BhNXxViLp/BJzKnw+30o8aCLRIrl/4vrm2GLgcMgX+DcQmtK9QF
WW6fBtolfdHYA3gFH7xC11IEZorY3JJwpcPOyjeT4JWiSVj95CQaEnVCkRBewl/Y
+Pww8czJ2nUnM4f2Kv8CA8qd98pUg7Ytt+8x8XcJFB4uKn9bto//LnUZ7mdAlXXM
vTLiDS3ZadgiovQiAD/OUDvf/Bk25LWGyFfN8PCRJY2CnyqjP/Z18awj+RqhpCrz
EdYVq3V4BU/O8GCmf8tuIA==
`protect END_PROTECTED
