`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MGL6aU8KMMNLbHMWaFZArCKc+BAfB5Rid8f32NyrUyM4ejxXzdaJB7eO7n8JFiZK
vjUrJatsslDsBRGJVoK0ybcSXUG3ZjXJMI+5/Yl/Ny2hdxxNxSNqY6oyt/EsSBTe
IADNPQ6BN49jMhQ2I6ZvaThdgq//ATRkR/P8l5DSh+H7+PPss5Xmpa1NGfYb2Daq
VHUCrJW8T0GC6ySr7yd5xfdZf95++2MUZGhrsKOajCTAgk0s7X+OZTYYSeiqRyeE
AGqX+3TuSy6tUBYUqAYJkwT0jtYZN+UtY1NEoBa6YFaYxFxoo7MXlZbrBgaYN/o6
ySZmfMSEyOtIUvDurXg67HbLCpR9tlBpHNyXAdV8J8tjvyus7Y79Oh6jM+O/rlmL
VtrXin+wAn3nSFqaat+t57Av6c00A25ZcDPOjb5Gdf7LLTPsko7U94aU8fpTxymO
DRF/muhs5iSd8roBlHoSlndLBnDpjkwVECIqLCLp4Z/FimMMBa+7f24M/Qz90/NU
+h98vXbW+9rw5Fy4eSKNwk1e4x44fShuBu8HbdAdTdxQOggVLz/q7Q/mGohet840
vMr70QaGE6Gi1cjqKV68XFYXCcuqbwYLjzFtLQG9pmn2goaIkV46BHgPXCGzdzAQ
OJjqhY3fPNe2KuvszAuMBZB28Tj4tzDLEMOjYtkcWvizeJyUU3yAGt480vuzFSuG
DPP+iEtINssu3565jCfk173NC4AxIP9BH/6OyN6ioye/sKk3GJ0qRbMVf8E3pzup
jBuhMxiaHkRtljB85bndJtcq9vvx7r2ai+oE2Feqh7DSn9x6n/3w2ecGtqdCrQ0W
LHMWwHSTsihTxUJTJPqPINivMdWaYsYczTYXuvXAsdN2ZZ3yqLKSAkOotoHpmUeN
4e/5NBZu6Hsv4at78ySN7ilYqlNNgni9IdF6cKHrFesuox7PtwYnHe0yb/ym+25Q
wEMfJVrxcHRB4EUbfoNyPiMptpUGJem2LHj5j3S9BazqN2PUNFAHcnHU6yQ3qIpZ
2ZNK32OlKbyE12hvk2WhjA==
`protect END_PROTECTED
