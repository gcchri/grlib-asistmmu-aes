`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3bkuCJFUhpyROXH2RXXfo/QXX18JWdLEEg5q7oTDVlDZTeDptboB0idbscpTfUs9
YkUzhHCwwsOSTJ8AngBcSUjBNya3CK29egkJKkTS+QY6GqmSTQKB5mPIGbbIuMmq
GztwEVb5wdloF7gGXjgpbht5vDzUSvw2FL2EvFDpFfAMxcXMNFumyhkYvQbda0bU
Z8Z2OORyhLqeLE/QOTn8Rg5yWQ1YJ1oLwjXezHKOL+AhxLEXwNZ63rxfnVecLatz
pr9Jn8lO2WQ/mcGySdpa4UUuMKTc7f7MtZ6OtRVwDNvfgKoWZBRX+/3bOfPtqN0f
+xl6CI/tshl9vtiHt0NjF+natWmSQDlZp+t8/atZZiPJ8/QM2sGW5ENe/74wFpwd
E36G5SY1QSh9dxgdFmSpBJeWC1RaTpvYN4aAMtNf7iZcmE44eQ+J84wR2hf2IXAt
uyh+uwIwnl0UGP2Ra7oaQNUhnclu+bFpG71Hn2RwhfhXIcbp/IKjuqGtAMUbRksi
AgDvp6gg02JP1pR/fowbCjWSlUX+rlkZ519D1v8LgmWQkGv9hGjFgxTqi0Pj1Rzt
9mCJFUInxjIwvtla+igNN2hRK27nTlXBX4V1iQFBsR9PMLoDTsPYhEmA9xN0upu2
MvUqYJQpOX6F9Cq9Q6rN9dBh2zp3LXdVAPG6ecryCoGTQnBbmdVjGB6kEhbcvbkZ
yycFQ2LXAVlQqLhrgTzSmYlos5X3gNVOFL5jfH7ersCek7vyxorJEgLeDaD0MZV7
amcoJ8TNaRQS4LDt6AUocAO83xyUeSJd3DUzY5JB50y6Ts2sOfRHFT2A1WTH6UKq
8yO3INHVgAUVB/DqN70RYBKkZYM44ZCk6Bbog4IKJFGkLA8Q5v8RilkQALq22TBP
W4uIjTkdYOZcGMB3q/xmiu6583/L/pDzPbQa6oJ+AoOwqtruLdF8wbdvCPaEV+9A
WasLlgOoeMSZvBel+Ww6mr8qP8lTldcAYWv154baUHOcvyMiy/nUVu7XiHWEGD0M
wpSp2mlJg4aW4QU3Fg4i8G8wQTDEc+3B6raTi3/pilMrFht8/RA41heMUroprcUF
KHIV9CVynnCXKsW8/oCd/OYIlWzaxMDSEUxrG4ETH7re7GtdndZm/mtTJF28PxLq
XeNO5my9/5zXAi2GX2c3wxQYYsBYPd/QV914bv2iluy6a7HHpEY2YHkmmW0ITQEm
uBJU7ECHYoUXL0CMXPoIWaSSnU9Y9ZqSj2iK58Q8wn6yqykwX+ZnkflCmIruNymn
4EX8FSHkvfsn0KnMLzN+/KRVS77gTxAMFXttS5lP9ofYJHKlY5LdbvAw8no91Q/N
o1DzqgcJF16TPG63CMOEqx25CPXWBJ5xV1/0aafmVR3PEwDiFarTbGCJusaEY7qm
rSAf7NYykfR5yQX8tw6/SUD50UFGkNs2nkQlAOF5b6koXE/Uy0MqQV9i0S+1/GW6
+8ZuecYg64ohfS7uC2NPzr+cc+9BNS1iXvsbXAWlj7nLFy2P0dKTy3tcrLjSb9iv
yFz6gH8TufTvuVBnzUBL13BxrUqLvj6meWiMEyOLeg8LQoxo1efrssT9Sy6Cqu7Q
IXI94O5hGvx6OYVbGwofY2oLQMf7IJ2uVUCwhFEtMRZIwRCy4Id7FjHNQiaOm+5o
Y5zezTFcHdCgh9Eq4RG15Fb1a6Ivrhk9sENeyu4L4p5wkEQ5UyDfG3STTwgnmTwg
ZOaPsXEi1bjl7jk+fbCu/QoLR+sbP2A6PlYY9J+mloOiSDLdwqoF7l3B3ev58fqk
1Q2tlS9iYhBL8hCzfBz5B7b4oZgEoz+msADOcvGqimL8VxbSM99WW/EpqTSDQ1MI
loBGPhhFdsRgw8YgyIYun4HX+AVIICa0VBHE2aKbCXlC7ED6GjVcwTZEvf5We7Ea
Em5auZ8ksrmzSU9ASQ5SVjKp0r9xJzDdaOecbc4OWEZdmOUWfenPeAY1ljT6ieoX
yUJKt2X/KHsVrJj9pgiFgZNV6/YMsLu19laLekNrUzT/xUQ8QLTf4i8q/5by6zq3
S4yA2IZUy39PDK6PQ5VgR3RuSGkZmog/NIPAfMP60OqkDa1aVfEP2eb21FUOCplP
NpORKUQyeDohWjYumfb75BXWpxpm5cYSpO2esmDXtybet0tFPYRcONEvQYYU3+Xd
yIsN07AAy1ELhSk04xsJCBJY5tbVYcBb/MyDrN1UkbbNk03Ww0ZQqQToH1i7puZE
6IMYWXhCMbjwlrnp2A6YWl+BiTS/y/uO0Xnfy4i6uptRVnhfTGsw5yHspReojqWC
IgWGyRGeTFlOamgxpzQOiDIhe0aVq2emINWzRF95ubmk/GBmT+6Up8EK7nU6I6Er
+C+daeiHfjulVw2Xkfpw+wem77ry3CENEdwu38V3qZtst8HBHzqFrrTgz9qaQkj9
SaUGb8Diu8lMvXWdRz77PtSU2QmbS2dDGYtL3qnDE1mAcSjoeSiT5EY8zEMSXXOp
Q5pDcuCyQ93qEDSuG4/8mplhy+FrITfSqKQgpcNmc98tGZqeuS1LYIvN0294VV8F
uA+jxHVmi+f0EF4310LJxjIs4sAjceRNKdyTwme7g3PcG7emboBQ7ZZULyCe75iA
JpNs29qwnXYPtFbNsjvRnILAB175S9TI2e/yH+fk+6RCJ27zyAcvISZU+1EAXSGd
kNqw/afQ6G2rPqFek2e0kbWLQgx/Dn0PUyMgBet2gNECVAxp7OkE7F5eCd/F5Vpv
410/0rwanj6GNu/rccqur/0zgv7kFlNfcGp7136cH9AwrVfsN1PgGk7UFmONHDg6
5j5s3XgXFdwp167fXqaUDniXO16V3byFGXOnrMKmGOnVt9VE5cg8xtru0VUpLfMZ
B5ZWtyl6D4uM2Een8w0AaYUXLokHkbwBt0eZcZ3dOM5O6JzNUlAflDlP3vIuOWqC
FiGOOUjRmRMCPl2u7+jSyftK7+HjGff10CiQeyw7EurALCFreIfSa4MgMmAOCy6N
g1p6GnuyM5Hv8rSO8J/reyctd3z99/NEr4Zg8g6QAhA+qnKZFvdi94riqYvbx3Dl
hwepd1I2/gIJg5SbiodjZ1/d3PzoqUymB3UQYNStskN29BjoIOormwIjGl+TE2aZ
H0FaloSdaWiaEIKQ/bCDOmsf5+rCmBql4pS8TKbHjtcpo7IqALOpiQaeZ3jzarz3
WTn7yMVJYlZpJ4yAeKkV6m+iPF0RSfQg/AIjOSPd37UqPfn3mwsCGMe7tdS+n4Z3
bKiMsVLBdL8DPa+ENB6U3EB0ML0/FXx9EEQglkSVf9+PLmGEL/uogOV9KrFlth8d
fTdgyl0tBxlsJFEYGXb3O7sjhEHPo/j1gqhlIvsZXu7DHxq5uA21cCzCxuCKLa/N
iUQrXAnAJ+FcdK6or6oiPy8Tv08FCPi26QWc+HjaNDrEIbU760XB+1vjYbqWaWCn
b2Iou/aaxcFQJm5yc0gu1CjwMC2MsLXoOaawHzZtIXzxkGtaCqWrnIuPviqljJpe
9jK+ZGWLqSBZ/m7sRqY+rUYk49zSgsGJWF4+lUAxZMv7i5ldUsGnBDvH8ZLCWlH3
9EQ105/hvxOtXgftz05LhVdnwxllKYuKACFS8hyVSvhWhgcI9Ic3kMQJenDUbdI1
+3GOh8BXnpZTtqPelJ8MMd14Ta93M9mPdTHR08vFYyJM6dThUgc96x9H3bsSFWfc
5PF/BwZ09J0UWUv//ZGp5q2qesFqhRnmTidfKRxbUrrjqUhBUWhROo5bGAVaVafE
E0efI980w2jpMfNQ41K4kRBEz4tDyO6iKIMkW6UhKW5t65pNPr+NcmPBWBisKtAz
twGo849RNH4cpvw/Eh2N989tV/osDrHeGCkBHndsIAnMAryl9cbn9vMshlY0KInT
qDscNI0i87emATMIrP2aQCr74bvcSe9hbthWt9tCxeTHJpQcdGWOAIVzF9Yhi8oW
2jFNkhy/dkqnlE8/7Y0NSk6LSh6F0igh/M6ZU7I+dT1ubHWR02G0sY8HK2tOLid7
l9mxgH+5V0vNj6dR1EO82oWv6yJIoHjWQ9NT7MGQJHMMWjFGKMHbKwuNXwyQ7Jbh
nhbqP02hEpk4tr5SJraHhHYNdjxMCHkyOHMzrYxVgTF8v3xu8jPkxioGsB5akNrA
YYnby/xLd15zTJqLQg2Y3kft0WsR8HZHKGCTlhgfjHBk9dYiFf4qra9i1ajRL4U3
2Hd8wGFlpJS6A3nnLiHmpclpvb1xM7Qw2zm3q+gL1npowixjCZy485pZ45QjMQbI
MzU4Sz8gRlMUF7CeKgyxRNySbBKR8ROBDCtXvzF9WLL7UCT2LLLpDYd0CUT1KLra
cEvGakdyVibtEOHeEtOCtCguR4eHfyY9T23HuKUPi/4YHcLGaxHe4VaymDCi4SoO
6o4f7+jaF3jNFX7yjmSSJOq4zmAbvU1eyCj0e9FZKuB/Aiy4lViAczLsb8tTYWhV
rXCuNZdu8B1Cvpyv8A9ri/5qOVAgve3KxmUA+vm56Y79NwNjYSnYmVLGB8GnOU25
Lp2asZ0sYujgOH4UB2TS48dDZnvrdsLHMHoOE9usGQJrwZvAmcqOfqg7U8yev0P3
NmHjjn4xdR51C/ZAaieboNhSO+d5V5pR8W4Yt6abxc0yrf4RU7Ix4/250CVH85Z3
hk+hkkJ60oUkkgFPXHH6kS9s5NP1C5LlVbpX2Rh/qAlxwnnXGedAPJswuhP7kvpi
uDsRba0Y1uX1OmF1Vk4rUj0Xx+fty4Z2khKTB7KU8WsNbPkW/LJEvlwBuAkbd8DB
JhDyFTSkjTXugZ+M/Q7bqIFCjlEe60GR8gpmkuQKQ8uOoayUHSRlQX8fxobUFyJ0
CGFneAz5wDnGnEFWdw1ogaTDSn++PbrtQbf3ZJxGePC7aoB0jKtTbvc0UayRqkZ4
nVRmy9yc6yM9HcdyStnhWhGcQ95/ivwyN+oAsYoZFJrL+Ck0ys2u4Nu4sDsvZQll
A1Wha6W7adu5XjsXLTRLOZYhY+qUAC35ZGScLLhqnpYHIUsMb5ih3Mm9spJO+xwA
S7t6Xwp05IThnbITgisc2hNwzAZmXAbUwXiVxtHTWWVpNtb9N9lHuosX12O7Bmpv
tULonwQgf0B7wuSPFSevTDfUCvJ8o36xs6T3h32hBJzbi4HyvyGkpMkIg36/xift
jtGv8TuM6YNbgXymN/+zKvZV3zoNugnUXNw3CqBkKZBQh5MaRhMs0Z3n0NLegC+4
ch2JN96/cwHehOfJS/hF8UXzXEnSAGguGqa+0M1sY3JDUS59N9P9cdV35n2gjVID
gwcr1vgSMlOkecswbj3Mpfpi1UuyggSzy34TTWVXMb2+etlkdtzmxzISkl4CP134
i+dphJX0PgzfefNBU/YhzWzvSaqj80nycLL3eTUoYcNmytmWH27iwBv5HP6upy8n
aaKWhzFZ/aZkADWrIm9om4QAf8GS0IncxxbDdX4D8766MUbwmw9Q/pqFHOut5Sf0
h6cDFmJS3npjZtqO2IZF87pcY1+46dPZbAgS9ALAL8CeV6WhFka8a74NjFjoWCps
uTmcokf3m4yzRk4eeT5W5UQpgmWAMnk0+brDvZjFWb/SchtTVsiAn5u3RkG2hKLK
9CCizO8foFCgQ0cyUjRmEA1Acc60mZ/ALC0rM9d3/Uw1FGD1c7RDuNN6NXddd4P+
xh99H6naBisP9Awr6xC81k4HZS+/Zcej0+UmMJ8IPLbOi3H8xSx1xAVPNIkf4csu
vEUGbNhzS2oDEeI6O6oAu83Uq/ufzu6DOrY1M9Ub5YbPHnS1u2gKjBabq/2BkbIm
pxZ9lL9ku7qH9OKw/z3aFwZpO3CQqPi7KvNEelOqGdBnruqv3uPfmverR1JDBuFu
Y311GW50G8tuhvjr+3+cFzmXTa8giRgCva684FVkazX1qeernrurRNRs0sLMbPMd
aN55khRPkoeQftVGPC1NodHhFAniWHOtb0hLXMm+0/tq8McJ1E4YUs+seG0pawGx
xBKMrJF81iwhh0FwciBRmWwoZDognarUK4iKlZij5mQH5g5J/LFLeMpD6xDInpGN
k5jD31pjWS/feveQbybu4cIR8I+8QqQoQKms0nonI8kZDr5AKuCQLKl6LOjPvPcQ
Quix7BpWnOox/kZArCZKQI6L1ot6BGuVJFI/BOE8N3/5aK0A0WBvzlJ6uPZHGmgY
0T+4gVOeHT/O5wFg9/gRcJhfrlHaE0jRMKKTzZh735YzcvIOYm0BCmybq9bkPaa9
Jnc+t27hIsUG9AOwRmtlKvgmlCGdKQmwXSsv/DLVMCXd8bZnFW7t21bo+RjHgYY+
LiTByX/fotvWLTSZbLLfrq85grurma/e5RpUXfs3a3EA7UpO5HdUOSjf6AM02Doc
D0xgranNCIWapPAWX6wZCbMIrltEcLZ6VE15cgs4Azaoh9ww29QtEdBt7+i763Qy
3GczU3dWrNsD/0y65rp051MSwPb5321jzOG6aM/oF/21qJNOyEFmVqpFsxKjrSqT
h6TYZv7/89lVJ001YLvpoZbCLPiVOWO/Z4Ud0PJ3SfqacI/pPxA8x7b7jVAxsXh5
oulFtL+aUYU3rZHuoUnZMH3ridIGSpk+YUOvy+KUXE3mzhZ9wme0FytwupGVUStQ
vCzyR+hG1NwMYRejDPYmghPDetb5OpV4hMavR7Qcnh9t4FxEqqRswyCIk2e174kU
reKw+aZBUhVPkimK5Uv6VBk0QvEeX+2SadGHnPa+6GYU/bz5xMX9DSTo97qSpaxL
FDkJVm4psVmF96nLS3NLqe8pmUkGoKB24CaIQaShV6EmBDsArN1KYCu4M+XDJjN2
MX5MmohyKBKLxzZFobyGVPxdpEjjmyKqngSQxKiSGTNKzpm3pgQWW3SmVsTRkO2w
dxNSeknA/bsYjhZELJss71+0XErsSF/2gJn4ty609KJgXXi3pzrwyFd60j1KoAtb
gPqcJcAla3HOgi1LC3NbkhqqO+wSMJYKaUcCMM3w2EjMkImWsPEvpSlMU+665wgw
jmcEpo7JmqcseAuklHaIdQmOEGuysNiKGzahmXrUiXVaMAERnPXzqZNriqxTdt8E
aJvl7/v8ipbrLisGzRyDt64Uzwa2LoG8sAC1EjkEzlBM3WJs0+HmZA0N9KjLlaM5
WbbRlUi0Z54TuwN8m1Rhjlx1g/vTxisx4jBfoH+AcqZLT8y2qygeBODZn48FtA9k
LHuH2+W7Jwp2TF82nijn69NE0fzUMqLG6R+/MZOOKXSlLez4aB9MTj+8zl0FyjMe
PFgJAj/JhxEfsCpUZg2cULZKaacqrFUVU/u06nbyae3NL/qZUZ2O959t66jvBrRe
X+YXX92TeHcbRuEejUbWyYyMuJR1nb2LzVujxMKc2BJihp4BBL+mbe/jnmlz//hI
RqSR4tQWPUDP6IUEeevSxr5s21744v64eS3lUeIK2xDtBoLpAlj08mT5v+12d/1R
WnaFyvwTu5odjsObPFzG6mTQGCN5DQPFM4Uf7VMmU/3YD6+++DMRJdginiigFq1L
xoxUS1sbmzlnNVUGN587RmUGkab3O249a02r/Vnd90P1qrRCBExVDmckO3vUaAGz
Lv7yZPJLtmeoEgUH5MsL33DoHn0ajiHY7CSKV60uTxn8dcrYUifl7yry2mwiCDVH
hmffX07ENHl8y5ApJAM6kUIZiu99LoB1Mw5BsmmjYaCURkHRssHF0y+2O0wn1Yit
lqSvPkAXWRhGGBz5zWf+931hxSLpSHqMHzyC10U7Dzj0q1EDMKmP/IgxFcJuOId6
748kk2Ew1W/SgBNU1nsUxF1cWJTaKYrTKnI9xdiV9C1yhhV6OeUFBlB3qBmtl6Fr
F4lqPD0b1JF6W0HKQIMPOia4fBGovYpAp89dHpcqAWKPTvgPfPBXSsVB+PouBo88
sESPyWMvyoixdIV3jhGFdf8sYlbdZRJgt2aaGDTlU9xL1a9zjU8VLI5GHTnNthJ2
9ODi8Af6d35iN+dJlggYR+w0egphaBSEN1bl3g3y9rcrZ5yOAQ7WZ10++Pwkl7+H
qA3FYapeFnGmtapT4NJ4iGpprHnoMuwBMvxYRECQO0AeVHKs2ve5P1qfoBjq8SZh
c6BPptVHHPygRNg7D4aVo44Wm09FhM/gNP22Gp+O1Cj8xBa5IledVo051ER/dpDe
S6FsY4Jm26dqjLfoYwXnXYJg7HEVrUzhzSualm0gIfcy8PANMZqq3/A+ajJ6STuW
lXHWgwcqSk5w+oo0W57QtZ/Q2AOC2vr/lf7uO/dSJDRyrfqfvukslz3IWoihsEvv
Qtek8Gmb6zEvskca+pr8F0E3OndVvLrP02yrdozqUfbwhwoljma5+Ph7R4usF5l6
lFSS12meGDtpRsL/fRuZGHv9irm2ZQZ4Z0KKNV78wutnTGaKVuvqKvW3lrQGlO1P
HcIwRD/vJ9MFM3jRGEeRocT+zz1tLfOQg5iNDJRfLzpZ2SC8w8XFthNrIRp3Yj4k
r4agUZs2OayumkL8hq7YFt1cmypmM32kV7qgdqU1eXU18J7m77qRmMhE5FOh8Axo
wawHzl8U018dfPdWnIgUbKObUXK23xei9zqOn9Hrk6b8jqWuCvSgh2QJzs8PzrWr
mB5S+fnBSSCMRlZYGBCcjNHxDeEWN7HVS2Hqt4sUz7ROd3agUV3vYoCWocseKS8r
GcnEk1s49kFrKl6r6Km0K6LHAAJMSn+TDWoV3J3j2a//OyG9ZLWcCRBzSQL1waD5
QD4OmJH7TFNNGiDiuWijylPxwBD3p98qBs3FnzAG6CD70GSzDSAkMjYCskPfsw52
kBrxPhSyCPdb7l9wa8Xx8DULHbyfDuR4WgRxe6hqzrkGhYcXSg5P9BsiW29nPP1G
zcg26Zxoz3aRLeM/IDAvqkEXpUET3nYpCKpqG6NJKxv9h0HOdmqhZwQ42S/lwX68
f7ukr0q4HqNW2oEwAc36rGnBNuX/FERJ3De6SX6hPboW7bjXaRyHPYIE9xCRkh7v
KJfgFvwIjt02UgGHGKmHlz7eBWTIFEViGJAjA2L86UDQnr10itS8M5YoUhwRxkBN
g1xg3u9Cag28SWyCBvv6OhemEWOefjE4T2uMZVFaeJACOFVN9p71Wzy17D8ik9NE
J2fqdUc/8hYjOVv57ViTQilOzYjTd+5NNSIk1iqA9ZMqNq5V8NJG3KPVKv52TQb3
OjMUKn3BIk+QAQh79SgAP5wCls3rsNvxPSP3M5U9vZh2kGQBKvnpyNuXw1GeC7P+
DSe7Jgi/i5ffXDtNRNa0MYmav9DPfeny4X16cLl6R/xdlmPYJazKAx7QFi9Q/+85
nfqLlL/iqlzHusUFBiWB3YNDagr1nOsYR6HoHSl+rsqLgQFRj82Jcaa/v+XIYMlK
gP0PHfi5DJj+poH0ol3m2aPam5sFQ0kcHv6LD2gI7e0PF1GB2e29EF6ufRGj9Sza
4TrKVuFQkBdV+Pj6kjmhFG+cvXU4R+Gj6oP+VdIwOSfNbZvhFNpTe6bV+F+ak/Ck
8fJ+OwBS/BfqckraNW5Ofh/eTtteEpzKiF+kWTHAM0OH8uYVa3nyedes2Z4SLpFe
ndqs0SLegRG7sFqTdrph2kCfgqawo7dxkyPCkMYpGwxPKd2v/hITnbmhO5CxRF13
CZKJ4fAvfrZ0WWAoBaD5ceBhMjmAI6a4tMLcW1/mYdaUukyc511tT6aGyZ0vhV8B
PlyqCYPjAqY8vYrztTM/Et9ycMcjbZzfKAxWXclI+KMhm9FzYZUHJBiREi6GVST4
bhoT+SZNVB064a2FeVlqmoA1uC2gJnpMfDg/cUjIqP+NVWQrp6p7qz7hw+ZsWDhu
VQNXxF53vVfgoXNvNBkU/RYjbcv/uUxU3YXVTnMtOGScqcx5J7wUiptsDnaOOtpj
tT3O5jQub1bBbaMyidJ/qiB6AXMj5P6grhQk0eRdrfAMQeSvIIaEYN8OdyfvGq9Q
N/ObK5WdBTt5QTQzFkA0HFJo5gdvkxpc3+BCH4Mf0qDXvdcrMVc0sIoNlHCkpNZ7
iK7q7Zq0pDyE84CQmKjnSGpS2J++TQ04a7viYaAd6owymIgLr+ie0kYDFJ2YRHhe
aKsx/167/Vi3v/EkoBwHcDkxwB8DNXLjSwYxGs65qhWIi/Eh7rf4ftMtqE+wP1mX
d+9DQMBDYJLO2PlkSalMyq/COHjspp5uJMg7kLJC0sMCzaTZvHkqwaDV70NMVOwR
J8zjZ/C2dNcF7CnmAr+IE37KQm+jF8hQ6V5NlFH10tclFYeunstD2c4OYUiWet4x
GMLYhWfdzqBHwv/BaqgrK6AjCdqEvpUGZX4t+WQj1RgZXxUVUsq48JJhmQ1K04Y3
VjhyY+NWPAXq001lnqDP/T8ZXVarEHQgpiXVZ1uQGCO9aHlBBM9u3F3/ZENrfBIf
LH7W8lxxpmaYJiEL8bdeC0idey9NrQ5ySVZhbXUoqKQihqEaLziokTgtvRyEqwHw
Pl4bJyt2H8QEud07X+iZGxj5rE50S5StkOmbNGcgc4VJ/xyO7zN4uXKYJ6TpEKvp
6EyuBEBvWAmskoEmICW1EMd4XSmdr7iErgN85Hzo6xsbYhBd+wgMt44HUdVC9GPx
WBP8e6lv2KSZ/GYXUmS57eFtAIHKxu/flYvK1byEaN/zSXkFdlvjGb0zSD5GAcLi
tK7Hd8K0cr45jaLEbtpR7azjrKij5P1pGEyoNwsrBc0a7PheurIC5xwLhdZyeu4/
E2cGtqAgco2O6cOuaGYtupV4MOI5UFp6za+3igmKyXH//i3FqEJzLmWSts23lh1m
i8G9D4wgvH4FBkpmjxjXjHh56VrdMpNSSCjLTxt/c/fa0pmM9px1y22dllfmXlDD
FacKA8rXgyiEN9kJKXYfP7bPL178Fp2PIbFgN2f5Y+UjFYfI66rBl6yD7LjgzXV5
7CqVNdscu8AjytSmQafXnfYlBSidANAyIxYGhK6z3Znq98u8MbiBW0SggC/KUGdj
aSl4SLNApNjAWb+/Fma7srlQg8scjM7Y4boBpW/n7iEvXplZ10OOiTFtdhez5W9B
qxoTwTUiBriGPmkyEE4JqWwzn6f+KwvGoE/bd5iLwkuBTDZ2f6Ait6RAIFiLria2
xZN7g1atSAT5kuzzfDf9O8f9ZOZOzAkUVGe4NygwTewjwN9aFFFrSSsOsVf+Be6R
RtI2taFqdZs8quPJuJ9DyEHkS8FQSYS1J+emF3lKINAqpdaFkNJFGivXL2DUPuEi
O2+26pai4sxGNz02IWbRD4eDtXBgAk7PQwgAgLdxRgc1Qaf3lBwXMahf0ncYFDnY
F8viPq2o8qCLLN9Uk7u2Nx2+0ScjIXHvaJAdlSQrDrv/1us3pG1PRy3khklav8R5
6thoLAL7/jDzWd61kG6ATVLk90vE7aI86roYcH4/bKN5Xx/uNhJjcJu4J5oFd7RO
PEbCEVNQM8JomrOY35CnAmfolP8knundD6z73UVzowOa7q7xkh0OW/U+Zyij0qyH
Xd5STothwoatHen234vfE8dO30t4sM+U4mqoAIc7BMURP609xaNlW8WCN5fQ1Mt9
pWMMsnkD8AfJxw5oMg9GeQwqi5V/fulCGeEaT1rGmmZ4Aestr+UfMj5tifU6f8NT
sQc2IgbH2Ekm8VB04BrdppGdnR7Dt4chwa+jKy0S8vgxxVSYo6rdrixoji/covw6
Z72f78llBugLuHR0wYvmKDm4vLxMQ6R3IW1QesoOI4WdA4Y3Vg/MuWa+lkaLSaFz
Fa8/QTSouxHmDsPChRoELkFQKAMfMcGsUkvqeFgafnq4vp1dxFciufTpDAHxURKg
GoseHyF75C0w171YnDi21go0cOP4ajMyhN/WQhbRYZLf/yJdhwGXkiitlc//Gspb
kRrQ5go8tC1KmcSBrLfm7iMWxOczz57MpVkMiy9yJbIhasVJD5cW+vMqDmfUG79Z
DWxtP9ml5ks3lJyJ8qJAKMPryKt39vXsQVyFPpbN8glN8IetOmY8e7AdL8DH9g+b
6WAEoHTNn6kV3NWHe80giEPeNAEBPtM88cj9/omCdGiuHj/M+2GaCiGwtl8UfGp4
YVmyJK7y2PP6ipCStBEAs3opqjf5OuG2xQidnzOXuiguyxRWSC+/wAZCAt3gxKA1
UeWUni3Hdy+DSYu6zEgWOmlW+EBkFF0Sj45zV5Q/OYqBjLrZTkIbHrntTPvcNQmh
59zaRsovQFty50z/M3VZrvuayiecoNVZ0rqwim0PE21zpC2uOqn1GjmBIENtKaYS
RdvUJFbl0NMakxNg40pXrk8EwxyzYeiNu8cJXryMo3bXZSANvqjd0/q/LVivce/r
BG21cAOuJJTo2yCKSAvtH2ohbZsb18Y/eRE9w4M4/AGfmCMlr8CpccUwUJ8CU6Gr
XgGgVafvvOwBcWSlzgHB4MCDLBlnhaES0HRwUcONk7GANbXjQ0VsS0b6t6MWki0g
JfT6KAMnL2TIOUGGmQ4bV7A60eZb/09C8gwxjKs13rN+3Hjlbqi+nJ9hDTd7aNZt
+EbP+EWYPPTNNzBjlU/AgQtBpUPGU5yEIxAa5zlPwhYKgiN+SfQFKtjCn/tffO8h
va925mMdikP5WxTC++esspNrRLDeQDYvRPEo6d7090X8gZN4wLadibVyaq7XgWLG
PCxYJCrpcxo6yMJMtOz6bLaSm2kwDeG5mAEWGdrMSHJmKsp0xgX6dQcnzH9UZJve
jkR6QIaPP8M2Q2lE5p0Lz2U71rYgApwpscybXcrHjTD3BnCdD56AxdZJuXHOXpBP
Hh7KrERn4PbCy1sxYXmTAxbjpvtqK+o0pBB1a7mxUeGWuzFqTmlstISPkJDr9/yi
h4RUJacrjzHdl1XdlnFIfns/SJGpShfRPzf5BSd/WeKv7VR2xb6JzFzDKS1/W0XE
VHPmw294VRc9GuWlkRcaM9HqaF8V9VA9Xj0hhElhdXEBHu5QbQ0Fvg+HqqNP9JMz
Kavob9YBaMyeeGyuZflRaA5ChJCUUUOH3AN8Kg+VwlwoaYFGGJyG4OjyQoVd+yNf
qBj2qywZA3iJbu4myxn7v23k6Jrc0qAWWivV+Rix+1FfWm3HvNQef13ZMMcAYS++
g0ZefSdm3fhgZ+gBz7YTghrWdnOpgwzMPPWXsCek25s5HKdPdd/XIKJKcAu4V6c9
Lv9lceV1lYlpQhZC24PgcGJSQHeX4xRahwrSURCUSDCCV99Eq7i9NAfxhYgxo4ez
b+RbSpm3WiBOB4oYC00E9pDqUZjLRjp49ASgbwYG7XPyJn0dOrq0KctQrEKSSGD7
/1jgn0pzWwtiTaFifmtJLwSU8mAUO1iyF5zrEY73BETvsWqbIRdbYcRfaJ9ZgTwj
mnRCzXVUyegu+Cwqt/fTCjVblPdZIDt/g23fHTELIdJ1okufvDmLPOFGYm//mWkJ
gCwWaheqv00rMfHKLGo0B+3lW3ePJL+aQre+qXaipiWOob5p4ubrE4zOJuIN0Roa
xtrQgDhO0d+LssOBPZKXBY0P4yvmK2HsH8YHiUumWoMp8hmg6Y/lOBP4TUjzWJWP
eAZlax3GUqaDyp7CtbzI1fNz/LSzWU721PdXp/4bQ9jryVqwdqGGz/qnqaN7hydZ
pItu3vluZoVke+7TTNEuA78YfRTH5bwG2qzN4wREcn/x1vCLuZc1arw52HRjXdGF
sE5Lw7DVzXWEV4O70aPA49JlDImk+sU/fTA405g8S6bZ5NAqTcxvOCkpcakL3tpj
HlacuhPsLd+FY7vrPu+d3m7t9aZiIkO4nF0Q9RydcEv2uCue+NJ/BWdu9WrHhzwi
mBmCGx4FrX2gf1plaNPBaTwBMJnqVo1M6YzZLw6K2esZRy90HbjWNfwTQorplAnM
VTngsoJTsTmaW8vUeaO0WZG3GgxbddnT1h2PIFTFtdyfrdu5tRPEGs/V3AF1YaP5
HQr/PusO5Z4QxKHbfRGq1+Z5hS/Oojb3ruHn0+OBo5t3mSr5mCh1OHVwxMPfcHB0
ONUbrUFS2XdJlHM7Kpcg51lHMjP1411wZJC3bwU8/KNJd0LVrKm8zdXyq9AeUZ7P
BophTDYQvlLqAYAyzN7cqNtWgHeAkcZl0yZpO4UUYn9X4k5EMRkkHj+aZgWLjVWF
ZewLDzrgnBXVJNvuP9fPWLl1rRTOyXxCpM0s1GnnwTGi6FP8Wl6+ZZKj0QXPxlLw
Z6ty/JjWWZmdp0JsDWJY3MGMdSeEb3BvPndB8qxvav0PVwAuzv+s7Ohw97CoF50E
tr19lLBSU5AG6IvJ8rx3lBcycyu1pvzClIe0/Zi+5ft36Ru7Nrl5XaxZzTZI4Nof
wyYeZ+wf+vRYda8oRgzbF5c189n7q0o1pb4aPXoqlYxXjxGGc+4Q7fLQ0FMC/ukQ
qoXIAvcAdqCEzFBzcf6SVMBsLc8rBteP2T4q9mVpTkFre2GOKEmayRyV/9BHR20A
kkXBWZXfR37yyv80z1lJv3hMImhkZEWR3LrJCb9W8s5wGFo9RDca9X/4I8PNJaAt
V4oihvz50KCmSX/oT/17IiuoE5JF9+PdfL7vU5ljj/m7TmFel/PyVx1WXdfzoyLB
8yO0jVloP+CcedXweTYL4e5LmolSEFoj8GHE3bp+bkuWYLAor975o9EfwkWsvTcf
pEt9CiJMEYegPIoQX7jGohpwku4CBaXpebId4K8QScDgkdOIDgdWql13psVDaGll
U1w5su6ojhM1evNIbDkwgGPH/xc5NkrHHv60fACK+qXm3d62MtsjhJAV7laIuSjz
fS2XFaFHXp6QjZRmaKSClxYaIxDgTJMmPnmdf876SYeCyklYsxGESLJWtT+wxprY
Li9YtV9vQhJtnKmAXipnUPaQEQY7en14nmg5Vsegg3S2bYSuefPoqMK0fdBnHgpb
Ai3hqn2wzyqAYhTrxo16uu5KgjB+mpSsg9qwvHThfJPg2gIEA342TpjQq+tf7x4S
+CGtqtyoJ5RhPTqK9hye23MMD9os4kZg72Iw2ilTdCMcAhiMmoYIoRypoOhVjfJR
aySIxFDaNxSZOKEymda/ZmDj9y0fLwyQ246maJEdtBgmGZlLQSFI7RLxxiMa+WXZ
Yo5PTE5px8gMMM7tAGlD+c9yhBQcyYEimSJa4Y40gMnia1Szh6nvXmP4uuPjctEN
JveJRkoyDE1EqVqjoo0cyghRe2hzVXm+NC34SeEAnl8WO+mM1OHFFYiWg0H0nWzJ
2PYvJDWJAwNo/SzZNaUGGMpSauW+SMISu71zCUbxj6V4G1zAx0JZymlJzyFIQ3+F
nmAIhEPwtQGD2GrjmaNGnp9X8NosS/XvhEJhrlTkrc1xT+/K7ktjjRvEXbajP/Fl
kIrv1hEcun1GxRx3KHGHEsLFNjTEPGjsg4i+HENImzlGF5wKxukRlopl55vrhN8f
ygUgVAItzjFKMe33L9ttCLIfygpy07uLcl06ix6g7T+4djlfhuqsMlMfZzadhJU9
XwcDqZr+/uwUQr6MAOnZn6HLFGheOPJWVAD7OYrjkEMOvnPYHKlo0Yh0ZGScKFIG
C0i25MctzKPyQikOBybYrXvN/4RTf45IEQzAagOIkWL0vPaOErbKMApu8VnhUxIk
7PrbTxG7WP3TNQGVUH2iF3vlD0V8FK0Zed9g0A74AwnK/S4x0D6MHbZjcto8jM8t
seN5jJfNsRQCxmOoLaDf00BLCGG3H4mUlin/PBCKhnYI9PYU/b7cMeBwE0uTZIy4
x7T0Gjug+SJzrWn1wpUH6bJ5xKezOXkv8CNsQM9QK6t7ySio792JFx8LVpYpQe6S
WW/pI6jg8PQVSTNF+1HycVhQaUhzo0HZRCI8Dk5RgC9veeQ9FT73OgHkoDZHozmS
obmAQhDJvvFgavTqPYQLcCzSUDdIIuwOFgFMHqW+SdL7rA76a5Q0fejBzWQl1qWN
6AnfUa/U0klIHlb/l7e9K+NHs3W1Yxy3C1OdrCC54nPCRkFe0FKpq4K2d5B+ztIE
dQcAgu8TC2m858KiY1urr0DjnL3H6MooRcXoaK1eLUUL+1WXbwrwTmqLatSQiJ88
UBod/0sbJMw5BeOuJpOBLCDDmDxcLU34M+M2JZ031CH52xcGpOmlyffP9aTs50vc
6dNwi0MaoIvrln1zGnzrdt+Xq4rACOkON1rNaRmav0A0VUzVhsO4R7X0t/Qe9TYn
d3mBqc2/l2bZRj81JemvVRb0VjgL+vhRHJ7OgxcvgNOyE1CDKKH4nm/HDWVVBk6f
nDJQb6j4zIx1k4dtUR2usI76qs3qtK26FSa1yWwwtMx7yY+3D6Gviomo/2QWn7gM
xEFUToVBq6yjebTSMn7YnPBl927T8zBgpG0gl79WCQYmwTwUAttUYTVBZOvFwkzQ
MWSpDY2oUhyWo4X06lv5UDnfjNRmOukDqunCkN/fgBgUnekjcDDEjXGuJ3e1yURY
Cqk8XWxYZb5i03SvbZ4CUs90lI1PrlbB+JzWfZj/XBP6K/24hDsi8dWeSa51iDKx
b+mN6HvVg2h2vuQB+AVPnNnJ8eb+nRC1EWGiMFFCCdr7DjmVXYYq79t7HQSBND8t
NGLq9t7rLnEpCDxadC3dnEtKeiEfcQ4xy2YhR5RBhE/Y6y3W57E0F6GtRnHY4MAh
l2NwXmjFbE0FU9q0r2jLCFf2ZCXk2DVrPJW/MknH9ONrPAxENpZ2AsqojOlDfWmm
gbYIvn2vvRRQ/jbR3rPTTosFTMfhCVDvE8jP9Q27DTtlMYd84TVoVkX4aGrUXvyy
BQaBBSne/9GI/x3gMmxIqU6GJemMeDtVMqWRkcnigYEsVMcHJXqBQ/ClQ6W0lq54
fBnFVjrQW4UBSOKg3r1jyB1pUbISrXMTw9J2cPkSAoLcAcZqE3rkcTZ9cQkTr+zI
1bSeRP8lcSV1kZ0NhmZV3BJQHW6ZkMM9gM6y3nCJfnVAgCwJTiZr/RWVIY94Lz4k
Yh8iJEMh6xMB4C6ADx0vgtdj3wHW/LygbApqAmc1pN6iykpo+7/hLaOzHktFFPzh
tglgO5mnl63WqnrqEzX9jDDf4VpbsGgzgiV9mSB4CCrqk8tyPWOSZXeMYjdlJrZC
ViYiSoWFpnIedizoy717Ph8NrsfDp9EQnKbPE2forD1f+K5qJwLGQKkzwMxYnZwS
6zrpua7ukuCobIv6yTFPDI19YQ0TQIlxigsoM1FSrYknF9LVdJg7zZoy695zeNPb
4iuez/fb5ytsnCU44WCMB+5qKzd1mvnfZOaL9UJfULoiCvf32HdW/J8f54wjrAga
FiAl3428lc2iKUHNf0z4d+MF7CLifAMVP2xRtstCuv8h12qg1c7K14UvFal68+DQ
ahXyxz74nLzUDfF6nliljKGYkyc7r0R6Cyzvcp5S3I1QWO6I5AQV3GbRmzsdXPyh
HzwomqaHB8kMPE9vATCrbfAJ6/r3s52Y8ArjhbwXVJWeF02ZN0m1jLkp6ZhbLU/A
iU8OlvWYNz455oLix0P9+cduqODtqkvKUuA+Vt5Dgyf3ayzgj3vakpztC+PaWp5j
NArTOvRtYIb2bdHYWf4VJJa1csQpqUZ5eg+CBTqtH4gcWthp7Ydm3JGwhVSztf6s
S28Hhg8X29YFlIPD+9QjmOlgiqnmRO0y7JuSdm5c8hDQKnelzxQk9P/glC5kmob5
dAAOGcwKYprO6ADYsIxA40bNH4QVNqA7g+iGtHNezmy7hIoDKOgUxTQ2BX1Ahhtt
Yg2+zlLi+1uetRhTweXsXgRTrTDWoH6S9YZIdozZyiN2jS9p5+0OtDJVk6seIXv2
GJgdQvuxgxy6Z7QOn/PW/03sisrtTI3uQx/BQaOj9P6KmGVkiW88pNxCiVeb/pWC
/YfuEOnSPmxNMquGLuXxdO2yRcmTHjAEih4pw8Z6aRBcTH0+g6JZYB/aMH1+NTJb
AN1xTZ0v7qHbLiAmEktbiuQTZa334dHMVMI25Khcgi1c+CDRBzOQNgHVMNd1GZZu
k+99mjXARiAjS0BpPUvkg7GMhS+EJXDdDkBETFQ/e5nQ0nbU+5QK90lLKG6ribEl
xKFxIr0MPsPDxIqB+CjsTZWcxrHTCNSoK5LTnVInAlRiGKB2aQQ7KR7jWK4WU81o
OqJUrNqTYW0W559AOLprhL8mZojWtwcWdSz79SJVI041H8K7XtzdyEBZpEp0qEss
JmOrct8Qz2Cyx4hr2cqx8P3YrTq49xoEx1PLwELLw0w0z8L3uHuDpdOzDcfLMdO0
Ok7RWTuB+ysKpzZKV8BhO92psL9z6Gw7eAbMi8P4UKWONdijANsGCoNsUNMy8xtN
piljaInpfI7icGz4tAsK/7PT6WQ8PMgVxVzSvT3MGbr9QS1pbA0i3dNmNcg/dtMz
VxwIo9q5Hc56C0aAKD1eCmqnPN6BhnSKbHf5BNBidA+2YD6KcY2Q+/lJ0T8YENFL
57qREYKpNN6eq0ya7YD+ng3WRVykYf6MNPLolX16vRF1cQu/NRHjenSdgrgALlBk
2QHNPdqTQPiCbqqjVAge2lkBEwR7qp+T97WmfoUvR3ySJhFIjNvj/4roWy3oeFdB
iQJJtPNw39oaG86iV0Ard6JJfcwrwFAPLDOvlfQvdhZdNSBH8389kwyv4nXsgPr7
RFzrfR4vCd6PGjaLC+4b44zO3f2ZozeW4gWUidcSWrACall05bl7s+xg9TdAZS3j
Dt3vY5q9NyMohEM+Nxt8ATVSABdwWFkpwiiJ02y/gr6gg0K701yvx8cZpu+U9c0q
ecl2YAA8okxnTCE9CCD68cK90qcl4f1OQl6h5N7x2Njh0dInkGr0tnCe4GWEohd7
Wmx+b6B0eit8zJzhvpMyB7uQkiJ+fu5aNRI5XAfY/A+V1SZ3WhYPt1Dlw1HprpFM
KcYqQVQwI7OCvoO38FQi6Kl7L8/h26/N4Uk+uLK2YHoNNE+ZQELadSP68MUER1sV
APlSR2fYcwxPD4YCKUy0WIaqQFCCnVABUa5eugg5swd+NyTty+Nc6KQ5N29z5A04
petYzdgK8g58cFW19lJjwxyoK3N9cmOmv2Y2fRqniJlcXIK10W4QF6ZBIYA0hMmf
1h9IvLPLYyaQjIe0SLM51aG0tzOoGgm126UO81BycFOlq9rcU2N+JzEgJKCZKqZh
bZqjnFftCrbLZjiEyHEmWm6nJ7AAqaQ67LkSVhhr/fLmmc4EQkBYuOW+UH8rDD45
y1MxGBvMBrVHTaw+D1Gu41LyfiM00YPx7VuR78engPphwj+sm8LrYNCh/vYx/V3o
m/4Wo8gp5GosTCC3VDZdn0UMuIFngy4ieq7pTA/S32IdpajnutwYyJhzkPXtiLbA
E5/xF1uNS2J3fc70pbOf6F/Bf/O2nCebZC+jJyo1fPLVybH1lljpnt0Yrfb8aA2g
UiTbLDjfZrL1NSfxEkL6H/JipHoqptrItO3UcLOKONblWaSdeBmvDF4lHhT8Nixu
gYEFXePLoK7s75/wLReTR/0Wc8wGMFGSyQyBOVmc+lrkjkthczlhnM+hELpqUAoL
0a5qt03vDfGLzcP8rZq7zE4mH6pBlL4VPIhzxUv82GIMqMHn6IRCAy1mFcXZX7R7
I82SNHnZ6AQsr3CKT/veW8eYHgItD8ybxx9NcjofPPnb424y0Z9xheEy2jgBwAei
SpSmXMXsbkuQsNtBLp2dfdOUFxh9qwOMVkdr2FXxGw9jPI4QL87vs+phSV/fsNZ4
cakHmDdpeHpN/GmzvOmcQMDKd7sMFyOyT7C8O+TNXzE6xCkKehKMo/Sh1xStNWnr
tdRIW3WDr1FfmSpuXhba4mCmcgKD7fCzr/s4o2kncEmEXTIOQJcgcdacHD3njJx6
3B+fb59xKE8hd4/nFQ9m24EnBTTQPcy2NowDPCZzdEuix+6gOFRdeEQFCHVDkflB
4RemvEV9mLdQdabwVxAGKg==
`protect END_PROTECTED
