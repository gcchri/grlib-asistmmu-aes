`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6r8alaNiJ8oyDQgPqzQ9AS3mVDkBNIHlL5vwJW3qetdH9Q4qxCmGAHH6AHsGaJoc
AQczfRN5Ucqj+wFaH37tUfOQ9TWghHsqSU6RdslVkW/g3sD3AxqULamnBWn6TEZr
gi+0nRauJFEeuJ4ZZ+QXj7nI/f39rBOU1zUlEhgtoiYiXYSTenBiUhQswpvH4y96
ehtmfEqi/2f7wV9IStIIY1F4rJbiKlWenrH507U+59C8jN+jzb4YscrANK1pHjgV
9oqbyGA7l5aW7msxsLn35H6cyARLK/Up/EMnrHq+wvuVgrCRUWwVFVIuD1YevNES
Cgqm1WGxPhxG/2yfQn+ipmwQpD3Ueg5v1hhZHjgOuEigjOu2/5RoJ2glLcS14DCG
7tj59nTufyqvQlIfWsaL1QJWPr9XarduGzC90+cJkFtgx7NS0UaANNe+20/TAlEr
`protect END_PROTECTED
