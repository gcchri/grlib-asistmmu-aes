`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NZ+X7XdQS3k/9zLkX57YHiShQC5rH8pu6dk5JyCCjI0VGufwk4m+zXnkASBLy/8n
dyNKO9FHu3pFNkHxACLLbpFtACrxXBOpQABll/1w7kOKPaAvei5ms1/Ma+vltgfy
nk8gKa0PyxI2cxkOZmuLNDxDtQidNMbV6BYr2dQM6xj2E0EOCMA0WGOgfTSosCLL
Av9oY6Kdyp18ZIHbVgvdka2+c1vg6bPxwM3sl83qG1SD8WbVd2Sb7vKu7qgE4OR1
Ecjdw0+u27o1ZXPyNbDaiXZFmcWAbq/4d4T9Lay3qqzer5lTJTklmjH3xDupGEOd
HDMoWPxGnHkuCRsi+Zey7VGLUo39CGyXPO1BVDtkao7cjjrlXzG2CacTvW1LEHs5
8T61EGdzVsVI4K3juwH3mG5OcUP4/Xr6W3QLT0J4mjkPcdgjPm7QydJNyLucmWXF
S8MI7cU5JHaiFgo3yfhv9B6sEIcEayFjgTQcdk9XNFOhMxMNjT15cfLQDFx/IQgN
mvIgxuGDe3FDs/IVa6RLnd/TS9zr+InuzW4PGHM2dXDUI/y1lcgEXxf3xwHHfCfd
NkxTxLN50ZpAS0SJghHkhkALszaIPzCGtVSWHz2IBm4hkSpv8ls5kx8JoGeCvZPo
fM7QXRkq2RzeZIbyzvl8U5BVsTHMPNAhlGdwYczScIA=
`protect END_PROTECTED
