`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ii02xygh3MfCctGYhd8Em0mdayKl8OxekpN8EYIwWDNIAexinfVWsHpDDSQSoxq
X0aEK6l8ase9Hj9NFfG7Ef6u/oxhqhOlLpeGIdTljkjI0Mh68TleOubvu5i92TTz
9VVPBDqYZsq7Ut7FGA1WjnJK9rGOt1JYoYKOLd561czER3SOpFJHIgHKg/jPau3K
yrztLC78EsniRTzly5E08amXu6I/G4UroJ9mZKa5xg2g1RkSrO++M/gzVgh2RQaK
uqkAzgvPbcWTjQn3Fe9WOV1unydLYcSJUnrHQHYGloX2kTSAta/9anoSE8tByK16
5lO5olWduh19ZUdUWducIGI81Mi0XKsOQPZUpBd4HZmPC1jS6pqLq9zLiP2a2LdB
Haz0lTKGdmhGpNrN6VV6fNGOvSZBPBDOKBqn2DNAXobNGtGNZsEPxST8sAWvoUsd
`protect END_PROTECTED
