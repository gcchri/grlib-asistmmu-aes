`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CywqaM7NbYKM1FoOG08poglsqazWQ0580PXrfveM6An943BfX9GfUOZ9F/jv995f
4325DqKQmsT/M3rEmptXSxBz//Oq9ozx3JDGWGh7ghrMz9bY+freOykQHjGOZXJw
ey6gcWKDKT0VG6VAI4UKuLrDs2T5TZ0FiQmYLGSlqUdC8O0j9Str5AhfxSlsuzEW
TDS/roHWaG4zlRTSe/vZjbUFmgIA54DNqV1ZMIUsLIUsZiQbP1d5Qxrij4xby5zI
coV9MbaWGUOqxDiPcHulgS14gbd99jRYOExsiBhICv6oZe0NBI+9rL2JiS91JEuR
YPKLmx9kHRjur7NT3/Komh08KmrXhb3yekGvtLHoYXuo5bB9TzHkIZowG6BM2Cu3
bbQ3dhzRFgQVtFyzQQW6e2c/o4XLFAryZwNi8btu4TzA0p59Of2Var02Rs6uc1oX
HL6pH4NQCJYtnEOSDRySnL26rQZS3h2ZCn33+AscfCI8RdftkxrJWplvjHaTDSNj
JZWbtDPT1Gs+cCTBvovaXisrE3XIjPZsSQMwRXORDdd6rPO7639ulZHxIxXxQHU7
+bRO5c08hRPPXrjimZPLIO1A2XqCNubvA1yderRVJI0G0S0zUgECMPE3Se0/QqHC
MHqmJnoaBDwMVS+30HcS1/S9neiROAWY5CNh8qptUPGJ3RBcCEc9jdAreUK/GS/+
7CN7ZT+FwniDHN74Lxq39t9ayDKhvdFM7wVbRXcSVyEkjFqW4UyePRWT+B7vAjZ8
w+ah4yOTuCY1EfF0Qg1pnxsNQrzTgih/JXckYIIqjyJmHh2qnAkWP2kVX+Fvq0kV
iPTAh2qLu4Rb2C7OhMfi2uDXXzS5Zcl8XDwAp4KROcCl6RE52erMmvIUmxkOB2sZ
j3KXSo4/uRnVQACN0IgOwu8AIsebK5AWwDMxcl6VrkkFWwqsl+oqJmwKeCdc8FHD
XhOE0rtN2KILGpsHcq7DVAagn/pattFfdxt5PyF3T0tiMohQCkCydLROi6L/mg3b
kn0K9vKoNciUfKQSdyir36idCOpFMLiDn47oSrb8M3waYNsnP4IPy5i2HS3+BE2b
YywDLvgBTndhjadudAWKnJznOQRJgy6Elnc5MHzseITkgcIhpaWh/Vl+cRm7KtfK
87JeInaxpuROIZ8JUfBlAKiRDBtaklDVODgkq0r8tyUiVlmCS350LD4bHnM7YNNL
Gq2Wc8ZxZ02t6xYC6cBQid5I4DQo7LBiBWqYvLjgkwYG7vhR7HPuW/XN8HlmPYai
IjBuwJbl7xZFepNBVei0k89avokhNHONKnuTkhBUCCpHupcksvonZffS2Mzjq5MA
B5AyNCF9O3H7tH37KGHBLXy9BVjG1d7joPeTC5prV3LzzQeQKCvPzSp8gVwad4zL
x7LB29bz++3lULL1cioHTczmVHV0acFLjG9OFrsTdkt1sUOzbCwus7dm9BdeWeD7
j5iLZ1CdZ6+Ha6VnKImJWbmMjpD1od2fYA10dgItWxtObouUcgSXAHObQ5leg+Or
PtWJ6XD5AiJrmdKs1oYmuFnRSei+Ja5CJRc7FCIlzD3R/d+T6yDLcZ4b6/XGVJnH
PX0EDeaa3A/PDj8WYps3N8UkHsCgvmYF0RHNSgIHYpGkQ2v9rUqr9tnFuolM9qof
4Zl9CjARFOYK3EEkRn2KQqyADJI4oWqrcoRbr6KhJIELgvehvbKGFPP8VO/ofmfA
5DMRcJMdLBf9hCFoDrZUZwrZqQxm5hVn4b7ZP8f5MNy9qbUYyWE02RsUwSbHbGP5
NGXXlwM9WR4lurUhLlyItp5kc1mVf/boRHoTqXa4+tLJ459kMD6LIP6KZSMwl9uq
IaqbnZVZKJ59lq53ADMfWcNXxCF2YzIPGJL/XV+icOUgd5UzYHtb8njQ5mkSdoVF
jRpza6wbrLb1HUXp3+Kw8HQ59xH52HpY7jS3YjsJ8Gg/xEKR3z5a9xwi48uG0JtD
479VWniotJY18FmM782pwYMV3qlNLAdlKTs5F6GlbOFBiz0P/lw2ItlCZoQnol6L
N9a32vMBrlkw0prGGXFN1KgHrflN/PDJ4ycl788C4f9Rgethfc40IUO0NLus86DS
zwB2UfLIpfm4tX9klsu5jT8Ac//zFU4wCPRPVmzKaSfOn2YkjEONiRtTfRjY95Gp
QqRTFKGW8VFEhGCd2HwzT+mnnMBhWnRBlIdcpYRHI+/PZPOwJ/XTg+bdTd2nOuME
cjc3HEbkeodQHM+7wF+QRvD9jMK0ncnJAigA5sDdn1XV0Vd4wASA2shYY1FUBwrq
X9tvl/f1VhEalFcRWrl123sMFuKjQBMoL1nqyoRTp4dgJ/LPyzXSZ2DInnZCVUJB
59dbyAfTsdKCwzaO8paVhaEmra9lW9PK54tdwF0FZIaKfJBueP0GJv22ftKV5Lf1
pdOybKwECMRQ2HGCNbHWRoVulQ1pB8X+6cL/181pgvsZUci6EkcIYWIIEnZZ2OAl
QoGcSHjqBqmsQRut43ncCXnIewCwM6xO31skDUM/cEuZAbwJkYSu91RVkoeAmCo5
wEToyC+ywLXNOtK3dN4+X/2ymBSw/2sU/IY+FWWnnZUBVVEmwTzY7Wp2gGrEraFx
DQNYePFeLn+FcPVJlsNRgT3wTpDQ3FnfayQN70F12XM0GAmr8ycEpYeZh6/smtNE
o30m1ECeFtNgUX+yD+OsCG2GsSH6gBX4nlrLB1xnBanw2cpZmCx3RAfgndvsfSN4
VK6idibquQEKo3+P3j2mFmh053MEg1Lj/J4j2HmiP1B1lU7YIWGthIqDjsrcTaby
fuPkqDMiHEKMs9RGnMZt5W5B2fTuI4wGmS0LbTwCl09ngvQwwtwV2lfpgIzBMvz5
M8d/6UU087bXmjMEjkXd8XlScpLWTqHv725uzXI+K1TzXDQ/QslKQ964XFUlP0qf
Rc456qIDZx6QHG0xsQucBNCE8hHk6bJL3JJetEJOAYHpbwCK0l8LMI6P5UqmptwA
9GdOmmEBhtXEtSG46Ge0Kks4fc9sR58gELEIChA5HWtml4MSP2GS4GqXSSLA5lA4
O9m1R/1UQ8WVXleWuObM6C0n3f+g8MnIJGDFQ3rDWFvtzWT7pV6zSP7BlmmaRCTH
BltLPD+8R5CbuHVcer6RpVK+77G22El9VCnOh1ER57hsRe/thialePrx2/SRND1E
QPy6W6N7uCrlPNrf9zqO/9rx2pjDN7MFZW1aGYtUpcU8eW/6Bq9iQeV9cEsQyXDl
/YQWf5CarW5VgIQOGdf2jeLFYCFEo11Y1RXktQoe8Ca4Fi1aUipBb1xITEmKDchL
AEhBSEB7GTyr5KbrRytqbOM6Bxw5DbwFtI4fyKkJ2Z1PWIk8LPF4aVbqmOZQxsG8
5R5r+bz7WDCtt0+j/pzg1vayjv3iUKRThC4fgFCGT7LwqDFYoIdOCkXSnfjOAvTN
A5Ty+gqLMD3ZU9nSmW4LoGdnkzhPftKUezqAz9IBbwkVmsSIIht4PuKG5FwAMgSz
s9295wJwHMe9rlMAafl3szwGxiljYNGBjvTntUCKQAXLfLLjZyGBIqLctBLajg5B
pehlSPkctuwIpxbBjvGberRUC7zFyDBTHKBfJvqTYbXDi21RH2f8Fis+ZMseF4RQ
uNCsDPmuSRwaH0XUlwHF37JLwKrD0et9QpIktDmI8UUV/EZ7938LznUaCWgxL0w2
u/sRRMxoLQgvQtpmM1pWTOLx9rq6yUh/kYHSHEN3Y1Lo8qfxsgZoOgK7oz5WaSZr
GRSE9QSEm6bDggDULNB860IgsNlkM6nO//510KLorHJIfkibi4y7b++5cgq2UraD
COccY+inD3flSF94vn9K940EIxsYeH2WNSU63GS7/tdDh3CfTp3OjYxr0nanhOYX
Yfxoi6f0ohwauU4BLe6zR6xvEiX49fPFImN7YKyE8iRkwPG9K8i2mRKrD7aAF0GT
9RS1KbV4RB40blNYgUVhJXRdYaP5G5GxjCL2+MDPjaZnZn5DOGHlW7hHrQ7AydJP
OJ9R9E0wTJT73NoTvGXQaKO0sxKH2CJgPdSIpd2tKqhJXBgjPkhgrCVFn/p1g/P5
nYS4D1Iv502FsZN/nXkDJzwAkYgbkhHDeTEItlQ8L3ajXJcEc7eUwnONhZvsaHdn
Rd+/C16ChrPQ2EEL5Q6JPbvb2dKsZ67v3D79YcjlpZTotiLytyzgl4eVhzkB7g1v
R13KEsjb4FMqXYDBwlvYKfc2U45zfTA95U2nuC/JplW6pgC8iQopmU/bRI/fVSQc
y/Lbm4KRYnX7MwiMF66LwheVGcn1Txja4YWRGtR8QSFCRcLCbcCAWlKuRRRlBwhQ
xZA5oOtJ6KD2yOngXhNne8+Z4eYO533rqbuy8h1WJx+GYqoNTEuA879JZ1pDUyrT
uOuC4QUKvBq1Qgcm+0OQqbFmKOhygiIrnLPYBFZ5qppJ/S95hiMpLay09p4okhYx
LaQnc2oPYbL19w9EqKpRLnuLbH8e0EC93HlertOiuyVu/pM3ID2lYnpdTQv8cXmG
MXfbvwDyRVEZAlCyXYjqoUNq5rMCo41V7V2XZ9WVJ/p6t0gTeoo0qZ/FqLfphIAE
zTeuM/uXO2oeV/1bZTXAIAnPlirbRAs5dFrEJZ6TXch4rD3opC06Hk3cAOFs84BT
rbQ8LJJloFfO034wgQMhMbapxZXJwYMuFNoPAYMsuZyOfuRh5u15otp4rYh75L0+
588kQesSLYJBFFkcjewTOliEF53wl4L/RDn0wS97MiPzK65Ry4jFZgAm2OYEkSPM
hkmAXRXVK0e3uB/BgVOPFFTfpCCSR2oOxBmYQM98PSmQjllWrPUiJBXmyPwKjfua
LKAVtc07BRBiH4eJRRGsjuAQr8VzBG9+25edRzI8c3YleWMH19cgT/zBnHDlOwnq
IZ46x5lIhTCJPHRQiVZwxJ8yJzrLLPR725Xetwu5FsbisFhxblYAe+PFIp6+w4H8
B33rZW92tlIGFvsfqjDw0WtcmBH0VoaPy17EZ5toCMPzTlGUjmw59O4tuj+PyCaZ
MKoaUUp4Bnl7gw4euN4LttInLzvpOpRcSNYffE9NGIbDB5jc1TXxO0aCJAmhD6Eu
KnZ6Fa29pQGZ+joaJ0TyLI5/xwktBNlK4PQ+MctbCBbbicTK6BfKggnLNxb2aQbG
5epNk97k5uqgmcD7Rqp2rn3OsZi2onwvCr8PR+yraS7pe8iicu6BjadUgy4ZTq+H
WTj2b42AXyfV3sqn57RUdTyq6ja910PFbg/bZJt48WbqD6hX5j6Ek5uDmWWYxUWM
MgDpV1j7ZMdwpqkL4KWXtcDFMATBZTHuv5oKy82/U3UNVGqJaUnGf9egZoQ8nfGB
kh2xBLaHTg3gMM6fTYAK4bWvQzuHOr7bSMePLok2g69mPCyrKxOT9DynVZTF13NN
yKzazNhZohazMdz11CUwFE9jG5Hz6Bm8RcwdUwRqV2VIve5WoLiBiLn9iOfR2TWK
/wBtS4QaMe4WYVhiM2MKymFYKCQ8EnJSmWyx/j3QymJT3WiK4vvT4C66TEbUyvHj
mabzjTDgO9+IKoNOvCbKsDLVf4EaIP6BISRGrdeqyrEL5eE90JKMRNPJ8sOEPDXA
mUdRaGBP7pbzsGRlOT3XtHAS11evIBrbQKs/EE3ZVBue9nrSwmdFV/jhfZhctmP5
oNT+0tIZmmreIFiGK/fZKokZaO8FS62wOE1LBOeME0U1bLuqfDNawtauCr09erY/
hBu6JvzfWubIyW3gVPfzv1+fstqOEHZLanDAfINWJtUesHPecWnwpkSjyYeRHhs4
jwVBL45055kmj5aGySJFg9TSVG+/Gk2lCloVWu9MUu9pZN+NNFJwNV4Rfy6YQmeS
dNytkDShutgWXYfGlgHg42lnDVnEckieRjMcH5bGzPyq57r0rDpfMWI8IPBhTK5X
XCFjcqptQwYXd9cD8G53Z+Im/vZT3vABKGo/ObqAy/9sVkwaI/MDK2jY4CcgDRt6
y5P9k67iefsFdYURoXwgZNXp3vTAYamweFL/2Fxv4QKiehl8fThzf9gOCD3EkQRv
zL7fQ3ZZuuZ+UqJ4z3lQJV411GCjFirO60CGVUHAIdFfYJL2mHkiRQLBSpUGtAnV
UqWbzxb6KC+o/V7dPfeJf0MtxyI55gGld3IKYHFZWFbacc2AQWfa66IvBj+Q8WV3
wSdONBfTJMTclR5sZk5P1zWhOucqdPm0STbx3nZ7dfBI6WDD+G91PATX0r452tKw
834/H53F+L1KrNSTAhOVgbe5MyQr7gLCqL+gEcYu/xwGV43rzmIQHK8GURDfzAPm
+v2zZ+7bEXyf/vEZOxNyCrSqUuaiMf8177v9p4TpbDw2y0Pgbmu+Jx1Fs45QpV5m
Y+Y5vXnPmcDcePvvssYbUlD5qi2NzDEoBMhc0q6U+hGGmRwLaFBIZyS+iiABilix
NUmvWwnXueFSdKaoWbkGXcoG9wXxV/lvYfP7TvMcFExZvuBf59OzZssKEbW2LFEa
UaXVyKt18cP9Ap3Hdg+y6sHRnSgVIsvWZLTzDEyOsOkudq0uIGB038xl1GglTG7Y
9rCj5bwevQN6RILbV/0u9NK6WrA1Zs7WphpBbNVtNP4cOzM6PKA+oZD3sv6W7Y/5
OfZrwVXQQPuiifk2mDlJzQCF5K3ZPttpbwN8p7/Sl7Y0C+92X/gADJ662llGCZM6
eCGZKodB3NlV7dZ0q8w4klvf4BuuooRF9Eula/iv/Qp4h6RAPsbllI4PZ8Jl810j
JStBciziOaqG94QOh5gOsgMUTtHeqTxtrK0JGG7ptZSqKn0RpR3AzN53Mam7y7gg
HFBxqAYjxEOFVHPm5CFhss/xzfyUvcJ1PVP87DbP8vllbZDWFw2JYBi9f/xtjzp2
bX8i4QHWIIgKCf/CEx0IJBGGNpXgb/JY4DXVuAkwrMZq0WK8ZumJqNrRr/1MIjee
P+JSs83PXYQdFf0wKsQ6AMcfyAZyYVT8e8DUPkmr2oqs+ciqkfmmIF6Ccw35dRzD
zIbGgHFR/Gx8sFJnD8Nws7dhXrfpvrURNcVztfzihOpwpa+zAFIMHKnEozwXuedy
tWLmUiQP0JyToh2ZDVyyfUZtQAXLRzITnWSRZ36xylFfAcW5mMurkB3Z34N+UhdL
jutOKCnmKRMyGvO9Ux+/bLGRFeERmWcT3y4gtpfghGnoCoMU9W1ouJxD0H8oAceQ
GV/0Evi7pNiFAVAbIqdXWM0b115ANUvHPDOO9C4sILoN3jWbsGQ+XPgYTjmXgsk0
Btmcq0QOKsACnCFAztY+GGwWnCYyCw+Elt1NiY8H2Gp9umOuLYhurnHMudfejmRn
xO8tAwGUXYPNnioMUCLwMiVeeUVWmAcrNR6GbqArVvb1vcsMEWPmwdYzcmP1OLD4
bAEP9Zk+2Pt05A8a0skPiJv5zbhnbtkEcCtMjvH2xMCARV3HJPPXc7dv6YMcw6cx
YbUHfutrhOhaWyaAV6p7Qj3gy54v5x3ydx7tttkDNV7i21wXKFd1lh21RIVBcYdS
Fr6bmPXnXPRhpvBkKCyl4+is8CqC+Jxex5jExn/+BZI28Q5YSs0xsBODOfyRRe3S
vjUilmDIXJBfnuQUCGUO9PFzyMuxJhnZAjkX7lxcpSTsEb+9gmpmJIwT8gSoPOQi
HCYvpZ0sHcnlmIJaLcrTgvo6T0lUySVbwZzDblw/R23BFsdaR/IggnBd3MOS2E//
mfsRsJUzWZYl57+JXGjHgTs/GgXcqwGBOc93s5eVNjoS0ViTxzPYBcs9WEXA8z57
JJSnp5VUBaoD+W0dFuOma+lZueS/xTw/RhQX+H+DdnZZcIUjUYtYeLUGG41xTHvQ
4ClFti+5bu8ZdJmh4p/trXDyLdLd/HTwbhq5TSg6TNEOC5C54ukBwmUc/HNUzFta
+qtVQ94cBDnZ375+nkocp1EIrBoJjxCeIpd0TLkRHYxWt1wDDWvvQVgn8tmkqSr3
1BhSVs324cghjqvXurmOdt8BDk8lSxcfPSb/jbA3J/kDQ/KnkSaGaOSGDIP9mWFV
MdFbCaMzma2u+O2MiI5tbRLaEJNL2oucuQHK9RlXQ+oC8S41gaBl7l7EO3tK4wzA
QIzomHDOPHOByOJaSaQjGvdsBvdloS104KBfeKKqOhQr6W3rJVp6whhmMyCkMjGf
/wtOGlGgDiBNhIRo02QMUg3S73E8CHeUPMk3cPl0klLx3fLGaRQqCtHQv1YiVPqA
YCjtYMtpUX/5hVSgCyOtl2VQa971xWZA0IPO7BwPC6hFB2VjHMuVXzi8VzCcKknT
ts7O94Ytf7DuodyEGxVMRFRtWdihkuV0G5YBAgUxuIqrwz3xXHsoZCNHa7zdLsco
Rfwkc/0LFZezJ7p9670dqI3+a+2VERzx45YmwC8zV8/Wn5C/YiL3rSvL58UxGAwJ
i4vK6aeTfvRVxeOc9JiRbZT7molcZZzuwAY+xbKZUFd26Vs/GUNOvAQn516hrOlY
tRvTpzWWXidOjMFxtcjH7fBJ3yzQDuIakgiLkeEAMmi5S6rxu6MjVfvV0DJDM6ka
Z0xE4vcVaJxtt0wHoEmswMW70QBByNFuuiip5gzGEnqhk3Klx/xXONMm9Oqe3ZIm
rM4E/7wfGwjUf3Ew5hK5+TjjVVRe5z6rtyGdceMFCZokpREXKO0Hsv83WjRfRrKF
xvn6OqIBSzPzGDz60N+F3ZO4M4VM9crMd4ZdtMcT8rS50liCI7SpuCLJuZ6loRzv
AMYZQ/hb1QeF+hu6SPrJ8gPkgyGF+T6WJZiUm+hdr48zwBo4s3W5VNXHctbVbbPf
UflhEkchrpkqTD/R+s7aaqa67msSMzHjZ54aCfBfaPPP7XoawC5mCerADjAwe5LM
zwFL/QC+VxGF6x8CHuZUuExDtJrrWKx59Ltdjtds72zckH+n7fTzEAzGqfKuRUj+
W0I656D9icozjhSxnOei4XVT5ueopshCSCSPONriCegX3TDSxQes8BbxKCd05ACM
ptyycTEEspvFt8zFutPJiDjvQeFXteDaD4yL8TVH8eqcA8M0v+lShFnMWCs3fF+h
LKi2Hs0cGyLOPaoqR70KlrOQ/cccHnDJKS4KLAfiKQgrfkB9Wm2qC5sMmp1Unr6+
umDQOTILoHtb882dUe9MRZyULkc35/ICG+cSGt4kgT4QP/yaPHYVIRijSjImuHNU
XLgnR84l0pHpcGrwKmbdQ6MUhboPxRSlG40wi3ML9YSeJ3nMkAilQw0h6uUkAGLR
5Io8MnPhaVbTeDhWJOoZ7QcJLN+Qsl6Rob8ShiGY42WcrZ12IFlFnNuHkVyFp9iJ
aqj3tFtwNYbb8hdD7nSkZHGIwkG3B3SY2wOke4uVABrdMzm+f6VgpX0dDFu11Ely
K1GbAWOaQAi+UFmRurZjEtNK2+AqeEWRSdCGnkKygDRr8Eyf+X5qI4RRvuZTAYLd
aQUah41SbyumBZfX5W4kXfJ1MMh2ki7hoxxBf7CAvCFDcumuBY2ZDzn+NtQR2yNr
fi0NtfQFwVWGKUR+GWavssxgYII+aZIAnm9fcquAINNbNlT+gq9m7pyXxHYpiuqD
gCW+P43yjC0YRPHx4jeRAmanRz7MH+0Q3jhnYOUHMHG8M5jDZ5gNrd4tDUhg209o
Nol/+FkaUy8u6S1EudLhg3vk62sS2CxIt9V+8vgCt5hTZDUMvM21kF7cZ+3m33Ww
Z3O7dU96lO8gUBEA8q2cHuHs94IvRjS+DGv+wlLhv+RxmO1/rWDbYsoZFjENhXnE
xOXgQlWrVf3JE2svRqU/Jb41vPXTV35Vtjh+WLqUK7iuMF+qAjG1yGlEfvyYL6QH
A4DH12qeBDbfIzLWWrZbwkgEX7vOuPoObMu+IRfQoW1lEPPjt3NaLYFs3obz2sAS
VNyb9D0Xrdn0mVQYMmPajlQOLCfdmHrARptAK9tt5CoeFujFeko9NZIKAUKYpuso
9EPa1ZqbGHDzKr/0WFtGIEd5VkH8Xo8VjHQlWOZNhianI1L9n5HWuPz0N2mTcucb
YFS4yhZl7FAsjnPSrD+tp7tG1XNYBER6OsqHkpODr+fJXwYDPQdznnIJmGQavaRz
xne1rvj3mUkPnqL92X/vYSnT6iEFn4+VW4jgN3mB6Y1n336rU40zN8RucGFc29xO
4qhRtfQcrY6xh3cCqFqcn2+WkeK/LEj5yp8L93sd0uc+gK6j87tPApLMWx4I1C4a
/oXE9Ir/DSadkDOAtjR3utDo0hN24aBvu3LL/MLSTaU4+3Y1cxUq6WE4gwNssdJB
oBrMeo40HuVrTAn58jVkYIBn8V8dlNfQuYydKrXjPo1810B5lq1kQe5PfLYGeq8a
btVGTUjwQ4vi3n94rDwsDs8gOYxA/jPWbqapiQX9XiPhUslIBGrBGNQ/wfg0hMV4
x/zei64Qk67P7/QQvo66vbNu4tCMYnc6y7WFu99KKiKnJLBLS3kLzWs/U/userJU
bZ98W6obhdnAf/30pghKq5OcUaiMPJcr2sVHePyfj7mwKSGDhhoxy1hnAqsLyFDF
a6c2TbFjZAN6cMMf+mElWpiUWpphBoGGSpv+T57DuUBWUv7XOBX423KjNvDztjPQ
HQxBVDrNtvt2vvutoAjCEq/dEqR8fhG2sp02yeWKaO0v20mFNJYRiL7Eu6/V5dXw
6CJKdIGNh5wXbbnymeopncIxzTcE1GGhSlpoR95kbmya4Wa07IEefSXfQvvqOlVA
WJOQ6DGK5utP9PwxU2X+0RMCNILU5nIFq+L2/6hoaRsRxgiqI+zLQ1j2zoKlxpyY
o6LxmRNT5gFlqB+iX4s7PmKbM3TzNTkQJ/NP3xgODYRR+3/TkJCYeZ1OZc3t548Q
mCgYTd80gYFG24ta0dGT3uDIRvjV6sdHBh1rCFT9MQtXLnU8jez8O89gY0z0wW8M
fuFSA1iOCZiYmy9gPPUDYEqnQ4Dqf2X/zSl2+uk8J8dfynPEXHhrBm4dHsIkCkqj
VWSvyGZ0AkxKk6mP3S1rz97kPQgZb9GO9S1eIYnlYSYXlURpUrDJSDNLz4Hl+8E8
H5RhM9iY19RDUTkV87YWamtCydcl2j8PX7XRtbBEv2xc4lXjxAJarOuqp13ElpBU
3oSUwYMRYVf0xruu8wUySiTR5njVc2CaT1I4emrhAJBFLLZJiUK5OgEaC1D19/5r
nrBfO2TEArulqpW2e07xKIACCxE8rD8BrlU21ya+g7IxA65ycJQgYl84elrkz8Do
VnpPJ4liTKHdqvDJP1SVr4U+wHCcVOdcLldf93L+EpLTG0Io9oJGudS50ep/enGu
enLOB4zP7/MqkpsbnTaMdJq8Tm81k/KGK0+vXlZ3tYZ9j75+z26gDgHCpyrFKmNg
5VsPUfleOMyIGNV4e01erhBsWyWEdHZqV6MT0ZIxWRNcbS6v3ieLTq+ozwnA0kp6
/+aGvyWOsP6MxM2QVfoDvKFNCrdfRdA7H9PpkkJTqSc36ZwHvrHRrjgElUQE/EzT
2sBtnW/jQqFxjj0mMmzSUGUok9z7szYYVUXmPbpSg3//e7ZHFvwakbYqyCJP+qz0
mnRezuCUMdsevUemCViypxRzO3TCXwtvwmWcvA4Gi2TqzUGwpJvAH6JuRoct/BKH
6NLfN7HqYR1Rb18nyEFSDzrTpEr6y0K+i5b5GoOtehLUNlc4WmxKmS4tDFOt1knB
WUBFAk6r0puht7mCIhSkMBAoEu3EhL2rGXq61C63TTmzHaYNgOSBFiTy3MnJ/Y2g
r2RFoqZz4NhyD/hS9tI1U2SujJmmGX6iiH2gD62vMHTPbCUr3AmGHzd1YAl9bUM7
lBUSxYcKUe+MspbKUAEBxV3Ukj9c8AvCrVOuhpF6OfNRV7RGR77jYt3uvFjyEoQm
M9rNC7bJw5vWU3datCzvqVkszZLcVVIjtLq+4QId4hvRVCs/0kJNsP8BthAmtdyP
3rIgDLDLlhd0ve+uQPIC5IPVXLWC4EzDlogiL16CcF6RdeO7Ux6HatpsJNbPnyXF
BKacoY9s+wVDnphgV7GIQiBpmcCpQXtHRiPygYrwhcfqG1Xclm/HkT8tG6sTAdkR
ScM80u7mP8Bn+YCXvwbUzEL22QYDHbT1YYTsWvguA1WyCKWkSsyTSXXoyctxqeAs
FWcUgF07X8x3iYoJOn1YqNhS6HLTmVAPXztxP50Q//13NuQnoFWy7S6hF7tgnWJR
866ELcnidXHXpXPoP4yH++iIGfW3BUaWlNeQkh6UGkD+t/5mvSfrwAqGFY9cHsUy
JIvtpt09V5irlMd1WVVoBCM9YXFCOjmpcE/z3OQV+wm6a1OjD7HEtgUlgctcHUzK
Hj36fY4MTWCGz0fU5tUVx7f1vkNkjBhdntPahsCI9ZtOg6k+eTND5UFkTuCHxp5z
YuG668FbFXoGs19/49oMXK8ONBmLPy0UstUkzdIqKTkEFAIoP/mSa+o/7EAC+8QG
9GIP7Te8R8eOLYd2H+CiB/XPcAvpD7i4E8LFBf2TvVNE5mF1GRQ88EPAnY8Wfe0v
CIL+yISc7h8b4nTN3+9nBvMjHlY/jt+WPVj3r8k1butzq08v5Y0R7ziN/E6glxv8
n2z2r7RBTMKjj0z+CE0VnUe/Zd2l3QSk86vgx/XLSIOi1zyrPx8DcH+Zkq9Zr0bK
m+982sb8FCUoLwxVtrXCuioJVLIsBPoN8EMRhVH0AWaZZbcu6164Tv4PlRVuAAd1
FOXGz8z+fgAUjZ6LMQag7WNA+JVORIl1oZWuOUxRoLc9rhaeuH3wVleEIHXmYl7f
OPnpW8P71xQ8AeG/UgTsdL0BZp+2HobKdqAqkadrBrFku1pRng7RJS6GzIdAxjBb
AUrmzw4KeoRtynmTlzRGSbq9ZTVthUm7b4wwg9T82211na86NTPffAptXJCBcoAQ
yt7HDbtZVfOZRY5H2c9aLmv5hzqfKXvUjU9QaW8+bBSkpDom9UPhBn4V27TOSTc2
iEoTv66DBfqymdfUsKmLykYwUpILKpWeUmiuagCoq8PH5STzPlYbsaydg6PKB0xp
Ne1gyFmyl+1jHAzOJyv5APo3965n8hA4gqHEm5NPt34iwgaQZcd7ziDFcbMkku+p
MzkDlfMcy5lEyzOYeKkfl8LFzCYQGUSUMxRdVjJexRQCSNowGGGg0YqZ960A/1HB
0kZq3loKq4K+6MI3WpLquBuPJdLJNyq3uO9eREpMrAjoffuv5CQBBw6iRS0Sq0aC
s96sGGGgZQ33zXiGU7d6utViq1hRjvVy8eAt8I4L+A63/Y1Phm5jNzzMfg8lZKyZ
YvxPRhqHKJti5tiV5fEg+USj+OtAIDCAK3Z/qvviLnYEAtmAW/i8eaD/rc6J4oxc
jidqQHNeRneamqCNAzIytY640GzrN6IMCv/7jfiKAV6qEQtlfh1qs42QhmiDXNSy
msBjEz+BF950u28RishDzkhqHRqkkjyhMuKrzimWht7EdNPqH41v1d54v3SOWpN0
L9eEd0ZK8JB/DG014a6SCL4YIWZDc71t8tE3xZ8UPlLkbhusbHH3GibNzMIshgvZ
E2DzkuppOSoz/CxnCVmooIu/zKqUV718kSRIJQ5dHRftTqFXv2aotFK62gO/qZ/J
G+QXZhZZSoy9RmQzR7ILhiyeM0nBeog0/AArUq++xBSMAz7TK7h/bXmJkOAoXy6O
OcxhOlhhsD+CS98YYP+IhNlwNj+nTp7OAHEdDJaeTZgL1YVFtd/phaKBbZmBv5Vp
xvmAfeVa5bXCUJua63/mn/yHkdTgaS08l/IObTbPu6s/41g23e5bdcQ9oCnmnVHR
4K1S9Y2zYchvOz3P3E49aKkCCgyJvKvYXlQ/1KhlEBMtrwxoC9kpTcLP16p2Hzye
e4+lAbVW01pPJ0Grll9q8ZNegQz8ij+SAzuLA3pJ0/P8XDjyYNjdx+WgH930PMyF
NbDxFoqnhfm2xonyAXtRcvuAd6bClbYYLmizY5pENHH0EH4EPTcQS5KTrnc4WX1D
HrDozzDTyGXQbnyejw09PPdQaRYYUXfDkyGXGY2I8wafauQVAF+RCNXGnrFn0Hqw
Cim1l0B1/3Krdj7fE3qB+53mcf5mxj3Bv6mwKGRz3pZGkdVSIDCfxwEASNBf6f5M
yHkMyEBctv+KaSQz/F7tDO8mbyx77pFG0wp0/SoBAgYky/LXS0y6JCbPogHubx9s
FMCBsXzwtEmu/mb7WcCElaj7mKCwqzcBPeX7PmDkqBji+rzAoJipxL6q3NKNcaUB
aliqHL1mMdsr5C/Xrz6kWewYuBij+C7pkZCjR0tcD/jRhCxQNsr94Z2POk405bPq
3oua5KppiPG0M3HdHojHMU5OV/bB9sZxTm53DWvbv54qECi55GWyNogQCqGiZJG3
DS1GVsBzvU3MXxaNzUgRGN+pA8tukM67sT8M8mSr8nwOxq1XpFd9JdCXITLHWrZd
j7cAGmHgy3Rn6tKQnb3+6vvgyuWK69HwUp7GPl9kmy+Id39Y1M4L0H8tw5GWlyS6
xPm+EG7lNziVmMPB/fOCrcKrqJMjtsvtIniiAoPnZ4hiloYFFxFW0zbgp+J+vYE+
fOYNXgb7tq6/B1RV6Yg1q5H/B9Z6vqdOpUyN2NVbnpRh7CCVqnffcOVGZ6pyWMbE
aTl/aOMn7NTCi+QPx2fhknHIqYa6gHBvXwbp/8Yttjy9QH6WW8BLZ2KSWqnoacL8
KL4Y8prs8qjtjVVixG/LJYcJot8N4THBcKNd66drIWJtEBUdXOvhvAs/r6NqxoWT
m28tDet5SNPjZ19rLjQE+3Op21lLnNKNw4C0yyzSPJBcGCTKY1jkQeZS6Y0iRcKe
+QtR985uVXHRTOZaV7jXW1qAzMyd9Tq/Bf/Z+xsuM4zrgnlFipiGWJcAfUMngySW
5mj4wFvtGbRxuUKa3y41sBMZG/5q07MBrhSab/o6USVxmL4cm4KMHSL6ACC5AIJh
hOtFBTtqTwbAL83PMOrPZ3vtrGoMvs2QEOlIhwIHitjlP96d70iDPgt1v+BmxyvI
I5bG3nkjOSgKSEiFDEGJBy8cR9hqFHC/g2DAJLyPqwPMaND1q2pxQ2TeI3mTtraK
RLqdm93XAhwyYoARwh7vDl9kQYvQa0O+iERz1W20FtmnYzkvOv8tG8jsA/CVvXFo
XTJWbW6t3cxaPxqZbyqyfnZCAvOY182R0Mr/MVyZp1R7z2Lf7hQObpk9TmCED4M1
UsvaJDr7gkcCZSYDQ6Oqwy4Kv9peAvVTgjcJybrKw8yvodXfb5kDdYfrD+wWjb6L
Y6R0vWCm/bQ3GQ/ORQgAe8QA08Z9D+J+yW/hLxJ/dzIguBKdLsQrvkwa3E0arp/l
DwePxX6HvTcWXByta/3M0QIoM54qvZAX+NrvSF7cOFkWfhho3x6dGhhcnU9gQ23h
eRugxh7cL/Ym7h8FNsaa5uCzP2ZW/7MeFs0TPzBx2CqTS7Sc6rTxhk6jU9UdS2Cd
B6jINddnno+oAp53rZW+6aFZUYpNe+Fu5O0HEZm8+CUA7ZlJmVkHPzt/bun8oebP
8qpaFFkXSljwPWTqKb0ZniKb7Nww2zxiepucICnQt5fYLjVx6TGC7/V1ACNAntPC
J0cpkPuTuDS6RDd88DUxmbY2Lb3QIsgon7wIw1fJVRdwgIpi5PsZsaKykpvmPXsL
KACBdrzlbLHCXMkMHhyBYFiNFenCqX7rQ7le8QNrfv0UQBa0nKI2No1WLGNhbxqJ
E2DjVGaLyUYsIRavAT1ts8+syX7tm56q1ko2sA9RruE0qVU9hjD123j1EZl+U6DZ
YavRqiPpKoobBK/KTbZ/02MRDaVOMENg1NjhsFVaL4rcZGIWI7xA6oOb8uNb3oCQ
vxIFEojqbpIYf6d4RUJhznTvsmCR/eJeZECgxXKw8abxFwh4OrZP4jZXLlHJZItw
ki4gypFVOKNFvKxFn56nI+7lX9kmYKMJrlJu5EE5PTEBjLsd2cizKqObpZf5nxnj
ObFdWBTLYxLlbmL3lWygH4iSC8g0b5hicQWC919Ws4DfOSmcPjtsgoc7SeS4/H1j
v9v5mUB23cVzmKMCR62AecXh+eqwsUBuF/9FsNLBk2piVY/FGu3n/xcdB3IkuZmc
zhtueawfSIE13/peXO9NNbVvWcsjXI5fkS8nZ8QGzPfFkXSyS7+2lei1FqEagk6Z
Y5QD7X/0qexmFUB0THxRr+9y0LpN53HIwqn9xVpLZrmYPuYltn3knf+ODGTiwOiR
ywFNQMxmJiVPeEj2zXbpBTv6KROGZ6cNM9SV/ZHO4fBnd8KA5qd2oTa+t4Unre9z
rqDPHRdZIcGOgcxCjHA6iB8HKVKzBa2Q0UcoNgnAFcVbTDwBHA7dB+glYN+7Iyr9
Q8iJTPQtQ50clnOIwdSaHIwR3lKwJfPzTN/9hYx/qxmcZ+El8hx3PWERZ68vW3dK
XUoi7+Pj6msS/7vAlu/+RqI5/jefkaXXOBdM4pp5MToJ7L6F1K/lOjyOsgTB46pJ
d29k6VMWi7tCBKJig+BoANgToOLJPyzQeb2TSg7U2OgljEBAWomSNnHU/UDNhnXI
y1AX8XMjTXC7qyh3ePt7+WrJCiIH3191o7D9xlyKFRy00lmV9x6vH6hK0E+n2o9Q
qTnZjXw/vD4TzeJP05orwtkTAUzs7f2MTrTXkrlYwFmtkE2JHsfac9KejwV+yTcy
yXJi3bk4a7WiKmFbAtAY4WKmNJFKq2mdQqNLrANWRM68miANRVQfGKAS5opYHHOA
WEdO5iJSzQsk3or49eCqgajI/jdY7h6CTLCltmAXHwsVr40UsW+pcBZjSf5txx7W
EYHtHjGIaXNYygpD9xWOMbVHxM4D6wGtSAa7+FZcrWN8kOowCttwqjGxfeDXzlyp
gyhIU//wZHFFFvkLNzMUglnx7CQMvOfb+D/Tq005M2rynUfM+2wZ8b1gaVY42dm0
UXAgO/5O2TTK5dL1Uw2C6BkV4wp7kLnqFEXL3bm9lLVWa2gIlD5gVMn82pYX8LiY
IUSy3Rh9OMa/M+Dz7xurtCvVnZlS7CS9ERLa7YeLPDndJCwidwVHloC5VADAuTcX
OoVy/9W3C+N3tsVNltwhlsPUNxq1OJMgRaCaOCChMNWzRpMby4X2EbNnDmw6c5WC
2i7Kx1ml72gambAJeRgFZJyRjGZ331zMgxyC/x84CVl1bypT57mtP9R5svJarglp
A+IWY0tOHDsbIljp+1XWZ+hnybxKoKZRqo84OtonNsdskaXPAk8QIuSXGJqZoICo
FdcYri/wS8Ff+BJgRHjn8KQ68x4AfM4YUim86TPIJIbm852Nnt7bUh+9usxaKHdG
mTAxZ1zug8BaJD1owdAeH/CK1DH2eEROdc26dE0Mz1DNbpu8SiYAG8HxUrPtzjX9
cQAG2Dsght9A3v3+FHAIBIlf2e0RvYGj1nBzBWDMMArbjvWdz+ER4YheCnc4vd8g
OaA3yxHknHTPvmS/PDwlk0UhhPEkTXFzNtNGdpKSVye3NuyRpw5Q2FqSZbT72TPq
86HZy9JeqG3x5XYF9VbnktRq/2uKJxCucsSC3YQepzDAyqqUScmJaDa9QTUoc8Ki
Tld+pADjmorz6wCPelRsnrHZGSwmiD5L8CEHHkmYTXe0Rru9MQciw5zOpN4+1O9u
LQfNuLJfSmqFGmwEOOT+Wl/YvcoiMgGMXHKK74Xs/ARMOTn/ELTBy69OtzjL+sCm
7Z33XH8dJjN/k9kQtwRJ0Q6QH1f5yYyiDkSL4/G78ppIRLrxeTLtnFJhoyKcDEsR
nJBQAro2rRtfLxHUFRjjz3zdw7Z/pW+FJswNItKXE7Z2K5N29FOQSCVUe2OZtmmS
wC6MHhi9Rlm34DUnGwrQS0nET6HisREG5IgZThkXxoghx1xdqN2Ke+naiAuL0fTX
VuatoNSxTTI6HJIHJbcOkdFMGnj3n0rRj/+ncg0peO7FSEPyhnrRpyM6HXUaWAjR
Nka6WwxX+3aucbMUiIfNXBgYWOeelzy7CXrgjbkpxqKWkQlsAv0ZzXce0n8SSrgM
fAUca5190L0HM/9nNP6WkA==
`protect END_PROTECTED
