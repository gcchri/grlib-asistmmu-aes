`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pq7SBE4hTcvee7Pbr6l3tD8zuWRyhn1POF/Eu5qV2JjZCY/1beABBISbN6z8ZQjx
XFuRBUUD8AKVgxA7h7fFFVFKWj2B6XW6il03DRATE3rNcYDUV9Fkm8ZNuhYcaq3z
ysOQsGvq98q5Okr7eXrx1rYa0xbwcF+Sg+qW4e5fmXwJOHm4mOMLWbsyoV1EVbsx
p4dUaZt3akOfFekBq3ozAJRvU8yfZdoRY8ff5sIBN0OITKZTCTeiZL0oqQSseXsV
X/iOLCqCsF2GixwBFnRi4b4qQ93abXPkr4BWtiFYGfjgBBdUBKsguHZEGTPCe/ka
ozuJTx05cKpYC059g8QkYYCSiajDLxhfsFs9Wl+xNCyE8gd8LMdR+aH2PlCUZ7L2
ArgHXPvXKGVRKfKod7D1wjDBR2M723pxlpATl7inzldx3M/SCwmVi0uvsSM5d+V9
QrFTob1acGU7IcXdoxEWytvFcNefSfP8kgZYWy5HwojWecTt17Fe9G3h5FLtk4yp
2Yrqgre52SqKK9RRgZ+43zhdb93eEP3K0s4Z1F6Gs+qKwiTGm1PK+adXzz0nVt5i
s2eKXiQ0/vo9PTBw3SVtHKwmH+ehCotYu/t09zO3+fLrDItrReIssayGZKS8gBFj
knMStLqwnOtsEx1h+jyQLGUHnBAmDa2igFy/hHFl5/qJu7KR1GIacWzpNWX9SMXP
VZ/o8Ss6ZAXJg/gOfToFde6Ij+TSxcwWeMUjwlAZ/5wVxY42xEb9NDVDkvCh00h4
1J8qS+fpxrIUzGWWGwIXLlIjTsDHusUS//mS2Ck8L8V/oM4J9/1HSrRPgwCcK5QN
uO8t1C/1sFhWyj2isEmUVHyhCNAel+Q6yU3LU+2WzGEGunWitBbzh/pT0eCi0goV
Kkp5MdTRrYFKYw51WD/4Efp+A+e094dySsZx3W1SCBk4JsFl1gOZ3sC1QkRCjacz
2gsIqtwvrYjfHY0k4V+9S/MHc+yFN835PghhM42YHO+KG3JVzfmC1mr5RS3ZnLJi
fNprubzJmQ23IbYBYkj8Z++xDSVEgdmyJ7TYSCeayy4y+KuSizk4X4UqNYic48cJ
QGR7QIK4O0rcBeW6nwGAP9Se2cQsuZrWbe+a6uv3CcK1RKCM/w3QiQCqICZ+I/xU
Ig2vhi54XtNrVWPsojdYQg3wt1mS2K7324mPOPbveLGi7h8bK3LkKJq4IxOMTEUY
7Cs1Tvy0MChsTN/ZMOZImVgXewnsTh684waAbxt7xSY1lobjDVD1xA9ALOduQGz6
ILRZm7y7LoCT/NlWrdCOFFJahFwGKVpBZ1WW//UmHHqyiJm5duyBOkcX+D0qEukr
/t+hWue76eAkPguEZTVZ+WBn6f0K6s+1e8kGF8mjLOjNc1tDE1f/cXgqYPEmk9xX
rRODxPQtfaORm3RDPYXvaMl6dSZZHUOjb4wf4CVZM2YG0uyvfx7/H8ljIHI+Frqd
2snojOgAYVSlTLtliNGBPeinQx403COwfV18voeIEWnOUbAuvbuBrp7f4NIeSMEm
IWNG1LxwHemNi0JcQH5nFYC4LxlE1PjYrKme3rDOrlaj1bmWaBpzoIwHqXkPyope
yDJcuTHU39sbmYde2cNDjPy5jGyQ048vYUcI2w5xQkS4r2rPYiwVIxAbbzTvXNGV
UxuBRcKVg9MfmgJQQJg9yKa+7xVA1YLFz6yHvMCqfKgM6agiipjOOVI7898q3V1m
KC/l3fsoeG0ezIRqzT9pzCA8W1aNkp3omGgJx/U3eB9BSwgQTCtjlVhXcTv859VW
zyM7LuBwuNvmHc8ZWkSFSZPgaQmNl8a7ROq7nEsj6HLxQ+loMj5Ya0duoM1MOb+E
hCipN3ZP1dDY8XDcQQYZifQvK2kOK4FGqAlW1qMP1JdLwDp8Tmhpwuns+eTwPepO
+739v643Jva9pRN/4Hs+OD5MrOIuQBzy3WGuJDpEPxUeFHU+mz4JNtrTYTdW4NxI
6bVmjwfMp0idHa6dQmvwESLPA/mQ7KUzw//sm0iNN/2qLWvsJ2EWq8KxqIB9VrAS
/hsE1WT7f+RHxpXSnb2LRd5nzMwpfMg3CYAOiOVoK1GJ8ZFcdtFY4tCtxMNpZiFM
hifCPkSEgcj9PaZCUO2/Ky5n37ZvWnzN4rHSpC83O6oA9OM2F3T9kBTeOd6zcYJL
MQkyRSPDtHBEelBCZHkM19kbgQpN4FJh1CUh8V4GVz3IzusLYjMJ2DMQvN6XjkVE
R6jZp073hC924y6QcjIMFShddMmtcC7KPPN9nlJVaOCYCvnMoCdaLSHKWaIWPAlJ
uTO86O9aRo5n7rXdXvVLT7m/z3QD9FFJh/BNyI+Lr/k4NwQ6PW2CFIP4vGPN61oU
8ircCPqIoO+z96RlB0kNB16p2UbC6bz/cg1lvy0N5xKgnXHTavtaWRxHvAel3mHb
HK4ArmS2UbAsRDtRDxi//QkjuwH4h3H+k9VztIafhZqTSXA9dC0NKgpSmISkDi42
ZOFzXk/TnfqL2CNrb/4n0D2Uqo+Nd5dxTnYhaKZQTEjGLIYL7vmVmxT/3aER37Rq
oJMuZ/x6zDakGIeSH7Qspp3BkFTNqx5mb2eXp/OvRGXlmrJQ7plniyoRTQUfKtTL
TH4+nr+mb2gDeseS3sRk7JDdILPiFX1D1y3Oi7LWJYSoOE2u1yNmVzLFgksbxS4I
5ESTa+3U+qWDUGz+kRPPt2zyp2wQZKtJba1QvMYdIGaJ0NHwCsOkzxQA7tDU+arh
hjAk5M11Kyqyk9MzTMob97yago/DfZfQi0J5+BcobtD3olJN5/PxPAmyxKnsUu7H
JZeF2IV4AE0n0EKlMtsqACetA/y9KPSr1mEnSActVfy6loQmS+zMOrowxK3TVSb7
0cCM5WUIYB1DSK/kr118GoIW58qez7vhlnpZ9+B6piBTtLC5Nkr91HioN+xvr0ev
BrG4Wo2GacWlshGtJfqMQwG3B9PSixEnNONezFugAF+7Did3QC+UeKbnPIA++c3C
up2RPK82IXue5Ignk1NwLVJde9jVnpOvaECo44IKEElttfWRYaIlk/HVOY/cbbWC
7CmTAxf54LBI4dL5Ea2O9rG9SCFtEp/APbYg0salXNGQr2c4+Bjqz7CWfMPi5UGZ
90ENh4QwfrGXN5aaTiJlUw==
`protect END_PROTECTED
