`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dOxFu6YJMsEGaES9zpAaSfNdczL5U36bvuExw7OCKsSbmnNOBI9PCOi9v1KDipcZ
mURVMvqLA09HWVC7XKUucDyS8v3SUA1HBdKj+YHazrRuWbu42VEpbidrSkwQd53k
BH7lP/7J9D3XvWJbwZI4qOJMZfY9GlqcV57GmOLH8u23qptyVFUNPRjEWdmDQcWh
gK8Ek8NBqpfj+tizaQkJEBhK7KDf6j+Au6xxpphJ8TSJNsyC1MtPBFhuuytXMN35
B/5fm75noIDbctHPPvTsI9IY/sO5QN4YX7/7ieO6YFHk5T/9Gb+7w7SFO2yKpW5Q
OTFGwuVu1Vds/XWMQyqAtxGc12VYthgwsSsOfL68AlzQdheAzfPdmI75mNXB5I3/
LV5FvuJRBI0shgpJ04HRE53v829fEtfekiHvrHWMAuEIXj1vp2hvo55EtUB1o67Y
NdXXXYi7qIwF9e90v3CHlWH2NabU7sWoDw2fQBYgmluO1rFmE4yPc4D4+TVcPwtU
ViH4q3Tp61Umxy1BjmmyF4j29EzJn78gQRn9vGJmpZzeOLhLY2UguQZK/VlZ3uPc
fATG5HMxaFS0GSE/ljGYEIDu7QCeooBfSSRNTK9N6SuWzwZ7fkjFddB5Yub33ijj
BvgA9oPlT1+0LFoH2qqP85c+RiU8vcp7iCuIaA8iEUIECY4dW9N9l33CXozb1TNX
FsIoFCujoHIxD9j8CC5UdRXW3S/0CYMmWHsEcMBNpEP3paoJrKaYoBXC1xvX0cOx
XyBu/kFAiLgRIo7oT8fNpFjt+rm+D0aGBrflMVv4JuPKCNyGUbvWtOWy7QTkfvYX
tErHZ+GVOZ2I6Xjjyeei2H/Ieyun9x1AOH8tK/7yoBWO6KqZI/oYgFeVAtbecO3K
btykMA4HK+wbOU8udVVTnelwK3HoLw4ky4daXvZ1gnmdppo63wWJngTHuFO8LRW6
PCa/Q3Asn2MaD8ZrPDjnyWf+Z/idQ5aY6EVGlnCPJwpVTa7L98HzBMdWDIGT8qys
sZ+tK2/jFUTaQkt1IXH1+j7TyEHwSxA6a6rQFes4kF4q8J+Kyt31uv8ABSYq/GXY
avhbBIDo+Spg0IIreCE9g1F67cTcJciZLOIdVwn0l0umQY11W2lohrDJ8dmS4+e+
+je8A7+Eeu6jp5sVhI1RdxbwO/Rj+ft9SQc4+MxnfPU3Fjlo6+I52qKnBkD6BJUo
+9R3jzknrUOVIvq+EWUqKdj7ds+a2B+QtlflUGkdrOd4s3tRasowOkNK/QVQjcLY
uoxCHj7ta8bC8oM6WV/llGQblPrW9OrD/ybnuOSz8zUB+EI5eCGhoJM+JddNNAFY
v4RJXLUbAyVYCJWzlAoyZw2LLaoAphPW2Z9O5HuE/UnNWwzlYO9a/h2eEZkfzdFa
9RmfzvLovG8e8kDbbVDerltN9j1EwJhLcYD3xboAY91faZ5n+XTrezkZVWYu8MYC
1UJc/8QjuIAneKkozVW0pkssmgJAcfprupgftZCIHr1/ktDa6VxqZQvbw+ALkm+U
7Mt4oZRCLgGIphlS7h1JUMeOm2RsB2EVydNLOvLQeHgC3/oQTAjyCBw8jOS8KrUm
TTENmc1gDfyAJihQHwcSeCXUSYDCEhMu8Vtbe66c4x1vviHl6uvoxD6wFglGG3kp
xoqrmxoAdaPeDQIkavXjyWagoErzdR5zouZd5qHyKH8eu1sD1QVEGyOiLY24lC66
rpEMrqzujUkW9D4+5VBA4pUvqiOTriqqWrm99vlhRhFRM+adBFrTc+au5FrB3Yud
gD6Nc6ZJCllWIBAZjwKF3PsTNCEmQ83UU2fG9M4giLgzHkQVKfr4owLe7PotlP7t
AfJLhVJXBJjlkVfitJGCMja2OJv2ItlUEkdLlmMz1Csrf19EF6N/dRoAuKeS9KiH
bPuml/wj4Cul+i88nlCTixvPAc++bb0jOLTUzMrYGJGnGcjxeK370aldfZyLiiK9
mVMV2ZZd+sGOYkjP0/lVXAwNvxkwD1fRYY+M+plGleF1ZsCD3VzJiRzCEUa9tP/9
W3kVJgy24gjsSlfCMIyqNZ3LeeePSVfjaoQT4ooZKjKVCeMCZomjwcGM2kPLmfoJ
GmAc4fqn35jnr31TiXcDXqLCkjg6HUJCDxFqzumVOc33gXr2V+TVgLmjqoA4L8Bm
oZKQxWSf4r7O9oYcDo6sYyAkI919aHpKDkn90fu/pajHzpPtZbgLaDn/1vhe+8A0
FxDrmod7C0UkY6/o/za8IPC9hX4CmbySCzltFcqap8zrJ6k94VmB24a6JhrmDbgR
bfYbUHku5DvuWLyY4UjYzmSkzhhblBNEUESh836Z+za1K1hLauzEQ26TndLDYRzB
PI8kTc9Mvf02r1VcoQxeGzCjhpeksHT0F5UUfOPjHY2EhfrTFbYiWn+svfvBHYq0
IT3ztXvFIHYEdjYyMOLz98e3QvuAUT+k9nAjfCOwA0tkDki0Uh0CJqpaOJ/PJx9v
eoCB3X0OUGJadm9ohjQIQY4qFnv+zsWh2dmgj3jk25VWILpa2UuMzF8g5w28Lwme
aydduPLYOjbrGCvPSnkcaStnweyz+bXE8kJDOK5xgNQ/dWn41G+6qb42Al32Y8vG
4la2Af0Ajf+kLA03aT9BvG7uZ2QAHUGB7MoQHrKawmS+OaYRB9B9zxkutUe7wOjQ
ikvAy+ymJ11199JjPN9F7V4n7XdXkGQ5HkJ/aCxqGU3u+lzKjkV0kozWUzZwDpq5
nBBusi9/CFBFquM+zdKB3V5F0mXln14CpXdvqn5wew2WPjKo1CtpP3gPXQsy4WoJ
384bovQFdQ+3tSmWS2fN9o6e1VfOg72k33amKOu+hEu89xqsLAiyR6Q4oKK+xuQC
3vcJkofw5eKKMXQPY3Nfk8fFj5flI4DwwQMr3J2lQG/mcll+oCQiZRJ+TeYu+51L
W2aoy7/jwDFEcVch6RKrzA==
`protect END_PROTECTED
