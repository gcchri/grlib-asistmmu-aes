`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
doqKq7oS+VF3qMydbb3BzXpYr6geClZdxD3JRvxCInd6JfFFueL6jaQphMeZUoZM
DWcTXY+BifWCYXpy5MPt0AgkOvSqZorOvCOJutL8kn+UwsGgY61rMKqlLyXP6kkl
PvgIfy46stF9e4S8sW+0M9VhfcK3Yp+Feb9a49u0aPSsz+hOI62fiS+YzFLzf8h/
xXKP4s4VVOqqqK4wKD0pf/oJKIu3VuYs65pgBS4HBefXDsAZ+lmyLqnhFOEi1GOb
vuFSrKtrduEfwFHPLjKHQCx3QWJtAJXledt+R0LU01yjAsTLbh31vMKuD61c1X6J
M7MwgMDlPUC/48+1SnhKR2ggC5LsmLaMdR6vclLGga+sUToZBQZAWCk+RLV/aQdo
P4GtGjTcSWEH903sMkr7OvAHeg3Rjye1RoDXa0x9T3U=
`protect END_PROTECTED
