`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ujwhSCBQouhZbKQAnXJE4goDU79YHy/QrzEGXPrFcUB3Suk8esF3PAEYUdQlnzy
qAueFtIMJ5eMSZcofg+vBUhfb9gI6xbzji/exeHPa2dOY3A7afKc9s8fp3zeFojb
vCxra3VlBUfxVzmPLxXIcMPxgyGk0//KuxR0JF+88MFSdcwbkayccLsx1F9DDAfY
4UPFnjvj6+U7i/nZsmhGnX2M7hUfm/neGEJAD+FdCOujh4Blnk9rxzfeQj8AUwsx
UMvymzUPm/Sr2lAi0zAH5NOx7trvp8N7sOonw49uws2lFhkPBSeEpajli9NbaHSM
`protect END_PROTECTED
