`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A6d4+K4er5vtdHEWHLxcFKeMc4IX/psQrDG4rO8PceH1vU9rn0WWDO0QrQ5UnJc0
pVIYskcpdX3nnGH6bL1IirBPiRaD7hFOmm7f6JuuUkuBZPbN6Io1j/WBqTw1NxcK
4pli4oMLm+q8hyeDo21XipR1EqotThUMeMIG1j6Ox/dpPA5fvttnIg/IMHF/ZBIU
8+Tq0uZJetxHsdhOEMshNRyKKlVlsFPjN/EpWrCmzQhSI9rBbm0iJ66h8oHPnpJI
io3nQ5InlIhxghF2FcMX54AxS8MT0fnZ9dWTTvRV97ckITPOTWzayoVPB8yWW6me
tFxsNBffICh94z9pGf6bkSiDEJAuwBvwHTzJpSF3q3w3yzOV1yNj+uAtPiNglBm6
vQGHyB0OuSiYpWkEGOt6TULOlV/OuMfHnY5ZROdnTrKDwVFA8ccVpC/CSN+TttWq
QvM71KmY9Gu08OHsUxz7vQ7BBdZQ7sbGM5vKmXsEMHHAsFbtp+C4mN55uRQynpq9
Jc3/dlvEOfsV1+wsUV6IkLG60I6zrtb5srq/dkEuZ8IeVY+7FfOjpUisyxiFOBfN
KMULiCIxrOdLPfzIW8tWOiJZTcL7evYz2bJ00XPXuh6jDjokQ1i0WPYvp8UQZvC+
IMX9Yrc0Ugt8QW4T3ZejqQUoHPCsvgd4Jyk2++2xQefGwLpRLPgEo0oloeToRm51
XGG7iT3pu6/SAORs9rLYyqYjQum3brxll5XnUqOk6Rj5NEF9g4BgiG3cDL5yeH1E
nn8gTsYAlMqY3+MaG62oW3wvjKC25QNh8162Kt/iqW+pPC8YbkN+X2XOzMECWv/O
kLHYQTZN/TF6wew8BgxZLg==
`protect END_PROTECTED
