`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JlGYRhsrTmfenRKKGMH1kcpMFBv0NGJCjr/3FN1Q7O9iR80WEr6JvAmSjleok4aX
d+Y2SKKuEjNo/pCGatlgNI3TvvHnoG1+02lAv62PME6Wp5iKnCO8/1EXpYIulFSJ
JkA0ByaQD+jsZobl2Ylh/lG8QTB1FLrpvy/oOGxU+0+ntGla2+E0kz3wu0FVJWYx
aQXecKM5qGNiS3/dEwVcKf3I5zJvvhq65r0D3SlBjuisfEmUx/cibs2yEaHgO6dy
VchTEThRivD+KrqMfhFIFA==
`protect END_PROTECTED
