`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7r3glPRiguMbmu9LEQyyLi0wZytJsdWsHW58m63FPYTBR3LJILGOAcapIT15u7G9
AOSmxN7FyIWPoa5uFGiVZaq9X/KeJ2RdlOGSeOgwkgs8BWHXbxtTqS1xxTIyucVc
lwQvAWe2vsjZQL7UJTC0kPWuU/gHjEm7o5K9eAxPuk19dFHWUSMNzploR69kru5A
z5l6bx0PgKBkRxFeRBIspK68/mZjBAkbCsSto6KBjmgbdsjXql7K+D5DG4kgxsLR
meOyIYBOLnUhglJYZrp1ZVwKAj/AoJR1GV63n6/ZPif1Q5bVDxon2uznp1KYsV0Z
MHuuMogRNIwl31E2D59cbSWn29GVvBvoMLTdaQoU0WLnRPTVPEOS6ZJD9NbvGyt7
ZXQuhKNyQR7yn24tfx1F9av7pUDI3i2RxDHMGWL97F3gPXSB/Hwlck70qN3oZfIT
ANZSzFTa5ERBl8xoCkmLwARZSOfiIOyg/LQvTGWLGbn8kJtJual0fp0jeCEwCNkr
1P2D3dzotVYq1AiWyHhWpyCyr/5tWMhn3zJO8USMZYU=
`protect END_PROTECTED
