`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qJ1vWq+RWfOXpuHcdhsiIex2NRUPbCLfmixXiCSut1AzAEwxTTvGMVIz29lSCYBw
u4RdCcDNGcZhWX1zcqqXfPrfcz3K/svm8Ra0wpzD7BzSfsiwMjuMxUkEWbcLSOeW
AAx9xFYXdMGRxKhCeG8vrzJ9/c75OaZnPrBPvxctbgDZwx8c/cbFdg2gLf/0ljTh
ltf8yv8AEaK0Vx3FdKi3RJXgBKpryOqDDwoyTOL9mkjpTHnSGPQpQECxfiRofCt8
6d2D51K+WofNQgClLS9tTXXwcSnfq1BHuSlAA2rO1zxpS/oM/cyt8cA6nno3B1oI
03ag9+7cqeXTpm3J/qmRkDbGjYGsfb8veK2KSyBHvoXeOabW0tfIGb9/8+O78ne5
+NxTKGc5UiErviuj6u3aKnqikOznbMG+kRCIw0WqMMkFy1bxaTU7ywhNcD7jaKpI
igXnZ9IrHxhfsEcm1qzFfYABRidjbf5KRBIry385tUECbNWVEs2aA5xsaQh62+Ew
CJtal5rJzRtC5btpHFOzxfyUvFh4YFfvRLrlNpz6gOGxFKMYkVNiNjNDjOXMOVfx
gqSCVBUgKJsCH03rslaNQimhOFI0N57SItkPZVqxjbt3e/iJMYL5w+TP5+rocyuy
s+lzE4VkGcBQOpOvgnEtPd7Z1K4akSzNtjUDfb5Db98Bbt2owJhJomkbtqscVT60
WAkpx3dAaasOAlTaQO2wvyDUr+WlZ71I2SAtvKl6zmiasfomBD9Wi3Qw5EUtHQf/
Mrqeddx7lypxDJHaGfsfMgbB9KUXg5mRCunPnv+KX21zD7qYVtR5bmdWryM075ua
OepCv3a5hydco1KuCT0X+DUz28OsvOGHf/vmYIOftEbAuH6rwFzHU4K0+TXmNovN
CXheB1EfR/JaivZRLf0A9N5INP4WhqnJJUZLe/ZWvp4oR+jYFXrU64tutgeCJjwD
wkZK2nTLcaVy1Dz70VD5GkKFnScjujoquWyAKTtsvKRer5DVmM47ZTnb9jTv1hAU
1h4/kpK8jpgZqkSjv+K8k+z2AVPavHOWlfZnPAf/qVLuScT7I9GMu/Wqb00XKqmm
VY5nkCOAtz6+mRWvtyCke29gbP9nd8UcuXjR7dnu/5XAXvvQC9jOzWg3UvgCdYop
SoKwxjhIhXnf+gKZDOZ0T3Qp1Y4Ndn9lyyPM3uRtXUw=
`protect END_PROTECTED
