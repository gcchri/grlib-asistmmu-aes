`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VNsXyCl5+1HDPbdaYY5FV2GU23QxluJKPZmWdc4P0NDf/NRMk1kGm/fx0AjaA18U
aWW8e243B5Es73jAWiGhy+D88SD7cJaEM/xyHIbQOINK7cHwJ2SB7NdfNlIsTWZ8
Uu94TE0zhHp7vIJIB6cnvb0HpUOA4fJqX17XweYrlOKxlKZmmgqk8jHL/e72jn4Z
7lzsneFC9iLINkbeiKjfyh5vBG3uOAXQoNmrj1vwPC6FBwd34e9JtEaSuipymXSd
8cZzORg2NbabSow+jdnnHundstGonwbmvo0iBb50UOhyjExAIqZhYtugJeiti1Fr
p5IgqyK+3jnmvRCK6qP83r1dgxTY/bO0fRri8boMD8xZ62Q739Vlw6SDELCbjkJ0
BOpltioVSVssd6hPLqs9RgooCO39L8dCLM9WgevGVfbDOqGV+3KdqS9dyBis0/wV
`protect END_PROTECTED
