`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UFwopGDI2FaUsy3GSpR37WlgtIWZzvSLY8BvV7COOqVV26NVBdKKL4cYqc6I+q+A
i7Fz5ydLUIQrw2SI2BTWArRzHlCW+1M/UFiitWOqMPDvaixg9F684puLqRDhHjK+
UacceWSgwKmMdjQ3a5gUZ6ZUeI+pQBbRrCgh5xcVFHIY/aK1rN3rX1k8k8dQFDT8
eTSz7TUaNDVb24HqmWa2e/BNAauiuVGG0+jJVkXafTN2q0xVhem+egb/N2/V9otV
UVPQeoAmbKqKto1v6eoHXzm8G1aXjW5riydkY/HIZA/3B/w9o+BCR4+Z/H8x54gW
2LxTyeoQQj8uUAVIyHxpS1it6pH3cEmHORaXAPNjTSBt+lGzHiQu2xc/bnRt97r2
tFY12PGMc0VusVk3LEYGNdu1iiSS5uM/+IIb8hgaimbRkYB1+OzEuU5vFv2P1Qfe
noJQ1f5VdpkgUGhGKs0vR8ulSdMbggZYJhu9TROb4PeJFSVFdhhzint0PQsCtBYY
nLAGxwWW6xCXF/NUsjxOalr2+CNVWpJfuDmT+ohaAMVpgPbCQ4oraUfQ+50B7uzH
QBo2+ZNdU6ofZvN0fNDSSnvY0aCn91IBRps0ClfzgyFZvNtIlguvdpe8UgEyWQYS
eJbrxNVAAkipAJhAxYUBtCReHLykv0qQCfEU9fTpgB1wTSWbfTy2Xatj1QE03+gX
m9qr+sodbGAL+Wd0RpKWWLwBx+QSfNUwbQpjiGBqW6xJWTU/4jqL19IEt/Bvj4Nb
VcS4KCqsMJo4WI611HFK8ekGkJWdJdJVTYdm3oD6kI/GCzEtmN1u2jWhAoWnFPkY
YLGianqNaQ9EOSPh9nGzb2/Aq6q/b+qpxy04SH6cqAGAnEJGvH2Woug5zd867/Wd
kdJRvbUYPIvHK4DRBFL+7V3wrhrm44ghT089fX+92XWpFjVhvQIFhHZdj1L0Y0Nt
09ilFRqpSqN3Y22xsT1/cop7kTjor8wowoR46KQssHin2RlgKgDSNKA0m0YMCwV0
NfDfgx6iw/T6Ext/uvAyqgKrczFfAj5VByIG9W39Mw3FcoNTWyQJ32gxvt2/uz6G
FNHvbZZb6tYurY9v8hNwLt9r24WmgLG5YQXORKk0KyYdy4qfH05Wq7msmUX68Rux
hBaZyUGSxXJKbK2/ZWkZESV31zOTr75AJ2U8IqSdPpaVvMhXX2NeTzU/zP6z1x7O
`protect END_PROTECTED
