`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oDmpgN27TlLmCXmlhZPBf/XBkXMjLjzy8ozJNUUj7DKDn1TglQZYuJ5h08zO5CdM
slMrDCBP1BFvzQWXuxDQVeSDqAjaJ1Vqjt4g7W82Lwer/gFdTlKCQfAMf8QzZDkU
iqks07b3rGVLz6z5+c1GGdrAgnrTUOdDhBrHTQVrlpZUGyyGtKjn/kC0emf6fWpk
UJX3aZmMf25KknVtPXMmurvUUF0C432S0Tz0jNhczz9w/CFpO3rN2rcygAbe6/0z
MycVVlRbYqS8DVuFI2hCnjO+krUHr7tqDbebXwiEQAM=
`protect END_PROTECTED
