`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lAL56ax7Ny577uBEDXiWC/hHCGB/3CLyzSAcqEXibuJRojbH9CalY9r9nvy/FpJF
kqtMuatm377GfoJBJXY04wtI2Zw9xY+W/OEa9Iu7otQb5pD8JMY3AJ0iy8P+/HPD
+yn3PkVKsH3CEmJbgQT8eDYda7TBhbkb/GkLrJtVOUnbuhBNY3sZSaxyKPxTGJOJ
I+u+6uTnPcH4bbGxam7veaXIzhwf619hva/hiwdD12kliQKKkBuVmzPg0Gy81MvA
BHCEc0eyWd2StZn6Kf3qQ5jkrvhnU3uoGBKdbofylX6B4LbBqKcvt5kAanmZUzZm
TQReHrdykoN9hANU8Uxhm3e143vPK8jkZjubSNLtLdEKGmzRR5nlF19vX5dzfbNT
cWCye0KLC9IKCo5uj2jweGsk3ICcvmwmWhi6rAnIbSJV1bifCJc8OSOCPNbbnIHZ
88MT/DccqhVGVF+OgISJhyifJX8QaCNJF0aZBHS/JYBMcMqlC1LInEamH0Oaif6z
`protect END_PROTECTED
