`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ppaTBoTaZOy8hGEj8BRGl4Slsybgcj4OyDXZtBd+HC4vZboGa16gzvpxXz5He5zU
gybaVAbhcKaB8V+iIGKoFKQ6ypqe3F99Y39LD0xD5XoyZn4/aHQnY12mm9bIaWna
TJCj17OJFYi7VUKV8jv2haX/55oX8QtigPRAQiHq9qUZ5Ts4MwpttNjSDZTfojgv
yprhcPNcrH6R8xwfAA3OyWP/YYpRgYiG8YxA8Hpc8IbIgt0kgVpNsCepwjST/a8z
w/heBAWWilSV34JIxCHAS41A1OGRdniKpZzNb0A0SiSDYzpNz9yYU6eCcFEO1KDu
mTObbIGg550kpV3kpJx4CLn0DB2NDHe3vYBAAalRwi09LQ2k7Dfxrpj9Kq65NCVi
`protect END_PROTECTED
