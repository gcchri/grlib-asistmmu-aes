`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hjfg0Va3Q1fqQgPobRBdvhNiYVQXqfB7HrM6ZjGGn6ZA6PoZT3YkvKQV6f5GovtZ
r0jJ6Ac+vniRJmuaBL2Ubh5LqjQWsdcyldqVY8xhJaikjLzg9AGacoYH/zHCxlr2
RfbYnc+9SvUc4JKh0O+CK0ekENtFGKcXbXqy9srFz9wCF9wyngFastNylecdTzJe
DZcPdIqsI1F87pwJk3zdyvAC5jfVtzYynQfujsrcjvbnCrT/nQN+JNGzjp6WGxkI
L+ljT8pDs0buWSLueMAQCNHYJV6egmOmrTjIN/X6euo8EiusGxBosemFbKw1C4nN
5AqXtzS0q+RzxlyUGdDEpY23I69ASfDrWiPallh3qQqyNf5TApqfhfKOpQEK6WUT
uFuYZZU71xI/UnFYjBDymx+M7kceNYN84V9OiuEVAGTrY+ncFYNVqtxkViIqaBOF
`protect END_PROTECTED
