`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Q+iN5cv4/n9nEKW2a97+11Ef/ys8HTC2UfrkdIM8fghDPowah3NN+45WKY+20n9
C+ImapGtojeVYu2/MBLEHSdacRmcWEShy7CyiBdQHrps8mwQ3xwBfSDYDVOP5lp4
vZMhgA+sXi819tJC/933ZgA/jWbwiLitjwD7gD3Zlnxo5vpjJpdQuVp5AhD/hkxt
qcAAo2cFUbNyxQ3udS9BY+YMMenwNuQBXeL7V5h4dm2KKngZQJxoPmQDxOBQoiuL
l4Oryeze9bOjdQB5l/Zm/iVp0dB83dUWy5mlIT2YsaxdHSxnSIir4zKjGR8X1I3w
NmEziAgEBIi9msKAEsAgba8Q5+WErjx0qRpt1e2Q+HwyZ04/rzoTSWC9cKRHH1ch
kWlumpouzZDyXcIkxhZs4jZxW0ooLeRvxhXj4S1yUMKWLt9mOtbc13uMa26eZ5xV
mNAXFR5p62r57D6AMB5H5/jUsK/rKJwouY4GHErJGSY=
`protect END_PROTECTED
