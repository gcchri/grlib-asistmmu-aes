`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PgoeaQQ5nAUdHhKWvaNhtbcBLsRvSDu/zqufgV3ZIeP9jEdjH5oFYv7JD35XyNgT
TLe7M4b5LWleTrmUMrk4utm4I+YzkkrULQ/pDhAIIZn0pe8A9Mp9yR2DsnHcpM8A
9BPg/hFeKuR3XLp3O6MGJ+fufpDKzLTpHKq6gs92vNj+doXHaAJ9vHB1P3ACPeCd
sjt8Fkc+fX8ycJmwHrdNszQXESsEyr4gkRPLh5ZQRXurhGuEadbblQ6EDtXyOmcn
Q3iyMmGuBNQt8LM3UDphxzGQqcNfJ9mjFlp6p8oqQRk0i1EKbEHotq812RjlcVZm
BwduboByxKVL3DCrthkcYOSh9d7r2xXUnoo++xoPk/ne/MV2h0E4NhzbgCGl8FJb
d8kharGtckldS1SRkGnjYWWkE+JgXXW7rF/0gU3xxSik9Fon4IRES5N65rRC4EvV
`protect END_PROTECTED
