`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PNSS+dAWJITAshoFX/V4MJduZGjgThMGyEn8YU5OfN2gOZTXIy0YbmC8r1seaXnp
9RtQkfUP7QpOEGHqrLkwx/iHe9JRL8L/ryjUu9dGBf/ptXLXADc1rtRgoKozJWNP
qoiZaZ4MGJLKWEaFxja4c3QyUGOKWb1CCFxGvCuOoQnodKL6ZhsxUEVteAB7vVF+
gZSo3kXVOR/ls6Geqs8n475MRhALKeu7sM8NsmXEe3StwnX9GOfTbOFt9SbuX2DZ
hrZtH6smu5yG3Jl+Axl6G456Hxdtv1QgHMUEd1UdHeaFZ+4OMCuOgejphKhAu2r3
5TjhrY7d/brH07rGBOZR+uXuUXPbdvu2IHBQymAc066zWFUq6zvnEULHRB0V1GyO
yBHAx2Hiuqk4cBJKYxpY4g==
`protect END_PROTECTED
