`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qfYjXSAMNRbKc2w2xG1yv19lBKvakMdXLNxTPFCW9fIpDk9+m9NXacmdXclsRNmX
VmysLGcVVJgAE0UVaBjkDcarBf5dCsnMquL8LI7W/OFzKjwXwShqkUD6+o4ftYwg
XMz1yYS6pDUD7eQcJ/5/nbrmrWDgKdYc8ELiHtSFCr+EqFJ+z2d5E5N8rmj5a2Xw
5Fz5W4CfGQuhFy6BP044Sz8ysr26jFx7fRW5w5ti/rTKJ7TOrFlvcA6ODwZoLyhG
qKYtSmyTvIIn3OveIi2472J6hDZafBIxsTwF9Vm0bZQ1hOz0nTbCRQlcjKNsxbBU
7mvdEqiOIAWack4a0risBvLJOjdcw/61HC6lVhPYYd9+0eiuYcI69qdNCuajryIO
mjgfz1zAPyg+EKIq0oS8OtTH5Zv0XlARQt9zP7m709O0/d8jRubhVrePCzHmsDqX
VgkN07JhD3di2VcvgLFi9JqgMjWqik7MO83r2XrVoiSX+8uPQxqIeMZJcHjVbd6e
`protect END_PROTECTED
