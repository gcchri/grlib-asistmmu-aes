`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A9TeEpO/SVSuNOYI8Qkbb4717Nd/LF+zHYmEkFIQoJo7cRZr/guaZB7E4DGElO83
z1XRSSGKb6oaOfdA46Z9qkV6MOS0OI2XkPDcsXSdg8vQX6+w4aR7dWOPTO/yt9sO
Z4cV3k82LmlMV/mRq7VUElsFTR6Q3Asdm39NVDfdxeYKNgVNXXjU4H5k/yhuu+tg
bo1IOcpofA6kZlOeXhmb1iXR7HcXr5tupNGuF/1+gwRcMNv0nsNldtX2JL3XWEz1
gRLHjb2hoTZRwc3teFqEaUaOg1hEn5E0nhas39+H1jw1U+WcVoQDjjupMr7uCfhj
n6CCblV2p7rBXW/heLPttPXibumhHg63CPFJ0wrPJDAxMiKg1g6PFPUKgn9BVd5w
efGY/wc7AHA+/1ePNuwu4RxK3wHnwEJ7O92WGz4HlHxumsZkldYk7D5XT8qGAtEz
`protect END_PROTECTED
