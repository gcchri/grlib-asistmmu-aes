`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yg48ptDMMwgTkajvQ5IXFyM7hfocOTp5GESPPwIRuvF2ZuiTGiBagAAeqLBg1R3/
KZeQ5RBITn6k4siLGv7n+kpI2yXmFIfgZlDYAs8hrA309DuPFjWcQKweVyU53/x6
h1+6m2AmhUg3CjDKjLjUn7S3O/ukaZlV6mGP/fVWWpsi8/Mm8rvEajbxJtbpTppl
HB9mJf7EDWSCxwbkpS293sdn5qIztE4Z3tHJ9bkHrjVg8PM/3Q8qVwhqemliHlVv
R5EIwR0hmSfK612RK5H2kpy06XCPGo3eAFjl9kjeLQ665NsEtgMzUWbeYmaCvbvu
mq0EZmRw/qJIq6qJOvJtl4nwMM+PO7aMZrc3ssM+FjiyermfAYy8sdcY2oi6iJtj
IKugTsrp7cMvvqG9cf3IQDjdS43PMoR1DlWwixlc3FS2nTRYU1+PjSiZle/mViF6
LIM6SMDZ7ekCuKSkgO+0ZP341wLBVetNGXCgypsKZt0jT6peBS92ywcedb32sQ5q
6Ev1V4D7C57yYG5LZbSZbZ4NO1TiR/XVgROaBiEtK5SzCsqoEtejhRyKhgLLtv0b
hYrdCKDXJ9zqSON/Roj6vdyOZJxTxJNQs/fWdYhXdiyAMQwbK4y6kwNkY59LQaYz
pfGRsUkbdkEXPm86Rfh2Cr2lJ3PF8GBxs8bgK1UTN1LlMb7kh6My5EHDdMMtVa+W
haREhi7y1TOuT3VONNxl4xPuj2Z3Um9MWvdqG2M4LI7rDhkUZaiP6WH7beKjEzM7
lKQxJ9/txbtQpUDrmn3Yf1M8Iu3dySK0F1Th8AFXOkL12SK5KnS2/RU/LyFWKs3a
8x9czCnoU3GbIHNflbcwfC2XFzJNilQi3HAQD/pUpQrPBd7jJxZL5kTSB6zecuA4
EOCeWh2RnUwoohJM9VTiemH6bYLdkBvmBMa685Tmt0Evl2mA9EmQYCpQrjLHyLYm
Vw6dYWdinhIbWg3M4JqcM1HrJc1F5vMGkQefRivQ57OthI5mmdengPPFEQz0Rdkz
zE1xN2rAzuLG8k25CiVUlzD1b0jqJvDhlltgjh4xFS6vK+BCIwMxp/gxmRepGiOI
ovY+RBbDEGcf3SR3PhDW8NqTmvrJlkMUyl3JcTqbdjXIlvTH+0jRnfbLYZ1Kao/d
SShf1w4B6vzq6pgMLHvf592FQdaa3NP5u2Tqhcr94ZmEJdocDTKuXLbDPF8mXdui
EQkKcZbE0CViKpXTrVlSwPEwzdRLxTm73j0cQDy1Ptk=
`protect END_PROTECTED
