`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CiJBS3JihBZw5yd9vQJnxmoqiDXPHYGCWEdjAA58ct6BY2ra3Dc7M/czYQVatJi2
VxFrJ5SwPf2TkKAh2H633s4JEkNmyORHy8leHP2C3MxblO2jypHNYwCKIFovcms+
W35m+FPrsqDXWa48lwzfkDwl3R96pgj2QkjBoRaFKVfPBSeTz85Y/10BXAC3dXFh
J97KoPgyM5x8V6ZR0AZUFyyn08HYr30vZhixgAqz/uSt0fBeKjbi0BQdrAGzpxBy
N4QOnpAczJSh2q+/cKNjAv64me9VcCykdmXWaFuL0Og4I18wxOpLhw4kT4BZCLuR
uFpNSiaTouYKOS0J8rEsQ1aYX9tx0ZlAIeiUiU5Y/LCWQ3i1Q2TqtUfiIA9YmBH8
/YzKzQE2utmwOBB/vNmIedCV4Ku4mWDS6UUpl81Wquyij6KcDgp7QTYhbmU2ef2+
FNfBuwUyo7QOKiFI8Du1jZxnel5HyVLJJD+X6vRrAheug3X0uPgkXNRa1bf/Zug2
5FaoXxL4eMUJerAkxAROgKHtFqs26YGfpb3290IwPg5VWE91+kIf4HU8ufXt9e3W
kiq5tU1yOq6Zfgej+vaeof/OjLpjf/81cdRlDoZDqVI+cyQxwoO165KAecdk8UVu
/PIQcb0ZNgeuEoeJwImp5Y3b+CwXzW8LZXWIJyt0w5mXemystuHpP/2L/Fu2R8vd
zBT4EHVX2XxWCTGLAnV3MCx61Dn2Rea2tviiuKRpVX98Hzps74XhxNAZs+OVTf8R
boGUenTffJGbm64jCeVPV0VpPOm0yDJKlnWULkpSrvk+GyTEX6JmfzboKHgYveWT
ynnI4L7CZdscKEAZFJBoHYaM1xIdmhEh3mkRpd+URj+FGgj3oAOa5ukN1PdGdpjJ
UvsxeZ/HjimGopqVUoVNLgv+HIkVvuY5n8dNMaXX7sn+QBOU4kSnIPzaKqm2QqMb
mtCOUm4gwBnIFRMYWd5Rchbhx9H4ayHlz+mJCJIbo0NlCNCo3BHosp/eVxvli5QL
M9FJFl0wImJJ6q26zpG5NEMje+878MydrP6Dw/PPVbpevIsCdLURK0Mvfxp1AMn8
9gJZgaFTiObSL5Y3zEOQm460OCr+DJGNGbN1X67AAy0aRIr8Fl7whdz2nEFt+t4o
swPzA3vmkfXGxlw77D1scfTS3HBMu2othLvxXOJxXA18FB8uf5s9OHiccMzxkWip
xKtkHHkZxAD1qfnmtUmupb8DAt+lcoGwIl0MbAxvAgT2Vu90Gt1AnhJsWuE7FXl9
j6btD8QZwXqqTaxGI6G0R2dL8pXLnF14Hde9ay3SGydfFTKo1/x2Qw3njjDUID16
0AjJalfwzbhn+eO/VV6pQdJ0FeR2KEy9rTKwcGUKOynJbRurBu8GAZ9YXS3u26LO
jkZ5mx1w7pp7yAvlIwxQvmSOX/r6TlXD9runte27PUXjIvavdj/qiKDa6pbk0AhT
KRBLQScbLBjGsSUVIFFbh5ULuGkADeQooLPKKCmoJjzXnfeAQE/aVu9OTZSEHXVz
H4nSkGL1BrZJk+yxOpnYBcEw0tG4IEOj4Ex6WvbgzkfgC30lWNm3fkfb0GUgZvXr
i3GUbGa0OU7W0nxegQQz10M629W+8hshSlDpClkmuojK9BRf5Umh/zhmBRYsWzzZ
/Z9cBAgeQ3j6HdrSYPidrZ/R31n612c2OMwj7n+EaeF5GzRUegrBD9vkuTneePWD
Jds2Fg/1RWb7PTBkrRn9B4UL4iyHKqh+j/lNM7XtzIE5BCZqFdfsmEmIojk1nvKa
p/ltQ+4sHraY8NEjj0UAUehDwNnBLsxUKPTvmFbyWEAPobNtTOJls7LDEf0lkEJ+
z+4/+bhNbluYiED9Yu4VCpwrM3E2O9+uPhOmVhETVfCg2XvI8iSSOPxMVKWSR+4Q
24EtFJRgCfT0+ZAD+sBHMetyMEX5GCARlS5G1qA787SK3taUdMNrcJZyMeKSFhil
Tikm8X7vh/A9hfgcFA3JQT0qLnlAto7E0NyVRFkkjd9oaD0ir50I05Dy2BxfRErS
7c52Tdv0IRci+fPOs2AIkesKCY/pT2jGLko5PXR/mF/quHm/TsCdNQVLI/6/VCpJ
zs4XE76Ios49gFOeMtEdDax88/II5VV4vedce+LwBhg=
`protect END_PROTECTED
