`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XFJMIW8Ctt1Xju7NeNHgHp0DKg+pG9c/hb8v7TzIXgGxqWQooxeKS/4eyyurmQOi
zH87MER7XLD2w+fjXpL7eXO1MDlFm7AUPGCCsNjF1YSjuZFoVay99rxiGKk4Z5xN
z/11a37YS/W+qLfuqNaRx/7e+bojedkT1VpiLiq+8FB+xO+vBDncl3AOslDnCXWc
i5tMVf+av+gIX3Dh3gBMv0x+wsWq4DdImpUEs/Ofy7LoGcX+hOTRHFvRyE8KyBMt
mv1bbVnuSJrAIXntfB7mc7Bv1PUWYZ5zSKThsbNItVrdVWZlFc6LJMHrb4PklzGo
N0u9gyU0MF62se390q1wRrlvcStvAfAH6WpXSVIq6pBc/obGRkRhazgfuglreWFJ
`protect END_PROTECTED
