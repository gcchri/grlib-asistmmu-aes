`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/36Swc/JNbePCRifc5QMVCvYQR6Ga828NqBhBly5ndagqt50btBBzkK5feCDuRTd
nd2oTuC8h4WeDfAsC7M6wT8AprYdqraJwWanZseIkBrxM9lS7Vf1wIeAGKSMh88I
oMt/z3/DEASVTnhopnhSI94hvv2KjflpyWU8K2w5rWgvvn5yhLgvrM+19U+seKlV
qFxcZTwQJhZkkRfCsVlZl2NgYrCRBWuX6oRQtU/B3uOMdyL6izaCnHWhCFxVCyy2
bsnlBqOzy/gn5kIF1Ytmks2GYJ27r9wjXks64iBwuj6pEuOoQep+Z9dUYKNgGOy8
c/9A5czfXbjH6K2EUhFEvNatItVWMrsbA4HqDTrCduU159iyJd7QKKmMbUCQ70hG
Yg0qS/45QENg/MDfxWthBnIV0l9zAM+ESL++6pYQqgmEpWnVMv2LXuziZVs2p0TN
Mp8Exc5zVIV8bFrE4L8Mjv9ziaCdjqIOBjrZ8NtnCTXqd7Y8vOphIZZmmabP0LbC
tQ/WsnTStpKJP0EIdojX855sM2yWNSzg2BmghIFkVn1G0XgxEQLcq5B75xChnM5B
Oc1snd+JXcF8gGg7mjZyV082aaYP7apR+yHYymlkA/lGtouHWCVZMB0USqOGROo+
srLa99vu++ngqV1iqU5PUxJcBKomOoD8CfTaJz99p5fsjtJBEvT2KSk4bAhWwi5p
Mw9XBbhYvio/HEaVrxNVuTyCaxvc4hPlla6YEhQ7mluolm2+PS5Pk78m3Whm4uAj
Tbv3QnFOolp8dE70JfAxdmBjbvGig/yZdw+uUp7k9VKF3feEAogAOn9U3J2mgSun
tiCOLnU4lmp7vj+GE0GWAJa66sf5gcF3wtBN5LYQ02V/xY60/5kOHocmAoJfQFNg
cJE+MmlqrWtrvTgsyirfAvImJUF32/zi72p8EnWImNf1j9/h2GZx98a9rm6hCn0F
LgLyrzYrfHkg/nS53CvKSh4R2ik1jtKUR4MraojnqaV2IIgSu0ds99VOHNE/UnX0
Mld2o1Wu0bHyPx5nwwkpAMkjoweKKa/0GhI7NUOvPpVePtpKCElWXNIQ1Xw2Xp1L
4ebO83n/zzGDZRPmRwzbH2LacTNS4F2FTypaixaXGdogIxffbdlbrFEW5JcRcTVB
DLmkLwb/NLT+/BnEuXrM1hYEAUPIj079zada66PIppHzYwhFXuHUjhiJDj3jpxb3
adDfhR7/RBlA0B+wVNI5mm5/ZS2y9jnwO5KI1+uvDF9tjStKAYrQswd2Fr4O7TDo
lhl/5NpdCH0wH92EDz3pPoPSA4QvtUKjuC+b95ovDlnTVUxVpG3XPriI4PZjW7NX
Y/QySA4QzM9Wvl01BOlazmdt00ZTGou6EksOhf0Pv6gh3ynLFQTEpZmtEecz2tBI
Wlg1rGUIARM3KHVzHKUoSCAhGTeWCJN+HhNXbOnhadCzYmu0wbHIQ4G0/bAyPRYR
9Nw0Dc/HH0rp5GlG/du7NS4/WF+dTk4rvuXs7tSc9GW8BIZTkosTyUgOwmRWG1i2
a5Uc4EjEhRd8mjtkI6apDa/D+frkSayouwB8tBUalOYkXwQJQdpzaBZjrkzPqD3U
xFZE3vVwQmWsztfKU+6SckNvyGvQfS/naZ4dIaYLR2oJ8M8uQfcgx6YCIt2FWctZ
k4AfrRWm2mVxnrJNeiEKBvm+vzuqdaQsmXZTkkBKELJcCjsVESavCI2wjQ9IYeCE
v6NJxCHPggb4XTnEODWxgxzN1csjKG00LEMevyT74KX1EJ4NapRdBwtNhgfll2yZ
Fq59U5G/5VYS6XQ6J8smU6vDfdzCVmuvG53D5j6Z1/RqXqOtozcxf7ZOGSwmYUzv
vG0FUAZg1fyQRvmPZBUm61/aq1zpLaJCLLFLWqXl6vxgtVAGRZlYN3QEfgkeLNw/
Ch3WZvkctAIlJzM7NLQ4L+vDKlkfhoQ/h2ScNCeuFKkxO8EeHsO5yRZ5A6kiZ02J
pIYUVEHwdznwD/b5bj6b81o5GO+9hnwPNLBUgM+4oNNK61Y3PMQR0cKOYyw4Oveu
SV6u0BARfl7ONnjZv7bBf6+UP7EvYO06Ju6mbYPzKgAEB0FoABxyHJbx/2aw7N9E
1b5Ai7dRHgb3/WsK5HRe4jfsOwVcZwtIDkV1PajPAYTCfOedeDZclyVPItWEXH+L
g5qpVdC19ZKVWTwX8VKWNxsyo5oVb5REpsYjvT6qGTXYHWFg1C6xFc5OyYt1PT+C
YTKtulWXAspb0Lt/2L6b8ngpWrxc2TMPT1OcN8T7j+PFPGrdvt4VzpXPqtHrTB5j
yMLBhSmxeMaGoupkxmLxhk7qqfDMJF7QnuAeFAEK7UUoI5TLbhaY5ArEGPsGkDBF
MGA6litCsryG75fb+MsH3NqjRzwyrIC+6RiFYsdYnSdSqbbRwA9ky5lyPW4+D+7g
UJvzA3EXNEQLlygyoLKPaRxvvl1jErrAaYMZWGFZ2BMUaLUo9nOB9n5SGCzVBzgm
rzfVpsEHxK3rkKnSmFskupvpiap7MOd8vnv0DcAZOh/TyJpSttPtGAS3WsCKEOnd
eEANlEVKaGJIgjGnuAUuezPSNhwrX2uAZiNgV5qHGhHhHaGFQ2hAiNAOeaD1TmwT
PxFQocEkCTcY5MraFnssLLTl+FMxoRgRfbtdqomK3/fNiZvaSgYq6QA+nHgeJBJK
+N7w1PQVlbjhYHc5Z3dDFlcjY14o2IpwPk7YE2WkyBXpC4tMyh/yMzfShQ2EjgCk
zdCZP8auMlpLQe78QcyujypEbUZU/U7DfE+Ez6X+vk5SyBcG8uRkrnkflqUUnStk
BuszoyRnhSXnmxgaIlTZIvmi++POpcUpcwlv7ZNWB2A=
`protect END_PROTECTED
