`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
15TXzCnz4ASJm3AgYQ/FQUGXDgMVmzp8Akiy1CBhsxIPtddZoUfrbo/23zK7D3UO
lP+V+/H+5FpzZUTZd0ckMyDCsYLY7Gh4iCmW3Kg6oWX6enZKZqOp8Fj1XytmRQ6L
f7LnMhFtTuUhNKf6HWPxIRe56CcUTEpPS3c+gNoRjMoRohcYN7nmRz2cgaSxYOeW
5EP0vpizPiRiu/7yGEfEXyxT990wa7SGH0ODJEQCQspTJfU1zuqnYO+0l/2ENrcJ
sjoOgrmd6OOsoaxNZ80CCg==
`protect END_PROTECTED
