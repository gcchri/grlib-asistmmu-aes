`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nwLmPaxk+gD4G5hF5tQ7f3jCebyiBPJXc7MUb0zuTR14qY060MX+I/51Fygvo6Vy
gm46GZMmo85MTBANRt4ricPrz3CHX5Tj5Da8/ktBTflq7ikBGSXDpQc+7FwJLahz
UVHsqWPUgBwkU1/+ePmGmTAo8VnMLhC9mDbJDvGd9mFwMqEVFhPvXBzwVoCAL1UL
7QP9Fig7TIUA3wT5V7151adwo2lVMEQmHpIJApI1+Nz4dVbDBoxH3POsR1XiawKr
FQX7He4smExalhk+3Cmqrwa/JUWLc0YUf6j15YbpCKtumH1usiG7I0l8XQXrui+c
Gj2Kt9FxVMxeDUgmS8vGuLiwnaDo8apoSl8PPHAYJLaG7UHw9ktTJlJDL5dwtAWd
SI5yFqE8j4pbGuIJB+2khHxD3Svwlt+3rh9hMpifPkahJSPEoaTg9+KjTAkcXIK2
GEQQM3efpIawJ8AINkNssvixFUBqm7mpDJUtDBWYazFxTxR1HUzxUMiVNrJtH92b
stAlvnlMExPX6i8O33s4dzUOtkVyrJVI33B/6D9xa1xZL3TRmORCThFhN+54oLUm
7rCk2nL3k4VPlewwkxaFwCAWBj3XSkYnQ0yx8MpKgXm1lnDibM3AjQJ1ipHMCwGJ
yROnH0VedypsZXzyf1DyknNUdRJy3mMoaVi+1M2irZyQZA11AO5kiM8G9euJLV/C
cC8sex++a5gbwchQ+ycyXt9YonQhWYPkaBestuyvHTe/Uy4ONlxxJnqAnO+RhTQX
y6umLd4P88Uk4+LRrIm+i00GK8G/6e4aHP4axY1iMNK6csrmE83hNAqBpQNGT0sD
3eloQBtn5ZAzCvMRYvcj+gLYuLj1m3IvEliY/1KJ14QqdDFOnyIhFA8u8nf0tcuF
ngy/MNtUaq7gdnfFqX0gda4T0V1rI9iQjgYejY3skW9CBpe7O5pIN5yQDwprYdPi
JxemAfkJAnKFQOWDDENt4ocsgA3lqVidzgKAim/zVSFOrhb3CHqFiOGc0EdwDMvQ
xkdrwXzuFEmk+NFjNB9uIanbLDSC9N3ihI83omHHnerPCMqkiSONYUX1Jy/WYmCA
qzS9wUt2pt23Bp2OTLRwPQkPbyrvynCLdgx2rmBWpvlpWhQfwep8f2wcggXXydEF
/KbbFnMryWTK7bnRjdYfcjNn25CY0vbh0r3PPQumkMpJTCU2IXQGb4ssScxYSMF5
OWDpRjnURTGpG7NJua6JXQ72H+zwMZtlpdYBFfeDeSE0WmAT0alN0pxzVEtyVkxC
XKnB1m0FYS6AUPWH+RxHpEDD9c8J1W55TVt8d5TL2asOY1/+6PLMaioHe/0bfu7k
R+SmDvcOcGIpDLzMQ+kk3ULi4K0IKKc6t+wlcK3M6m456oLgBE37Glx1DlfoRgXb
p0RmVCIh9X95/XlMA2s4BaTNsVWJOcGUaQ95sTTLFxCI33PFplOUkf6/fuXaVwQm
1/voT6wyt8jzpB5QkrfaV27ki5vD3eVdZCtZvqTQNucUSHeAkeCgrjCLdCxwnCJi
IetazF+Kl8t9f0hbI+GXzIRlvG2vDJkUuSlr6/Heh+w+A13CrGx0QIoSXjaS5gcb
FUGDRaJamYfPsYhhtrksjg48jZ+NUNteyBWMx3D+T43jR1ZLtk4N9B4si2WmTWjA
SUgipVAdwwPtpwvgbphJYYi8c+89IVHm0Vv3lqxfYjDGRRWmjywBsxD6ae76nQ8u
dDTKMrwmrlplplBx1ntt4EErLVpgW79LqB2zrrjAD5GMkzEjM5GHzeM9xdAttaej
NyZz+df9a2HLeAldKJy2jUZPfNc0BRaJzHOiAHMyaBqQstOPSVWnOIlnkmMVdbBq
0v7Kc7KWN0swaZJxE/k7bAZWlxxU55iMwXdX+qDc0k1lrsIYI+MzRsFj4AIdPkjs
`protect END_PROTECTED
