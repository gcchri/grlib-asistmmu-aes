`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rwBtDW4R9z4QMe+eQy/1ubxicuerQ6kAi2dlBvYDfj7QIxn95naUhVbTQXtaH0ZQ
FO32owEq4+m+rn4uyiSXV20m1mr1Y4z4+i8O8lfFG1wG1i4xBdqYXUqGJeOvTKAT
f+OB0GSch8I4rSLz9WBO1axLJfJs30LkK+tIUG6BUG8kOxbvAjCK2n/gt74GKOBP
YdM6pmPQ5/A9TcN53WLhAQWxfCO3kEvkOFjTusiNrZS+quxBWwwDrgVoEXq28u4W
zK5IbdAnurCCm/Ut6Caf1osRJOyVUpOBb6qEriBkpjZYY346FOky+rOx2G8iPWO6
AxtgNZufzHqRnsOomO3QHcIWPI3wLL+kyAUWkWYhgwYAS1/Js5JopkTFFvJ7nPwc
sw3vfO3/PCAM2OkdoilZjgIz2ejh486b0ClCaEWmiHtne/JKV91hHVz0M4BF4UbA
`protect END_PROTECTED
