`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jv/rTs64JyPHq+zUNU1LCrMYvkLIwjq7U7YgUUGfG+5pl6+ATW7+FLg4Hm9lUuhJ
W1nxbl90a/2I8T4338HhwjkvtrGXHfbx5H0XWB4YXODBC0BE+wuvVs12KxGO7Sl/
ob1aPc4YCXBLj/OXUINwFWKTZBxighnkEhD3xAHWnjCPT/Xw9O7hSyQ5c3g1lv6N
PJLjhFsoZwi///SqedN0L+2cpbuASqIhrl++6ZDcC8kCZbeMtswWXzUonTMYg4/z
6aDBvZxGPamYJ3J8WRnltsmDNkWOlhL7aS9NhEBr0DLpvsnGAWgl4xJIrMXpjH6n
3ZsI2nwkL9sA6+mMhe6yNAoZRE2KUrYJAY0jj1F4CnFJKoTiV/3jpSmv321afOfy
eDOnCJzFV1K7ORmCv3bh/juMq6K8oJ4U9crn0ptjXWA=
`protect END_PROTECTED
