`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JcdBGI8J/nkMsRZ3wew6ZjSVY5k49yyn+nB2anvMkVEx9ZeNW4isAwmpKxMUJPrW
nxNScz/EiKrJgVLWdGlMrqcQsQeg6MXZu6MZnma/EEwg+kj9glJMq6ODjj7anVyn
3oswkHlX3X2DiFhn8qg6blCiE2v7PeVPNVsEV1Ol4RmhPNS+UgnRwj3qIxEeFRxU
KxE3hXt3iiyEh6zPtgydi8hGwS2f+Lfs0Plf2smdeWFcIe530YNG0JkLMWD1IcHx
AunQWV6hx1S5hn35Pf5qWYA5YiWfB2QnFYn6Bw45xEzEkx0oi++mBVYCRcHSf4pk
kF2/qNFvDrhLyJHiV7p3Lg==
`protect END_PROTECTED
