`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JqjgOjJ7DKd61w+NneF/zQsPnhw51688WIEHqpuIJJT46TESeYKnN32i6+SXt6RY
pim4myFkXORk8zFf5CYG1IdGP14pCbH3DjCiKnTf7nAIxAuEesnLM+5Z6bRueu9h
r/11oYdieI4GZAWqZM2/0eCHl/LJp1Yl6h2zodb4DDACnNjvctaFCmeKZSc8mNsl
8KmQDsdgTa94ZFnZWnXmWEv7qSQdGmtZ70azXKYkCGDFgh5JPT3EmETZRNnhzdiI
h+dqTtPcMshh0IAeuS1cfMR7zwPeNrFEfljM+5w3oOF+yrp7qU9D83vab1fL+cR3
LOepTtSEmb1NOwglo+12+85VIU2fWxcBow4dFoL2RI2HGapp7Y/fl4QXEb1Gejdc
eh9ZZw3GjN/+9/q0Ed9n7cfX9Bm+rB7K8Ka5nLQoBMCrrNxCN/9dDwMijxuLpU9J
xJkBe7ODBriqTchp6qa45aL8ew3eWLf/IKKGVUxIP1AotJWKC6pZ5QxLPUjQ92Ue
854GinAh8d5064oXEKV1O4NEwXcAQaeRmSfVntrUvlUUucH9iSEv2VP6Euj+gMo4
PMLLKrJtsUisU8DN1HJCxwWTxz0BKDpVy0jAqEqagvrmNHJpRO1grCqdHE1jhmRs
YQxG6Uty1DOSlECUFIfqwjmUdsrUAU0F2IwzwfqFOERpPX/Nei0Kz22I2XEwZKB3
3g9+QfSbcTZiIl5zGMyUIuBgnvtwrwb2z3EjTaJK49PpKQXlspGoCiCHw70d+9Wc
hBix6+xskfNHY/FMs05P9xYDJYmlhWpHxKSgOSRouMC28SnefQmTER2y9FFAEPT6
VM+8K0Vch+cPQK8BiW5SCF8WJdaG8NGIfo4Ik5cM2zQGG+FGdEdWplxA5UiNY2uV
j6P+BVhzK6Pf8ZhhfloTpB9gM/IvLU9DXo50d53JXD8D+jGvkUj+ohnOtf+Rn+3R
MvLLyM/my/t8WkuEuXefqMXUUFW9+KJBo5q9ZCA/Lbkmu/EqSE3cE+PbCrGeA2Ep
InzThhSwsgS+23QAbfG2/YWnsfWhia9pB/ikZ3JXweZUuPv2UWdyi/qFZ+Tmwje0
aoNUQx2OEXkP9U9e5A7eM9+7mh38MDCla1VG6Gh89xo=
`protect END_PROTECTED
