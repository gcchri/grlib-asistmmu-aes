`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sOgMRv93XhMHL5QJizpe2QKkix6RTqAHst7LDrzBHxrdmyWUOW8B5o0fEnPbASw8
8vyGOoCh6GNQmNAPfjIQIdy4D/Ovd0KUG34xl0/OlIsB1NCB08/8vmpqjx/FRmb9
frN8t7ZMMuJpl9h/LFy1Yl9dbZcxARG/4bqUL9fKr+b4WwDfH/xyNrZMzJGzADyJ
2Sa7DjtTCzy6uzg/t6ra9yjjwA7eB4bg31v/rfo0h3dfSUXr4pyqzZdV/782twlD
9+NuYIsvqjWkmd1yZVbTiBzbNBvGiO7Jr0acYhkoOJVZ9g03MLnwgyzp3OH1H+e8
BDiFXOoo6sV8dIgQMvuV4HYELHBrLpgof2ICXxDE0p4IJ+whNGCJovUEgM2p3LWz
AKB9SdhRzv6tLX4hm8qFWGy1pCvQa1/NPlomejN9dTVdb9mUWEgwyXuRtKtn2qjU
PjqrodSuKfryczLSIDfTBERHEDkqXtkjA5xgdTEtBqbMmPWaelW5mRvlJdVvGr4e
qU4uaudWVTvSh2MYfS7DcZergHzuVK+iKvg3qqL8FlFO8RphQnSmk0EYpzWRh3xu
CvUxuu2VeT/5DnhC0XYkBORbzaMLco1It+9lsZVECkQ=
`protect END_PROTECTED
