`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zs4RXTT4myOUDU1SHamR8d4wxR9+1dsMBF3mLsFBSqCzk7FI09XM+VwrguD3umWv
cXlMR3F0SoRs5gl28sNPPJ7ZHNwHOzmxOe/q64FW4/trJeVem4B4LD2UA+uhcrTd
ST4i2Tp9pUUbDAdigV/HEIp6IddwFVP0nd9RJOsp+0issuDHQdOFkmLkjsi4uek5
CkO3OQEEKDF0ZGYP4e0hSbkikhHMEROn7X9wtfdq6De0sIBfgJCaiqTEu3H25NTE
xAddgvXcZMUl3N4ZPcnUR0vJp8hBcaLJ0cTlgAbX/srezShcjxdGWhSgsnpPICS4
YGGLbc3IAn6/Z51JTu7gAOz5ug9myOur+4Lkm1NKQwGYL4Xt3SxnrBga1+1hpYw4
/cfMrJdqZA31NE4QVMwPGzmX5vH7/ykinDHfeHGVNqbSqQaqFFeZiEt/UVMHG2WL
+98In2oCjqU5UBiVoh8v7HjYgrAaAWidJOR1TnAUCErv7A3oc+Fu9rRy0mkFsKeb
kv67omYhMm3JOnoo39BgWJzXQMF24kzGAXyudnwxyUaSewDxEAv+oa9ZFYHAd/zh
83mzzCaYbL2TUenBpT2cmnmU+HNOZ2Tq6KNj3SI7Q0B2Uck3hWOdLm5+y2YGF1Oz
3NpaDXgNnwkj9R5l3ed8IXbUPIUIC4bTCJaajBeuoS0JEb/BLDfzE6fo4TaNgAOc
ZmeOpGzddtDwOJyyo3C4ch9iEccXWnG4+JCrRCBbZn37r8wsBpIr7I/dm/xA6qDh
xFYvqK9oIobeU2U0Mgm/D/wB2Rx4G6CULDyPJxk0dOKcObGdo0WA+tIirfg7nxjZ
ndEqlAVod0NgOwskVx+8JCXOxt9rRiNa3EB9tw+HAKNXYAC4HXaEy5jcxRgHPAFb
SnODmYL72KvlZWFyYFvF03psPIX1hg4OjOcHQRrVArpCT+WW4lyTNrbgBt44aNVN
n3RmShruRIzkBn+NIg/yPaDKG25RF47wR0H6E1zzu7HJwmu219XoKNl7nrspkKoC
yCXTbVDpWiZBIwVS1YHFnJDvUkI3r5YviyDqvPaDekk8vrXQxmC8Xgq17n8NHl9x
NW8R8qzKq8r8fSg6sWyVtIGu0yoovvgiEQ/nHWxqb0b9skosHtLlJV7DZ7DfZLaL
rkEcPyMs0EFqo4BkfHHPrmMp/vHc8Yps+xiMzolXo3qv9mc2MN3/At7gYz8U29Sd
LvWtDYvkvfQijgzmeQocgyuCuf6QT73q1pj8AmQwuCzf/QtgdoRfkjStPGPEiFYd
zuYHjap/tGmwHOzCsJVMNRXPXZIjzOdcXmiOpHajRz2EuxMXRP6+MojAH24Xm1d1
l4BvUeu8HX6ftwR4cZOVY6btBAisMaYk3GgfS4IjBXCp2tc+7RpbDEzm6SkLIiBb
7zIv/5u0ed8yKDTfL5YuRvbJk9yOnEI8cudD1D1fupVniy2XWu/bU9VD2V/IlvGL
lVJkabZMXiwNK2KbDR3yGypAaiaSO2lqAgphT/tqXz9zm0zs5A20MRnw2nERZlkT
s5O16t2rz6wupfUCUGRIGOW13BKRK/aJUJb4EjrldxwDW28GIKsdSoZsmds4ZvYs
FiMaa6ax1ZmsU1c9H9Nrg1sPxuRG9GXOZUr0ZC9vePrF2nw5H11Uecsysag0i7WJ
tjsQGWCsOZzDuBTEF1gx84HqptFKFJng5RXOO7UJ8M7JhU7IqHIA2ic9b3Y43cWd
aFsriL7P3tarLN0TkgNayd1oLmVyLFaseYimoIj5ft0QOc/gHvVx6r01ojnUZeZZ
PzreBm3YL9WZuFJyL76ZV2Kt+i9nlIc1J5ZvMx2zNIxwcvrBj3Sob9dsfOO64/NI
ftLI8sEtuteFpZgfcYkHCjeGs5y+RiIJKJ74tMaZ8ts=
`protect END_PROTECTED
