`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GSzJOARfliediHoRYrgm+k+2j/ExfCFO/xG1DtHH90m2VJF2DwRGnGxGtxc2zmCE
kb4+J+GdRqSccIBEeUx3rNT7uwRzwxiCHNzXKwZJzBKegyuv/LZ8FaYqxSgiKEqx
u9RTn6zCmb6vxLem7HzkQqinNNM6cqUBtsaVYMGGoqJFfRbBagTo5OMpn+apkxRp
sTKm0fRGq/CNh/WHPFTAgN6UrfQpInPO2ni16BmTt0WpADd/drCY1lWtEh/aY+Ld
LBCmB7WbngToSYTh/oja7Bt3ifl48qQoQ/8aApjTc/6bp3s6O4ciVvyzCBf23cGo
fwra2VOOaMibL5mBhk1246pEnFVXonE68iS51MLIfD3eJeepW2sYpcW71D/3rvTp
3rU4ReuEJchm1ogNtXl46c1uZ18SX+jWVccB8KSZFfsAUFEbsVq/Wzyj1t8sG756
`protect END_PROTECTED
