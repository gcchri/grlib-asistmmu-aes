`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQFq8Di/05ehchTHbpPxbabex0/S3+jhYpwSA2qWNphrKNjqsJvLCBCFCqWxz6w6
GDM+dyg57GG2UoRLdInyQxJ3L9/ews2d1p1aNCCkoioYWgmPuBNWimoe/oS39ZjE
ghYVvEB4mJdki65IE778re+E1DEn9VrSlMrw2H95sbl+3FRyTR1Dx/gBVtqVNSCq
9fyrB1SsHOQjcDaOoKDiBxd6r8RCU0sOzxllfQbXgt8I7mKrp1s8j1PyXz81FtSg
xK0+7Q01KRuo5e4YzyE/MHQjRCcmUeFMKQrcx/CYkjHyrfrSPuQ0HeGCtPMV0MpP
s9OLWuVqem+q8pQK4+rnlEggZOzYspoAPprcSuCBxI5S/Iqh6BIGZBOAUgA6Hd9s
Zmde2cboFd7JT4av+rFuItm4SfBDNMDBQPWn0X8JkFLHYPF6cznuob/yVxtCs9Aj
0BsajSCuN6tcD6vZE/hSGyRDpmSvVETRcWVCT9V7ZCE2uXqb7YFbWW376fNYUMV9
sR7aQZPLyn+KgthCCrj67QEEKfjsvgLov4M1s45dOnwQdMXpgtnaOthqZsw8aDva
9K5P/FFE3MXn8f4bZ539SVOp5EUo740bYKSwpevX9hy1EgUMFk/XBRUqv42lfBFM
0W4lP+c24Rf7hnR81DmEVue6uDftac8GnEXKK2bmbyId7PV/GcLpPh+En1kyVSdm
+6wmV171So/0ao4TQ1lz5kF/cWvOHBfYTg2grmuiRC6v4iDOZAcgzxElVQHARuJ8
+YHO/4qm58l8t/DUCI2Cgi34YZHsNyfD6mdt12H80iieDhbC2XnBNRsroy5hOUX9
c3R/RnxsTmv7/sgK2yCu0A==
`protect END_PROTECTED
