`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
58A3smLdOxjIrBcd5akuMttWiietf8rIaj0fwo7EY+on0K2rJ/mTad9KE2JWrFA6
VgdDXC+EjVNttljDI4ot+zRqjVIbi6oUA9VPijcNiclPM6fXhAGfvkc95xmq5xQe
OyF1S2o9wVlKoLzCE48CCw7JCM5csqEnG837sp8Umy9Bpx5ZxDZjakZseEfe6zaz
2+raqt4snifm/ePDJEiIhh636Hifa06L264Xp1v6Y+u9ERYGsarXLiuA1FJORwiy
mXQ29udtumaqevo1jEeeS84/waHlcSmnp2O4qvx6+lst3VBC6tVXh1e/peCXtLwc
diDuzoH4APMgcBX1L5YouXONqvJJKYWVzPV9T5xsaJJx6hkBTTZZIDI6BdlTdh0z
`protect END_PROTECTED
