`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WofsMNJfTeFqZbMWqxsDXg4Qx0KtfoLXWqwGl3hTGx3TywPPi+RrLPQ7HDpU3rcT
igJhrQ2Xi48oCixlERw+lZJfHOydllWbdxGinK2hu2IpnAgu++paEm4gzgTnSSCs
8FSZUvc0GN5/n1cqMdxmC3KU1eYlksO0bBjgGkCKkwmz4To62zZGwwEKRBpLpeuy
MW4QJQlQUHqXQU6sfLTn8yHgi49GEPMQizaEspfVk/v0XRmk1kGqGTfE0TaLLh1J
f2UWZ9CEXy44ESjagYT55cLr0VAMv/tiwrAw6/cTpwTuBRmutXZJ//ZnMWH6dQXV
jWD/v5YKbdVI9EzWhMwVMw==
`protect END_PROTECTED
