`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jf7cTorQ+yXhqvQ61lvweJRarU2hVKZI0qcltyGEDePfITinvnBMxxwP5jwKZH1S
/ZyxfJT7ahbmMuOfPVk0/pk7t85l7ZH4dYNTlhyTQSnSDWMk69oYXNg5R5EgQKqY
yUSx0zW17foCW4cXEoguTs52Zmx6pzvjzG1W5nP2oqI/zxpmyCbK3jpUhmFLoeIh
f+L0QUO98Y4ragsUzQbludHHAtNG9lCJ4RdIVwvR9Ov5bwA8muwdS2FZaiWtaaC6
Vo3bQUdP0obRlmGmDx2y2tF7ey4E3sp7qzZntxklcBVGKZYzkLUMmCOGuSGrQxsG
qoIjKETXffeKP72HDU1ysyqyBoQiff8xHCPBHRWesQhogjpeMSQFe0J/7O4QY/Dg
SF9NYPN97p3ZiMyaERJ1dQ==
`protect END_PROTECTED
