`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1wov/KR0FxLiwQ0n83DTePEfUMCc09vJmCIJhO5hl/ya384OEUAotApQAa40SPfu
nO1cvpt7VlkGpDsDfKawWxJAZm02ezfi7Tfj95xd5PE0EnwzdFbSbVDMOBXwNwM3
2H/d4V77sOgW3geNtn4q0bLw7GIsGY0jBaFu+4Wan3XuZjqtQNGPAE/3PPcdl5Je
D2vTECqAkVkiyp9Yjm5gSKlPX+vl0/Ugc8IG6GOzCYt3Bu0UOhPCFtZ0HGkvk657
/ZFFTwKCgafv5xrj9qzYfgYKizVq2gSbnurlg+1YhfiRpiFeGUriSlQBFx2qaVag
2Wgu3XtYLvLJp6Sfc6xWdpKt1ZghPwqloPxJ6qaQyeGdGFx4u3+5FCUH1+B2McCN
Td8JGVwaMsHn3uLvbWZoRoo5BdZNGx8yFwGJT4OcSpY9iwK5Fmn2XNisucoH1FHX
sdcb1eYnLdSJjkUFyyhErJfizeAhiKcxeWYCtlfKnOfMRQeS1ZsDJNWBjGYIaLnN
UpwhIqqDbYIPZPYnlTu46VRD9VRhUU+cerLD54KW130rvE7pk92QoupxgEFXNHOx
ADqb4WYWPDpsDGFxI0DRv+PPJ+Kd5m3rGN9bLlYavFpJ5R9zejFf4qgwQtOAK/5V
lFuhnJixtAuHbtHmBhyiomNsk86FDTQKyVMS57VSzwc=
`protect END_PROTECTED
