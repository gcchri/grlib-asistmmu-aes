`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/OEnKNK6Z/L5U0hYI+MzUvQhqckP7qIUCe57mI75gS7vDic1MUBvpKttl7HUp86s
iRtBRvrIbrjqAEYbNhmoTyRpIYwD57/O80vOAB16mnFRTOk6yj6pebLvSP/1nJg1
bnfteH0bTM81s3ljK3ByTJQuw6Dz1WA5dfCRC8A+c2Snfp/vVodXRVNbX3s7Xtvv
zqpQZ+hpQCRozU3ppXveThli+WGo5VjaG39KU67s1ZI2Gqz1+j3bipYYBteHn3FU
TSY0KSvaPnLfFXprHVAV6JmYsXFIrSwVyAJhArd0LCMD8u5RMvLLH+whx5qZeRlC
ROGevgn46LuTqS/tzPC15ACbekUACH5f1btpoKVMuWlkPTeaeWvrcQ+bBV8FPZPd
inbaoh2UiowG2OJhe2b1XNFQDfDcY2VeqdIEyj4TupO1kr4xzd0GESVR0SpknydY
cUfCosCijinDkKKSDKO5nAKoKeTDjJNdxe4jnYasFsAp6B/oNjOaUGN8WFbmxYSY
3WFPZma5nqtpGsaEg8gpVKJGS48rEx/y1CzRYJ7w0GPbc/0qwzQ+Uv2m4NPfaZiW
/Jpe+ZDKAuCrU4gwHVTxDWJdGPBk9g2n4VNPXhguwFH9VJQw8rVHdExCU4dKuoEZ
uA6MOIKzC0Wj+hYyvXGrgK1TSjvlHP8Mvmdajsbj7u3oBg0kNVsME6GNymyMpkNX
NQPR44xLPUGe2hVtgRBlH8u7Go2kQoknuG+vy/9/LnrfKQZRRjf9QC8VBbM3/fyX
qI/7cSJtdcuSHT+oz49jlLtf3DSJw3H41XzG0Fj5oekxUSHR/SHPRKYTYojZMabc
onbSgJNkADZXU5OvV2z96FWyV4dcsfBujkPTpIMCSLQcje07SYf8eAnFhj4aGYap
oJdJtJb8g/1Jvx1cgqZ8z7vuze/KBxBqIu2Wt4QGJ06NKaI6yAyLTHwlUCt/kEw8
cTkSjwbcI12nPPNfoJAzFV4+t7c/nR4PFwEP0Jccql6H3mz3JUpe/ici/rIn9J6f
SI7ZeylPimzzuiiffafjJFQmNVJPjvAESZfXbuTrCrfpfFYU7bzepCqlgIqmn3kX
9PqrONf8vsdmML2uSiu5GSZaznSq8FEqHJe1O893zTjkkl1ofJbRXFzKYiwPGxU0
pAKHJI2nJoh9uvRMfX3W8qxQXbbCiKBDqFLDHMduG9Hy9AodISEIOQwQ7mENAetc
ro5026tQpCxr1RQPyVaB9w==
`protect END_PROTECTED
