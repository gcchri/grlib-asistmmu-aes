`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ugvlPto8Yf5iXZVv4SPLhmS1bQBgj0g3sWLrYjBJopB6/hIJfYFZ308abSjNri7J
m6Ejn7sGKzCx3xGo+kyZFDjgpGbXRyZDJ3PHfbCSgNmhYP4Hk9C7n+vYSHktXXy6
D5c+ruUn2vPbjMZhfDjyITKe5KdZy1VEpij4TfdQi4SVjHMTMjLU6Nvukaha+GZM
EgiRSu0GzTgyA9k7ilNmAWBtaBrNxDcvrrmHTlWwljv0qEAkniRMZYKu6Z/ySZlR
OFRoRU1+Mw7BUFqRWr0UzLNJ+fFWfDV6hZZmJ4bWYHliuPXtUHV5OA0U2Ffbsgsy
vtTqZUXJV50PBVe9znXMcDKANoCnHcpFeGwEjzOPbfycQzSNqxvpx1OOMkrjm2jj
nAWDs+HQ6NbZfz31a9dUnUNbFvAiLKWjsoo7MNY76zQ=
`protect END_PROTECTED
