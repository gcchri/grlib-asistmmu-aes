`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pxFNNFXteFJdk1u5ZKPJWDDn1iCteRgqIKLbqtx71GlJX1Su3FqRh3qusFDCo7j2
eDOsvZwPqFW9ZYmyAheav8JfDTbvafYLtYvq7rXuEt8Zy4jyDL2mktYwHHi7EGIQ
dFY8ekV31KD/+GNC7sBk8X3/Xqw+jaBt+qAUEIxBrbYZXvvjY6Rbme5t1Lt6WkgD
HrqXv+ZRAUEWB/crCYza4ypMIPe+fYgFIaLjkkIigFYWpltHC1RWh9fQ2BDbzdIA
LWlfyBUzv7MGIdEMqFo2bUVuoXBW9+7Lk1SPMEALojD//xSTKKVKVgManDdemOfo
Vf4V5M82eMMlDCAvwR5dDL/lY3KrBk/KY1Q8IGvFx6UKsLS2nf9fmbvO60M0RYTt
KVTDByNra6Y39HWrZpKlfyyi4nMx7VnthZ9p935NYbQvDkB1q4e8W0RpNx2UTet6
wXgxvB6Tj6a3xKXcCchXb1+pAY0Dy7/uzo7mGbHbnfzAE0DPjnYhEJcE+rHa4O7K
Y5vKcGmM/hEGgp03glctxyLuojcdYajmQHS3kDjsoZxMP4+i+iSn4yY6T3INwJeD
0k9zSvPvq2ARHqOIlMTfDdTtouxlbn80n1RHmo6xo2jD6oz31r+IlIJ7GVTQK0Tu
xJhYOGDaL+BM0FVXSN720QkhUZzvfT/gvqAr0DATbeu/i1sEni7UWNk7wB6sJh3x
DuAmXmblyI2eBO8VzAqwXcI/ogN+1jowygSTohzFPjs0fud4wxMJLVtKtTljifNc
Ia+M0XDzndDvEYnfH/05l3dPl0L2NM6gqwQxjCw++a9GXa9GB+Du256WSOGb+XpL
6paevvKwWxKs9KSrTUjrF4o86Nv893piGp7tAi7ImSNBivmZI2ODDilIZ1ECgsvk
`protect END_PROTECTED
