`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BEP6gFRbmOvyGvUpvRBycOJwI9VpPZFZVBqvHtZySzTN4+ThS6DMPAqSS49ckMGL
iee9IFb1ymhhAga0b/e2WH5oKw74BjbHjwzui7DCN8Sj6rOAFpQNCki25L6Xkkb3
YkcF/k9Hx9HZmr87G3vYIg9hrv5HPyua0HntgGEbAq8K7wvi8v3kTJHlIOm+OibI
u57+kzTRdTmmRflMR4x4a8kfDDFS6xzSTeUKbQlh1dqdAYBZn52IK0ELCrY5/SY1
fUACJt0ePZkAv4xd0V6d4SW9RyjHkCczwp7+AvZtI2+iVjnx8MX/DXCWLZE74Bei
5w9EFDeGRSpKmqMlTl48RNwpn/ctIVtl13QxESWCiHLJN4ZGrZcMu90bjtswWa5h
yNp8kosRON8Aw9KPvKUQkcn528qB6hy4TxskWXNHIZc0ahsgrt2KNiWYEICqjgtj
T2n56Amch3K3qsEOUQQjLm251q6sKk77MoRTFITTX+m0btGRa2i4R8TIyStJUXlH
kli4rVGyVqF/c8Nl9PsN/d9LTYjxgCF1o8nO4031lx1+CaqTUtgBZUYp2+ky4Yin
aKDC0ye2L+G4UNWNxVeuHlMExGWdVmm39MutegGFLspsGPOzABgJEGFMrRsciZ+r
losdcyrWWzeBSsE6kB6Yi4nRfRlQdbTzqjug4SMxNjNY69bxmqy3evtom+XrC/0+
tBXA5T36GsLL4Nh02jTkmA==
`protect END_PROTECTED
