`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Li3MavphiA4Xvheh6Ro1FWv9aVtPtei2BCS0SltkyK3tBXzmgcz8RSS19X9WWv7f
d6zZsCkmAxebOaBPNBDIMxvbU2fGeKPhAHGSZV8Io1qvu/xCc0IPIKdtJEtRbV5q
j3kH5yKAygQ9tAyHSxqhUkXyK+ZhCG8TbLHeIetKfiYf/MlRcq6IqKowxo22Whf+
uhclhjbi5yBN3rLDv2mTt7kIn4hw4rohXqXsbNppzTQPb9l0b4hqnJQluBFpu4be
wSftgV1d1W9mPtwVGY3KnhXtRdPiFYjMaRuyaJivLxe85wTakPB0UShODHaaN2kI
MOecwaVq8oJGJ1sBDKfcu4L/80LBjB9eiR65Z2g1CdeVEbJhY0B0G+6jQPlN9rPT
7K666CTovz4RrbmK+wH2Dq6/Jtj5KlwE8UqCpwdBtSYXwM6329ewaUKkTOPvEZzS
j+AiEPRpD1Lxe3v3+ktbWryTjnY8yHUScMrFpaoOU6/d2ZMTH/alpTwjN3/zyduH
bO3l/boOYbhlxSVDKfSVcoLqq+e5Gn8hb5AQjiKKRF7zbj9YVHZNVqmPPP2sEUBV
cGnnzffKgFNBc/tH/tyLD6O2C/ovY0qQ9nb7eQMOF3ounoR9TzkCWx82GatUUJyP
0lIQtrwTA43GvHWfa/ZHcl3qVb4qvrXVjnq0z64Gxh0=
`protect END_PROTECTED
