`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VDt5LpnsvhOCtLCkOVliR7nlRoSUUuTXL7P6DP/v2011wPUyxiE5Z2plqiniHr1w
jFpYFWIyjdaj97/+Seti2gJtqi/TwdBjsfdvN7nS/g0cxpo4ibK0gW7y26OcF03L
baU2p8t/m3exStJ8fIesrJ3yzFCkkzZzOLWcNQzOjwqtyt0+sBrPpSmk0n7h2boB
8LNwn0ZknFAA6XuOOAa6tieVnN5U7zxpIQZVRNK+mI/22831YW5QAS5SlWJt2kvK
UykV2gpoAmyAYNGaf/z55yZAV8WJdvu9whhYhlqzkvosZ81FFozd0N0Ne6fkcsJo
igiDnKJ49277Z0t6t5xl26GXHGdjrsrJfGLfqTN0KNvfHDn4XF/cBt21qs+0n0or
2DdZt0WoLboDEMh2RFOsqRhUL3O6drBuqDpKTW5UbfEnqhZYfqFDgHHMfPbqE9XL
rOQTh33vKRsVJLi/GdhaTw==
`protect END_PROTECTED
