`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9/dClh7d7oTC/nGgD/KLRAfv4xoUvPO8AJL8wMCnKRlK/tjIgBwJUcR9wJb/CYZy
dHZZwYAaFYLJlVDaenFBbusge9RK1JDcLnzScd+08pGmfJ2/QvUzdQJiG9Ko/maI
ZDxlGdhGqVqvaWw2Fw+UtJ4fhgZAxi9mkP/7qzWHjcz4NnI7ABzZYes0KIxYkkAD
QZZbw/DYu95+pg/j5Dwo1IFbfNFCgjQrkhuix7zFnymrIC5afkGsh6UbwsZ+C6pa
SOpdLe+vHKt6UX09EKbw1m13NPFhhTnPtLgDhiSrYua8xqPInpiHziDgRDZ8Gpmi
i+68BsGgzO+4U56c4Ff8hzLc2anDZo+pK6wiSprWzcoYhSHkCP/TbSKuGYTdQNYy
JiW4cDl7ququAXSnErv6Pc0Odm3aHPJB/eEATP6hDDpogLBSuwcM2ZxHkyJZvyoC
5qlh5TlRV7lsr31ilitibIetMm023H0V54n6iFf51lmlx6qvYJYUhytxx6SJas+V
KQZ/HNRELeYXTgYec/8nCkk/L+FlDGuohInaqLPLJv0565bcH+Hg4aAAxbaqMyiR
t0PWbZJdUu4e6H3iVCXONdYO0e/awsaIqFkINsYrjdYyBcvIpqWJdeApz/19BSEy
IjP+wnPWSLT9arWpSBWZI9nAS4wpJ/4MsajWgXT/e0UjCsvg8bkUl3iVM2mtSF6M
1y5UpNhPj3BqIEblPJNS57MXjpLtalznO8M4OqgwCjTc6IBH6QcVk/V77yLRp5ll
3TQQZC+4bImHfyPwgKCgZ+zrOFI4osxMrYTzrswtAOEkqfetMklYPOOzjHjDkYRX
/8+EbMkat4NpkoHwxGDXNWI34QIR1/HTDFM85HsiHYSrp/9PdjownAdpUFkoyEdH
`protect END_PROTECTED
