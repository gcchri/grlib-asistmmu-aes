`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hwlAntD3JqKGhpXdbLciIGm2hVlYpmZkj+lkYA50I1nC4b4dI60duUUKjNYiXBax
M3JzG1bYUJWHZ0FjZIa4q01UHv60Nh+te5JdosaXHdIu14fAlgprCetQmBglIzsJ
fCouChhcaQyjl/Xif1A6cgjoklPqJnzK3N6KGMr937DpMZJF8wc4B29urL6yoUC0
xK8acQUbMr4UtQPzNeBSacCrSZdYQwcAF+RNn7i0xAoUfzJR+zOF05DQGusdBea5
W5eKCAyjakiTbDQ1Jp47U2eMUJl6xy1XoFR9DvyKe6Q9pAvuTn7D75E0tcfqxAN6
1549cZhXPfJMKSSk7DgcK+buYXtev4FmYjwmdNnu7H/POAyEAH29HMA8kI5Y7GGm
2GLNJ6+eL2TtxGUEfO8EXkmdVg32/lWaeA705gGA9+9pgO7LzqWABZqzk2byAY/x
KYtz/l8+5XCYQczwc+DeGSQ2mnkWU4p77U8VQDZNUYUoySkuO3NGinUyeXMYIbzZ
7zYsya8z+MKhBJyuAqsIa94h2jPZyPTmo+WWBSyCpiwAf9hr1q1ShEcMZeSWhnp/
4f7RYh/as73AQ1T8PZvxfmahCXDr9Vph/fB0Zt4xdwoV/qTuvlqEdpmsUQUYhcRp
2g7990nC22jzFnDlcomIKsP8C7h7/LNEKdYKwmtckT4=
`protect END_PROTECTED
