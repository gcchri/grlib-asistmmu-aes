`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bpkZalpLA+RgfZHr44dtOoy4t6Bml5cGMDkAOuYpyhBURno8xy2Xags1Q9WKTTxY
9eM24n09yYdO+L1swzSsOZwRpUE3B9gHJGGIJ2cm8D1/OYFPMzynXv8vnGUGRtA5
7I7lWDS/KE7BY3IN391JAAA0uz4yYBFCexxmOH1TOChYf3lkn/6OtMaQx11DFi8V
U8FmPD0PwZEx57JEqTzFpEdE+UMlEzfvb/mD9UpZoCw/qC1jQJdSA3FSEcZtzwdt
c++TA9Ofvkiz/xB4TpeMiPS/yei4wr6ailIee5mZNMjFdajF2SK/T2Z1N/dYuTb1
yuqyca+O/aI1q9J3ddBXLTTszJo6itZKoWLglY0ES41rbFYkUdHVp1MdMvBc0KHC
AShUI2nf9f1Ri3uK/8UWHz5EzxZpZycB1Bk5hhJ7r7KQ4ZfXrU+NfxKzvQxmwWwx
vur6gzgQsrDjOeBlOr/2jy/Vcs27TN9Yvv8xF7rkF3ZkfuOqLsKzVUc09b3fFAlL
0Te2iJGuW4T+RJHGytI93xyo33MrK8/33pm7Wi31y/LktdRuZXXkT+Ut9Ix4z52d
sZFQLTW5hQjbPbgmmgYmA/64dAh4yNIV++4Vt1qVqLLlAmr+jMZ8ZqWEreL7FNau
/lGYuYA9rVcTXKBaPzx5pzDXq4K6PhUouGk3mXl/5QSjDPX5lXWRDN1eTBe/TEJi
rKQQlRu1vJq3dbulF6piCDye//UWWpYe4/vF5HPrY0BqJsXqoFnKkgGHbgryqy1S
csRGeI4ukq8bkXdhKYYN5KaU/Vrhj/bZraqc0XhUCzuNfMMj7DmX3nz7oEJhHAga
fkHvGhQCz4ARMGClTUZGX4zFCTm+iD5SnkG2VqiaseVBOQvldyYP+myYr3LnK9XK
tjin4gKTZo6tQ+CvGDNc6ulh5NDqI/nMnD3XDUOky2wB9JOVUZGQO163vO9THZWu
Eq4GEOdgu6w0j5se+cXxzjz1WGbwEDPkYV8cTyO/syIosFhI/S028UVnFnh7P/9T
9g6/ZFkQj7oWe6YeEAfSb4CnZ++VD+AloeyMrqQ/S/Oj/K2ta8T9t5OME7+5x37Q
idgtQWAkd43UNasyjhgRlg==
`protect END_PROTECTED
