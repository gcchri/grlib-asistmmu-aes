`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LhfEUCeWBVkTXJtzzza9uQC8g9AZNfkhqczWtR0yyxyekUIzH4K9dmWssTMkvlLm
6QRHFFzwalta+TbngSEdWYfecABT7NHLEhfu1qAfMugtexsAqqLsuLIRZfoXAh2B
NIILpVTrm9A2Na0o4IfYafxPzjhz85sDWFsS7a6PLHmubyAGaUF/Jd18F9YmzYZv
r50Rh8mo4GrlmQ/CF6ywPvyiGyAvpsP/N5xEuPJ+4BvATeuiNpGbToJsxbJNzAYU
eoUJx9BsOTvYgVawCTWlYJf7WIZCXUSUPgrESOGVQmBqIWlEdaJNp+7G8038qFWx
h0Et5ZxmcSHQL0eSZpZ8jlVCX6B5s4tXMfrJRIwQkALQBnBALWatUX3nuniYNIR6
1Vhjg/PNdfCVv97FdMPbiIj2Xfqhv2UfAwGi0SGGN57TWua1nJBAD0b/7MjDqbPM
ofD2bkV4HTxkDxNlaSIUDH6oPPjtSRJVrISIo7jSlrxboWJEEwk4wpYBWyXGlhG+
ePy4AXlx0zvfU/+VTM03Dt0jHlmuUW7w48i0NP8XyZ9Nu9LRy1IckmLk9SnTWRRK
8Hh5xMSiJ8mtnlWeWZSbuunZ30JO+NO9SBoUTBUE39QhD2SL6PPkdYY+tmSraofH
xL+aafwe4o7DAjMDa4Yfiw==
`protect END_PROTECTED
