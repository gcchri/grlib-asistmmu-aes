`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gupkvy/90fuLaKH/IXuQA77Er2dEz21qYfIrQzOilWmPDD7plgFxKs0STL7GZs8d
jFvmgMJQzia5Yzx+F9zgDclpGkkTlYJlXfMIXl2gPGTazFgmWqyqZWMNoiqtkIoq
/oNW111Ih1ZUzCcXIs9dOi+PB9ClxWddHGKPPzSjjSWtuzdr0LzhjECK8QrH1UxM
dN4E3Ao1HOqHZyV2akz1DS90a6mY9XNhdBOx9JbmbsooJ3dgCzImUjcWROpCvRxB
F4PPxWCmgHGtb9w9NKEzrhDvY86D37JboPCczr9l3/cX+xhxKXMNSU9pauuvCJqo
dnB/2PLCgHegs4Upv3/5aTElJmyoZrqC8nTRLJfTpGbZUQy0hP+6fUKVSGorUQnV
FDxv5GfCFSV3pLLpuqAtVYEj5icoG+fbokAt4CUcgaHi9I2Snog7C5emjFnUQ+9Y
qSTN3J/wQ/+MQdJKk4/RYOn7D6WStRJi5rIYsZkLMwDV1rhSHMFALCK7L12Fhybz
UZKkTgYsAo/OB14sh1/Aosmqyf5wSCo40BDMN6TEgHEnR/W059M/Scv5mGwr59u/
alFQi//r3+3aFns3pbGj5ffDZ1coyZAOiWXSskIb0x93QzQH1x+nZNXUdOAz2zmX
Q4wBdYcgUHyvjW0Kt11Q3g==
`protect END_PROTECTED
