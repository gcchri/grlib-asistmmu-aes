`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B4fm+6dpHe1akSVFGrd9RfmcSsPX/VWjWparqoS3zxF4Boo5qoWMC9PluDmsruhl
ck9+XcEjLLw04UJ/rlJuB+zV7xtnLMxMsTSdMbIKq1PhJur33QAznbi5LDWEfOXJ
2jfyj8m+C29LlWL4+LzSytQsMmOG0UZ8MiXDUSMnol/ez0N9tXYJzNumzVxMnV9c
ed0t1W/Bk8re1XfJDq4tg7n17XFVx2S5JCxPGoh2uKUbu4kyCEMPmgW+2q0PHOLP
XbRUiZ0kKX3nCqcKr1fj1lVLnAAx8k7PQvFmJz2u3SukAVaG6oHJ13UaV9yhkkCI
3NOBd4r4fce3pbmze5pWpqo8Iomg3GHPKgLzT2RV/Uu8BqtD1oYrplpAsbswgCMG
ebEbrel85NkEcJxEl3gCPrN741Uv4ejUvrAuTUJHz/AisES4Wpy89RMRSXPaa7Dx
khMdvR7Mr/5WLYsqF5nZsLRcFqSmr3MzPJxLHJ3q/bI=
`protect END_PROTECTED
