`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
17hMZ2dR1FYqH0K25DbJyhvRoiQ1gRjLyPcH8ci7OEXV8R3thpaQeQbUVnoyXQ+H
nH8IVf7V9sEQ/KAeXtzbqJ1iplrPPkznK9tiYeEVsfwUCkvzLg3Brirx5MTjytHh
pkW5DYm9cqxBym2G++rSUw1+SYzQqKLlJ6uM9Jz9SjKPVGgum5NoqqnHK6pwGOIx
ayg0qnlDl3x7T2Rtov8LBnztZ5bR4NhjonwuwQFuokVZjX1qKUegHGmKNd3skyjQ
jMCfgtOvvn44LMJcqcjrAkla6aCo9JIoHwj2XGiD6KIs7Q7wxHP7vQ//Rblm/FVO
zzs2yIFqVpeULq97FxiAFFdmQaLIGqKK/RMRClB1VnBPUpewPzDAeyqbBs/4SaR8
Xvu6CatEg5JE0dS87R9lSZrzcpDnsdXjmlol2NlNzCHv+M9zkrQ7SyQD4TBS1ZTy
h9cbYAGOm2K/AZVK/qZ7qGjDcEF7avR/NcRK+fQGmPuFj/OYiNrGN84r6tjWbOnZ
POA3EgKWiHx+zzzzA5vxdVFHWrJS30+KWKajEXPfGPUKLpgWVIJo3+S6U2ZQXQOt
U92+GGusC/9smIAcBLsfoL7Yu03CAsKpSnlv5B8tRhYFlwCRyKckkE2QpAyJdqKZ
cWG4xJWrSi/wLyWz6ZidSJ9QgYbrLTvBk9ezc1qLYtscxb336YZKdbI4uIKPx3nG
RxkqCx8VxXQSjq7wi5GCP4kdleEpGuJHZtfB1qn5G5r30+IZxWuCWN/jfQJQPO6I
FB9pe0pRdE3LnHZrLpqK/RbIX5iIkSwisWGNBGiqZ1yAFXDRTqvoQW9APBT0rEB4
j+FIox+1j08OIGd899YTZSe1Jw8GlWftKAOmKdju4EC7uBtbQzgpWiqY6tJOkTJa
H5KyEH4uxltt23H8nsnWQSkONYFHE0KIEwzjeD9YfTtYj6hpk80PlbYPxEh2MS4e
mPtJrsMTZExfe7a1QAaYgr1hN1oO0Fbmt+ibdwIXsefZXwWY7wIluPaZGc74NB5A
rDaxck+1qiwZUSNKlBxCPsXDt3cHZvYe/fIbd8vCudaUgSKKTDcTh4A71QNEF4cD
pHJwiAYNa6ncrESea+4c7RqkWulVVzl4c66GAqKbc1B+EScEvLNpG/lObA/63yNb
aBdkiNnm7V+Xi2ccc6BtnWMJmM8FrDc1zp1mDiiUEp1oubKaM7juPU0LMV9sNs5z
2NRR4zrD0wJZHT3jAaaHQMGsDpzZjqNPEvK42Jb5zF/gcilorj36Eulys/JEtCJF
pOjvLfxeX+HG8TGShWjtV5TUGGcoMjViO9zHOGYj1q0Y6dvk7AN/cwC8H7EWCcGP
oOYm8aTMAhrqFpLiJESkaZ6r0ofSuq6GlUalsOYqaaB8ag38Nih8zjQPX3BoN5JT
IPfLAlk8J0aQqpYdiTU/o8TFY+XN+IUG5yOOinLJg9lesl6NLpH6vxOpjddf/+sp
oE1vbHMOa+ltv7zrg0Zhy9jOru8UMGN8FMj3/FDt3fXaBFASGtfLkEyBbhSW6Sau
V5vnGf9eFXmfIT7OjFAsdp/rXAHRhL0oc6UdCFgyqGxqgWumvqem23vyev+i6c88
9IzLNsHyEkD8zxUL2f2kh5Yfbp7bZNZ2wdunViAXvCiodkJMfvE0+wDkF2ayfOWA
+W59bgx3Eek6R/PKzNpOU/jB+DTg0z5czq5Aj/0XlenUr0g2RWMcIwHWsqejNJ5V
NLSnj1aPhXToaW16REf14c9GBNZUjbYjoSklzzr5NMPYlsL4dBdeJiJsoyAaNVKG
r9kpacCdF00gvbQ/jAlhA0FSNYwCmGdX0O7utuSgEW+DRFkZKhW5ywAGMeI91y4T
ucWypv8m/ylVS6NtO4Xr+92lhwqJ9yVynu3qMQvZl84=
`protect END_PROTECTED
