`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3IpkbrCIgF5shJwV7RSPApA4tp/W6hosJUHRaf+ObIm6MvHxcysZMfV396T0HjM2
Yt5FGQgiZPZxMLi7YC5bK21gw34AgTb3+ZHbnBayyZIAHcFMKa28W3gPzej+pzP7
CFqjXu0b0hzZnPXHSMpGOV+EyFbimRVfJw/IaVjWHMEa9NBHl4IMCoIWhUCZJ7DR
xM+4Y0G6leZphEGsAHKrtyh9cdLrS+T3t3SCuypmA2LnQCHf3TDuPIFi6NrsCJrt
vU1Au3/8PviELNA19L6xMHP7Hj6L76uv//ve9k4TU3N6YRv/Q27yn9mXOmjIeVyk
qmTQ+CKp4+JJKou2RK2FH/lMsJObxaiZ0tkgx6LHp7zCP6Goz9hHgw2r46VkPMIy
NBoKYeRgxZRPJYkNEGwem0G8yizZ3r7buTtOavJwke9ravOt4uBD5CR+FGMyHg1Q
FSjFgKtgGdzXq5iLMpsuhly7XUaMpccQRtc/GVmL1e1+nTrhrGgxL0jCUkuRWfZP
6N0pluZ+CaErMkhS2rwNyaKDP6FpTKbtJlw3C9wTNyBYlt2mMZax+aziQUk43g5q
/mBa/1M0vlvP+OpOtUJvDd+WgBdl7un0hj9MPh6u/uD3SMbLLFkdPl2LWgayIqM+
V5/gKYyxEtvJyJThAIB1bcdmE9s1odxv54fMu8ccPsMH75iPKK5Zc4vumtv0mu4Q
X6roQ5pUT+DJDzFKCw9KlV5I+pIEutgsQkiMsHsL7fM=
`protect END_PROTECTED
