`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y1WQNHAVcLgqkrxCG1SiZbkSM6t2gIwoaiLAbPyj1VJXX6cugezMb3GVPjs9TrF1
O6rWCcA/62bPXVmibvwMqdW5JmpHCOI9g6cZbnYKKpA+cKL7/u6uCxFekQsYsyoP
bmcvPHDAl2a+p5mxg5PiQzTnlq5cgeaQsk6qL5b5yrTOeiUdrRTdkyPYB4BnQMYk
HK6t7RQdd5wOXU831epqIkNUIM1uQd35u3xT415ka7jYQ50Fsovs5TuV9ANd4lv7
3HPYr3AgQYL1ZdiWRm9QErVNVKJcoSPsc/yE0JJnNQb02Mk27pTZqb7E2tvnG2Ir
+0YyR9gOfNicPfqif5mlIj/RnzMcytrlP8RKisZhRaT9KW3PT0qgyWRLGgYOq0rD
gQzwgpgiy/u6FaSJ++t6TQ==
`protect END_PROTECTED
