`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tQt8w8zxZltZJwPk/MhFlhWV2BW0FBH2WXwtO7b39GJGXYeMR3erHwRvKFkBBarS
UcIcF4jv2F5J6lsgAZ/Pm1ddJs9p/PBDE4kcl0EFV5Dbbtrr+rXNxnD0owVzMAv1
/pHKvi+a9sIksDllHU/DNYjcp+X/mQl8YwpJs00xUr2wQq6/N3n3i8/cARIEVOQW
3UaMfixW8rmrcMUUnzxR9XrdyPe7Gma0SDAPt7WmiOs8nLcmIPlgrqR1ljVYjyjN
p237Pl/dg1APEk9epRq3rEW+zS8i283fzAp13BWO+rR+SjfX8K+6knGowDO7kVGH
xZ4iFV7vzyzmhnp771MvSpnIRAofDm66m4VI7MLcLzUP5QplV+miLDHmjQ7wRP2q
`protect END_PROTECTED
