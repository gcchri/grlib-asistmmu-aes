`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bMm20ybTVaHlprAKdYQr7KXd0iBXudWUCqLRb9AcY2Cgf9HzL3q8tBB0iTheElAZ
QjBrCvvtGhPOohJfom7wHODIdjA6MK6izTdKkFH1R5tx4QRfXtB5uD8q/SK2Bgbu
wtnRaiOZn1bIqave5PuQAvTkHV+o192Gj7nnDZbJEAjYRQs3sIZSBQjWOr91Scck
Y9x7Tq0KOFG4d4OEeAFwFX2v+4JaL95aOf+wgzgHs/kYbn0yBxU1Z2yqnVwMO+rj
sVVjk3EyKs2NKgpdoMzNArkYGgYibdPA2uPk2louueJti3nkOXXFy6ikWuGKkE2q
0DXPFwLgfxEEgZjUDZPstZA1+HShoszRHr7/gGjFQUnknDrxZr6jxiFIbPK/s8YE
qDcbTK3TnaJ3DKEmT3Okcw==
`protect END_PROTECTED
