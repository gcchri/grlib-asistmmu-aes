`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jhvMu5vDxzv3vdeMXUuL5bOdAWep6XRxNLS1pmtwDR0G2nuEfuOAYW2BBV0gxyMa
bGkjg+I7uPIoDchSbeGiAth08zQSiYpJygIt5XrRmDHPsMJq+7hlJeG056F6BNIK
mpXViNnXZPwl7841tQpxWBUYDU9tq7XK9Z5sZndHn0I+9JH/CuxfyuJ22qUOSIkx
bGWH7XH49JSki+5xK5Sc8Hjo1iAoIE/vRKtNatNaJhUVYaKXfoSLvKKGL5ZAoeKx
S1NLb2txh0iu3qP6NaO7znA9iPmq9j9Rx0X4gnAIscVdwFPD+QFUG2mt6XRChUSZ
YvfS+u8C1C4cA/cxJcNlXjevaP/56Cy/AnrWTAJ5QUl5ulKmLfey1ym6fGh/b1/a
K3Z20AkkmIziw8ksGI1CGFP/B2Wj5vFF+JZKH7JAoSuFeYFL0sWMYuviWC1NcJy5
aHheRSD6efEQLwmNTOOeJOmY4FpUf0s+s8KHFagoUl74DgnC3JXhKXWqSixQqR20
3q83C/BSUBUGYG14aMoeHqoZdY0m767P8tof6pgbTBI2JMftJD5P+vgiEHUWIyU1
xZJf8jLhopR0Fgbm49Z7h5SXREKaoZ13Xm6YlQyefAIhjhYgZmRPo3wiFcpLno3E
u4Frb8eGQhQEnlL5bgl//MQAXD4hLeYPZWGJGxmPi81+f7XBc6bH8sCn1aaoe/aO
C9+/FtF9UtsV2iur19QXwTgvhckXEQ+WXcsGaOuvjuqjXmQ4X9qSXXUHIKJMR1D1
4m5DusQ/7Ux8qZ347YyoJCJyG2peYdCLrQYnDnvvxqrZqlVwt82JFLAQIBJcyCDi
d4qNLPd0ITK64PfmnVvhSA==
`protect END_PROTECTED
