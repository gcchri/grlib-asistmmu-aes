`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QVeJc6uA4P0Z9KJLIAUZC0/aG2l0hJJddBeT70tkCFxE9DtkdbGayoTF8g4vZOWS
Yp15MuB/6dapeFGx19FyBIBzKfVZwkd2NebgR1Nur8uMt8E9ij07jlBb0KZlMwMQ
JVmJIox2zq3LCCY6CNsSXhwmx8viTbNIeA5Uh4FrOnhyJsGVX2exThK3ybuKffxH
/MiomwbTbU4KDOikmI6N18HM4dvJtv4n2B+hocHEa7F4NHcFbqXSSRuPF6owUyFo
KSUqgu6cdZysDxzmZ6mga9nqpr6YWD0o1SsnQL7a0gRoRWalVpp2tO8czLtbX/Hz
8zb1lnUT2I87h4V80c+FE0AI2X9ROAzQpo+v2r4K9V/4ik3GKT7/dmZK5EbKBaoz
COXHRbylGHF+tiAzn3F7O0tmhrDRnQoF7zvB6pA7lk+0KKbbIG/Qca+KZsQAOTH5
VfdiGRoyvek6UgdMTmOnIVFfv4PFnBeySGe0TvT5tnk1bLRtG3y1rbUd7jcPAsu0
2qmRswrbiePHpTvir+fiqgOL5k0I02slxb1rOHaCOJEw/eSqAY4NyuVLXk1fzxfg
rik+Rn4BjJKAYnX/4Axq3fJkNhSW+TKzcbvJUcelEM0weiWlRGjk4mxA0U30oBgm
B/Mh42ANdwodVPG2NWWHFQX7m6iKNCIPMukhQTGcfciS7hq7r2huIo+5mnd+5eTX
CksB9ADBrAM+L1VSn9Rp2DGIwZmaixukYobbwoSQQ+41TtwBnP43IKZ8IxTat//s
LuiUB7vIKuI8ep/BQCEgb+OVAKvxvlUz9uDFlt6blyOSiYedEo/isCKQPStuqVVR
YIB2VFrA+44DMDjUfUyJRBH5iQGc93LE3EQqscbUCTcHYPAmRIuyhn8JsNjnCOo7
cjTWsIXc3moHDNjQTqhobeWCwUdf5o9RIIhhrwRQIjh8rP8eO5wWJrlosTRZlP4B
Rp2vUd2ZKxX2xr7j2Dw/GTtpR0Q79zwKWqbD8R5tgfjzj0xrNAM8vSeyxb8Ci0Xb
molN/FckaBMV89vfOn6rDXvDRFclmAFlyHPwJpAUabEDpwPVVooqoYTn3X39f8Ev
FvwxN6g4HtEl7b8B0IC3gB77gI6oynm9HpkX5gjix1L1tufwN84YbuR/h12VPKYZ
iUNNZDTzcY+yVKur8DpLI6M41PtvDIQhicT+glkf00H2VbnnBTqmmycX+Exco30F
J38reH5egfLfG/c10awUes4O7PT+lZF8clvbse3CGqBoM5RdzG0xR4RljhE9Jabi
a8t9TXBbJaezOAY/QRl1U/BFhLSEWglaEuw+M6MBCM/Uu8sctl+QCClF7rewfc+F
O40q1CucUVCUQzrlB/Rn+9ejGuqxGFz/jwLuN7fycB8dhokwSMgM+3lgS8ZcFrNQ
mxMkNMcPDVcTrsJNMfgmBcF2+cK0fqUXlRavApLbOMWnBvGlgSJhhKYTQ2G1BhHd
txjG4/0gHkCsO010xV3sb0x8g4cLQHJF5/Z1+LdlEUMJqzrxbi0zJXx9wUXfMu5H
i1AH6qfjQ5wAhuPk4DybOVaAYOk1kJ79mL42hsvnKi8yZ82xPlo+jtPMKo0ePxE0
s22+auJLFz5RcI4chH8ni3LIrmI17Mk5wRaSz92ZzEj9LpQn+KY5N7ZmkACk4HLw
X3nW/zGDdRJWSbaPH/sSeC3dh43tZx8VhlZo5zYX3ophB6rL3zi4/J6jtaO4YF4b
gCrZVDLlbdl4y+L3SCcWtaAnmTiIu6mZWgeQFBbDzh1/35Bk5JNNom05KMlGeBVJ
i3zsHVTmf5ZXRF4tqvoUtv0mrtutNkdt3oobwo2GxVdSfTbikHER3DGpSzznloCz
RtqsSYCOKbYrQ2+bYyUxyOqOlH3sRtVnhSeV6WH8DbVI9Z3XlNDWx3DQVmrVov2x
OO09y0wRHlpAgZSSZ2Lur1poCxcSrbJNmAYxXdRCJJmj2D0+s1HoJiKxL08cHEp/
QDCRsClL3KUg0gwBXgjK0FUIF9AgFF/z5StIlmSVT9wySCl75k/pDgcjfLw97db3
d/v2EwIHZlrF9eeC5CEhRhExXpgLEigB9Ebbwi7WauX9jlPcGKOgBjePavafSxqS
oyzU2USSf2yVjhk/K5y8DlUwBbqIgmCFbyQGJWI5Z9q3qE1H0Sftkle137k/bkLY
ci3cGdSdaxxgTUSdOTVZgOboZ0n1iwt/ukyr3QViX9i9keKLT1bmgLrxEiCdW4Ra
N+NSzbnrVGoUGaXBR1JxOcqaIFLgVHzRA9B4UfPQex6M6LPao9NMv/iNwdc9mdSY
yZ6caHlROWcAUWFm6szh+ph7SxDQ2cBz2FPdgpP69X50YuqyNkHOGODkkN9IRRW4
`protect END_PROTECTED
