`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Aizc+SwEIMQ4PXJttBNYxI2bTdEG2bm6i4UGoCUbSTUHlN53ldm6uzAh5bEIcsH0
AEW3xUEz2cdArh7GUARPRL1ecP6kt/EhHAOqZakZeT1z+d7nvFBopMJ/90rAWPLt
FjB8K/knIiFz4yzuZRMVt+yhsGa4ObF9INQTFswNxHxJmYIX74i2CuIs8jdm8XyS
kkmvMkGhj58ujEip/JrUD5kBK/9aGnKsmAxlLmSqZ/H5FGCbGafzTnG6KpWp1m+0
kzvUFSbmsyR94Ebo+3GFhISp5BNa/Yap2w7Am2FrRWELYwbDrLU2H0MiL6Bh+ZV4
TFkCMO0hDCpTlTCtiAH46Twt/kGyOAvSemjcULvBOfRdJDawuTPC0+Sdo3VDw4UZ
5QshL5JkTl7CK+aWYnE6vaxCCKoZzgXz48TG3SxcBaJMUblORLWgoyHxFURAZHe9
CCF2G//kTMV8oM64HsV/+wafIc1P8fs3euTOXB1h8sCxgTjGLVp+lPSAELog6oD9
/5gngVOuoynT/mlJd/LD1CLdho964e/b/1faMV+TdQN0dZBu8hmvGX2z4OBCVKlj
4GveC14wCuRklu1LwbPVyUuCNuGC95u/5kvPKu/2GAI8kwE/LQL/IRS61j6frw/U
MC+DoIKAIgGljIuzZPhxIy0G74uTugfsJfd9gNAx7/2NCYQF6asySp6BOkAq5vjw
M7uCLnQ6ja4xrxNl9V28a1AnNBw6RHJt5a8Aa4hQK155bkqUPtoHssDvZKXEywae
EZLU97tMLdUqDKk3Hrikj66nZGrV6GDHN8ZHyoXxrFZp6L3w+oAif1j4KPNA1N0X
+NU0/YfQ6kd3uGotHkqFbI1qWVi6ciXWl5ycN9/DP6gNFfN5NNSNpVRAWbeONiy+
rONY9HJBt0f48x9hrjggt/6TlepF/K24znbTTZugIxqkDzgBAyV3jZp5fIArr0vG
aBtBtQ4Mq07iPEhGCSVtJA==
`protect END_PROTECTED
