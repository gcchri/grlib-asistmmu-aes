`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rgzXsKAFFF8AE1au+ksKjx0me3wGGAd6hitXvk1xpcZlWQHGcEfXzriE+WelKNNe
74OSUKmwzNvG7NSMSH9JCgWcPL7Vt55If4oEEZnqxM4ymFQjKLQjteG1QYG9vrgI
IvdJBemn0xsvCnJovE4GFC/Xmc4IWvCqSOGU7VEMhgzYpsMBRIJK9Cg87mD6KB2X
ES4/NIMVaF3l4MaKHoWUHofXuBIBScsv+3oDzgvXdnEgO6g882Ys063f/JM70TgL
jzrpBsM+JkXmE/jZhTnytF7O8i9F9hFA7whyWQyHVSy8lUaMM3s2mIFkILXsS8Th
e0KPfJf/lw8JiB458hVtDvYOg7KZIxUQVxsAEEWoaTY04ykLK8ikpmLEllL+yjbk
+vt+OJNlUnwsRO+9lHPqrG2/8tm0IWej9tDtRHdGYTaL5k79CjrCmj8MkgAciIYw
GpZ7Qk0X60Ry6z2tNIzwtkSK1kASkVBGCHLUefOEW++ZVOm6V+eO9GqChB5y4Dxd
TxsFRIiu3+JAxMgd08petTNntHHy6mD0XO8RJ+dpGqUDrOQU3naz5QmF4ZIcBUUf
/2yIgSxJ3M8ThI04ZsHLcvrIU0tS5BF37zvrx8fkkCrqVwc4CToSu9BaILZmY423
sRj5eNxr2UGCFe0DNJPiDvbtp+tXo3wJiB/ZcLcZbcIxtKrY5W8s1HAc6CKItJ81
zgNyBZyfDeWA6uCcmVnp+3Jx4IKzcsLAv9zXsCVlKNpMeH6fy8aORVhQlDD11T+k
pouZuOTOTDWFCEMnuc18BrN+9NSxe7lKZ3F0WMcPrAIL7D6xk0eZHGWhcptafmO9
EQztH/0RbviUkbJpEQ/PVNbTZmx4AjH27AtWxH/Tn34KII0jIrRtEFJKhmkrWWsP
zbIa2LT3EUUKATA8V4OwguCZ3mUSqvUGUhoZskEHKZo0MhpJXgQdle1hF1AA+c0E
znkdtIni+O7lNK9A2iK+dKXv0qbtzA030SGRZwDv1hc=
`protect END_PROTECTED
