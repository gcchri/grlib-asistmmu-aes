`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
esKMoLwil4Zh6Y31F2aGGue0wHkYHzae73nmQ7HR73E18mVVO0RHohZEGAK9b00m
+bYV8XCLi36jDcabmi6eQEUd3rAk8J7svox8TkdX8nYhHrkw5dkuiDfnJchMpOt7
phflUijKfG+nDfpBkGYoM4IxwXCQ9xqKUQc3+mTxH1b4A9/WbfgK0u7r4MCooGpC
ALRgZBTAbwjfG8060MfwBTklP3RsuK4H03hLZ7LA0fc+wLQFe/XYGtX0IYbK/NDQ
f+zhi33JvBAgGwlb5DQc3hV2di0uvW3OcaGulfXaxoIwSBQ7j6VlLrUY20APNQlX
xNBlVwzwJHxmRbtlFEEuT43FiiL5ItsbhtGSHsELUJt5rzHXT3FOoPVTtHQ3wu4t
RU/8lXKDsfr0u27UWqUqP66OS+jyA68t70x/fWXobe+I4KwYnYu1w9f5SFFWhpUz
csPNShKLHgVyxRyivYgMiTHWpS9md4GQ+k6ifzDwoTrMB8WW1QpqXlPU/ZzJCA4x
PIhCY+BgMRykLPMSY6WuoPk83funiQ20UCdPpyQpobTra3yB8p70odQRlf8oa8Jp
sFNEH1ZUscCv6XreDX8T/TnqmreWMGYrxTDoIO9CQO8=
`protect END_PROTECTED
