`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i41fhXyJVZ1ucY1PFf7/tUM5opzmP2MFv7ZZ6uYgdddJpZ0+qZCaELGs5rzT1H07
FeaFjjyCbjQ3RHqHrbAF5pUnKrRp8qF2agNDF7kxVgVUuziuwQVDkBylJbvxp/Un
n88XrR/J/WBiQEN8SPcacvmaTbWmzabZqeqY5kFcSF4yjiN9upZAH0qB4md60bqY
hI8/B7xqz/8lWZO61qxdOW/R0hEX1I9tXhU0tiJpwmiGFYWFhklfHwPPchzEDQnr
WHfzn7GoWXnfm1ee8D3AecWB159ZBem8pRNVE2nd6IQ0iOaekzT3L2FT7qUrz0nE
YmjfiQgs8Gw0U0dX2DzZePE1LIC4kIyYrELx4+Hsi/olEGsQ1Q1XtdIgvTKqHSfA
0QgCT+XiPi8egZIZK7cnpmlW33mdXGwxvBeCgqWVLfLYPp7pLstS6HH517F+9kfn
CmrgBQQkbeA0jDJXCEk9ghwsuTGEFZET7IJBnMHDiETXZPvHOFx3Gg6dnIVm1usv
KZA3BNRHSXzllX/Wr2FEeKEhus1G7jjekkvem3UOlosiWbjiTKFkAZo4B7cfDjLy
GHaEals9hxZ+1pS1s2KHzS3S1u44sekcaOdgFsPJhikI+vVJDZA+7X7kqiR0TfEG
5TIlftAc514J7OVIFoJT+JCCHMB/yW6XxlGAG5x9HrT7JpQcxHA7DY6OZ5++IITR
o+DbU+skAS/GCyRsYabVHfsDmLE9LAcDBR/k+ptrafh3U24+lijU2mxq8n8DfbKb
viSBIsIZFHeHkIppsz3vj03siJU3YZI1OD7uSQ9xA0wOQBeV4/wGALKgBpeiXhhg
11vdgDyNZHoroeqxKviz8MVjwpbJSlD8+JdXfxNCf66dRVBEtwFH1drWwkvpGVQV
xqzu3wc3zWgnrSt/1zMzD8sSeO/mUL4xFijpfgYkU4/ApnNCFN6rh7s6mNavETYi
RmgmVvdv+56mT7EpV0qCgcabnlqQ1ydE+lTWuhnZ6TE4u3Tdo/ajB0nrZWEfxP1W
9sjwaNKAC3yjidVtmpoWCsZq1FvSkaPKmhoO1J5NLL/PtjrnW1fnQIb7kPXMo412
lMJXhWA09uyRelBypBTME4Ce0cAUQY7P458sE90ORDXDBEBbgZsNhUajAOTqzJIP
kR2JDutKKGqdUGo64CkApUZD27f+zEU4RiGUDxFELUjaEQSBCZCYnpt2nTXjLc8k
58X9aH1f6lh7JHEAU0NrVL3nfPZvhCUIMlvoiZZmWE+pfmPxOWvyx4oZMtiqo2Dl
uo5zIYQtKjX/kFJYr7gMjY6PojIr4wdilmZX9UQHY2T8r16+r9lM6gk4/oY2Cfnt
ce30ylBEwnx1Xp+6nVYqFOyw34UebjxpTy3HApO5QumbjCLUORzB2JoPiHT9Z9hI
aTx3t2mGQm37YBD6lXXrbUd8+TTOz0vPtr0aetK8TnFzTH5RU1JOURX+VPnnHExB
T2BXxEn5GAvlkJM4PzbKhqYq5eANHOjI/5DM5liPRfskynh7cynaR8att3Jc3T/6
8P+OlP/uxeZRGrLmh9+1KVqz02GxgI2R6kGY9FVR77fCemN0r1YWtHIHiGPwEnYe
+HNBNZw60PyaNNEGYEb/OPc1SGVQZ2ncpNXNn3sp532DKQtzLrwYJTlbNQnicA4z
`protect END_PROTECTED
