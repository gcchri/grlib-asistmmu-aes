`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ip2eNw6EbaQtEbCBbWq2pqJcg2psm5DoCqNbsSX/HONPjtFbW5tAgrw3FXNxnQqD
VoXEZnd+h30vSTWesBpQMhfiFgLXvBpbekXFeA9ublT4O3FhpADRuoxJIqA5Ock0
fUSxVxO1G1KOPK0D1ErWeXB5nJTz7AcEuZRRleb/Rw4HtQUx2QIdjbKE+eT+2zz1
h+Do5Mm8G8MPGX9Kukbs7UJRv6xi+sMOQ4VtUJ8ji/hDpW1+cbrPPZgAcRxGKqaW
KmJYJhDTdsWDQrQ67syeF91X6J5I4ggtPIDvEupqVNTkKy8oNJU/zMOD5eVKmK7x
OBdYReekshMh5UjJkl/vAwTiv7ym/XDPV4WsZCWrjWhuchxfTh8dc+8eDeqWNu0E
8inwWWUUraLZPpVwAFkf5g==
`protect END_PROTECTED
