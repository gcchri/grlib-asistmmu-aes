`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eb+/2FOMYrSeq9JFjlm1zOaU2GuPVr3J3SwXKfn6mQp9klz69yuhtdwtriOJ3N5I
zOhcz6wuMOZa75bMYZZ+MQW0NzM+5QG3x2NoM7LWGIlbree0AmUq3Ktue6PhTLpK
1jFH0Dr4DIEBuGg37zcrUe0zfpuTGmlv/YnYcP/iGJsas/46AGVaVqRRE8HntkTb
+/zVHsuVe+gB78ebW017FO5WIlcy1Dcayn40ytLUQ6KNoduv+8nbGTILgysGI/ma
wDqSh1VPTmW4hMgYk3v9W1nnLf4OaNcK3LM0todQFeUJ9pP1nPLlieoh7KRaSUCf
dhufJ3HPAj1mP5rxctCWLgVPf0wUf0N7QmbylFQQpdYA43jyXF6LtD+gpSHIStQG
oojJB5LffPj+bHg3WrxX0mAYdi8rmGuiwg6Dq/aH5jt92svrzxl0rZtZCWtHeach
gOwoX6ZzftGS7qSZR+3Oj9aL21L1hYpz/G3/m5VaGy9Ru4tuRZjNjW9YKZzObvEy
7Fb7Sx+aw7dfvlO8xueox0MnQW9eSwIjYslxVTyWwVDIjkXOeSYFFguT6IoQQNQo
jqTWwCQ2hdSTU1PKok10eFeZ0ME1CpOWODx6B1xNZAXnK3AxHB+rQxwdLh09RH3J
fYuD+VrPCdQaQXgEa+vgHS1AXysD2yWYY7gf+RGqYnyiMR85DENdvcdLxQ27MEyw
Uxuq+Iks7FSKSefJ4dlZ0g==
`protect END_PROTECTED
