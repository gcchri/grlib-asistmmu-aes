`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ckJ15GuzZU8dcFwZymi4z5FOUwwh6r/ePU+3klpAK54Vj9bZFF0fcfJBt8MSVt9w
Qv6OAhKQeOYEMsYGjCsS2t+pxibd0TmN0rC65bicYLkeoYj95isXuIzBbjB9+ksZ
qhQfE79LtDMeaUbd+SRpqA==
`protect END_PROTECTED
