`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G8CpXtio7yV9kBqeSTsLtVGGuxZ7+vCENq+Y42DUBumI/+K8+CBn83pz2wAEFGxS
wB8gOJYQEhDUs6+yvCMZt/oIHXv6maLMMS5kh44BUr67KQYVfVCY3vGhEpEZORSP
SHpMsdeWGf3tmk6b8oDbqrK32JJHwZjaI43Y9wPrKhYQLiNsVgaemV3aaIY43pVT
LGdJXIutm7FC8APhtjcZyLbPwH7xeBwRyTh+twqMaEr/NO7gapHjAQW0ZQ9MJlLF
doHvj6j70E0ciaa8/+A68HitQSkQyrUPtPqVt25EYDJYIuI6D5CmqQNGbLTi609q
a17+NKi6c7QQfvPudUJzZ5k4RMQ8VYnJiW2UKKRoHWNHNyWhBZDyiAaQN1G82/Yt
pkM5lVetPOdqfOOjyHZkiT+Y7HKA1w5iZVbgbhcKl/WltNKQjd5GJkygxqKJ/KOM
vyozoRopB13A/QqziF1cH7X0uXI5fL0tMk8lPzlFiBElaH2IK9TZ/3tcZg2FoSZm
NihTr3tmxwuvk1yJz4dHoZTmmS+QlYlKyEMbjVmD4b+LAkDLyXHw3Zx0B4vMZkEj
GGIe7gvfYdB+aeQKdwDgvmGTYgualCMAsxUDD1ZOZeE8taH7yqZUih7FrB6YiTC3
/43pO3tHCoQUcKmCZYNaddp0yow3t+Lo4bk9+hPEXwpV13QK6maxH5mL+C1QRGtG
EQ8E7fXJy+MXBECu95/hsAag3efHumaQXtC/kCRa8rDXj9HO74KNv+CL3XMfpGBz
O0P8ua7ucLPOb9+DTk3delXuFL9eGsYAB9Fd2fhW9kdZVIBkNkoVhcwgFqlLZDVE
JyyJBbAPo4Le9fs4jo2cOBCqFU6/eijIfFjwRpZEq6rvQA4aV/tb7JzUxXp1EG+g
RSPYz2eR6zg+DY3ZYCwa+1XeamXEbKpt/yW2AYaxaR6uBus4Ls2AnizpIjnOXEO+
I017Dj8RiE7O44bnGE392OmvQ4EpAhHRI3XHsU378VK8LDSSl/nxIfptQJqx2ljg
gYcHHmZoTVm679U9xQ7d284+r20OjJq7ju9bLIg0IXai8t8QUdnWId01U8xbL4oS
FCa1z3QnsuhJu7Y+bOsMLlgq2RMpmKAvyU4QgfXogV634snU2LoDI+9ANYcHlcez
NWcAaSd/5rc3QUDPE9PMZ8IzHStDFQZ9+87LPAk3cKouGY2McEkxoLOXe1l5l5Xl
C8IaU4DTiRm4ARQTY8dXwZYeFdE3nKiexv4LRS2as7/BldZzzWyP4TgfjeVKJv8U
dXmGbovIRZdt9djtlPTUaq6qBVAqjzYEoJ75nkGMbGjUhx+WuRT6HLyKzTwruEv7
wxXOmAbhs6ye0a5XbykB5nSZFcJG5B6gaxKn4rddpLlMyQZZY+oMXbIJP9fhJEN3
ga1mNiYmu39z9GgSMpMU5FVw7J4jf07zC9p/R2zC5sQK3EfxcFn7axBs1Me5+8Fi
JUZmWFeClVu2NdYXUTeXrhd3cWJISV5yE5ZR68yFTMC2qsTZHWu6pkfMlGmRkDhL
cEnpFIQ0um5M4yNhnRMUGEJEl6ueHzc0R0DeqkMZBE3PflLCxOoGD4LFc4BbDPyJ
SFeUcUFVJKtI/zMMRK4J9rXrl8bNlSaOHzj+M21FGRO0oq3IKGgMRVv9kcko7f48
gRuMNmHM0ZaqDY/HMRZc/TcJ/uNakvQaHbubWO5hlvvOdClNmTZbFf49CUNaP25P
zHm+ZXVUYTNpBP6zlvazhiEvfCt5mrQ0nBPsttuIVkhbKS3ixpJHvDLTjFXOmxgV
okF//NBdrgTxajx0JqPqFJ1/bCwxAhAxnRTyaKOkQS6by2dgNW+jPtZNCYDKWM+w
Hg6RD6/Nqdi1HyF9iykXEXe41D4XpcAm4J8fB0BxGHId542IJbOgfMgNFykDWwMD
j38mwAwoUCd1kEkyfignYO32kQE9UVIa3fgBUiVbcnPrgbHVYDQFa+49MdxulBA6
MSNQcOgiepsWO5EOcbKlFqAXwk6jgBnBeioADYa2dHzc792wu04SAGnHMQJKqFhl
dW0j+D9cpnYqeVZcMxmOC9SYUpl28XeTr7sA6P5OQSjX0ErYXwF8di/lok/r919j
TtVji6p9HE5VxUaGKgSEF2gHgA3tBiFz9j0WGWLss1xNPSaz9waNrr3c0Pav0oGA
mBnsUyeTmJ+6bi2MC20LC2d8VlNQSkT93s7sfvxwbi941mSECrVJV54BMvU2ePzj
+h3VTeQMoc39lKd0iRSdhHSgyf+b5+n49Ga5nXB9r//PxYlMdk/X/SZL3KXtEHEr
DzMUixlMZiGNzpnaNBzXbJgiKRtQ94UWm/xFkWQ7re4661hf+NPCv/PvW+ijEfBQ
VHLbED2uxGl7uN+F3tr5a1yeDRrndYMgkpY3FzPB8T75gnPeVNkgSvMW7yADOozz
Y9tMVQ/YF8v6lNOeOmE73PQ8Sn/gUPhMV5DT9gZ8dnur71DwnGBqngZNZdb55iV4
g1dTvzd8UJ1untkSJyVTxEi12AKYLFPImU5dtroN36ewiUwVpNWUE2iSe6TRr1e7
jK/qERV3aR2uZOtLhKQ5Jz5AHsZxP3LjHvwBgnVwm4zL/ap5n18TogGvSfuGUfxb
x3Qyo/4KJHVVAITepTD5KczCvCJdr45mxWciwywWq1Y=
`protect END_PROTECTED
