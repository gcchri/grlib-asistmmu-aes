`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sokOl47GXYRYbwTXfYTKY4dz5XDktTjWBHj35sPNGxoGd7midyAXbUZKyobznxfV
JsdQauGUQ0zDJzpo3ELdkYvHehbQd0gKCHbQWJNNxcbwX4BwxA3vQ/LebxKak3KN
LwMOrHqlTtRjrXam6NFvQoVHFr/Nsnn2uuOANcmCCFEyHNkwSvRSh8IYhMsHmU0d
RYGxFN0d3b+RipkNRNlJmln0gmzsLiNP6RLO2zZdTod5QP9bq//EvVGsvfOjEqtH
3r+VK6BzsuFY/MF++DWV5DRg0uNLPA5TZPHYF1jLVRAqbVAIhKs+Z+fKsEjx1eNP
crCuzLpDWMkgTHKz8SA1UJ47aIpnBdIC10YeA59vfYCHnKDr2J/7qg5LBQSFMu6l
/BBLA+j9Yh7GSmWDwCV2ULR2i53BAGKW08m8jsGm36CgTlCNuLd+1HngGg6R1mrm
nVsaZVpnV9dLxDvCMVXevwWTWIeNWCfTigOs1FnHMaBn+N55mYuUFUXAL0cN3PcJ
0v2zj5DPhWpVqgy53okUQqn02CwcpInLmiwN+PHSqwmKA+9lse2vSBrVpHJMrHWp
UB5gZRW86E6nijQEB1wKzZI3CN95dGIGqAVl33QrFLTgDFYgyiC/wADHncO7SNfh
Sq/NCKFnFHl9SDvrp0c76vM0c0kNvCQShi+OAJGrBCWg4MtVfHqujmvaSnkGZmit
l47pydXjYohvsMnW+o6YRO3CLf5xVMVpUAdLA6fmQX4=
`protect END_PROTECTED
