`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dYeLzmSMnys0j0QPVHGht62gQXCfa2+LcG3/vsIQTpKab3RBOSxFUa1m4pLQlx/2
+FAdYAhZx3hY8ED5gjt9OnyaiQTXc/ZgCMlGccdKfIcFXd8elg00whOWfFHRlY/a
QNKsy+N6X1fuM7NsqoqQkwIMJx8l2IgPPrLscxQKh7sntp7QXEnTZrA/QJQ/WnB1
ySAFcdzVQ4e7ISDAr9+OsWpa8d1JfA67u+AQn64PuHzvNRpbmLxgtcnozHg8hzQc
2M1+B+ROGLbz9DP2ebOxu77ppaOIPkviuhNBMXAj33p2CD1OR/uFGmGmMrYNaDz3
ww78jiXzXCwmP+HEXCGk//XFsMDugkWvzux32t1+2XZYExkfs36zyfu54X3cg27N
o1KPimoaqtSi/DewNedZCto17emeNtsIXxdFPi9Y8/8LJeO/l1h8fyh6o5jF0cEF
BgSQmJ10moQ4ZEiKsn/70tQrbv0LOgLqm9y4H2D0NY/efumltjuqvxmHE0tKUhwi
OPfAcBF1dB+VQlY9W1p6xsFLJncHREQq7mpzAvDdeSeNmYdRksKZWXzGYUVOFW3E
J1OpU8uYMSpOKuRDf027Dy/oS9N6VTM+xLYXXNnjUtzSea6STuh6YwjwjNcGtpIY
oG+G24XSA1yvPkJYTH7VTgpd6/YtokfvWAC7pUzvG0YF1/QGR78TWjy9UzPO2PKb
7SL/+tr1zq4o352qBooCtTLj0khX7CxahrIds/I8jM5m6/eYzYucMV/sMwa6FjTg
7YrD3ddshWA+EdTEYuHtBhu+1qP9uuYnxwnKyqLCIPQTIn1oFuYzwUgz34APoByC
06UQqgBADokSWbh+uxkEGMpFlJ8aN+xLlYiwDaZfRcWEEPx8nCG9DCVrdQaF+Gbs
Uluj/gsTeYJBBeQ1rLQw7UgEMm4/X2SIjp9XYC3k5aEDLAf7/D/1F1nm7DYt4fR0
3JWrtgfhDsFtwxlazt7CpGMd1CI5OvmEevLvUeCnfcCKsl8SSdpB+1VWw3v2rHzx
tHsrYDF9ccguiBQnR+frbxcaCp/1aOODewQU6EuWDhyrZteRjBMj1YjEMZm0YOwj
vMe3ksd/gCrJamW7nM+glx5NSU4fiAUbNi27EbvxDngdaYD+G8zd5KkFyqrW46CV
Fe6OkxdAughnaWxeZa1VazYiDaX3tumZEP6afFKHsqXqpTPZ9dybh8Z7fyi/aFE2
nfwAbd7puBKT7tJNLTU20+/fUsy6JAk0pDZAh8YEDQ607KrYtBc0bRzlIUmwyoaK
zdMzXor73VYBhc+ZxriQ7W+mClVuTu0oI8EWEgJKZDc6pS7BnzolXq4IiHDTJvww
X2MwssclshRjEq7o0MX4vC0pxfIPywl/USaS0Awep6Nw0sXWuF9sZi6Lp8swsdUQ
gEUrvqC7yZlGHHCx6NJtOywSz3XdngF6oLZ1A7+WdNPViTGEg3E4o6pODvBCCIKr
/N+kWgapa9N/vv0A4rtxIlQv+Bc7iKtF3/J292M9SAyHMqxOoliJxTHfv5XASqZu
gpFgfA454cA+tQvXnaj4eZS9T4yl8vmZ09a2AD4fKF9ALBw2hWpFPQg+yaveHX1L
VI6qKzlbjcfA7vj8QWvhe8h+vYk1Q+fozgXxCv57MLL8S5FcP5KGQS5/AZJWpGiy
gknD97oNba9oTJ26ywZqi4rh02wGva7OthP1sNs/A6Fya7rmsqyz8eUDag1oIAZr
OivMLMEin3Lr388sDMNSrRubFU04DjpF+wl30Pgdchcu/hxqrJSVFtHVgR1LhnT9
uJvfqDVJmy08Ook5D+041tSBKEMcbdilbi0+A1giQITXchFhVPdbS9BXYNoYhBc+
CXEGeHCTQFfcfdRkZYYQ5I5pl7c90fhhfrp/zvoV8Ab96wrcCIWc2GaoMhBlNDj0
o+bU4kiCX1Gxs3AQFHRhxZL6F/UX7E2vh63jXm3f44S1JdTU9fdvaG67sdQLwqGg
1VGvHfD0GKpZvdSAGjLA8ukFcUCGXwfDIflwBbY2qqetv78G2KFYuefdkw+sPLPf
OKX4TtMKIzYxl3dCxkPT0vYMYyvTY0Wi5fdK+MznWSTCzMG70PS4RiCNimOmARCA
97j433rpn0PzZZBqWq4/zoSWDkK3CEeqy4lqzsNtQcXTGOpEZhK0rSZlULHQeGn7
oR9hArn2cbnI0vPPoj2l09y3PE1fvI0rBXN3EJhsVJfzJiZb3DU6RVck1USLRlzs
MsrjeZSrJA8FKqSCHMv8BXzMoJbaZ0wGwOH0tb4KZ7aMrTTkLKyM8xn0LU/pLp6a
H+TbfcxgdN7kzb4OgfjKmDN2Yf/MrhQaTECZPt9zRJCl5NCWfbGRM1ZprGsVAjbM
CtSdT/q9KuBBjF7BKl+XuduXpKUP00O43iXyqkpfgDOgrp6FkjI/YzspHAz9uY74
Btw7dyElkbVERaO0J9IDOuIg/hbhO9M87DZFCslERpqxsyQnJffSjDczvEboGOkF
h3482PE4vkcabKZpIF3vtIgSY/mN+iVB/E3z9nXYgdOM8ng1fwp3M+kXVkzp0RUR
m5ief4a60VKpCNyMQ4Q87B5+buvP0L0sMH/K01HjyVIGxXBKh0hbXWs3Oxs8y9ex
3RTa4CUq19eEbT7QhgUHVDreirfQY3SCiTNchMomEoNwG8Psg3NKHbzu4gJx8lgW
TY91F59x6c3JXlp0fQ5h2ooInJfV/HA4Qoag6WBcnlMZy4j8v5VAAdUiffvnAcXJ
srTNn/oc4a362vUpMr1rAFJ9Gaw456WxpQVPKhntnPL8oyQ5icJwgSPA4T86p2xk
0IehE57R8GU7LPCUqoKpNanGDrw+y6Q6l24jiVOd9BD9ASrR+lCzTgyfoXKreUZX
NWpimt1iNGmX9azihsSNOXwj9si4nteQ514P9Unvu/D8y64NKHuwWe781uNpagCN
iUnw+QKEhmukU8FVKMK89wDl2PddcVUOz9JB25vxxyCfQTk9QiiyRuQmr3sireQX
IVVZK3Y3pidnLX9jqepFj1jb8YDoUZ1B6OPOygrXOa1tjsCpqw95m8z84R05yGrf
ovCxuJSSDwYrwEBjK4Qg3J70jrWjrHCjZsOnBvUaJekXNq/pchJaQo3vYeoiHcay
bn0YYCHMcK9D9HEPj6cXRJPjFObtI9uz0u4FOG19Nb7NoFDQp1fv7TEsJ4adh2Sz
TgybMw0IQ9w35RET+a9xCMj4ycKgUx6whrojJlxTWJPbNcGb1VrclbK2I2QgNdiz
xdoxTX3k8ahN02pTVOMJ0nDcldoOLAy34pg/v3CNGm3z2CDgoEiY5jDV8NuOode9
v6hLi75zYuxnn0oSL/Qwd6t2Hy46a81XWVtFvFE0d8Mql+cOvBWrJxjyKsTlrr9f
TxDMq6PXVHaM1H/LP+px/1KObiizX3iT+ZCUVv8sjzEp5sKnHhEV0QWaCML4i+1N
J2p0tb0vOh5XlXVSaKDP61LbadKxctc68nJClL0rzineCbvonoW1W9oCn4crjsVO
Kf/2/L1uugPxdrwQfQOuQ9nDwOpsP5+qoau9YZczkvDKPf/3c0S6iZmi7VTSoVbp
ALytQxKWHbaYxue47abcGrWhUl6iKRXGTYD77oBQPAlCPPo8A7ays6zMNaUV50uc
tKNKtn5iVDsA5CS0QaJnZL4CzcP7S20wtYrmBKUMZNEo4c4fjJelphjl5EBEiuu5
kqHqwz2Stv6PMK2nWXY2kA66CiJsOxnlI6xUnGNiOiZc5LrMo7lyQxUuHL7vvFD7
FbubhzHFJrUFtV702zsbUEglU/vcM5dnXtRyn3jBsTbpKt6aPpW34t/+yODSWXmw
trDiKZyKkfSZqh4OpOgau0v/tO1DL24DhTip21p4JxBS98DuTlk2Az4M1nZUmcGB
8jw6OSaiX0GTGRzLpV9fOcMMEHrBhIUgt9n7/R3tBRXJhwlazRr2glONiQW5khrV
fFhDOgko/M3t7xkNnB6/soV0jW8wtLjfZBGJiAkryfvzGLjEUAM34QKqAv2e14Xc
K+jnKObKnerPU2YuJMhDG19A0TPhqV+BWbSClzS9M+rmnIuhAigNjXiqqR0Iu36c
iYK7dT5Sx07vs6u1HdqLt3cWWZxzmZXuo/NK38uU2EEP7xGYJKNfdznKH3KwZ3Tw
l/FCOZSwTPdn+9/ZcQw7JHklxuCgYzAdLtGyYgL17gPceknyX+7CcPk09UBOsuIa
AGQVyrK8squ8U55Qqq8qeSZ4NwhmICP8A3AmvzMdoh3ANJEntfT9f8dv0KMd67vK
72upI0bBZwd1mrCNfN2OJP2S7tl8vhsFXn5F5ebzihBEH9mrTzdyiT04dt0nibgH
2kC/r2hjI9tAA3++3a1TVc6F2QOuok6FrA8vCB3av0GtF4bviWYI5Z8iLotj+Q9e
+ULeBepMFjKJFVzaSn+7BMmsPqW8h7mtpNKGZdrFHb/VPq7c07CGu4btjphT4RYh
nOXnUv16r2xAj3e045eXiJ5qUC/s0a3fSnNyWOy40ZKT6rfv0k6PuoBFw+mcc5rI
4xqq0SzGX68DLMEbyWP9b6vKEbfzul3bWmU26ts4+69YhPxN6hLh3kb0pPlzFNOY
P9nefC/l0X8D4DpJcooLxNc95YWAGXPIG2PFvM5kmDbbu4gadXu63gsVngeng++g
QpHLMQXshwiIAYg5/YQwSbTEdo7zVaD9Ekftaq1P4NDUAOLWxX97MPPlO+Z8n41B
kMo7Y4TaiMBwFQfOZvY29JdhickxP570p+TMuAJh3hwmKRW0bD93L9P3ZS8imIYo
/yj87FY6+5lCYwIuAo1AoEigAKsK52r18VGqGyt9MXv5WAtjRBYFpRkqB4Q4E/eI
BaCYGiWm3S+nmmfspH+WGpdc44xh8XbS5udaPor7AAV6LlROYtd8QZWsfs7WBZwQ
ihBDrqphu/RKhqKETC94G117TFcDCgPK7N6hAISqDIcee7pNaZFjFVniZtYTQg6F
C/zE4MkRo/tUO29O9B1t/E3ITMwBsu+HqrgwxHloJ4SBHOGe1lhYt+0gRRFbyJ5u
0MHK+opwFQrpWg9ZuRUQoEpRZk8ctJwAKbun9jr2L+kX4oanaeMh+8YQeGn7wmAy
hmEV2KjG+tCaAFIbiULcM3zmHkG/Vf/K9vSVqVwImVhrxpzAnBMYSeLHxS6ljiCs
56RG4BNEsgIB0iB4AihVoNlPodfZ7VivODJBU26P01HFoo7+RDKApcu2W0qnAGkC
H4ZSAPabukKYx2xR4yrPKcr1NKDxSTxlLluueCxijXD5s4dltyKVXtpq/ZjlP6hS
waLo6+KTwC3FXkwqDQd7SCxYqlMxhvricsuddHu+myp92ygMM8z6cdilpmxf0jk6
imWL/h1JuidJ0lJdM/4ctuUrE5CpqJDkjzTV2gwSSj77FF0pdxeMHqI40YkSdkQF
5c992dMwoFv9FJiIpeidz7w+VFdkECQS+OvAbgGXYvLWyj8hPKcOa1/nDoSOp2NQ
qOELvq3UUcqQ1mhOLwuhY0zf+dlvI/9ZTIMzZBLTycPZmEevybIHwmzwXIeUvb5A
hHbytlXP3s0TUl/HndRSYvDxbdZBCsSq1/KhAN3pgcnm9rrCewOvCoIwQZvs4yIJ
1Gr+70v30BEhnhEsnDjwTgxNmaL2GOq9fjVK1epRay5txZ+MdS0VeOUJ4goynM8O
YFHOo9yz2VJMR7aHp+/SCjiF6UkvHKOgCe5oMOijOvBbzWc4EHgyWXTv9s2UA1+q
6kAz4JUDtNS5s5yjXIjNk5ZW4+eG1HzT6P4OqYWTeBmsloDg74Hdwjy8nOmRAP2D
2rHYxQtq8IuPXMLGsQNGM9Ce+/f++ax0X61R8eugSP/UllwNsy7KHjl47up48NdC
KLx6HEwaDEK7n81Z/WFkdY9Eq8X4TSov68CYixT1uSsgUJsDWuoN4VnUNS5wG4Hh
Mr8P9kEjcEJO4t6cI6RYvn5QAw3IA6EWvFSbiJTVMjo6MY6GgsX9SKL1eRxNCCa5
cMvmgNT5QeFTSaL4LV5wXRjaLtZRyG5s+t0+WHpm3X+hkagVpTxLtBw2WP6k4LhN
UU2SdPshTwk52lY2bCnrVnt93Cb1tC3wfRxLOf+FA2TCF75C4sP/ic5xqXLJZd6N
uiqf2gyKZY9m1d24NbUcV2EnpZJY26tTQ6IPaWs6kHUGaHS0zgcKGVvL47kG+kWZ
D2ud098muXMpsLoPc/pC1B19kwTTEdg6spqYeXWWt5nzf8NpJgfyJGgF3qQa8HqX
uf7A/Kub67VDIJWLj6DxH4A/UivrHlF0So1/inhe/ai/RibIk46ukQQykvmBQd4M
ICQjKis3+P8eAB77MCauDdqykLPNr+b5wfYg+Qx3dmxr1boW63+c/Zmgc6FNzl+f
N92Is2caIzToGmlnYc/MMPWgFJDIgZiJJQwyC7qmCGDD1Nfxs+duL+OfAONBf1mW
k9xMOal1s+DwdBIi3oI5wvXBaGs4eTHai0ZxHVC2PykN7X21GhSzKK3FH3feqgdb
ugETjNkKs4mvgk3CBP8Q4C6LDi4Ov3rGGdVQGt927su4ggTpTgo/e7t87nHjqUoD
aYVROWHsvCJq6gpQCC0xPG83O99566h3iFAeGmWQqGsOkUFxp9RVg6Ky5Ig120jk
ouKa9DBtHqNeBbKTjme2tOraEiIGWk06V6r1T0vwOKsOYoVtvAPj7PUxN8xo/Z9T
B6OvBON6ppIeA/MV2WgA6c4tW5LzxX7pbQQGQR/qBzPZZHsTtMKCuQVR/Nt3CPfM
Dhfj5jPEdfwxMCC+t9+4RqMSTkJZnT2ijVgZlS0oARCWvU1WZtE6A11dH4d5HIK/
naqZOv8HMSoUDhzEDNn0t4BNBlIPm81fZldBaCQiqXNmjsRQ1c83kXWOIRMcar9P
zkFuiIu5dsS4Wk2zGriZO34ePOQKvPMj9gHjHgMHAN3jKH/GiNYXhQqfcl7KMIMz
bTReHBdD5N9aEuKuiXXy3ELcEZj3/PqPJJbkBoSUJwF7u3rMFuHaUJlR54qb/LEc
LghzYQ5rhBK8xSjXOBqs3AESVijrx0NSBqvBD3Uq/ohk+4ott7tzR2jig46GMKgZ
cnq5reJjHZyiTxkv8vFzPXi14dSaRwJma3obnSVVO00hPYr+DVRW/TsFTZsXWJgs
qfbvFeuHT57wS+wQLPZdYNqnXwutmgM3se3Ajcs9GuladCuV0dBtjmwl5hzN81Dc
YNH105M9J1+A3reswOZd26Mw4U/MnLoERkw3ogGlF3vhcfeZEYT2idhMCC2rjaOc
oEYUY/WV+FxXnRz3M+8D2mCf6gmf40282BQRWNyKuwvAiwWWYfY68+tanyBIxvbp
N4TjED2vD/V1dLd8vE4K6d9NUO1cpmqGTDxdUoWC6ViLH4LrFgHRPgbwUOOaMQri
Jnt7mDIfJloPmLTFjsKhvO/+C8V7/kADj9rCRp52kq/cMJefGPmN0NtFwWN18fkn
leh1Ow3s85iFpz24etCdKfVRCe3MHD0E/7PWGgQuW+zhow6DMHuOF3PAJN+j3KFr
V98LAJDoYcVlfx8A0xHKxq7kP6AhESEeGOYb+QA8lvbRTuwTQanek5sVMYUVs2V7
6o5dUjM0kvbbR/fjDXYBt55QgLJbPxtGg+CLKfUjW/o0HKcBJihs8o5xnHaqdYfv
EhLBKdadw8pcohv9U7QRUTpO45fdFD3iEkDgZEZO2slWxIV/nUqtY5ioCbDExlQd
87MtOEX9MM8XCFp+GR9sdT2t71wszGbhwVVxDYbDQGwGFMWVSFpNl+PF/AfwjrUY
3aWKXylMH2VizdXkQsf5E1Dj6jHuAKqGcsn5M+C9K7LKZLv41whDw6+OUdyi4YgZ
cCJO9uiW4OTpXzqlCvHAKWL+YEA8TN01R2Q/gfjTarRbbsgNay23Zh59naNslv86
nRu1H4d8ZZVcVzo1J5njvuO4Hb5kzusDlwJ0DB1t/XMMGWq1toq6Ez7pENWTH3b+
K4mcvcL/Q+7ZBUIh2WrXTQcExkMnt6a1olv1c0tmYcl3YkUL08IDWRoDNOrFMPvF
SEqXC1iYr++4qBfzZe5DXZVZbRRYEVuORJKIcjQL0oz6U7uwmQS9BtJYeKG6x0gc
2b8KgOms6f1UxW62lActjs45mAX8Qy9C3DD2LUWARlEW/gcRlbisF0rOOspqfYeg
29U/jiejzYwDYvo3w1iRvfknSfmcmN1mTbmAoM4aZLBd9RvKeXJp/TIm9ca7cdYU
LbOKG5VPXkDKbQZ3DZ8y58dX8yzajrCG57u7JiYSNlAldbDQCzW1AJq/ZNx62xC2
EYFxRuuRKrZCf4UdBA6o6T7NQCZunQ8fr0CmtLw1QnRNTObYXswSivYxyidvBixc
oIK7ENl2MpgTSKqyrRXBPi4QbGFcDfzbig3z5AyFs+V8x0zKC2UxSwQ8kRjKkwm5
hhlTiXxBK5soI7V81e1ZCVSFiM7x7KN7UHGaVyy0zHjpM39ZP/p+oz4YsV1q9Av5
cl3CnVKKKaXg8o/tuuEuor81vgNXY5QI5AwBSUm9qJGBrfml4TbY54UhF9r9sA8r
AXteoCyMnay1dqDXBxeS34X9f+bzzGDcIb52i8iH5gj5x37YCgzTJoFrGoqwqilI
HmB54puKILK5Y3erMUA/7RCkU694Yn5ScTts9C15UyaPl81bMvpLW8t/FB5eD46d
9TS7Y07NPoS4c5kUjbr+G6NRLxt6/sLPm5opH5YvlcGHMSqlZLQg4u7Up84dg+KP
Ug+tzfepqR2JCXEvEmcLHsAmHu8BN02bHI1AbcZS+tDwYg33Lcfp3Gq42ycrjCLN
kZ64nHIJdNCF5/BTwtIOJdCbKhgT4zGFqZtSjZX6oaqQe3ayPfb7ATXc/aBClO2C
+4f/B87XIKyE2Crb1thgrrEFhOyxlOSnN7e/TqZMxBhC89jfzuHhJvy7VUbb/ErP
Dv90ZXXAUlxv7XG3qKpRdiabCxJIVYKW68D5KQ7gawFc7fFm0/HekUhbIGhpVxFr
JWKkIb+Xw8vYL3JruKQQd4LwHa6dZtNLMmqsPCJOTb78NGmQpbWSGYciNoEG/6BM
2IyL4khKHIPfUu98jZ0lC18dnuVWGv7BRnnzolBaYDEaQS/H1EiFOxq5Y1UCwaGE
zyHwY6CkhB2cEDWhXE2Wc2EcL832Jedr359tZFmCbUO0kav/IaBbFZHYq+qjLuT/
QUdryj1r0nqSNFmWYAVhoC87AKUxIl9P8zKQXqMKz4gnNTJPs9SCtSscfsem2azd
PxfYcDoqkXfp1UvKkj6ktIEQg1DdrZzA+/b/VZhdBsoY6WWMNIRFedySkBWYjmOd
eyuJCoqP5w8d64FkwO0ROmT9a9ZzTskoklitkK3KNpj0v9iRNsZA4eLRBSzgQyQX
0wcR/NbNoY4rG6UqlQx/Xu9Q9zgOBfhpsCLSISadr06rCPQ4dJFZFNV+528WKrvL
HjV3d9+9pooKfsna+f5nbB5Xpf1iWhg1WrJQXRdHXfokxhyqv1Db8TOLnxZhHz1Q
UvKFCBTxOFkv0/MSFaJcm7iJ55HSnbJ0iSM9hpT5z08fSyqHxHSETW0k5AAnnHO8
qE7lZxbaWZk1xBvWdLzc6GEjbCFZDGmdSls4XMqJOunTi2vlqPhGivhfNU3GPobC
DrK+hz1i3PvIoUdiYc/DWyHTHqs2e8Ln4U+BakTkPX7FsbatNsHoXW7yi3i4KarX
iBQiwv0I1aylJN9yNBRzA30COKskc0U7dxEr4x/9cYHRP/b739HKQh4vD1hSsvu8
yDASgW9vs0h4j6WuC7QnlEr4AD/HxS3giFb128b7iF2ZXMtcRaXXXhgPpSXxvc61
inP4VhK4+hnCEhpzrRWeNSsc4UOj7Kl7Fnd30QLhIQGc/HVEdnJkPjxqjKdNNUoJ
unmjKiVMQD+eRFM8gzhlwqI0w6SslQx5M7FRX+2yRfrcdeBIUQ5ZEep/RNo00MWG
2bUFLgOGFqP7g60SoDjqyXroWD3x1cquK8f/uQpC6aWlraKU6+oC2lGvahcl5diP
1PT4KHjlFtlQNivunsjaBZ7HIy/po4LdzpQ8ybH0GxeiOoByraYrmJB6q73XSBzT
vQsvR5+L279yExNBAg2gzJGeeVqUXqrIdU11FqcF8Ogm9O1Dv+QcrcpXo5CFsXWq
zepTqgb960ySvdhD6cQ8I0cFO6dxqgEy9wyl5yhoGdDepck4v9wL0pBwwtBabTIY
ax8U9kYLVSXyYyslMMRKtP3ULQzwe2+QUNz12l6EnyTrW+yVqmHnyRBwoYUvEcpF
qHo59MqlOGlMYv2FKZ0l2mLv0yNStiqMqSIOG0qOd6G8OZC0iWWjiyWVX2o+V/Vk
jQT+DzsIGOU77gaHAC4zbghAFAeRiHJYS+7LE/egXIaJaLG7T1NDIHaf7PA3ssSy
M2KhhQ4eoJPmZeE9FjEB199jjoHoD0XMXHtxlDgsMeqUnUIgstA16djTt8OWmx3/
ZshbI+qV+toKj1AoIRmCvjkoYYPZkofV7rOfZjlQICEsgoOQE+1fPb17kGbexplY
AVFLW334m+ILbeKHP87sg+03KOewdCfzTS0exGSywUXDoo+1A8PZuc0NZCXCBO/c
s+v6mlH+6WSz775IwfaEE2V2mZIE4YNARQjlPO7vJJTX+DoqweiSRuQLHvX0ply+
KrxHoofhOIDgutTHy4R4/2400MHmXo2HA9NYS8tyydyh2tz0UK/ynCBsgiSptkn9
p6Nhj3CcaDxKOOxZNBG1dOhNEM9OnIN124Xf+II3fa3+GMLYaunLCTIsQPNbo4ig
/Q7wHltBx1uX9gTh+BKsLP3JS3e/HZ3F4uJkjYC3pPs8DySBjJMFbAkz7pPHw1wS
4ovzcnrxsft7sUBzEw56bW/Za9Z0vJSBe+TxA1RYXfY8dB/S3qB0kD38jaiH03r/
H9frNo7e1TSecssJBh/vhfNTvSSerqjdQuozzcF8A1FpFSWPlDe5ngrKqWYNfCwJ
WSCB+BwVrGxseK43NE1JvOUb3v2a+r3DvoVOCVBKkJLGZbtKH23LkClwc0ojR4ul
la0Px2m5Q7JG3/iLZQv+rZnvJjeFbJVuPPNwEEPtuDsqFJCqUdNudygaqtXyeoyd
CdURKIkz08ocMa/w+QvD6YUcA46vC/NYy9HQnMWpTVAJWwh4Ff0M5Phu3MwczJdx
d1t8UIPJp3TPsPA7R3wi2LmmcN0cg2N7oTRLO4iUhHFBZe3UnKKbEMYtekgzCDvl
SgIHS5v+eP8Xiby3ICn1VMYTM6aj+1i52YmRFR94rTFJ959vUaZdD9VUHH/H3UXW
DdtVlubc0GRbHuYa0OPvpx4WW0ru71hJJWsOYj6fNMr4qiyDQP9HD8NGR3Cu1H0T
Ke6pSiAuGs0XWlaT7aOlLgf70Qc5XBSCSukm0EBRmCxXFP8gvhnuWw4KmKIXOo2L
oTUckKTRq/gT6atKtx2g37nISA3weXUgYflon8tqAL428aillwdMRdavMMEWUWG+
hG/FyoBhH8eE9KqNlva8b7sZOLz7QWhAKIia0j4NzK/coDm5UNYpPyYoC/zyf19l
c3y+8Z3BTfsVZnh52dnBheOdGARj3GeuCiGyY8lEAmRGCnv+0i2MLgJ+uQ2HZPQe
JGYJBE/IL6cH1o65v67KZygf2TTZ16/DLhDfIfS/+NHl9X7RisUnN8R9kDb6WHB4
oqGcG5nJQ1rWbz4xrmCqrGyafyfzp6h5H4rrmeNusnWiBAfV3SawVJJY5Q3VFkJ9
41AYVEkSYWaC7x4VAwGZGuOF8D4ZL03EDuLErHIIxsy9Idqb9s1dKbsiDwa9Ukyu
Kf7ouyRyGlFlZg4FXYBkw00jNxKLJ1kSOPDW7/9suDIRQhjKspjiO+nEF7yKLpzL
nbJdrodsA3MtlM2ihCibvb0eE6u5bmTfrH418xLStc9adeBWvPRpiTtICGiw4C+u
4wXnRjGSMi2+E7J7/wvv6hORBldyRoBKTt6UVfYOcO8AmnYXUCiJLyaTpd5FsbR1
6OKXO8+/8bJGEUxSB7JpXpWOBC+LEihoiCYbp6lmHL+ZQr6Lo55r4IH3Qkj6XfCB
GnifyLIBweqUEQld/Ijc946emvH6YFbf6ibT5uTMUSfpOxNfEuCbzyicKIDk3rAv
l26EMJA4Nd2upxZYxHiELvMZJkUhZBSa9ssqeFkxJoAkAMjrMDKBeHsU+8xLU1r/
18lf1JrN5aR2eSTXRiuLbVLU2ozueIJ7TGL1FfaYJc5/exCokzjHVu5iDMjLY5Dp
n64AHrCqQOHvSIroqr3uucF7CymYZnYA1jraXQyOhy9bTIP9FtK8+envpPmqLxYl
ZHdvc5b+vbEcj+h98CbIwis/5596h6HCVfggzeMPP3T677wPqY5a3twetXB5Hk4z
CctkXzmXxfdjw/jjW/TrJ9yQGzNY8GnGXbetRtgcwk5uM31H+CtJFRd5mssveVE9
lwMdjPCkVrtNKUnoNUlIHZaRYAPmvWrRvSD1N9/L8k4MzvBLlyFxc9XtQAWwqJ/l
+rB7yykxpTjsqgRpwA93lEv7DsYx6x9qAtqq+9IwQJISzSU5cC9BrrE3Zdsl1Dl3
mS8/YKsehGF1H04APYu4XiO+wQ+MiXbnq0Rb54ENmJD5XCQ+7LT/4cAB6k2I+D8H
VgYONSqErpU+KZc5gebB5cAV7yyOCdOI9Uyrh/FAITzxyG0w4ZCtNHcvNg8lQafw
QTy5u+gNVIwZ9MG/I1faxFq+B0a/XVdsJfmw4Yogia+RCdjhLa9qOgHLytEqN3ri
qpfWh4inE5ufMQyepnVWJp2TNYtBUzuSCfvRsNKtJOSTtiULL4CRWBPPj8Ks+SpH
zKZgTX8jTWblH4HhAQSgMCLNy0rbWoNqhI1QnLTf+OQ/ruH4PjaUsXN4Cp1O3ia9
OwE+4+Re6908L55djYb/XLgHXRZZMOXhh0jkAkUwpvOY7e6VpIkDs2XKoFG3xmHx
G154SPIB5coNFvmW/6qya5vD7nbGVa6JP6XnY7EU9J6pMX/004i5pCLpQi9DM9Sw
UgZzoYvzZ2Bb1insltMpYIpJ5nlA5ya4K0XSK4sBOtIP5k5PYb6OyCE2iYF9ApVS
fcSqGxMVpyUvl07zt4WFQQpFiw6Exhyf1CRWV75NcxUY0CVh5DXU4c4c2sZ/lcgk
lhHa2KkULIclWylDVnfqsDazkI91EcdtDaLZE5fvxFRT9JgfJJMiUHrlAlqGOu/H
WD+1qZ+sD0cu0/Q7HymMaaMqwAKhLulU2lHT8rWLEMpXTXwGqzCMTcjbi5Xertkk
tYKp9CI5KQbOtEMqvBZuyZRF0L8GKeULys7RiGfxBcHoJ6TEfU/+QjzaSZVu4YdQ
HRruW4N89QFGmIN3QQWF1f5rNmg2PSDxdWhyndJE/tmwSdEk9fphFQe8craMNKLj
Jk2ceUrk52/c+r2bAkIsCnT5OHAg4STZ1Zt/lOxHInLAQkRk5GESzMj5JV5mHWQj
um4/BqHUKYjCx2ANiM5lczy6tCWn1DZtnErQDsez8/kTSpFanuRzSkdmlqVP030A
aWeCBrRmAlxCyHLxZcaZ2CefrkEFtcOEQBHivJrs/0XVw1fxZ6uVCenTFtp5J1cI
9cFSIAFj1blfTaLWKCdtrMxf+KVvjYcIiLXr2WRsXy73wH2N/1U2kSLSCsjH/foB
w44srW8/h87Hl186RnIcdLsPlkRB5XLdwGnkArCKpGK0tgxTi+Cu/3aH4PlL7SGM
ni9Q7W1ynnZX0tuGWsIzX7nG4YRckVRiJv3rrJxObjiUwEb2/UrSDZHmqJj1BIOV
jkxB3obOIC39ckJQ4G+BFE3yzueNlj9qeroPAFw+LTZ696760oA1CvbMDMa9qaFo
HbDCdLtMg6iEqytC91fCfysXzCP1VeBYhJAFtKNsyKpNP+kbki7KmOfIQPrcs74o
553P9AHfO96PddnfGELrkg08M16yKTdDRlabpBBtIn5H2ys9srjOviWmFkk7HlMX
mbmB1bI9kg1eqL4qQ2BWjPLIFhy4/42k90S2sPr/s0MvT0BmO7ZINMC8QFQl3DLk
AY0bBfDpsbfxGivyGFwnLqRhgmuH5DpgHbxIi+uuUom6M6i6VPR67EcX0W7fVSOb
QGPTXUzNl+N6DjyitjzItFnOjyVpP8ZV+Gf2hR9vzAPholqCpNPyBPxCST9V+eL5
F1ZMtN1+7BgsRbSfQ/AHg5vTjRbiEO2pLBfTbHidLmbE/OuroLNGceIr5s5r+P8Y
PsdTMN4Xx3fb5acvU6jhoayubKPzQoO1TKYhXcgGLOmls5FD2U4Bv8zN5KLsDAGk
IgloBzxlnLUckPLxgsnqj39qoTeNeRwtvLt+6vh4jgCgG6CIpcZ68GNkK63kXSLc
Ykq8vH2SefPRih+Sa6zI1OeturIzCiQfto09i62kKh2Lt5/zi9VPkC24OW52KwDv
d1JlEPKoWkAgC6Gc8SWgpK8rRrgdZTBWUX3edNEZkx4uxhb5kE7Rcm2B9rECM0Tr
xTVOjNw7JTfhXFcZkNNZAlQnqh/YA+XcKTS421oC6kBKNcBHAdUYXr1cGRRhPwnY
b6vMPDNzsEzaMaJVYzBCSsrZJRCi/TucY/GNXXhi8B6p+jQiBNuxzJg4EiEqT2HX
3GLRluROeNgz8qqnLZcWNtuUZRGa+tfF2EZlx6xNqvFkYfGFrGyluYDm5kGXtCnB
IOJEF4A0HHj7AEZCIWiLZVJWuj3eeI7aaNQaP1QV+/APaiWsZPT8M8IhK/4AOIhx
Kf5SK9bpvP9Dyo78TFWVLvO+UzSFwpi6Izew++MMQpIYsoK+ybQyI6MuHqnpz08h
TcV+5rLxnSODcYljAxqsxYKbWuGNO1g93VJzAW+9xSR49ZSdbaiU7ISbToCmJOCm
2dRVhbL3IPSrFu58Egm44Cn0QSW8Xly6CLcTgxf+HAVU7bGcffKkICoqxj39q/Zx
MvNgrfSGCCDDKjPn4SSwcl68oe8lLCkfNryFBYKfc74uyQhPPwuFCuMKhdQmKXDf
TTAvXq8gdY4vhlEuYh4cqk/Ws3tsPTflRzFmJL2Ilk6j6jeZfiluwFvKPHOkGOw7
r9ZEA4JavpbNiK69YwmddQflmr6YozG+aNAOaj9OFXw6yIYIdrZUFLYiSzyQaWvD
ZlRQjHhGzmsi3O8roItHdbXQpk2HNu5hnfffvpQDdgzFl4+hfzKfrTjFLaxc8pla
7rC0IzjTHbyY16tWLso+9bECAJe7bD2QNqNjEhFz5Ijz92h7Z1Wd3NDCPJFZhA7t
CFAfIIEx8SPzrlyQL1NFWGeCSVZRAzYTqBCkPb4KuEF6HkAvnonBKjSiCUVFTRyZ
IAO0QYa7nkjsQkA+cMMOo+0fbRZMXRV+Etj/sicUlPyMkpexBCJZASUlhEH5Suw4
AAXcZUXKNbDovHLYfQ0CY+oRPq3Cc25YTRZOsJr6OFignKNqa8fFxSu5qCOwNtAU
itFaSiP3wTL3nR/wV5mWA20uTqFy+g01UR8g7W+EZc7P8o9mSdvHxkooJDe5ds8S
a1iWJGuSutk14cLdbIVBKM3Qy47JVVIJ7a7NXw/qMdXFV1+y5ZGB+TT/U79yz+US
mNgaCDJGqEHX4SjOD1B339zwncdkBd+sb6vHe7CgBYiTJ1iLg03MNx1Z2Ieptq/5
j3u97odovXmxAo1+CFzOA+bjKQnE6VUpYQ4DzgPeIyykfs3l1L9WhXNopAcm9nb3
dMhSsAfmysWpZkOpgTSHFqbXT2InCw4r7JTHFvl0P4rBSueoGkSdzzaB7fSrMTf5
iJRXkTImObYOpVO6M65MsvAEmVjzjWgM3Sq0NZOJ3Le7GkScprAvz8VHnqr+qSWF
m6JBgvF1xG4gGXGXaB23xQG06oA2SUHlK+h+2Va13DvR6yVF36SDc719S8r2N2go
vkdq3l2WAyPega1OOlQCIduZN58AZ31r+t3lJ132p2k+YJUXTDxYWUKPKZR60uUu
wAMnKoZwDCW7P8dHUCE7EmKZg6+L26BoIMqFMiPpn+rx7WUesLNLU/p40jPHvG5E
FoSWxWVZQ42PinJmphavqPiSRvS9e95WEAdTmeoFbBbOj54khEj5vH4uoc2EQ8SX
BpgB6VWDD5IMFifiFiZ3EjhilMn1/2hKqpZb0N0RbgmgS3/YqF7yhgTlYauK+9kP
w5AEOh8b16Z2HZSqBcYDASM6glV3b/Z5bdU/e5H8HOhkTp+sERc58rggnmiSXcWh
yxmTpg/wjER9NAy3vFovk1X3xy8RsLLmMTeTUggYtb0vS15HamJcYcPJJ0UP+JUX
25Fnfzsm11WEq8da6K2mGSVgzFjFF3HE7OtSOmZlNtdwr+tWgSGWh15azyiYBP8F
B7UnpVZSVFwA+DHxWc/0UQwmR9zSKyhDUYaFXc3In79IEDMxLk2aPP7iyjuId4hw
gkMiv+LIMALDog+3Lw7uysaY0ytAbCDA3SQd7ukryCV1wVSbRiLCacee+il1ZwLG
WKNCTLEJmjo3H60zdpRZwXoLj9KWDTbFnj7+z2w5D7zUUTKbLkrc57SL1We0jEpq
BiCsWqr7rqZjslzmcIotMbM+WFDPLObN6ZJA+NGtmvuh2AigdS5QhBEB+trEp4Jj
yUPADBbtIQL0RCydpZJLPuYwhRBJ1Edq2le/44WQz4q8sLXXS7QCS+tSGX5uuWc/
or6IVGbXOyQ962OuPgVZD10IN3XA1ZcLi0JJwB4818mDHpGRUIbumXss+b6MaE4h
o6bXhu+liweBmuiCcdv28oUmu3CFX3Q+VGdkGtxCO0aZrJOfXKWta1ipDyRXpcTT
gFq+UAkt23l3JTgvtO8GtQ0TFWEAB3mpZdNw6BrPIco0WNeuHR9DPk8dbpU7tYMj
VB3e5KCLbXxpRkB9jA2JRpYw67m+Cl2JMHpqqromqoUgBUaYEcq8kHX1jnAgmCAZ
t/bIHnvAg6F6oDtMi8L/3YlkXQcrFa0Sorr1Klu0KM5deR6yO0s9IZetgOVewqmR
GmjWspl8N6gderX8xIcuFyFcDJWo/6c+nt8LfQHsZix8M4GSIBOcxD4Rho/BXUS4
InSSe4eZ/khqqTaXG09VMKLXDSxvjnHmLHFa6GonioUIztr9LGGzoeqiggBI7e0Z
3b1vioeaGp5MUvh5RWyE40rfWzmgYFuZ2gnO7wtmg//ZxAH9n3nytT057xIrnkTL
COYehr1VFg0epSzPgdqfy/4A3HinuFMBPR9svkZZR7UHn4EtJbcbGr9+pKANGPVQ
Lpg8g0GioqFpKKQYTybvvwrFoR8gcf7txK3F+3hyXSuBolFP20NT1ecI23Xr1yhG
iP4gqBUGj11tSfoPjqYbkofFzGXOVXmBvmWQrkmeQdoJpAeHzOWPDZYsBUj9ac2Z
jh33tjZTHe7x+ubnuNEqlOpxDg7MJa/GX3srgCZHjUxPM/rcWYRAROS4oujOlnL3
ELaG5MOhMxtIQFenTJki55yqCUj/ZPYh+Syo9EV21mYXaRnuqY7t8IZ1wtWdDIGj
hB2vl8+Y8w1f2AuAKNNRcYyAEHdOgAJXJBxH4lTGl5BkQHlvFmbnWlj3jF4Hf2PX
CQ/yEZyGnBv4LujCFcjHdciKWh6P00PrFZioM2dVGF3gY0U0M41CZPAJKrBHNFd8
dN4Ke5X4IEJQOoX+RcBIF3weksvDS785MJTJtWmE7QhFU353cPsi6lNke5pv79Hr
8i+nlrQy5BM+DW+IM0TVt6ANK7AH+5EClphuXUDXgUbBT11fsT6OFmOHnFRY89bA
3pp2vEn/xi8wX4a75OjKmrkTy8/UCiVnGrO0M0dBsietFf051YMEYtuGvdMp2pto
Q/UGgROwksHHq+gu/2YQRcK1sFexPdWX0AvSogH+bx0RiIzxKIyQB95BTcPIlMMs
xa0HfngAi4tOb52s0OpYFl0nJAFpgeVvKrVR4wXWi/FUUSpdYhxugBImtWPYyXIS
aNhHkFmwClWsJx0pdcNaE9WkFTgDKq9PmUThMPK04QOG3FQT2INJIEqcDL3oFSbf
UaAbNu26fy4jI5Wpqj5A75Yg2f/bUQrsHSpQgVAoz4neeqbGLxomD481J9ttz75L
qyiIwaHwV0itmWeKFTHW5MGx/rxLKsOXNIkBMbl/vONtiTiD9LKd2x20+qUxuU4l
5znPlYFX6wdKl/J9io9V3mJkUS4rBWfNG+MbiSzQVX3fFrdbrBmBfbkkMqXBAgLx
+w474JHUNK0JcmE+CD+7Xa13J3mTbITQLbPWjyqZDliATxiniqGuQowUa8Rc6QY2
OB0guO4SouzSTbjKUMtEA2sbbJoD16YTRMTnCRYFNtO/ILSAlOFkZqFwjC95EBl1
z4Ew3buvq/k9Yg5qUw0rkHwP8oJhldvpPq+kwH/bt+BYJCfK3/ICaa6YTa0uaXrg
byNKc586zR6p5gVzh9lZHcda1lQjqRaW2UQBu30H95sD8khYuyxb2MsnSSpSJfff
FYxVa9sQ43slRHUF9QnxItRiseU0TQwZOkhf2gqCMe21w/Lov2TuHR8QhPxfHPW6
CuIjSlT34dUmf4Yx8NtOiJ0nufxPvM9H2bE755i6fX3cOL27tBITuON93dG7O2bo
SC7LPEvzrpVvnvZtONblROKqc9g30ociwebyXWzoh1+W/do2yoawSFT4HDidS1Cj
YPRC+UxD9/9pwE3zO4LvrMcy9lm4s5tBBGtMGyvH8FcsDIlGCThdeRtCRTfTUHhg
kKT9oajXGa+3WLV2AWlrwpNmmML6/Not0Lqnam0e7NHYZu6VtV8CZ5rXU180Ya9S
DvXoopHISMqo0apcum+sFBH38zx0hl66otuliDiypbd1OP1AbWg/bcjiRA2Ijej3
+2DdKuwUz+qvjFv8rUgvj0ESsa/FSsfvYtLhCpcnYDY9qLSLXxbd7mwj+/5MKH44
89G3tUGH+zw/skdU6kSsCaMSMV47lfB8tBPff8gOQ8aloVhZrEycHRazX6XmjfAz
qHb5cr5vpG4oDzlvcdRzQTftknoApdDV3iGSnrvKLsjJawZd49Vr6zeeCgL9GI3S
rhFPXDfbo4V3mLFeXrbHkGCrXumTDKSLq77DpdVRafaI/naJhYwjsx4Yw43DX0tP
ZYNXKfc4DzlVK07b6YBHjYF8NRzGtnxz2NSt04mne4p+IQo/sfW3MjExPp6YCe2v
NmMwVMhJulHxpYHGppzmEfUMtFqz6St236ICqkRFC8tKRFg7F8g32bEhcgt0huGG
puNE6RfL/wYmcTPnc23eKrUpwj3YxKHIE47wnHmuA8d2V8afw9zPmPpy1iXHqxuW
3DwISwlCmNBnTZry7eZFu6PhAHCB7atjXtagM1ALBXnGy3PE3cbB3Pzk5mHG6uzB
dps0WXj2UsGNdh4V447nKZKXrz1Di8N4ELZuL+nkTlE59cKmChYVocqtuvQF2jmm
gmIAn0olmEfBVisAisrDzvS8gXMsFJBzJXtlU7EcVE0KDo5QPRoKJQeSnDRabiOw
e5jTbJIiBNuL9lMPsoaGyQdXG+9//QNSNHHxEzGtCIa2KngayheonS4auirPpbc6
9BcRyb0guVoOkJdqAUl3r20ID9BO0jaeqSc0RHEyT7orBb+GTqcUYtwebskJcOim
OTq0fyBQSw0F/aCu3Xac1EKk0R3j3hAV905YmSvldZL9/ysjb4wP6zNy904FVUJ+
awGwR/ZmpocJyxqoLUyw2uEgEANF+WdPqkdthVq+aXzD5rhrGyXkADW2/MkCvcML
RB5LJ4CHoIOZ/1yzN4BWdMZEAC955AuHj2qa46aVRhl7QUFXkT5VOipGuaeK/Uk7
UVHN0V5ZV+GrIwSjUbmckCB3xHiRgSVe2Iu3LzWLFv7b0jgEWyZCS6cquxFC/ipM
jMPnRSTdH+iGLmqtHxdG9pKiVfMzickHcE7jxbaQFfIzz0oAWk/w9hcUH4OSQSXB
vx11/p/Jk8uaJk3YhrU2+PUfsB+nADuwUmxRDHQuFtEGQRUI0uRHhKJsD6GtM5jx
Ct4lHjVPXUbC1bpedaNeLTDtdVUwLffW01W8bZbzIMQIu/swwO1eE0B1UEAgD9vJ
+NL8egthKszGYmgtgF6S8p9qRQu9FxfrNGJdG67X7HrYBejRl0zVbBq/dcugOomk
Hkli7ti5QLAkz0xWvtcAoYNpSWUnHYu0EIrl8Ik35wUkaTl6/vhsSMm6md81j8X7
1qX2Kqn1zQ5N57Bt8y+V7XGjTZ2FsRv+aqPFZIG2HCeQOQiTByTl/V6EAvghnYtE
RDh6kV/v/wFsGwJwESleK1NpfYtZoXXH7C+lsdBcLIi5tzCiyKEwEbpzPnoNeWCA
UpUXntpde4RnGxd/E1MXr/XUGW5vqO1b0fLFqQKBqfFebWOo1/fsNoqycZU3fpDx
zNDVvZQ4qMKGYTkgbLnLJMcWw3JVsjApkFbufKFHpRHSBUNFEfVjqhvPKI1YsAMe
L1r+2hpSJ7SKseRL8ZF15IH9ddH0hYQICkfaOhMNaoeoG1AuvA98C15smtLS5qbs
1A9cN9vaCgZTOQPstKDCY3cDE8mUMuKUI9E0IswAaa0dLiPARXJNkqulqM5rpd8Z
Tjbw6o8wpAvwBetbEjKyZ81ycChuVsHI0/q6XL6GTDNaCvV5XQmwEnne/ttdWreV
ohCFy9AbkzICBmmzxRzVGsxMwGyBbq5Zd+AzIJR2zAvxgmKfcBgdg35FmKMNNpDP
R8dOKVMQfpcET6B1stoIJq0pQ+3U/x3OskVaLktVL80iwM1a77sQc9/INs6E3hNV
RFjAqRVcxDLJ/SR7vTKABil2lvDHPwqpYoGSnakhhcjbWUVx7fp7qs4aKAXbA0Ob
P9mbTnPAup4sNJS4vS2WDDHu/1TLDuN8RpnoEs7sP5yppRJXat1EWRqwuIyqrQ2g
B7CFH48l+3vna8LriaIvLb31joIBRV3dJKNzuiFRpLUWDuOKgvveS2ZqB8sptFkd
UYF3O7Tn3pjIRL4s2G2eh0bI95YbkLKV7w/FRX4kM+dzoBae7N9JjeXNC//pUGZ/
Z29A7D8xSZMbBOhQ94SVFft63TZVzbX7NsL2v3yv00aIMp90epZpqUAPFpGYt4RH
s+iaUJhrne2XhQiW8m2indNSmO6fYdoC0cZQRYnMnS247mSpiNx06mKYT3caOn+E
pMfJKRHJ9VLqo8jLq2mjPevVbxAImgDSqUr+4exiNJ1X1UOJo6tJyUHkYY9fVGZY
btv7D2TXqhoLEAy6CTc72FMLLl+3Vx4lKTQvfgM+PCDYymgNLC92znCRfhCa/qIx
LLOeP2jrsVyhBpbVgZ2zAk7FtbS5/Gt61sNVoKU9URVlmPtdDaDg+jKx+zCeiI3I
6lY8jiAMh8qihKIlwxwKXjIFvkpXzPTDe+Z3cwZkJs9OfRBZ6q4/gp1Csd/e0LUr
qOhKXMtJ3OXRSq3hbpsPq0HT8dXHTy0+aq9+ayFmNYj9YBf1C1yNhLK5jL22Uvsv
IPtnLIcjQaXEMy7JCf/WvjKHwMQOAz5lb1kMy+0ItASn77YJ+O6pSugNjH2u5iXq
iK/shECyXfnvIk7lcGAKab+2yaZwNlB8jVDmeRQf9jGpqAGvW2ffO96fzT/ZcYv2
+udabopgtu+C/wPMu2tVrlO+BexHf7wwYp9zYL7O+RQqKNcHcc60sQF4bq4pych5
1TBprChRP2gjw7z+JP5VZXS9jbGGDovRJQtOZq0fTp52rUdU79CJAyp1jCUMOPB5
jL3BDyv6rZGB+3TUxUmnM/DGKN79NgcdcIqSD1t75YPloDuuvE/KQvrOih0CBTNj
NpNGJcjr1AS77EPWtoSHYHPtFwKZL34eH7SplfSkgz70Hs57RIZjC+LWl7J+lcAu
aWHz3qpw3n+1aNgi2qZ+d5nNbefImtofDAIw6yfVS88fXVz2k4gBfw1zywO33pX/
d+DvZEO03iIGkmvAsyi1geqMVM1kWOp0kM61msdt5XLP60mubL6feKAl25Jq8lTp
bsWNJqDn1Z56bHcOJgasp6s+Go+wYmcnwgqsLbFndR5EAPqXZs6ihw/NtuGewYLr
m7esiSOmiTQ5Du7UNkY3BXUK0HubZyGHilpW7LYqzve6aF8kFmcidMwmt9az/LmS
3xO7EXoWMYIDmPdx+KPGAO272Ofhm2rsqUPaKe3S9oyLre/RFCXMJhxpq2OQC2k0
JB0O+CzhN3H3gEQsN8rrhl7EesBi0eFUlLpyqV4G58VbS+M+m2Sg2KcHpTV1QqbI
A7P1nVxxghCezYGhSZXzqvccCFF27G6UHtdnejMNnrpUjW+fkH/wrVuXTXHjL2+o
87XZ2sjvEIPdFUb9rASpchc2ewcCIdcEKaaRl0dEoGtiZ+S9Ejw55MO65/aN5OMd
rdJqUPLjdgFocmW2UwbcqrXTR83qys7JQ78RuH4vkVdRwOqjk0ot4XtWmns5JU3t
A4Aw/QH7s/MtMTU5vrITwH66SCZ+KlbVGXGV9eVU04aKy00Rcpx8/dCfMIdmEEbc
YDYLDmB0qLrN5MoWURzIpdHwtRVR/NWgOOJtmeI7djznAlt2MAT/Ei1I08OYBC09
sEQG1AeUpFK1mG+AnfzAP4/B9RYrd/nikjcGuIoDxjsKAJfd4O8SVdRpxF7dfl3o
uwQiCAM4h+ThWD4fBq8U8+C1e1MobPHuIqkJtBgAlKqy0UyVxj+qBcViHyjXAIgl
EtoZv/cLLUldvhDjd0xDbX8Bak7FzGcbsHE+mF0ROPA20Eg4KvKldZOUFMHscRRx
FH9+Lr8NlqUKQqDAYWASMATtnIfdsO3r0ozpT0wTzzTqb1ojs5cFHqHMHEnIS2Et
iFWCGCkmzM6LU6vAA+ufM6df0Q0koHKNL6fvJ9hfeXfxPAg/TW+hugcyRYTRiD+1
uU3wDDtMMS0YtX1lkt59VsnugE65bVyZj1mgFRa2COon9F4juGNSdMzTUckU0cRx
qXzM6MKp9UJbtnPYP3Uz8NFDyS/u5/FX6yehpXujEfR7wrVyAQ+h4J/oLqSGpAYp
peu9bF1msDM6kInWgfTnAVOU7yBRYlP1VM81IWkhPuFvElQTA++4aapG9tsQifwE
JnQM1jxTts5o5+dDmUl6GEv/NfQkqsgMUKwl/bjANaonMLu1OoXcpR6lfFtwNgmB
Euua+DJC7sU+loUN53s9qGT4NI8+2SPtY0jOQFG6DlRAYgVrictXrKNpoq9U0vc5
SGJ+0eIyK59ttkm8CrPsVf+ZhLIS8HXK/VX9QSkOO9Ko1jLP3mgbT1x/Ff335fjW
dhl72KN03SBn9fCgZ6lWsaMUSJ7SBegL5ISgxNgnpnv2nUAMMddmRKZXoSL2hhnM
Z3n8G4Nl3glYAU4Uu/U8FzRskS5xDOxPTkUvDLypPy4lRBfXKge/RIVv0WyUfDPO
FgBenRV5MnhmcaMnzigf3E6F156tSN1N5Le1MyKshVLb2+V9LgKrE0yGa7iWWj9H
yruYTD7e8hLz7+F49nxUm3dXCesIhVYDLspybIXqM+WtNgLsGg2hsTN16fVHWGZu
JzXoSYDgmzzm2aZSyzYQwph1yD6wiKwtLSqxtblgEFYe28QmtbYQIrF11BKLuYHU
TkCA17ENKLT0+npexObsp8xbgWaBwfjAv1oyDtjzyaRq9rshsXvutcWFo2emcid9
jtT8SRM+cQJuaKvyN33tMO/QTicLRAWbZyaLbUtd0w5MnmcgZhxThFy/GgfqQjZc
ax/cnMN9OF2/gnHhJOLUUj4ynkdmIa8bxk6OJhl2ZI6Figj/Kl0KEG9Gl0lVsUB9
Z3zIToccKJPBCpooyRJsmQykjGYPxZR9bV/jkZ/lIDpL7K8HXGkRQaohgDPSJgPq
OvM8oXUyExI82QPIP/tKszlUCx6QgVG5vlUGzFNZienMACqHJMARbVaSkHDw+vAH
PhX4m8lLgSdVFsWZ4QDmGOeLMsanm057oiMRLlNhg2GCPtAdNDBy5K7ZE1ZuJCh6
rF4tM5AuLKqnx9Ftvsp+GvJKwVwC11D+Fc5oG7NHlpmRkT5DLas7aBko4jwUGkvd
d0GA0J4XbaRrXF9P/xIpxm/RWKVm2mDd1pFYJqww4J/+uNW/Xkim8OpFXsxGxutE
Jg4XhPWsP/D+GuLPknWk8InHankTT/SgLe475G7WzOA8m4wGLks6gnrXYx9NWuvu
6PJPLSAueZg1BFoiEetdx32Sd2HP96JeAGeaRhvGqAJMEsqZSfzPkwpnQoqGR8y4
Fh9AVMYWR4ZCJeOcTT9fhyfl/glbRllckxs/cgXTL5BdPGvpoE7Dt8CiTINjsfnH
scQ4O6+rZEIpUMjgmfooYoJhWLHlju/ug4H+dg9iJ7SZmOynCJs59gmZyM5ScTa4
kTkU21Bz+IwnwaBWRXOAQzYnXeUEl08ehWk4wla8NdtaLDlOrUxd2b6flR+jwh/k
bkddcyO4bbiTaJzymL6oKihapS9RLVvbjHhLGuHQS5IenzlAL1vWs13RtlDlFlwK
YzG/IrIVASJQc1SKN4KG78EY65MVi3bO4MzqJPoAglw7nsqczASJ/61PUwXKh5xZ
aHa00k8uuDYrAY06k9+d00elFcYsPElP3tATJNaq4Widljs9kyhYLqLkecsk7yBi
oQ/eCMGlsTiUuJrRSBs+fxbMUbxpCksjy7qPrT1Mal/rDw4QfceoYmPjZj7ff1Lm
5/OcG85u+J/P0RhT4PWS2WU/dAkz+NkhhqsMhN/WR3RzdVDnzT5LWn5E5g3Ywvml
ym844as1BeRBcbJPG0WFNzQ/oaYQY8xu3YB8+sHAh2B+n5QIokdlu7P72WwTr+md
rDJengaEN2IEZzoSRT3TT2zAMUPmV1hlUUuN7x/jZ/rEwXSxxnpntpyYoqNYQt63
7VzxEn4dBm3E5XLnvrwifqyl3RkU7dPh2dt0Wnb2wXeo/40Bw1jm56B8HqZpmJqh
DYh8jeYK1eME/ibgIA84yHQDzqOUBM81mXK6zXlHgA/iJ0+4m9RNVbZMcnRxy73i
NY5dWqFp+mdWBgQ+aeerICD7Ej05NDmp9+Tw5YLUqtOcRhgd070QFjAbVJ8TkZzX
0DAz3vzvdwyqLwV+WKgYVBdWmCkWl0VJTRtbK1IrZjqXJkCBm6F3BYvTe7hH70e9
9nXU2F3i9joG3DX82v4gQ7a6Jwchfxuo5OXRYlRjlb+V15824VA95CV/SXL/9SnK
Oce+eEe09y+aPXUwT1SF6APKBf+BFq8uNmJio3IOp1R8Ana69L8xBDKjCe8TWbwz
j4kEEMkvpqiv6yBwE1arxx23reSxtJ7Jc5+AZPO/TxbNXK0vYMGACjFJi+ictw0C
7HIp+KabgKsMCZA9xYGtUNvyK7TLs0L3hmAPGXqqJ8pwTVLl/56NZ0LfL6vbktry
n5481srR/whUAWmKwiqDnFbwg/ZSq7cPYWlvsjp7thtXQ4VSCsixoHpuG4lGPc6E
MQpUX03z6XUydWuuQIsI60RxdVKU2nvf72iBn3tIAFOa9bFKT0tlnxnssFKbweyi
yjjGn/KR9TZLFipbRzbDDeZwip4hhUYMf89bfoE3ulKeTceuSchWYpfquUJhPQXE
itcfa1yShgyF+HPsj9qRYMS/sjRESuJLPBjDRc8s0lC+06KGH3qT1vQwOnFg/Akb
M+mZl2xGZYXGzgMDTo3aNM32M+FvxOy/OWsNxAu3AVxPPMb0BYZLHYxkhCuJgevY
QMVrEjghF58rBJrQs6YsBSQ2+mABZsfHm7GhY+bkV/e5HYoUEoQwYbSUzBS/N729
LlT3pO/eMvGxzi1DYNqAaSZevikY+xBhJQVD6dG8fQLUuVsq6eWV1MPmVtjxhEvw
oq5t5M1WmqAvazhySIpa9oBkZD7noLwc/1yxa3UvRALzJm4UYb3oQPrpP67tFAqQ
y5H+FFRiS/UiIvl1RdZtVJNBfd/lMqPzLQjySz9cGl1C0mylNp55Quhv5UqeNXeQ
LSFkWXtxRqjpLo3N9bNDO5qG4NaJZvh98vgBXC4O4ErUP02ynChdAPeheq7+Qn3D
tB3gMnI3sROXCQk+aEQO9IxLvNukx8zBQYQisjwreqzERN7jWCU8/ykiZUuuRy+9
ft19i5CefE44ET8CQB0ctPoEYL/FpGxzkZ/0R6LfVxGNRNq66HEzT8DBddS43/gn
OdwWO0XY0ezi477PYXWf201jzES0oTIfwWT1ceLtraps7CYI2xngDXdz/8mSg/+m
S5j8Z6o1mIpPkNmBrDy/QZTihCK22DIJHIeVGCDxjwpp6AlQKXOxK06D/N8LWKH0
RGt2VvVoioGC/pPAmvpHbW9nq0T6K8e5lSDvBiA/vVjE1gF7U7/LIqEqgoSY8cEP
IbG8yRab0S9LuPL/QVjyACFsgFHHVUuVb5WzYk4sQvejh6VuliOBWjUeFQzMNInM
51jncErr/9MBjdffKNCTZJGJc+bC8nT0Io9YAN/OyAlSqA1RXSjCuI1YUJFyZUyZ
pyxiwlpTcRYB025zq0i44nAIDFmz+rQIL0o96kxssV978GEdpxdPkilIdSC2W03H
ABrYmATFdzNR2Q3iPPcoqOHnoM62INdeOxIylj/c1XvmOeKITgurdm02iQ1JfKze
ZW56arw3iz1XFzfhFU8DK2MUWD4Ae/MkLU/HdojtRqNe9Axa+W/XmGtHZ/PhsyZI
M2fusMXN3HM6nYaYKlB9WG37C/sXijw69ABJH2xEptcHSZ/7cx0XqcQQNYxQCX2a
4XAbR2jaNmQ3veblSELlFtu/qr0rrSM/DR3rrirynXRPa4cO2u436fSyiDLczVDe
4yPUjwWswsGFKABIL+bXnYtBcyR6hPzYyG3s0wdWYzYGBC46ZIThPQFSiNc4IXHP
ivqN3wXrQa9n8IcBRpixTxRor5xsTABBNHV2vmVk8DvGN/sws7lGOmQjJ8LqAW8t
hFwkZvFleJZ2LftWW+eUqcHZodLhwAk54H8M40iZMvBLF24fvYj5Ae88SCSvDYa8
R5LjOwG9KhS8KKV8H+KDfVdf+Ci9VTgoN/l2o1O5qdCL8YxdAOD4tmVu/BUl0XS+
5ClonStuuU6BZLKLXISHoxqfQyTTLwQx2vpZDJ8AC/6TMSsjw2jM8gtt6m93Wcjr
ToMBTLYcMLWBCkKAYcND+Jt5OvdhiHgXBxWsZg7s5bKT7QBXwGMCysK4wp4l5rAj
pvfZFquazge/ANOB83Z0lkCNZbtIxxlZeHkLUitcg2Vt03bZSJJs1h2rOWdzVNBB
EQEu7h3prA8VrEOIU5qXB4/Sc4a2FltNmMzpS/LcCGT6rb3Og+wAHc5qye1n5vnu
UVNwMKppFqIkyPvGLHylwkqbcbdc6Sdh2qZ8AnCBK2nyffSsqsKNH9UWY+1GGxew
Q7+/5etY7g4wjiz+u3P4YQ8h5bpWcfwIcOuEqM78t+5g9Fgwr2M4VUcJEy1Wqf8B
lT0/nK9adpY5okwNGaSYgZbr21zcwzkb5MR6ultt5bvMClIRNPSRRcYbrVodRyGb
cnjVb0ZWMl/Raqm8UmVpKE67pmvpunlB4TLKr3uZyoHwJxQDiCUFZ/mw/0pJVA7I
EUbnprQV0ecZ0zFo93sDYe623PfOONukUERZoJ7WIIU9/Ep52yy6vdrezjiUOpTi
W5V1wLjGGWWRi66UTQugcRM/YNS8gtdmrpBNDBYS5eqJr0PVVVcEiEygZgioniUE
e47BoIgBGGVeovWNjlE4cnP+GcXsUKDW/hDF3bE+huijUcedVI5uY/M3ZNI2Bhx5
9IjsEdQWdV2kVg/vYtfInpF2nNXQzQ3GSttWoCVSA+pe5GzN4nXkWl/Ws1q/mEBB
aXWyCDPbPimbIUOByBs44Oh5g0waH7Eil1J/tkETE9VpbZkonIeITy061WxL0nKW
+T3EgpksDqBsf5HRpVF7ei5gBss64MlO79vvaAVWVLLE8B711etfHfy71hGvFqr7
cZOzsvREBZKlluhczy4rn3SF3FGTAZ/ogdZEG4XaL9xKhQ7EQ9/lnUCMKVgvkO01
VoeeeyMq+aXCxGtZbF5lICRgZLGbYWgSp2wdhkIarJIRJk2PEfOrBiLrOxXNgJTg
94qExaov59GvB1XM8yf4bBLPK7ZvOpApCM7RH4n2De/DduUgA2icrZWo2QnHE2Tg
sTqpsq0Qm6i36UkxwJcsT7pyXZV40IXd8Qev/4KQ09J9sYsSRauBsC9v95TLElj4
LAd9Fa9NSB4uBbACISizVt5Fi4ZdxYDpFnCNxl7EBczsjBCb05AR5iLEVtiwECna
bccJybvwTdUbrzoincHNTwRpZ3rmWXOjz/WYtfndHewb5Ys8iK2JbUFqM5KCuy1e
mP0tGJpjXjazMkT84dalE+GRAx1Orze0ilOVYOkTFIJ0Ed3g2/s6qOyjJr6TncEC
WrVDZP/zc57VVuAAUI4zKmX0a1jkObBqzHoaDsevOnz1rW+Wz487ZRPy/Db/OK/8
xLbf/IBdkSrli6zhIVDzfh0qDtNbDpS8drok2ZkSyoyT9RvAjsqlKLqBN+uKyudE
2hxhSmRRFJimj3sEUtb8h0MFtufqZFEXZBljkfoymySYIzNC1vPKQKOHs5E2zJH9
UevSP8H5zV3q85N1ruL2cDGcZavnrz/q3XOaNKQeD2x837+F3a+6M4i8W84T3f6J
E7ZGYeih3oIXkkhRhmx7rzIWGlP4OtL9jXnHzfSXp19x5KR6rrRSNFZF/vHHChGf
/9KAxd8xTWfSxO4mkvGmvtl5P7wiqSJrmQcOHu7L2NAtokQ9SMlYKz2JCz0PDI8v
vwxs4FLsgCea/19ynQVsURboX5Wm7typdB5QEPoNLDBX8Uh7oaVinFfVfr2h0Q9O
diBBqTrl8U9M6l4D0YjYm3R64JK11eYPWpdhyZFp52lMu8SSDu8MqtWfB+LTg3fR
S3YiVOZ/grJmXusg3EqTvQ19DQJqg60jG6h0bYvu0ZI09N52E+tNpVTRw4gZVEmc
jJsLubcK0Na1vtdXBslaja1oqmUZuUR8/p3nhfRZgWLckY6w0axJZJZzndmL65Ap
vGarmW3Rej66uhhL2c32MqfW47CpRdXtZ2mFThes2mKLyMNvmYO7KKLKuaMrhVEj
e805Ixv6wmiA0+sflHq2hOXyVaQtyxOA3+E5h45DIOmd5xFKCTBkEQyRPBsPQnBs
iJfDLFuTDuLdRwJOcts9ht/1vtiI+n5aCUuG7GDSK5ynqx7F/XAQTNYSpnApMOOH
rJ8eGVqJH/09jEncw8eVNko4UqgEysAPMzR7w4UIOY/9GIKudpEK+KAFFcf1tYQP
WxUIeJqqNdzpc8PgjAiPXArWLiXRHNXV3MTsGzG/d3Tv44Qk5J+27JBdIJ7I8J3i
1jhNshdSC894HT2qwoz7ag==
`protect END_PROTECTED
