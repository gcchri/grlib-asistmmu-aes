`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sOE34y/hk19S0V2sfzSWptPhxcnDpKsjNQw48YHbDfpEHeChY5hZZILrCqjtYfKj
A4uxzawJohS3W50wWZE3HztE8ty0DTN3Zz46LG7d4u+yM5Mz/CBKGvVqR3io5NE6
Bi+l4zP0PzKdtDDt+yZmxDKg6cAMBlEUZB5mqkevJBqLLkV+i3bye+7rKb6nJ5nN
UQgyLNygdZdUad3bgmISm2O5jR37d6wIIe8m/+0Cz5NJZeyzJ+Xmj7lV1h2aY5Q5
`protect END_PROTECTED
