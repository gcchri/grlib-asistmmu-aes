`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3lQ5QS9Y/lIqn2kr1dVZoBN9ia5fdVsJc1RKTRvZ5+PV2NVryQHgLzQD+Q3Cst/L
/YuYhPBqxIC7/oKvABn/iok6sqdKE1OLhan8Wl3vSf+G1+jhbb3xuPlrK5N95E5a
wG8nFb+hUAAjNZFBIg1zEwfcc6to/7J/HV3IFCTqsNRB/8KIPpatR99jxnobdkDW
D3DwBd9wEF5Xm+LUa2wftwqNOtQ6Yi0m2Rfzhlw9dKhL/haTZVftpL119ybVkh8/
s0+u+o4PmEyRLzE+uVLv2xSaAR/Do7QQFwgxzLtRH6M=
`protect END_PROTECTED
