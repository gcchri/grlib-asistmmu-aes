`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pulF2jpg4Fn3Mvqmtf2IDPCGJQVmXfr/Hq7jKNGovbOpoiy6t6BMrqT7qnQRjwOG
Ybp73idCa+85zwmsw459APHJ5KDft8VUzL6HxucRfZBPNrLQctxlR3iePji0QaXV
7w6i05NjvL/Fkk3RJZzibvjHnCrvU65ohv5Tb0gv8aKHUQnbg7f/VxsZWG9i4pZ/
UKSe/aKzdRn2fsSTVrp9crDVtdvM3UJkywBTUi3JhlrKbsRc8xFX+IhmE4IuZIe3
bcNtXUWuNsfEQmsIPoO21uNk7+bT/S8bzvJjpCdhtBgYCREa1QECBeJGS++yvZQJ
Xnkd0MVOZP+I9H6c4+BPwVWszmkRlrUXqVWUWJJCic6zZh1uKrWnAVgiuSobHk/3
`protect END_PROTECTED
