`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Aj9SMyI9uaTHe6Bo3xrBEcHvdvNzOH3XN3cXwfH5Pg7kRFXFIjD4/a9TGwRxGR0
mK8seo0W3ZTosaUvjNfszLeVn3SA55r37wyAcjXQx5+jmWBVTZ/pbWiW7w87M8ki
glylPi16oLxP6O6j7OjagCKFbZFm0WF45yFOGHdfucRSi+0i4KkLzurBPJVKdsWs
Og+xtwtu1sGh83jajFxdusG1muoT8Csahy7L6KUj8QswVyoGTLYrLuOb1MGtMmSk
9pFJNVG5aLJviVlipasJ5A==
`protect END_PROTECTED
