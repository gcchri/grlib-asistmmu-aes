`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6GQXkRRadZiKM0rEv7ULsft7a5qu0PjlfGSsyHr1jqksV/v1bL6tGqaM7GvOzJlV
vA7LACWH1hZnxnBIKMLJejpVlBrQ0TvdmaJE5U9phQxHuWn3nkMgHxGhN5eD4iyd
0Hkx2LQP0CYK/3cPpURt57v/0jf90qm9pXPU85iwYhU92HQQAU5s/t7ZqDQK+kia
N4IMOezwTwBDujXMWlvWwc7utbR+yNI/e62THNf4dziUyHEGJ0QOvkVp3Bj0aJxy
8kpvRWsZxaKzW5ge6W08wpBbjkHH48fQQcHW1zovK5jtj1PXaT0eGtzL0m/V4clP
Hu2pEOzjozvntR1XN9vpbZmkSgirgb5POeKUvJPRIujKrBtpmo4gASQlwmH4GBUq
`protect END_PROTECTED
