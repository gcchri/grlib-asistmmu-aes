`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vFb4XBtccQMbSe3TSgW1vASQhJ4TMJC5dtwk1LXu1U7Y3g+fYGlQLCocPv76k8Jw
A1XLKCWBbj9B1L12IbwAsNhfUr2/6UXufhQAkRR1dlm1UhSKK+JDl0B4Ooi3Yysx
eKze8I8fQeDgn9CQR3iUTWCTyIbxSp5hEqmkAi7TbVWTbOemXL6hyYHebmniR2LQ
GUOvuzAAtdD/iohK2S6soj+AusuiL3w/MdWtZFUpFd48b8SnWOOjNCiiWB32klKO
fpeMDbAkOag9ewk0SOs6XTv+Wf9OHakUQY3VEUCUH9XV4Xa+aOgodE/DgoOkjQY2
NSr9Z4SkCTsMzBM3aK/TNrd/6PCto3m6lLZtZC5tR8M0tu1I1Yq+HsCeBK7kukp4
43a9MKv0tTeloTe4bgfu0cpZlpwYDPFSM9FAL5Lu0riMpa74CeZzYaKW9CtbNo0D
y2kJNiSXmBtYp6eqmfgop4WLi/mZuZkqLXGqYpPHsA5TIfMKiq0DM6oz6GntPlMK
`protect END_PROTECTED
