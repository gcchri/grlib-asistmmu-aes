`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DA+XvkfDJt+ktRiQ8TMWAy5EEASWQ4Fnl+Q4UV6Yf43Pop4q6rvSSr6kS1iJbjMv
H4km5h6SguCHAB97H0rhIJ7YsDyqPMR72UWYsmtzw8J6kUJhdNJYqaKdpW0F9CT/
nIhEzuabTvblRXE6+ottsVi3Fso/JAQuDdKlhtn42I+jU2QTYQ5NTxhHqhykCWk0
YbSJLtVUPIBGy6M5bTsI4SCKEOC2K7h0XfGCbA4Wceh3eX4gNtliUsRkPW+kRes7
8WgqUezE8st6FU6gu843V22JJZtcQ588Pnbu3fczTpwIfSKBocHcHQICU5+xTMTH
Ajmv2SgVtynd6q5EDN7qdRjyE2gP9HYYvQZKurZrx5hOOmM3ClvXMVsl88RuB25Q
U5YRd5pTx82CI2epbykSdeuW+ikLGRp/bzHgzMGiuLhnQWcqppM8M0kUUF4KkwKA
5HlhZp/wjEF2u4V/YZjmdCOHo7YLMluz8GHFOWnp9Lu/DJPyrm2SJNQAzLoKbXAy
`protect END_PROTECTED
