`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nb9441tyuR0H8B5NsZ7BxcPvQwT+Odi5N33WlBTlUzoeh6Qn1veqeiQPe3kgnbBd
d9dMl4wWMT+vRNCeJzuWb23WYhllEjuGKkX0WfCwB4LjnIfHXokEKGxOh3SIz/ZB
hFOYq6RnF+/7PFoRq/zcs2DC0vto6fNruUxfasLpJUTeiS7C3MAWHsicqrB0VQ4/
R8ozJWA9uoI+4wKL4EiSM/2DfWpoT9dHqnE3FV1Yb9ms1JTohD25g34ISo45pc5b
az+htrDHzjge6DS7rZg/vmSRjmFtmbLSYUJWOEAwiJiK7Uhco2fC9CIPbR9ssmkJ
ojojBO73k3z7Mm87nBKCCY7rhLgZWREvlD62qu4eNaUCy5yWBLUN2RHjASCvncCM
wxP+DNLCTd8UnAJz6JJP83i1BL5FcrVCvE016q5TJAUwkFXMSm1jHofwYgyQGtoX
9h+OcHvHMrKMDi+wgsB1QSj4UiAJ4e3GFldY1NA6mCoz9gN446Ynu3yhhdgtNAnK
Jj8NoljRCibJaMEU1+SpvTUlRFDeRnK50q5pQs9HxRrFz/23QLp70Ff9w4vTsy3d
smvmszj9E/el4gt0mlVTU0omyRkqQWE67UFlXypJwJLB0rYjyVRhJE9sSXfme4af
LexRl8gUvIKm9myptx6yrmJGlPAXtSQWUmFr1E0uO+I3Ot7gYGp54WBZWju2b0QU
zl2b/ib5CMyG5jsoRu7xYrym1Q87OkGlD64sPLsbrdDWmAblDyiIKsU+teHniSH2
JaCiBO2CQVlhCbhhmzGBFozuxgwcR/L96zpUEthUMnAEifMMNumfTfUN4V/89VDE
CLAkuRTt6axvJMXiH7mpR3payDU2fYhe9lCGkyEAF6Jz3yvJfSkuSaxR8KGZn/hR
FqNrDiwtSTaG0HWAc295Vha83mJLtLeQ0gb0ppyKCN8tjcd4f28dTaTBse//wARS
sdDcH7hkmnRZLAQeOMC4XeOKD3R0bMqtXsuY1BP+zgezqkNe9kxWQMHdMV0QhmVR
FJ1IxFhrw21PfvTKK7EtKPYLwUYeql3VHBvtzlhUteyXBJ9e0ssmUEQsXChcWjgD
C5K0fl8LbRIjb4Nw1x4rgq4lju8HVn+Y5FiKDjngF6scYyNQR2/kMfQAgss43smA
zbEYNoaXRzNM/jdqBeilFpCXvADIhEcMezjmD6eBhigLWpTvPeDE85sOQrbDEGki
ZJ6DYw9XA52baeUB/TNYmK0N9n3PATC1Tql/oaqPYBpz540766qocA6/XEbyLEaK
M0GN9XIXDOkn2COVBvbMaY/4pDXPVVU58qXTWSYSp0lDaUCXUFndvAGLmr3hNCf5
0JM2fW/Pbwkv8a4XQlqxyGbNrIWAoLXiQvSzpIEX0HjSyhhlyZcncjpIAmeR/UCi
s84ZYv5gJQEePA4kIb+DZL1AbM2JrdfMgjg0iz4TdOoI6SRs/jIDkPQZVHfe7cUI
XCtIygSygCUKEZobO/uUhxRu1Lf9xjrH3D4o460qA7q2sutc9Y1Nxgbhz0AcG6JK
Jl9oHru4QMR/bmhadBN+/QPuBKwYrtOIU+PhCpsxdB9srCAHiHJ00slTR+uaS+8w
aeIWA4UWluNJMggm+6Zp7cT6gbsM24nt0Ri9q6xit05M3lOvaJhLODv+U7SoqGMp
x6KpPE8U+ymLtcXwUhn4LjOhNUy/i21ZvwrF+2VZkFC0ceWXFylSuc9YjTCU8ojK
`protect END_PROTECTED
