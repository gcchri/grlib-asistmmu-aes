`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uOQyhbMf7eHts0OKjxK0NSaLoku1OLpZomVE61ogFc17tqXG8+kl+BJt0BygdMEP
AfeH2mbns9zXaxSx2bFCbSo7ZmhCMrHF55titLWvxom4KcdFYTN6OmPtsERDU7Ex
z7PFo2xoZ4QYeQvealg5oBxz1UCkl1oe5wl+dkvA4Da5hcWHjTdnAJLLhxmv7jGW
OZ8FPRXyaNI0YB5GYMJ/kifm8ghdV32pjpTA4B1YEfs31LbO1rWW5xU5ljTaGprF
mjP9UxkeA1aq8C2mFQv56ibLV+sadAilod3VXhRuXa25FV76MNYZA93pYgxavlty
ZFGJHEyJEbEXIZ87fqs1FnQgQwPBDF1e8OL+7ioVucEOMcn8DZOa8OE99B/T9C/k
6t1eHexRwgfbLj10CuHVU9t+bTPL/KFBmUsTwyQI+CBVdrQ9BVlpe4YBq0xLwBVN
YK8mmFpPdBZIEGBdWb2YD7ceDEuTIGZj1NiXVGwcQEutnLRKn0c+utZpizV9tP4P
DcsiyK8ofi1ErZ9ShOLQZD2W4na3tUqS35ScduPzKB43ULWVg3cYXsLeauNVj/MQ
`protect END_PROTECTED
