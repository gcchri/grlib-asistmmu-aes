`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
On7BrQBwXAjERc5gP2pJAoicdXhW5jNRBp1rMBK+AOSw2CZnB7TgnZr6zynduonE
2sNC6HejVRAT1pjmlXiTepjovMMIU+Odx3MEV14ceewGV7OLkE7Fu6O13QbKPUcB
wYjknCDLBvJaSspl/HDzSetdLJKui0G7C9p3xcw+D0ouegCeS/s3I9dx8X+LYHI+
HPNYLTxB14hB37xRml/G1GcCsm3BZ3gkzfexgGWavm2dfRfBJm+Cm2dcc9bXksd5
Gs19N9a4UQ5EFUEnTB2DW2fdtWHJZNxY8/APPBwEHcXlOmJ3rc/5li7jFEZCwqri
cJl3Oy2atfZbADLJSa+YbMku2iTl2/Nm7PpQAtL1KrxmuxUNwRjeXMUAJLTyfk7J
/nV6Nkt5IozZkGNTKgolU9XYrjU9tDiU4S4RLkXnwdKAEPfkoSK6sOwTJm4F58cG
+dnTRKXzAuIdCpgbqGFvDUJyUs3y2Duo12tK8k7TmI0qAPn2s721t4sZkjON+Eix
JgM5P3VVxwHbhQWb4PfXnMu33WyEuCEPEJ/3LRZyg+sX4EVkPqm0yI/tTuf7X6Cr
gCR1W3Sv/MggWJ6LQ70GEJycFFVv3JNPQyoTRr4/OjrKoxcwLg0TDdfDGOlaaXYr
cahcyPDdJqxfC6glKALaZ/tGZ+HdoJ7ACti03zvYw5o1N7A5lCYc39VLVsGU6DbP
p/T7HcsrtoqqVKUP3xjtnhbQzNcKj9cUME/8fAHNlhk/C6oCgQTPiftaHyyIyfc8
f3bpaj2t1yYlK9jzrKMTgrfm0o+UqN5rdldczlQIZAklEB4/JEWqk0ied/4yKOGQ
kexWltxDQrRc0aaRxl17MEW7JSQLP5w8KYlDzl0mrIAdYqUdQ+qSPzVfC2GH2ch5
uYV4zfBT6yqaHelnrbEep6qeag41CrFbx+TivY6p67bg1CZtGTPI+lbpBV/IEBzF
+W4C5/5bN6r/E67yfYqd5NXnEJoKnFWvOHzmh+yhzzC9YXLkcDhuyZY3jgIqVB1M
`protect END_PROTECTED
