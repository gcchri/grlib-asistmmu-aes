`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LgIl0N8l6UZzOMeKcBgi0HPAn/3K6PlcB7nv43SEwlrqdF5N6VBTLCglzGEhIqvs
VDp/ZrqM9fFR3iYTvAzKw9ptQK+luxB+DeQLWbkE7LRuoEGcVfSTd6abldtAj+Vb
opL8uMF3Bn0CnTx5OWc3jeWCLn7elCG0ll0t4eY+xocyO4XIDljrepp0XonKH97J
IIguZ0wReD1LKwinQOYYEYsgxfwjXshjwQDYqllTDN0fg5Xzbyr63SKYwBx1AT9m
ZlAkFp4Nqmq6AxWc5FXkfjefUWJbQ3QScY42zqnSQuUyUaaQlCqtcIMvtDrF3ZFy
BmtGmxHt7r8A9HSg3s0b5p1z8jj05RhzpDa30Cigr/kt1RAXjX0aB5Y9Kn3jxrCG
`protect END_PROTECTED
