`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e31rCvX3n+59k1BPpoB606UYfHKix7JD91Q3mPOmZqo4nYoWTmMdaMraDbayyrLD
gia5WzD90orEM5Yle7MJm8PGOxVS1w2Dx9cfRbr9haaxOInoBO3ETjXylg9fs0j+
BKOdrVmXw5yXpi695L90828OXgFeAZ5GeDauCV6Mdl4UU6aIC0I3X29zUG2463F2
5ERUVY32YeVk0lFvydjnmUeCpl9xZgVPSAcklLsZ7336/ZOlH520HtWg//0i4Obo
4VjSfAlzdEjKW0kvvjwnp3AXyYxHWusSYv4KCMql4EkG5dedfs8je8ErbAek10PA
wVXddUesaQG6z6OaOMXo9otPuwY4D2iePopiTj2l01sBPMQ22B7m43h3kazDvA6i
50jCDqok08xDYIkeHm/ueXq6RgBGFplbKccZWrM7k2yg4eOce0Nw//fCxjXUKmy/
QTTStoitl7wnUfhNJrkgsmruzRrUSNhm68N3swfbZI2ttlZcJu/r8p3aVqXxxrHQ
IKJc1eEdPUw26GksMUfhdkOkmtW5Za4Mdw4j7bES8ub5L3AvKS+rJGgRl/vXBVIA
qMEVavQ5KkFgWKCyagtMj7U2w8jHGZLEQ2WeyWyhVzv8hqLxObotwHKL1HZ5nFIk
zo3rR7tuj+Titlcs57VvJaGBCG+MOkKOuus+xDNq/TmsHeDiElMVu9daVi7Skr/Z
`protect END_PROTECTED
