`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fTcBpmRgnKDtcgWQbCufUUeVcilaUOoWr13rR6S4o2rv27+pgPbEHNnVxT0ZT9Oy
eH2KYHXaZt+zAb1hdkrAq6goFHbPOGf48mIrNf9a3qPHifnxbR7qBGzSzqI9QWZE
KT3Z5vJ+RVkGi58Pgpeft2U45rZIb2jvg8xEW6lMXjz4pLP5aC0jRC/C7+PBknW1
fSiB+TEiQpEGjI765Saa4vUeHOFi2FrTf6vgsQfMMiRsqzqe1glawS0kjCL7yKS0
soAnZVcPkMTFQOXDqqYbhslj4Wh9PEtS3LOijqzXV83xy+O+7Dwc/oirqhvOaMPf
5zMRQqEzN4wXEe/BDRR6sULbSKmfnZDKNi+9CH0Ci2vaOF+dTy++d1zfv7zH3cl4
tNHp1aynr8moRd/GCapfscM1/QzlqtBOyxVIuqDO9c0WQrQOHyxge2VICtowX4IQ
2Pqn7GIuKPGdXSHcAUOFy0ovcXzKTcCAMkc24GwPzvFwW1GK++SfrLcPGj6tFwsv
f9n3QQed6XUfz+o6Bk2hrVTJgQVqdMvtJNqbSajfWqMsPOmOqPOhlibIjqp7lpCn
fZfq4N293d7FTMwcXLDEhNb+YTNfEdgYHN2dF/QM9i++yRNvHi78iHr05GQLGVJc
jN9vyUkdxPs0ZdHjw0DOfY4X43hhCPkvTyNIFAYE/mOLaFz492MZQF2Zx/rv7sCt
cyWuAVuAumGa1wEce5FOESI9ETjoFksyXsPLMyQynio6uyuJLtq+7do/WpeDhjcv
gAI/cl1eszev1Uw2vZDzIHSDuVcn+OH93bomhm3ulPxqaGavdyxBqTbAdvFhVo8Z
8N3saHIMH0Ow1ZLf8v9kbtuJnAJ8vcjxdCKLQEmCBtAn6gZo20w5MdCH9oo55SBV
20nQth/DBWx5ILQkBYd8rButTNfUP7uB64r7mqmuYPQ3zruXUcnzIXR8F/I9KPn7
ZSku7s7m7EDKp9S3qZxeSUioRcz7lOuCTbqB2vYv7gCgzdRkE9tWt/XDlwKfcFN3
/P8hu2HALNdMlT86OrrIgYXWfN6RMkPWtUjU4J9Q9wzTJyKGTMZbF47k92zj3OTl
m9IzmMDnTYf/JrqBuGRqAkyEh2igVKZ5cwF0rNocw0zuq4qzRFMyasmKIYVJog/J
JvDknpBqpCfvxe6Ga5yMUIxu2JT2BUWdvLZ0pZygLvS8dzZYyOyUCO/AetZ8zzQ1
JmnqqutxuPIgaJlqHeQUH1Trt4+vmK0KcXSFifVulJvnJ0Sfg+wXYUcWy0YlRbsB
Ls/cgzA63K8GJ9jmQVP8Dg5g6rlFXddV29staoXQSwsm+rcmjticZmnkoM+ndjKG
`protect END_PROTECTED
