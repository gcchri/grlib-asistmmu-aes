`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iYsrOBoucbdAUgKGcE0RvR/LnkriQIIqI7e1b2gfqe8NO5FPASL2g8x4S7cXKyeA
Nk/okSvDMyB4T6qTSyW9b4O0gTVoIOutu8k4vdivKiQNGcAGv4b+pXmRolyo6Rtt
sNpMOJGiMFFvRML9LBOggEvRZwbMApADD+q7r+c02VnrMYUa94WM2GBniTUjWam2
TzFCYVhDljtnT5ah1CiI0SSjzIhZfy65CqD+VmbcHV6mSwhYmV4t7ddKvWMMUP9T
dnM7OpKvn2kjGwbe0CtM/ztu7YqOaRceCn3XLw0LERT8KnY5apJ3EosP5iyTvY6R
dDD/hheGO/iACYo/ZWLWmPOVbP0h5TsTHjGs6Bck+ihX56YTkY7NJK56f3DwiMPE
JGQYSpeQk5/2VXlavwiUbLsFv5JDapgbadGcZXccK3bEsFuWxHBCQuaQhYLBP/Ls
8ErFVCZUskKJza/uHmqEr3ShG+0LpDiEZy81JwW+19POxuqeV8zhPeNr9kiljTYZ
qH9+B0tGEgbNC1Rp/Us+AIs5T65P3puRht/CtcUAVZ4X2zPQHTxmBTMOsdMl9Nhi
6pqAux/lhBGxNN7tkep8Mg==
`protect END_PROTECTED
