`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NXJUfFsNTJrK6l1Y35LjjOVqlo76jLpyh7ofts0EcikhcWNPAI43JRY7/DvxYwyp
472uPaIk7w7LIwwyev5CJQf56JHEYLEMMXR9VX86yzZRzdmSlNEKPj3cBnE6/dYj
o4AFRl+Lwdsva4ffhMxpBP3zlF2ruZ216D6OoodFiPJchArtlUXqFvSiQeSP7LlS
Uo+DyI6MQIg3usLobVwwuuRn5gt2LUUP9z07PTGn/ZWsFYDkglEK7mZrnLONFfEN
AQpK5+8EgU4+BOF+89Czj9I0VPfpEvjJ4j3mBhvSkIUqh8rSuGHAntQmk8+lKNNI
H1u8QXMzehAvWkBKH88gaKu0gsl618edf2EVqBIQwnzfmE3Iy9A4nr5/ns0kqjTK
JNMtnvwIbvA1dzF0Q+vhOJp19xmrJl49mJsasVS+lR1sQ/6RNEWtAp6xBDPhecRF
9d74cNOGW5xJu9HkcS2b0E3olOHpTdy0+Qq9L/WIeZmNador7VKiL/ZPMxXO4C3D
2esG96xqa6EiO8ZnV2d+7q4KoT2rGqzll9HrRMQZYCf30i05v6l3EXkdrq+6riGj
Hp8WIrNM9PD7PCPPEHfVI39p8ifp+/c4V6dj9tTA7aSILi50C0cfHBy0nPhjXiVq
deZlrrNIREkrtq5dLmjcYU62zfofiv6NMb2mKTrpQouxSbeFSAyHN53Eo3DNyKrM
4tsBqMvmKTCt0Bgmwia/Cjv4kGObso2aePPhP0LUP8qjGYtWr05FQogrXTIA3uH4
dQMw3imudDyNMxXh/GlaS/oQNCDqLWbh2As9Cg156noAFF2+5Co8/4sCZY0t59qt
JIfCmjF4Pwm8DZUiOBPqMQk52hwV2AqeT4wMic5/R9+SHY1cwrH0eXt2XI5crCIi
pwP+pbzjfQM4wFH6y4+68upEIJWTTCv/1fE8EzaqF2UKo3GEipXcAsr1TXKfPGU7
BqDy6U/yuqXj1axPuaPb0xbVgaMBAY62KT++/yOLKnl1w+uNt+KoXjsMcLWxjAPv
br7cjytEejz4MGldu4hW/apuk3X3MzhKwezyXK2EslFS2sjIPGEJ7S5fUVmO6J2t
2m4c6AqfA7wrWbWD/fR6NholuPE124KcOtgt+z43Dhp3wPyE1HINErX1ujK/NTrU
Ref4mALknpXGLvS36a8xjXYodN2JyL5NYesaJ00sWGrhFB+LU+q8H11TIuLcnxwc
d7DFkosIXytUQa9rL0Re8kooi8a+eTGTqxl/62otQVXn5DyS808vzjRCNISU4xuh
0IPsWIU/YljbTuMGe9s1MvBjKDYMknOj2FA//bic2xO3ieKpqUkRycLXSbATvpLi
nKrAVJD7XsrwDgfzdHL0FNaHEwXuJr7PQtt1L6HRjF9Mg/MYF5Vcq75N6Wd6RHsX
qVF4EPly5qU6XpdF1eoFKyT+dHdVHCce3NnCivvaGnxAewCAbY/tfJs4Mzw1UMyb
AI8BAcbtw6RgvKbwMWQ7bJJ5uiNVvUlna15Tvrg2fc6zExIS6iQV6rqkM/nvrN13
FCy+C6wO+pRE5FMWTzvXT+mxLBWALPOLsb+f9l4dv8H0CqdDhDASBDesA8sujcgB
qDjf5vaZ+mU8cLv2j65UtsmjksowokFwdgNfrck3TknKMCCWXOpgYQ2l6o9t+fmd
NHhVaceZmnYTrPNZZYOWZJZlTRag3EYGW+Hw7CrUAuAd+P7WPZmr20+XyI/0Ai2u
761T70QwxEHXEcs3e0eyqmYWhRXjbuNdpBy0Kn1eOqEwmTBOdZZatM7967n1zSOK
x7DM2nXSU/O8oNy7bdNgBFXS82WE5347HXdJkRgaMBUfQbt8O+08gYQsnmx5+mQ5
NnX9guCK4FtMdLreBt5Qyl49PHq1VPGS/gZjUQBmuylBPiRmZUyyUng0eyffYEEs
Wl6CF0TcufjjyAXl/P6/AlknsmHkO+XI+KkpoeNLha6/nz7gzRXJK44NriyY3mBJ
ovBI/KDZATRmQZg1uUSwO9MG6iD4eswe9bEVQPGKXC4nxGoUkh+GELLx8nek5kJG
n9m6kajmQOJ8vy3W+NQKpzzC6+AZaFBbFva0vr3abqK7qORMn7iqfMV6wsf4leFY
GoMQje2DvPIs6WbMaCZjwny/o67KK3XDWdqBx5SOoZ9EQ7IykJGoeFVDau/l+oaB
vmisS+AXH6IQ1RIOPI9IBBxUHNmtSFnkGbhZ4b6bkVCCxgBKom6BaQWtOR4kq1Ia
+QVhcWhDB5DhYzv6N5nFdqhvZlCcqQw5oJrQU0yp79aj6bKXUN25mWcKJe8skjac
nVl7yE608NM+o+/hWH6yV+Gn/8s04qYRsAzpm/DwnkXw/Y7WzofpAxyARxxnaRsS
mZ0ZaFjfbXts39J802XZ/P/sLXu0wCd630n35Rvqv04SFGNtlifRJ9sIFy2E3gnY
0H79OFy9+U074S4M6iFy9VWgRSCxxZ+OjymehjYWrRS7b3N/qn9W2ZVDMhSb7nQb
ZWYREvD86lX0/cmJzQ1n/+/qLRJ2cz/sQJ/CwESHhfN/esDoMDUtLrmmJ+yJP2eh
Vs8io8wlXk6No0dgCVf8n1ix8hvZk9OSRwXTLIYapMrP1R/0af/grGBgu9WL9sRF
Q/NRRjxcepitk8uHmWbeZi6SvnCMzTD+gYC+lwCdFBYHoBWXlaHrlleTRRPZhtEz
+uY/3HT25YAJmNofj1J3G2MMdXB9BEUSuUojKAyCpti6NMCxuZlE0DIzW0KTru/E
axFT0D2jNt08znJGvkhbhA6fNJnCqDtX81naaDkCYNBXFexKa9eTeQmiF/0tdptA
3ZfBZ8QkHF8jdBeFzTXq/9bB4WEZdyJ7CCkE2ytdZjqzdeaZLrmuIXEKZ4BKWu01
K5eHdn8FvC7AeiwKVjFlBDB4bv7s1Y5XKFuazgnWqHyAXLUes/j1p6dofni4p+1/
uLK65+laOWLMMMz/5vOiE6m5XAsXxoFncSaLTDMEGoNgyGINkgm5Cj/wMs7wRPq6
mlWi/FLHBrq3Sy2grZJ8f5s8Z8pC3JqANMu+nt1R5NLFBpH9j5V7k+4/AV+23NK3
6F/lfOQz6LX7aVvmd+9FjfRW5tqgtaGUQiCi38mFFMHRGlvZFcQ9Y4mAZYUsvSau
Z/80nRQMBy5MYC/hI8eAMYeeN6kAewcOnwAh5r8jCWbIRuNwBH9y2l2I6XGXcFav
DYnAmYO6wNMLdl5qv26gMsQNwUEl9ZfVcY8e15tILnbo0HI3LQDjHdDZT8xBTTm9
HvSeVGFSOJ6ztrLmgUZ3Y2MAGRrVV2OaJFjUZgIf3aCWGJhRsASawTvPn84gt99N
JYpSKdoLERib3qg3L9OmnINemyg9a5vETLnmtAu1VvmJlcWUDDCg7NGzwtoCSCfS
6JvzBrBapFyyocWgfaqqwF+MbagypTDr7H9gM9Q6iNcYfw5LWXZ370DGdpu9fafM
d2MDf+yb69CCbRVuY3Kp8xITn0Jxz0Uej4fAHqWovXaU6vUa8DTy5DTgaGPoFFUh
6We0frrGtqthXay/tdwB06omW+GLpy1UwzPKZ66atrNTmhA13pOyWbhzOwMx08kN
DE9yF+7dKIPbpw/SuROlg7zsXKMAgOti2oilPkPCKNQ=
`protect END_PROTECTED
