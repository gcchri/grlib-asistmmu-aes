`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jgmUk2A/p3foMyvfYnVcE6zk/kIdSFNH+fkvzE97ZqvFDuAZrMowmdCrSg9RU1uo
Ua+KASE3iBgdtEBdBBivd89jWJjOutPHZ6TQr4qGadkCyA6BZxzmhdrAqWwhYm2n
Td3e9aWazDSBS2+jEVHGyglkEd0DQEF6TuPihpeKRS6EYkck4lCIlr4jKriHRBNe
hGxtffRVGpe6iGQ51mZarHTXxzLoJIUJNTKsXKysLjmj/qjZALVnfmNKTE8iScXO
w4Zo+6scJTzvthXq2aiI2kp+4KpCSyHLGyiamlu5dsCMQF500OkJ/tJnAeqAZdon
sXDKsklGUMCxn6nq6HvMz41hiNhqVxzBwG9xf1/L/WqurA/IfB96GIZKjRcTaq9Z
ZQF7MrmYIxVAuH25e6xhIZ4HMYXK+NmK7IJOFohgqdc=
`protect END_PROTECTED
