`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jf7KAFH5VEnN1cK+fDMseVhfusRraxGzk4Z6AXUrbufxetLkv+m9BAkMn8FleSEy
lt0B1HcIaIfovWleRK5U12F3FO45VCB9XqdVXnUVRhkcHy2LaUYPwBV6a6RyHWB8
Pg1D0wosDmzJSBZZNNecVY9IwlWFW4tG+nomcfFPp8PZPUlVQY7B4qLW17+trEPq
JB0AgLKmV+y1JplVy1IayYl60QGRXi7YUg6KA2jfR1h5Xu9ddzGtkAuaeRTsBkGV
91w6MtAYFfZsiAIM2eG62446AE2dAmh1cVmDts33CRby6XUOCFIejppM/sF76W3/
SYqD5xdo7hhBpgNttCNtkkcIUfiKVbKtA7H/cUuS3GNIFjPFJuWJVSdV+wTf3+ye
Q+X2PF5vB5GzPb04vGu4ItlHj6erm2i/JTf4QdRj6ugrminCAJ4wUQBMRbQcTzJu
kiTaY1F9iMMY026X+QEvWHfGkCAxndovyBMHO1v9H47c7jJW1SkreJqV6DrUvV4x
ExrsqciYVZfOk/cPhJdvisx0eZPCE1eeyJJgT9UKtuFajLHrvvtpB5EMl7FEnd0U
rS5hJ4VyFHNxwcvz+xP2XeNZb79Jegyl/YVi1n+0keYV0UWQt9bIDT8f8/PDGgzq
MTENza/4Nul9nqdMdW4cyrbxt41htExkmomNfHHsOobnIcp9K/3w596j5YmAW+cM
8v52T1psApX4A+52+78mCi7KdK21X++aAscR990yPF4rz/yHUfbsR9+utcACPELS
+MhDhkKAqodPUB46eM+/9M6PLx5TO7m9lq/KV86oVlCuMnkyYc7Gg41Z+MMoHKfI
xEELBgXtFdpVjDASLz7d5P5E1bv71SUFP0BoCSK1VJWqMUKGCf5eGqW+Lz//D0fQ
QBd4GmXZ+jRv43CB387nkDX63ue37Mb05SZKyjaj+kY2AFxtcq18wgq05i242e58
Ofz/5CTOlMzp0fgUdgc5vutC3M+z9JnZHPltYFvoZ99cTMKC1+f9muQ21QArOnpM
nWTcojhxl/XiaJjwSzihN+9GyWiUL658xcCwcMK2rnPp9aSHm4xvYc2L4yFCylGs
HNoRS5ILvbBeG4XCUqZ8jA9IeTIkNg2McvQT0xn/M+qlReDwOM4lRa9TEIJ2+a/I
FhVRqDVfsS5cEtRhe32e/HA+wtSPHFjwa5YUyCqfDQvhzMSuYwT4h5buvVRHD+S3
tydncb5SEeoSH1ZFoMdfR1U+3t1r+spYf+uicnCd5mYQXAxlpEKYEsI6S/iQIdfI
vOz7AT61uow/tSemvDkJwKCQtEP6wh92QnELTa/XTEEka3QoztBDDRWwtQu6lL0O
uGPlIN9qXDL4B0bKyHW9YweOwB+VhPekLsIaL9MA1+bxbmss//kGGCnMFmSGHgk3
HoDuVee/WIEbOWuvNYWsWbP+yiyQoAkeS5CKjKdH7JA6Tvezsxe9s/qCHhRnEjVS
VGfRMhbOKx1Fc6SNBJEMrViGst30AmgpurVjfBKcjy/E1ZvdOJHLznqydDaD5d0Z
olu70dRw8u8TzAW2TACBOAXievxdZxVGqnQPwy0B6fI5PneWBgViCo4zUFZCOIxH
VbWD223+tbtOoDDVObzRzBw70iNB4cPy1l0Q2g5xJwLc4mdIQYgU/GYa/F2Z4jGI
2hPCoeUos77JR1pU/zf4JbshLkqy2bTqfGm/xlfv9rJeKFS8tEumzfdudWFXliLd
z9zp9T2C+gdftH1/p2nvcHYKnfCdjMjkAM0mDkFOnwI8ngFI/N7/whb5RsNQbneD
V/MKEgEQUbfqCGiBYj6bf4BHZrvfebY+v3T0kWNoq3ijVZraoTMbHjBg7O9UUecZ
6LemxmKAW8o3AkGcfqEhXDDtlRV5w52pyO8f+GdP8N0Jy3Xc4dB3ylpE5E1TLPkS
6bmC78t4sjrW//ObhcvO+e9LpA4YEqI7AOpzQNqUpjKEm9sv0kccY/gkE0YfJnA+
ippYd07giO2FwLAJrRWhLmvfCeOchT9JzpMmZAFunKPO+F9K4w4v9L/wWTK91iTH
d9viz9e81tqo2hoI08c0nvlwm2IzRXCqhuDe9xbHKkJGsTQM6zYvcMKXmobntsGJ
Z9gKPVwU82atI3GOFxyklbMF2jSKCKAIUuZM+PpZyz3/a4zMJqMTH9+fBThHUjDp
6+cNz7GIX5NmDSSIICcm+2ct3pIiTXWSUochzgRcl78IbbSVpoZa/Knekx4Q7dUB
Mj0ad3HLjM45MDh7JbppNIZuiyT5bpDsUE4VyFoDKl+SNfVPZFbwiBigeSsj6lOd
aD6ENymlRFA0IBHAkGUTPQ==
`protect END_PROTECTED
