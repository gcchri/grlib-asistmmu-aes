`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k04Js8Y1tO9glC5MNV4JChv7rnPngw15lmu6+XamOUK/h0n3jeVjxhdOOXcsDKeN
mRcomGy9if+4NSfCRo3tJXXieTeP9R+K4q1KCOTy30/VVlJXp61iS/KCoXmANCzS
BeVAdzm1u4/DELWcxH68jweELPssmmRoHRWwVY5xc4XOEyL87xbyGRCM8bFa/ruM
0NN3bke8tLba9q1eRCqdGzHxZGKyAUx5UgYNODjiC+yR1qa7WCASqxtFhYpc6BVe
+R4SCv1mX8znDgRiEg8OkRoQikeeQHQAlYuhT9PdKZANgQfD9OAin/O+WrX1O5PM
7Ym9xcCsZ26dw6ENLOXhxWzIfJ4T9YfxjEK8FCwgMSRZwU3DvU1V6Bizi0n9r4Vj
i54YstK4iAvGJl7TWZ1SeWTu1o49QFzTjlWNNmPaZdAiMqeT2zLOaCcHa998BuPD
nvu63x7NNAnrRRsYdo3xih8pnlYugQKhnnSHUrpsVWybeLgVHzTDBixiQ64Lx4D4
h0G9scsBsTmXcEdffCq0y97xbEE0ksAGO9Qy3y4dXz64oVOm/ExxDmoOC60Xj4gQ
dZN9AcZSZ7LfKLXpHk7+1mvPN8Pt5a3oOMUtJc2d9HY=
`protect END_PROTECTED
