`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GHYyn44SB4v/9b9YMR6k+ZdrWil2VyMqhZdv/Tn24wIa3WCLaAdXLuQL8vVlGRhk
3lOSgAFnhEgNsKvm33hfKBlzwO3+pgMKKKT1O05M5cCLU51QiPBeL/iJFbEfFSCC
yKJTrMx5wsFQic/iKBWTEnEWOAXZ1wv0QU3CwoXEinjPW8mbRsxRgbpUmBGwIQ/q
ijCps7oakZKVSEktopRSRhivD4jwwhsi0V/95LZc2bErUM0T+DNZ7uEGVMeAWtPK
hj11WId31Bj1ECQnOlQwivsvU/k1iQooAuwUdTHzy3lhirgRFG1NcgM66GyRWWzA
LwnwU2yUXn9UbCm4ov0gXDnED5wrIswCLQlCZyy93a4=
`protect END_PROTECTED
