`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dt7mJLQc7GXIWjf3XkthvkCTaw0SL1kjfaoBeceWoArieJXd7zHSOB22w/dblSvp
vdrQpqVGT3GR/T0Tl9HScluvidzFbWtXomV+gBXXQJ+N24e8Bdsz+wPz7kPNp9xt
anjL+o3BRK7Cnmt5a8+J6GMB47zx1HQmEttQKcdNXjuE2vyqmrVLl9MiaVH4jMJZ
gwf99Lc28ktRLKBumWE0USIS+gb1jmNPMU3OQQJYR6khtopz7CA1pJEL4Sryww57
E4r20it1NLV4MjdT8mmkB8gfJXo6q9PKkCTx8eUISYutaHjT6Doh5T7zRyedGSyX
+eAYI9e8lj6eqoXRo39UtPxkj9qrxgB9xXkVLHDluXufyOtOs3QtghA/U1r1nwof
UyIhMRk0X+1lY5Nlh89/DEKZYmZGCd0Jky7qBB/ytHb8d00+Qx8cX57GIED9/Uyc
v32iBobPzMaqlynFu8+2XYuWLOszV2xvRN5+pknyMhQfHV+kUCvLGIAxm0hETNf8
3KfzCUGtUeqV1/ugWwxbrtguoZdj/Ja/Is9TvMf+ADua/isIE4DzG7FAsCW/HhlQ
bVoMQ59cQJPQyhRGGR8cEi5Xdfnj7PMlAmxoY8zMmDvF9jricugmA6Tmhivj3E49
HLoA0qln3yRmy42fs77Ko1EgE3fpgIw2o71jvdU9+CF4DZL/qXn0odZQjZDJtyCx
qxIZvD1yoqpx759YxMx89rSNf1TlxlP9Dkp2vNi9r99tKdc+gXpE/UcPUfWoB4x3
oSj/FTCTcZoq5d1KIkm6zd6CWgboiThqBJJxuMYoihAOunXdklw+8B7vKY+yVMCt
glSNzhoJfKYao4WXaW+MMEU1Cs867AsssQqPWBbzvUHVLIRH4+owbrpY8b5HjKx6
8TLArBAb3mL/Jk0D7E+HSmEOuQSlNXnG0krWHBV80FE3y6dQa1tN6Q4XuSZgE/Wp
5DLvVKWscEWNIPLkQV27PhGdXXpqAG1im+QNAWvnJ9R+O6aeQq3kyMUFwlcNapBq
wWhRy8gzNlWGgz3ocgsXHLGejrUzYk7Adk2L0HD/fLeoWRFgo7ipu3u8C14gVvak
ZDz0irCSKnn6PidfVWj2M5DApBe8ACJGz39++A2AmqpPaeA9wYqkxqCA5vzwD3iC
Ktgo9fzpc4Y3YnpyV37JHwUMtuFFo4lsmdyg6o8jE78aZhe7xRPbNpUXSCkt9gwc
+gqLZMZ/1ruuf6imhEIAgWDwJ0nOO1kQ15nlBmXrzi3V1KpyieP848f1crlAHK/T
2MChEeEQeAEAapXarc6RxU6ANxv8InBBz+o+85sAFWGqBsiMUL2T+hVbY7u0WunM
Gymtv1jfxyPyEuPKDaiXAihTi4OWg7Bj7SA6J8CGdDpXfCivDqz5yK6HRHrWGy9M
+iUEiRc3WNcoQjW//d/iCWoOESWdYgGh7LlGgw2DfrraWLmbD6JNCK550ke48270
EfAT4mhJxXNJbIZB7hdqUvJ2YIL3+7ehuOJ46Get39Vth14tHBG1ynYX8az6oWFk
6JIFc7BTcdmBAeUt0r29vM/9JjhFcIett11F+DPKpi5IyiGWxI4cCWK2EQ5SeldJ
42TlB9GfoNwprQWxAmSn+eL4ziLva538DyYIBl51lmHVrrX9mw2G8T8gnLYqH8KV
ffi79qGT5L3LVpg7b3yBmyyYg4r7xxLP3emcIvHbRccs5/I3HnpfAM+ybC49U22q
gelz5MWVzOO5fGftDydTXUu3vtYAZXUHzjLj5WuQVRF/qMaVsz8/yum07XWTn3KQ
+RBf35WCnwp9SbHICt3n2OKuJhyAx+A5CDI7emiHLK8Ja94eFLm76DPjctsWvfhC
bHX3DPtJNqfpQIJdziVYdf5eN8t/MpWTPgmcJa11mZKdVMufH978qtFPr7ybEK6X
/6YMhmxV1Jj4I480B8hsazcJ3smvCZcTHR4cB4jxtuiU1+ZMWofiZQ4y2YqrzR2o
utmhX7n+mNAX6MuBdJdJB+P2AC7MYBgFQiIfG7tCOUF3HPM4PgvHeZQuCymP2gPP
Pl3j1otaAVZH0cMezuegcQ==
`protect END_PROTECTED
