`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vNe2r0eRR/5PMpNQWurPo9r7LW8CuYgL7m2JSL3iLTBYMhZZ9+aCmzArmErMJt8Z
g/9HK3dviJfZCeYyq0u6a01241N7hA2xEsEeTWbM2+jneo8IncITzuAPb2bgjVGh
aUxcXf78/3cXpp+9OcqOvStMrhpAPvlBfv8D7g7N+xyWkcOEcVgHO2C0qgG+9LJa
XI6jkzeyfh48YybcpPu9+S7MLwPL2syOFelFIf6WWRLBVXAtf+qMemt2GeZktjHn
Y94fsrdDWU78vPTF0xe+/GsjtipHI/Y5fY2NlNcn9DL21H4XRcLHitootXcVgJby
G45xiBkBU0jznGbHwLvPPBagZMs0+RfbJg1adu8sJ84ch6GwW5yXkdJPjbBnIGz9
wFI9ntfIpAs78jenTMf1kYMRYDtxSl2iFSdiC3nhTCleYR/yzAt4CchSvetKW/ln
riz98Clpmojoa4nMgLxL0M85dVs/xYS9rB+Ex4PjEh+fIEcHUebI8VkLWKkynm6v
`protect END_PROTECTED
