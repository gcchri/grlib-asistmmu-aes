`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a0E/rDyprCX1D9OKEZ9vviIzD8rRqufhSUQgZHcKQAN0AfxC6NzykagdgjGLm9Xe
ntjppwZ8g5JSL+nK/sqyrdYJFxk5VsGgQXzLkrlb6thterHVHh+e0nc3NP1EHmi+
frB8b6AOfA7E8lAQZWbpNqnlVx4aP7yx8xL+xITJs4XLFYUTpSjwXxXwA8roS70g
TWckt+DwYycDCGIOUNi+Ea9UebWOXzee6SwA3OMYnSkbyXB802ZmMeQ+9lvW3l15
JKU3l+OSV9n4l/r3ued14QDmbEg5Xc1BM+jr6BKhbdQCFcib+NWbvrqp0TS7XjWh
ePvzN23vs4HTiGI2IPa7TQ==
`protect END_PROTECTED
