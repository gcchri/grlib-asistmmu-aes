`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
47LAQIRjbTjrh+BSEurb9Dk50miQViU2qNGOhr/j5RXeYar02kJXVLtPIvWf7Ezw
LpZ8aL9b0a/npcpBE3yT2CfgLWy5Q2AxHYLUGb+xB5dMnc47N8juDOqRHPc7anM0
nypjTsRuNeEWy+Rdy4+uWLKOoSuG1VSFuIbTt+bDIUA1GR4Mg55MF4ip39Teq6kH
ASrqaB/wf/N1wt/TTKOf5OunwYdhvZHlmbotpelLPNRRzTum0LMXOlGi8lTMKzHK
tuNhjOowX0jBsCYha/8hlxCtOwHg9UpQRaL1sGW/8bhFha3VHnhMYVJhvRM2Sy9X
Pi7JrT4zb0mkUU6Gmg132t3+O1XVxdTXwSeLhxOM4/w=
`protect END_PROTECTED
