`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G3xq+Zuu9JJmmUPmGUdXjynQ06M/k56KyH3q66RR6pi3dyYkdl6W1GyCkuEsjIsa
kjpgEd7RLpE7w/pG9EoV+arZgIP6y1fWHVA8iY9rHKfkhL7s8NPFQYu+NN5snA0j
RweGwzCfpzUKJm7TZSFLLkmdaWxFrWNVRYMqqnKvo7SqVTqMTeRJgzIJ7fd9Zw2M
HgWB8OzjzxCBemdIsEE8DRqtBkOuQp0B4bIa1FM34nxdrhi9vC3slZzz0jqv0r+H
Vq9SE+4sc5oRtZjjbV3bPIitxOVYVIMn8MVDduBkRNe8yDGdaizC5/oqbcQsJI6h
GZ4GGo16TLL06z7zLUiJECY+cqQT4JAiTBVISQML2KS58h7VgR2Sq//vQvhoLCUa
bzzkBQCy1EVriDBIVy6raA==
`protect END_PROTECTED
