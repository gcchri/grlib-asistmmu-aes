`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j+OBtYotba7rjLn8GlM49XilNnD+MB2Q+razrRJrlsP2NUoLRYQxLQG+I4uGixk1
y0w+2DPXoc7md3L5S2dH+jH4F7TfsLw1hoJ8+cCyC3mHaU7SJkLnW8LP5UaQUMn1
WZvpEwZWU4FQNiiHPJExhe34zWWnYRf18hFBFe44DbpAYciLUu2cLsd5mLk+ku1P
kMinJOBI/59QRblE6/iqlDG+M8YgAPEph4+Pu3wo/+Ejy3M2Uzr3mjTtqJsFIBwO
o2EGpXu0ECon88vCbAyknugNLYtnxJc1uy9UrEQwV5MRw4ArjYDm7OOKDq/m6K5P
J39YbW74aC37gIb3v2gQqFfSBw2beKUfxt+fYCv0CvU8jrGtOLY4w3oBLaKrPzs6
q0bAt01BX9v9kwaHnX88+g==
`protect END_PROTECTED
