`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZRZFZwlKf0FhttEHsORt481cVwU+wnymqG/kZ/mWPj0P5AByE7keidaUH/CUC9QA
4xLog0vnSbC2JbUpTd11kz4j7m1aTwp49416Ku1QS52LdoIPon3/Ew+QH2QfxjCr
MsA4PLqOnFzzmlajFSCMO//m/AI+Z2a9G8NdvmfQSC8Hr768np2K97mSkjfNSDpR
dBBcb6biEyHK6PN0REqaSib4AaQZWHYUgZew9ChWVoh1gS8piRoU0yqaiToyevbm
P/kbqlso3EnI8p9vPhgd8nHLkmUMObZ4EYzAI7GpICGhHoaR4cWjZCag5zJaJZz/
xWeBk1YDK0IKbjyBbA4bhj4G41aRxQlET4uSHJCYWxpd4SDuDzKNV8jxGMzo1Zdg
qN26bMM50Iz+VhKv7BCEzHiqQ30IgpoRrKKAa0a7WXsYaKsvqTe1LVu3jOCVbOVH
2VBl5qV5fOTs6CNGpeeSOA1haq9HWGwjNFgUtXjgM5KDluYlAb9cnjH3lcGFcZhN
A11sPrKhupzT6XwheJdJXgdn8JFiPiDa6/LHjF04W07RQwaHzwTIHk+AeT/C5qwz
gqaoepJkXPyvhU0WLOr3FZhmEBDcgpP71roTk6d2CWGtlSYorQ3uLuLMk+/1Fyjs
lD58oRd7v3ue+A9dyAs6L9GbUWZMyuCw9NjyeEt7qY2BYvi37ZrjjGzUWEFm78Ke
`protect END_PROTECTED
