`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k9X1mHUu9VSqZN8ciJO0kjB7mDh0XrHj0QfkRCdQd5lpIBeSEau4qw0W8sDO29BW
nDBqJ12iMIQBku+jQnDydfgbnq9BQvb0i2Zyr6/PzusCRIHK+wsGw6hSIbHuW3kF
NxLpfblJhIgRTpQsPg4RTb9gYywt7QF59Og9bCr9OPUQDGYf4WnCLFHyeDtRFieh
Fj/2H1qkcr/XqoZJxRCZBBitUf0rQ100Cz/Y3tvfMXF9nc/f1hPf39OBYXZwaw5Q
QcdJunXNve0Ma+5CDB0mj2ZYlOSszUUppZNYzoLmBs/iSj/JsTr9mCZouxJ47XKJ
UgJyCEpDJPWv/0/6ZuvuMn0xwXADHq4Gw7aGt3F35joACq5ZNqKWlmWZV5fqT4uk
zh4mFhLokQt4vP91n1HvMujPLhdL/0NAZg76rxQhkja/N+zAvzHjaN7BTj+bXvrO
VfLSUv9CUXhXr47MzfWSbknMmyu58qjW7jHYSowPTQrEQVnNyaAM3eYBfxW28xMa
M3hkL2LRj6VmzqdTcovwnIOB87kToGF/BxJ5UBrKUeBlMANNBrx2ah0OJjw4HgZ0
3ZLJfgjGYexf1wIsycr8HsI2NyXY91rdl3BiVOtvCUoR2SGhkcjhdxhLLfv/C2sK
UN7txMBOEDMj6k6L0hUPbOFvLNREmpeeDcclmlTe/1LBY7ntNhhrH+W8dDkDMPmC
sarohoRlSOvj3x98SE3hUK7w8j4Ww6Z3gJw0RgPGZwUKhiqUrTEiZZmaI0Hd8arb
zbdprWrXI0Sss1Lp5NcxfsJ/QV4yPkIToqJYqj/Wkyj2EHHuZyYlgKBe+CzVLYn+
pA5WUfyyCxliJXgrBmU3ntx/AdblS/CGnx1KfKejHxIx4HSaWVOiIp7YQ4A1gZ0M
FIhTx57odMVPrgRnceruW/V/6W0mf6IIEh63bbIA0w0uJ93noim9qmRjQHsu6QIx
Me8YNxK/ROkGxW5QUOlppcr+2TAhagu2nK1qzc0bobpDxxpuXYzbPM3ZGT0PTX51
Zn1f0QPAH8XbIz5QmUdXgUCjnNLmjepeZ4I1o3BH4CON6vSTid5djkii2rOFifen
13O+ezJuJyN5/Jecw+G1R0rxKAsj1HtdkvLIP4+rPU9StV9iGMD1rAicdRWnHzDh
32s5IIogKcr0iWq1vo105zSf2bewF1XbewdFFvFkXK8eyHqZBxSxQDfqOjP4Ad4H
6kdOH0I7pyzR9sYlFZHmjq3D9fMuH58RembyO1n9ysBJDN4U6adyF0TbY/cFov42
HNxpSDHCqkUAp1+2okqAs/H5QtAowDPMeeCpIZXyg1aVyQ/dl+W37JBi503z+7eV
RyAZzXjSjDxiPo7qbMe994MpCEZ0k9x5YykEy1uo9ZO4shtwZV89pipY7gSSZ6Ct
TrjO0FHbc9ngUKj5JaD3YbDoQZpBiKHOj4JLh89edyPcHETrdbeybapWsuGjLpoq
JRcESBgm85QpDFPw9g1n3oYpViQCWGor3oUDqZZGzmY4iRCj6/ZVM8nwrGUyQuRN
CCUmdCscv5h1rVx/Cqhj4VFwNC5zZ1sdQ8sxg1RsO4OKAM2bqBZLTIWjt7aERd6d
dfcm/28trfMR6wKw00JSAIEfD6nngD7pAwdEaFC+B5qRowVZid5Qd6Bay7bI3yrw
L3UQYM2bFHs1G6t+Y1IdpJ0fY5zhnnha80QvyJOxOLffrGAnSFBpNDLvyi3zlcEU
YS/ovKDUe015qwE3MW7dLIkfKuvU6pAVfuBlprUxJRx7stWxIEnauhlh0kA6wA5V
ezgk8pHTXjk4h5cWyvkERisQ8tN/2dKcpp19Jq+U0KbdWN3USfhQdfcU2oZUY2oL
L+nXLmGczL0dmb1qz/aoDYL/ycAzs7p2vtQnSM40qypzlQxNAiILGY6zlYmqclo9
7PgGub/er4PeETwjaJsjTIBYimjuWQmzxkEB66TKk8afwIZrjkPsALxz7H3Y5Rgg
A4NeyAd3XOOHeXv3SbA2Bq3Z8KasbSzIaae+FBMOgwGDBVFWcS33BNzE9rSPVVdQ
48MjDUcEksnFxt6kTk8UsznkF/HEWABD8qmpYVcn/0exy4SjEDZi4M3lTTIeGsSr
x0f49/2he9EO07ZFAfzhhJptd0VkxBe9jCWp5qyRcsQKqrsQJBxLQeh+6ghSpmrJ
IH1ZpzUhkP5fvZxmp/2S3XK1qTgbP51HxPfX/sEfCEUndspgdT0ax4Q3hT3xVvzq
5QvGlBrcz2wvp4sjdOWqs6sJBbEBgcut5ZaMDewcRmixL1zrJkTJf8Hiw0YzdT8e
aO0o0cm/hOW4+7eH+sKRHhmHyuRclpTfXRnc8ei2lZj3Ajco+Lg2A4eVLIr6VFIm
Ys1+/YE1hY/MEG382dzjbc0VGbxhtP2MXkqaM17zV+q0ADcuM2hKDaTM7cIhK8im
tLfQb4ZyEH18pnenYOjZxXxHZHTT+XLnCQUzio8FXZN2vVpOZtu6a+wbWwhAQdOL
nLTsxRuDjGzOGO7zOaIRGl0q/3mAmXKIQQb2vkZPV1EHRkVEW3ZAeEREE+/jVgt0
uIqGkMApAkrQI2O/fXMJdvO/gFM+o8QuVonQNX8wGf8taonOY6dgpo8l9+UPPRtu
vXidW2GLudgVX4MhIeMPt0yBfd+sB1e5b8QN9L9lG3gf9yHmZTIcFwXVDtmBmNHJ
isQr1NoNg2iPdayECPNOGWo0vMVx/qq3javyYuOsV4b2L16usYwJ4oR0PvPKbQ/P
HV1jWf1iI1EjP+Me/ItpsS0MBufnuOOSDM62F0cWrvD68Lu9q5fcZ4FYY99M1jgd
GZm9Qi20dJIOEUfF31nBjtSP7nJP6KXPhQnEQrrVPUPQ3mi9xZLPLG32Fq0Ih+w7
sGtsoIjfA7nfRo+sWApox9l6dHr3B4Z6vfNtC+s0cL0tTlidBix0nrRfwN+0zoc2
p1//0mrXVRS9UlJUpsm6aaie3lFd9e98f3el5gDt7P4EMqGhEgZh7Vrpbtq9YP66
I+4bFXXZcxoutWZjXEET1SbTgvz3MxI4dqPv1LyxnGsk6jIoBgsmxtgRBJeKG+F3
BjTsuT52LOE2NDTxlpHFG00Hw9G6XugQQJA1LLxpZWRdTexal6N2C48KZgnJ8S3j
qwjnFA2HzlLE6Vo3NIqlCaL+a7KsScGC6MNssq3bkuV6lgtknORns8+yY9kQwXZr
Sl7zF6Utzde2WV/sP0tdykXeOlpVhGxY+vDyNFlMUFGAXpPsExIMO/J4kREHPoYX
f0hmycL98UdPF2ZUcX3cc3EU62Y+cPBCD7WEpVTZgiG79Tksea1zxMhM8wPKk7IN
4bTy6U52sXtdli8IhyyWrIr/gSSlxUFnZsozv+xBtog5lNSqUzdyLeqPY8ITqLMT
++hDvAnHZJOTCOwgFfbpk4u3F6RE9gIfuI0TpMqrwajMLMOYudoSOd2QEKqcN46n
6+Mt9IiYh2UOPXpQsDD8DGvNTn32BDi5YWnDbg3OS5lgw803LZADF5Ceg1xTaUIx
jYUVcittxExv9nDTwfUxBji/PiTGIVPecpuj9CvHkvHQM9Be7C3oYui7Va90Qgqd
7lfIbT5iH9T5WFDlsVkphjmN8zCv4adTzC4/HIFU3szicTDRM6e48/G3l3dnqiLa
+WBcK6JhOY2IVa82Mhu8Pdwo3gJBd+CZt0shPjUAH6s5H4EorDmO4qDnQ08BLZkp
WIo7/aXsolMf595Ig92yFJlVkTqq9d+ZRT5Tqj+LBbbZrXrhmktSVGwjh4geN4UY
nOWgixWXA1dtz1XA+8fWHvuPIrun7IhWsUX4/Em+9K7hZfYMEX9H54o21xGkX7br
EX7WA/JQjuB6smBfVWP/dIiVDSjKu/qVYlU4rk8a0PcN8ODxdwJ1M3adKIacTtRk
saZaopQt6cPfmNFgyyO9o0kmYf1Qe13yLAZishDpcJt+7Y0HQ0j7l1eATviWePoB
6pj3X84jgT+iSE6vctGtD/Qm6Oh/ko3xOu4zSp7Ym2/kef/1lKRCJxh2jO0auqE4
R7nqXQTogakgRxSOavVMfQdq9bRGEFy/k6cn7HiTu8BRizBzgpTdtBgPKZH8l2dR
6vA+Ads4GM1Ohq0Qa9N1ekWB6KLIq4w3y7Gx/htlYCPISk9c/FZdgiWy7siApfc3
pzh/thoVnIO7BL4oWlueGumzUppC889hjM9tDFw6xuhaNWzqIv4UeU6BsPe+LbbW
zkUGgkEPsdcuyo3Ix9AePz8ptMv61YSy+fBTxU1gJoTyRYtizICEEiEwyxA7pf76
lNIoXI/Vzl806FjjKw7QfqEv/PkUkzaU6lhVdO2g7Z5eTJe9FxZby2J4ElcyXxkk
g6kKMl508PBMFeuzeIOOdUL0PDERl8YiMmgqdXliVqkUOGPLk+TJ+wpqYEjXqPUl
Yvurpm1xdiROx/A5pc2eKhcegenI4/vMl91ugTRP4BE=
`protect END_PROTECTED
