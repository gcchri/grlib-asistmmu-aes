`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4XSVY99g11MH9zqxyTFPyV7emWHseoxkIVGN46ThDexviPMe4g1csycoluwfW+E0
ajrEAQcKtigrYoKIopKbpLylWGPt5y0tvGNuFrgxV0fG8NBErJRONp5KsSn6Ta34
HJqfE1hTEjdhNHmrEOeufOlTR5nnpEdK2XnEkrSgZ67uWv+iTlY1TQU2yCkaMrQx
+u6M62mwD0sHiNuZ/X53R8QGgvC37RPIph1nog1mdbHDwnOTfw0638DGtw0KTYUG
pCdzro+DMp66nbqCjI3fD84ycWRL7vDU43y4uc2EgQs/1k4gXxgzim5ycFovfdpi
uhStzftvX4IDNJy2AAeIJ+S6b43c22uq2L1XdTvJF3gI7Bc7amBTohiVb8oqIToK
pa9EV2i4SOI/ZZrWk2IvqYpteaW67qkUTHB6OMwOHPN3RXfeQXievNvvVdjlWhWM
cvftWFSI33HjGMYDowm9zSxLrgfOzGIsQSSs4gfYqtoMfPQ6+3yPXCTdkq5VK52H
LRYwjpYJUqa0HdwJsj5AC5l0lGMCt2byk711OknZ5GhUYX98T0WrsCEln81ab2WF
qGq6A/hkAQEmDC+epfLpsoXuGuUAG7Ggk94rz2zBdBnWsPgJh3LAsk8cdUGhCtBz
sQzyIkgjqr+lXBm5sGyAw2z5CINKlH7td2xWEUnbeN/q/vXijnrH87qI+5WP8jll
3t2zFTXvjEg2PDFV2Uy4KSRjY/7X/F72QLm0V3GJPUSVudyF8XkBYImLzHYlqmK2
ySX5bqZiwnqhLP5h5uWZnrYXRXXRhn/hQHIfLcKxcId8uvGvG2ITJXpgQsFj1AQd
IxnV136de/kh+AoI2HHW5Oz/xE5h+UnvEWYWI9yU+wB38GapcIgyAvFPOOVCs9aS
ZXyfHWmcprm6cCatVF/nIcbRHLL6GCTSEMSuoBzsZEzOESrLOfexCPd/nnXQ081k
swXPuy93tHqTcEhlOaKg3BAQw7I/sCICF/rT+xAoM1JqPolejg6qrOC//ZcFA3+O
p6dcWMmsMe1wMj0SFvI70dPaKVh30TJDJQGk+9tM6UWhsRBieBAjviKFPwNJpBbY
DurRBUqpASBl7gHrPLcCg47ZITIJIfwRd5jkmW2kf4b1VwdxsjsyQ0wpzNWS4deQ
IzXv+utHHU57RHCEZZAqx1KjuaMdAcIrjszTDmV035BMFTwkjkeR60GCCTwCAPZe
/674DRlC20aZE9Js2AlkWWQqYRvE9SYJLryPikcd/y4HruBGKvD6wrPIalCnVb2F
C7IBG0BbVJHRYoNNxc1gmY5KkmeIKXsPhBTfsuPKlrDBKZDK5UxITN6kcVJqYNPh
n4svDIRohvmKPtqaea0lx7BKvHmQ4t6T2f4aoFTFGTytuslO+sDKG5NdrVQTQIvt
/XXsDOiIp8xIUbpykSVsaC1RhXDUY7Py+jrX4BIItwbF8OKWeOrprw5q7RU69Kbz
uH8WpTsambRTcndgoIZlLOU5i6Q5oxHCjRBOKyUzNzskodXvSQvL7NbZGuWmohXt
Ekw89gqsTbr/2eS08M5vS58HAC1hBPKsd1b5A1/rZC5aCMnQQaicGcD7E5Y5AjCO
CvSqYoYL1iy+R/fzsPh9549/3myWCEhpYInKx5gm8/P2q9HB+ZK4BUpHhmHyF2l9
ePmwERMd1QMMscV84bAkiGjtdcchxMS1y+zzcXTm3dpmUcdZzAq5J0TG6c301OQx
I8/tMJfolWpB2RGEUSp9OYAY0XwvNW/xJZlrAjuJO2Fdb2hUlU3fyOY/no0+hncS
l6OATieCs6L9Mi0snpjGPzMjtdYxhv5mQddKtjoKVwtjFQB/R0Vvun5deA1e15DI
JOqntGX7Di8x1oW2ei3lD37vzmAgHvviwYykkCMVimhCTc6xEMdsYgFEyDi3/4JD
aLUY6mWgHa+ZNiQAk/LOxfGKWT2M8TvfWC9EaoQcXjBGXEfNl8ENke+EOojCSSox
xDp3nZlZ3VrcyCjaSY2mQMnyx8knlGmIWo0iR1WG5XMMX1z5YuoZw8z093MHTlhB
`protect END_PROTECTED
