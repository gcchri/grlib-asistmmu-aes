`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a8kT1zYyZaqxVOZKoZW+P/8k31K9KUOIXjze4Y6tK9bFdfsIghAJa44a2BJ6quMM
mAuszxEXwP3uG/DDI12GbMapdHZS2Y0dCQtQ+ZBgnbkyhQ+dVOKtgdvm4fd50fTz
CpD3y2luDoMJGDHB6ifBTaRlYWy4ArWJegHmqGBcktJpMP7YkVbVN8luli7KCunu
zLV9K4WtF1VX6BcReuIXvI+dnWVucEz7jX43ZlaDGFcjoYslAuXBeDiAkBCpDbde
OOISPi+nZc4WRpoHn/b9cqkOJK65DDD0DRq3uFS8csMTa5kbj9pJmW3cUJPaOS1E
HbBxuGPQ9OoCcHLpU12eYJg6qwLKDFOlZPdZb9yitTG102FS7EGmPkDJGMvDug9W
hyxwSO0w/q/C4yQVXyoqJi7rSvoHI6qhMGrACm5rAzGXhvgJtzK/4gs086FgDvCp
WaS5xeiJ1LRD9qgiVjvGU+fQahaSIDOG0CJ7P2f0l/zwi+Z4KCp6Y87oxf86+q7T
+wjBP3KMWEAZyW00a6xxCjRQ7TH1xSvVFmnU/mb3MGpWwt9aXie9RkT22RSx371l
rcCBzHid/ngLWkp9mfMEg/L7XEuwCd7b5Y1XLVkQzJcWLojtyoD0NKfEYfSxzD4z
ALx2G6CxAVn57UReq0fNhJ1fvVAU4nhp6F7IgSSNPBJ4pnvqU1vuw0qX961lsS7U
zDEmzJ+KNZPMfih2pG3dRgY6Tmnf/gigsqB6pR6Fv/BvfjXgIyYIzvqZt8CXJ4pD
stgHtZVjNnVL9eSw36zKq6fw8FEenXytNoCdPCJUeIxvBhNEl6Cj+efHQXwCYsSZ
utI922K+zdq0sb/qI0MTcQ==
`protect END_PROTECTED
