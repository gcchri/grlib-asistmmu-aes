`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BJX4qd2dcCws3eRofLKZ5p0JJiPoHQ5Z1GTCf6w3E685G/Is5/fz1tIgstpU7b/M
fXykKqkigDOgA/Dq75mrHnKlQvkx4dE0KDIslDbSpKEFgpyoQnNXcqiJ48sMcDzp
9mhHxY/Cjt4YO+Obtxn6vpqE8LySru7YW535sET+bfWVKMLR/rQO1Nqy9OCDfRsj
lDb3W3PCQpayc3Zt8cKAhFhzTdy61GUx1YtogqcMcQJfozCoySQ8cngnedqF+sQR
YQLRYFjCTdf/zm3MCyoO1PtnWyIgGQ3cID7sLPeIMjsidUYjdjPwB1Ib7zgFPOpZ
DP+/H6wQ9YnDjjr7MMPTuwW4bSZBU2oN3qX5rwO1HzGOpzVBnIWd6200V1EKNgLa
`protect END_PROTECTED
