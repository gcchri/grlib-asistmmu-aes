`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y+50Evlp18vbI/nYxK1OTcZ3PZxWBK8ebQKrRokxgVcfCD8Oh10uyhfk81gfHMv2
DPX5KxQFvgBSuH0MHW8mFYzQ8huHPAuZMKCPNd8D443Vv6OSMqkU38cv1qiWGE4X
2aQgTS64eIHE93Vkfw/JBum1LdrKCvJPYyb0eGdgtoiHcWJtCJGLtlvFeqctZseF
rZyIeshj2x6eR2wE0+BB/ezj0jPq5zjV4OL6BAOM1kgPGemdWUV46K5E8kPVVMbD
Z6qslcctXWOJGjWNIDLlV0D1pv1JzvoLWVMK7Z4MaawvaIkdNPIhh0GddHBLfxaI
c1a5C6t1f2gX1SAmWfULFJWX+Vk+zuIcztwGLwexDJ8eeru21JOoOWLWNDoAUfeG
FstSWuPb/G4VhHnacnWq3LJVZEUdqXoqFCVgA6rH1x5d7rlZlX9WG7vC7x1F/+KC
UlNvv+goV8agVE9pFDvVW4UszB5qoBSEwh7oS21HlSS2EqEqSrOo8SFUJpybgdhi
uE6NLVtJnh0xAEsODe17NbBozh6uqk61IjnFzgmjtHpHvR54aNumxuIFqyRY6O4B
rqyDhTZcMgs9WT760vZ4AYvp54/a3sxGHRLKTyXNx6sAdC4aG7R6BlJpfheLnPUe
dUrPBmHY0A9ybzX5oyhrr6mQ27plrrXGB4bADXlUHxnMoGSp1zpRIzg1LNAPkG0c
Aly9pDTw73EtvZfrAaep0wwrbRQg2IzCJUAPJGNIyhG+0wW/CLiTE4erY3m+Z5/6
1yN6iMGryl7ZJljCinEjmNtnKrBMHu8JhYzBF+RItJM+9AedT0ed9Sgpc6qGGNZw
7J4D9u6wFd5S+YtnG8+2dvIe+IWtyK22jK9iuHkWKXekzeITFq5cQoxiRFohcZBO
+QxSTxO+kVMcD/TVZpzEOHcJSH44LCH40fOWfY8SNkoMm+X/s6v73GNfHkyodzbQ
MyPhI9PABazJ9eTNtN/kLxA7bJRzD//6rdvYvVj35H4qgh1qrZFI5dRNClXXS1wJ
0fjoHyTSrlmpP71p99/2/hZCTrSTIeSYCn/i80qKus0CEXZguf9zDtxExA49cJe1
MFPo3oYxmXZJ+XUiyFpus9w0DIJXTlvbe/qF5IHcAwVd1SpS/jq88/3mNmHHO4Es
jySrYzulZx14jOuZzEidHUvFPP/opf3yMTHAoRdohxSOxVobkZ9P/pIvcycV0IOH
2g85FHA5h/eHBpqTagfouHcyzQuQ3qWU+s2hwWHftdCbGaCkFEdP8E2Ql1geWNsX
l2Ghr+MkXGtdIwf5jgIjaSSFwYRciSHNi9EjT+Ub8GgK7gLo97MFMY6bKrGHKjZ3
vdsiBTZBHuNHJl1+kK8AeyIhDvEvXF9LB7CUm22Btf+2HetWHZHC0bLm/8dYMDKi
0U7EE+NXV2OPGrAv7CQyiHv1pJPuYr8nx4yLFnxwtBu0Yt80TZt8GfOrIri8C1+K
EI3pMFSBQIIXlos2XcQKetHK5qMVIPmkzqrlHaEljhQs1ME77Z47G3nVXMAjjJD9
713idy3zNfjbOBOSho4wZEGIWS566pl0a0RyggOO/SmqgWziEOGIbqRASJOxu8i5
ME3JhXfivQTltzTNc9WDTlx0a2PBVL2x/5VltSNceKq2ZFOnJ0SXSJXoBxlQwfCt
RJLy29bXb1qfsE2XEwMgFzT9tA5y2JUnT9gI4+ZkBaO2ljJCQNXhAk+frqCKG/A/
YI5UWrx3POESV8rBTomDLOZG8l+HvS4Y4yJ3CqJohX4M9Ot+SPiW+CCMqM4SjzEW
P2Bh7s8DUFc1s+8FkfAq9zY9P52/zsIaW0/MF/7se858SjQg6MLlMXyQ6VgwZI/o
M9QEPw+czcnKvPz974jXMiMhaVva/7jIfbKNxoZiF4XzB+D0J/wJWYu2An4YJK4j
nlpFOirjZWuibAxPMZtFZG26czL3J8fIyqj0eqfQovWE7PzmJ8CTisJxDmnQ7mGf
JkyC28nDky5rIpvMCIDujANT3c7mdVMK3bdo+zqS/sXzXCJ0sm63xnQ+BSucl8ZO
4eMtW/Koq9Y3JQRb7lJoWXHU73dC9wQOFYP54jnXUelHrb/lnSQKIDf3ydu+2W4p
U5kPxX+B+ZrMgbDTOA9Xw7j6yCZUoDzfOIPO/Td/zpofW0pwhmM4L0kofc9koF4s
CohUqT+FEeKjnlEVTwwvC4RVf9MN/yQceakX0XQv56fUECpconI4pFln74Gu7Oiv
ZBZZlCW5ljWEz7gudcfTPkcwesojoaDT08fJAHVBiuTtPL2gyJwtOsPdEkhzE1oy
x9nMZc6nmdUxPiQOh2Bm1e3lR28yPzl4JinbEkNrpG/eipWsI9CGvP6aggLKQOub
z/lj4eNCzuqAj9ZENW8Qy2tN8olmml+E4htU53oWerJzX/bBXZJckMXt8VzZSJbh
oIRsJwkqpaZYTk7RhwjPCVmAq0n3R4/HdMHaXPs+JBYNCW+RbEPgnAoTWfCKlPTG
Bo99+lV8bRC9zHPXjGo9dPuhl4D9AT1AQBNHMbCHBbYH3sD1Rco1mVL/cGKh+LM7
YzkI1sKIKC9VkQZrisCvHE5JJfi7pKlZbluEWJBhJpLOB+grf9Ng683Ib9OonMba
kDBtRnWUImICt7H+yAQjlzvsXpZquKrL49SDbnpVTz2BxXVLZW9lV5zfLjeeQs7F
R97NcIVw977r7AYx45pT/EWtWFb0Hu3VLUAXhQ5xpQUB6ywvoiTmNm19TL49aGne
4ST1rS/pUeciLWgwV4zg+3HVIoSj1cgJPj7QH5uctRctzBYNT8zLPqXmWdjPyydX
cWaap6pQclX4ZVdzpMaqi7YB1QCGy4nPKjWnrje2Zq85FMVf3K6gdx+bw2xbiBz3
V1UG94/u8EjtGWFl3qqWWkkx8zlMUA6IIHRwz4OL50XUocrFmy+pSCNpzg2olfMv
/DcWpWHhdWjLjSAwFjvHkLNFcoBHkPwe+xqlqhas6Gu04fW6UtXuLfzw7lJk6PGI
y5MOr3WzIFpKYy2ff9Yvl8dRyvlyTjttQEHdKCvZWLP2GSgvuJfhJzbvTZa4V7dF
+5WdvZYUAhxSNQvvUekM+Rff4T9n4Mpt7zbZqmDbsH/97ZLFBVetiGuj/r/k62oH
gcouFwZMQ9knB11LuwPTj63+oaRc9mupXb8/sVdUCIneHnC7mQF4xIGje/iYBfDa
DXtfxnccRM4dWvJsKLpxxzLXbPfScgMdL6aMmY7wloSzDRAgzVP1iZ3tbc+xSzE7
7jalScLylZcDKh9SmaPGnr2Wjd83aIUbugkuwr697iHCZTOl2M+HIFESLzzErbvG
4mEAXzjhkUTCHICkgj3j+W2HnAuwR62a0XgsuZ2WdUy1oj04uLF4mRpeAJUHQX/C
ouDz05Tl7JuQdIh198obLFS2ogY6KQwEk9/gfsSMeW/sb6bRpsyj4CH2UdI6ZWs2
aBcAuasBo59pl1jXu5j4l0Tjwp/wLSTyGCZi07QWJxj0zjT5pXANxPfOUUa4Ise6
1QQSlfXvt17etDjRlRGHkEbnwUC+9AiEuCQo5yg3SSs26DzEDJUqqtuU4kSNQQl4
IRfnwzpzYWylYlen91mdQV57CH7HQ4ALvFlbGlsN/ViAvBQkuTPV5p0cKvOqG8HF
iEJ9RJInLrobdcn6jjDyVG2CXvqMdXWUrSaf92/89ZISc7ZNArc0RwZivdyZIf+k
3B7FJsiurH7aQwu+DnOqrxuh+IX/VU2azbXv2qbRZtz6kQF7DOd6TQf2Rm/DkAE6
MsEnScg7yNTcLWETitigemsg8q+qdfCS1g5CQufYZBXIOrzs8n26TkOtanzL/X2p
xvoeaFUe4ZRaf0dqHkyacc9RKUgH2po3jyNQ0amPy2gaWfoW9l4UNCbt5q8c6qDn
eH6BT2/y23yJKgMkhCGcK77RBPIycmW5LBNLuHmmYEjBhX/b8/T7efKytBKwTsii
DfmvFKswp/BtqVrUy2Cq9wUSyq9tlYhl27O9w/oK84h0156XdWl2QhcJp02hVZB4
NDDcc7N9LPkzwJYvqi5DaSAar4VKqjoGEMYqffzMmRfKzApUEU0yIzShzd90j+kW
gA7R1XrnrRYj2WuJou2SP1kyiQdz0bxuhkSM4VXasGQJV5uyKQMTWanvf30MR/H5
I8Mq9RyozGUDiudBQKB2EVJtZltW6epFOFt+I/Hp6ZmVDniCPoeLy68zk0LGLDJC
hN1KcaFh8rcUT3apo80T5u4vGclS9Nkuv9Lj5efE+VNH8NDsCiKYjEufBfVanJnp
PXgKX/JxR4xBd5rE0n2Gjx+tvMOQOQ94hZ6Vl0JfN+ja0eSTV4KcMFLDcVXpRQqA
uVo7k2mTeBswzr72q/9QzeyZBobyo+yeLwK4v2m0goGxlPJ4QUOs//eyJ6/QBtD7
gMU0DjPheBlV3a3PnvKNIUDVBj0ALokNMS6nxk1Zg6qtcGSLC/IqjIf0WuYcQmHj
r7OkeFI/4AY+muC7iK/4AWzXyuu4dpGpDatt3NN2WdH18vqt1N+o/m4Hu/PsbT0E
noAQ63aJv7bRxIzIMy16GcqCmwEoJHE1Q+pgT7HevSq5Tuoq+MVWoaCt65Q8Mc1l
hHZCvtE/3T0pPiGdGYnPzwBRVSOYQSlECCWBx6gD2mALzvq7A2jjAuocEU03ayMC
F7XCQFw9Ldhq3SUvwU0xbB7tPZDuTvisvmGR0YxY1qfucFfiy6E5Qe7Cn1SSffl4
wZ/Rva3CRulCgHAQCIaZIHAA4vs/lAInSjBkYHYG2hwqyf5dntl9fwdEHPw92HAt
crhoxz7yLas7OtCiUmy0JCTpFMA+Kom7d2ggXVee/cGhEkZftTRpnh5UgKkHQzAV
hu3BekrvJlFm5hquCvocoYrOW4HAsLUrRBgkRERT7fkUedxfvvEXHJjimKRewvTp
Sj9d5olLTPPsga3RwFvw3UJFsRE/qGtYqVHjLRsbpYTlyltqKdErSVGHkZfd6vWq
+VTGUwF3l145TEU6PKoakZktT6/GQkQjFYFzuxGdyK5dOqSXQQmNXrE9QrZTkTB0
3N3OJDQfqJkIDgxTjH1Ia11yVOi2rG9EZrs6d+SxjA5V/E0H2KKTvYjqQ3rrusEf
OgNky9catlbgFsv0rlcl8XzgE1si9N6hhVA1vY9GQG86G6qcMvGOjbtOLXl7YCoz
hKx/T+eGlR2QpRrdrYqsEqZB2hwFPxmscS/c1aoVuVzdScN17pGPqXegUt1WYAWv
8uzHD+5PtTlU9VAqQ9ThW2gEl+KTvt1Adpn7Crsj9nwUx2trQ4gRfbeKdisdC4uC
hTsJhaOOVvDQrBRs/ftS7GXUoxaojBKiqTDp73k5wUfjgXtESRkcgjNRWm0Ht/1F
g0zBRLjrq0ElD16BwMe0dZcXl1kpSP8G/51QswQblj/sPYbbq6Rwbi8ew/ZFouhd
hUKr/QN7Yam/WUi+/7wL7lzy1qf8tjnPgwQSt77tJqojxOMwtLkUD9bxj+4tiwpp
mpwrqDsc/fwycUUioKpcS1Amx6mONuhL2jffd4GLeVZpRS2nqzpgBKMhL1UUfRmu
7GWMxL4ABaz+4AkTgE9/L87vnRHwYI21BNJbfKOW4M25JB/VLDvfmkfVVZ/dgAjr
fXTfSVXjet9JUhqwyvaAVI3wjl0fVytNyqmTRjx6yzvUF9+hO3Zl1OZS3cFlNfst
xT71pDzODGvQwZ8iPiGQatkgZTjApl04QDGHC7y/88nCS0n1Ecjix61dVEhTow9Z
aPeSNK66T6IhTZgOjlL4HVZzGg6SsYnKScmDPAN83rou5TxYNofYeBFr7ZYgYefS
fU8efW3BzNI73JX5r93gTYrK3B9TleGt82gbhANLgl/QrK6dwUdDfp/s44G9HF0R
wwJ7Ju9JF199YVetafKpM+VbeNKxNpakCYbmW04dohxUPq5rZx8EEixTBa8TjRGC
OWqTXLE5rlUfsvf346BRYOaBfj4dji0KzUM0JAponIazpCJ2uBIHRy3Gv+59klSC
LMscof9eXe/P6IQifcPkc7xujbUT9GNqFrrj0fqPro9Naom52VWHfLEcDSWImrgu
ofCzGS17O8tpiJVfWvF5RILfv5TRlmlBR5dx8b/7SfOAY33Z/zObur82Hw9x1o9E
BSF7rl6CmlmT94/lgCszzVvb9RKEQUtlaSJkgtnKcfITqb9VcrzdXPOMkwtqqq9s
b73UhRHIEiSxiPyyqOb22NAFuYcQ0zmr59nCey8GjnE8NXZ8fDKWejasJltIaOAn
2iSfzbdEWruRbYXyijy2xkltUKIFnM9Yt41ZDChdLcjzqlPBsZ3H/8BIvnzy59c9
0Ul4rYRCtKGMkeA0bvrrkn1TeNPEfDldVwr+Ia9ovR5XFLkrQbvdJK1CvlIxSJbs
JbSFIrmlsKbrkSDI2AyX2A/DhiFTOeFqPqdV9Vwu3P4INicv6XqkqPnXtQpfV93Z
fUpweAqyx9HtVzpcl0qKP6Z9CSpXTAXUTb6maabAnrPeRRNuQGi5tLCVuWrgF4ha
gkQp2sYfyqXx4YWaYHphXUjK0xickO0/+9J+frGYtQ+5WJd8krEIrXR+XCXQ9WKc
HWR65n/2uKBa7EbDAgrTgbY2hmk1Ivj8Ti37MIcWFGmRY3ICs2+s39tCT/I+qdur
6r/lb+Dag6fyt4JHLh/bEC0UwKc97TNw+M7QtOfUbqcyJMYZ5FHiA9UiEqC/NGYJ
u7wMiQklcyX+TY57fIQQMNNYIphjDo2uPDE/zIOr5ltuTC725csXUfCdsyPNTTXf
QNaWB/xLQMEx+TXLIijYwpc0VD6kFOy3WxCHkq1JbJZxBgoRPjjQRz9lUeTt88yp
xhsQQq4DhcHRIZVOCrmrDYW9TWMnMcxpjXyCrA1/m1wnqBzXcX+Ztqsu8UbzmU8D
oI8LtHzpZN4GS5sujvGl1adDcW18Xq3JZylJnbz4ASuB1Wbuc5N3vKnIxoSmVmnN
hDPLiuxE7H0rpxufYVxmPnG4HulqQWO2fSe8cL67LSdeMIVzMvgIg+NbUO6dcKB+
k7i+F/ksA2SRCeUMCeSe7lFeHAQGxC4wU3/eB4fxQnZ2TUOJ3wSLQxgRHUI/gNtm
uz/odmZo/GY9f2vrAD6wYj4GFf7T1CNQvBKQJsRKZowdOoNqSvf+v02FStEYDkYO
Y3JUiYt3KC054pm4e0Wp9PSBQRSivlyJDgU4M+IFzHS5oCOMEeUGVQ4Y6OoVEtRD
P6uqLPLndYwJ4OBSqwTVl/Gh0rwYhICtNjJ+1iAMYVxd9TCMyV6Dsw8+qy6GfVyV
TB0ICPLj3jSGyamPYBV2KAML08U3gjJbla+mtkmBliQ5fuwZIKQrlqXneaM/BKdT
3thNBTM7u7zc5MIVkhkgF+tEST3YfGOADPExmS7ZtHO//q4JBoy3KCj55eta7w2Y
7FOKG3RdUccUOzvl6cQxnPT8gynlEvriQ7Ve44P8ZxkhjcLrGbMEBbBr7S2gHEzd
XVmG9mK5OXIYuC9LncrLeaxkZFMaEECPJIzwIPCGiHLhfg83qu9BhmjCDLvUIvNL
Q5nc3J4V4mLF0VSNrQ0RMqEcbXRUQXDXxpgKzZlEszCnfLj4NmSTYlv8bru+9UDd
X7ea8OgEiUVMkV+3Z7XxZzgZoY9IgXvLLGllx23v1SABTI2Wr57zgIBX+12m0yDR
wRq9AM6wsJWeTf1nDg/guS9qGchZV6kPnzlTZnxSt89jHEUk+iz8ZGjMKSZw0XIt
SEqSExpB6MOgb0LNsJ7ckGUtk2KvnU4bcnaxu6LC3KKu3shRapFSbdjpqrj8ojMg
EjKNvGMpXhXQqMf+Hpx/IIEN6bznckFEar7LO2hzDBt+0yJNK/GO4vXd0IrcwEDI
wS/6OqsEz27eujo1eUmemZKOEiH9Q74iBEggsWLYZstPP5YrXMRVabl3RyckXVyE
f3SaK7GtlyCP1pYoaLEhb0hPKrFisqE6jocTE4G+1SzDx5QnTj1dhJ26Xj77fNWj
limVZi/seh3KgOpoQ0BqiLjtFXW4BzJumPUdEmQ6CPF++mQFeDXi/4x2uIGBN9/a
GzrVhEbq2fTGJWxZT3mmQCNIxKwrXKdPf/5jpI3l1eXj0Pt/7mH6y+gsnLrBf415
ps6JItYSrI7d82Pv4rMVQy9DyXgdbE3Ze063bjENq615tRUd3el46vZUQ+3zM5A0
4iV2ELbtHA5HiJoq90ye1pAc/ScjmINy4gu4hVksBrvZgGVTF4vz6tE8+XTsgLiq
gAWbGZdY3dHFyLFyB5Nn8N3y7fd6EQLbWCDZ2TIwwNtM3BBsr99/H4uu4piUhP7q
xdxGZ+DRC8OZ3miF83mWP3pRjC/cXfnxAbwT4E17q3I8YoGbZ8Cr1yinUsD7aKlW
1LJIr4KuKebJPmv6ztP8CzkOJwov6DtcYk07FXxyr/jz6AyiuXRZ0P1n3T4wTfrV
ZoRoSvRy2GRWz2aQGcAe97e2qNVbME6npn5ClzclDI5Ve9lImcXzm2RlDYpqbliQ
bg4UyZy2XD5sIZS+TYx0ScAisY0VgVfmMYmUnHLP6K5VwaBG7HCLkQW0PDiXTRG7
AH9pKn2LFZ36s+EnPVaRNTiwEr2ZY1aL4J9Aw/xxA13kOSaqBRwDm0F0dvmSdnOC
yp5M1b1s3EDw6ZG+wE0jS4U5RWt6SrSY9ivTDeozMLydLeb2RnHFYAko6SYf0+nH
Xytp/L3cphF6smaaESYb2DtoM4typ5E1Y4ytvlnZo7zbD2Mu3RfWl62KSkmHfiev
hhNcRlkZjSzZPiiyahua+HKnHcVAn4bV9fryYzxg5R3cSXpr22dUFRaAM+PuHMyi
/0XJcF9N3B+2TBieU1AOdEpXPoR1uXFWOMC2cauHDXbRgmYNE1hUUjLk+PQUfxR0
ZdIJfN3mVKprSR4b80lZDpqg1dPGvA6f1WO28AL4BQQKjxF3NuFYE2pbhwPdYDfm
nXLVEexTNrvq9QhMo3krRwVBF1aaxn1WDfZ097MJmKABvwCR52ftUvYUNncLq3k6
f2RWztUqT0OY0AAGwfkdM1WUgTZoqM95p3wse0daxk3grLQWJjpSzEJ11oq+Iz3j
SiaZgMCNaJM0lDfTyWZxANi8yCStVKBrSGmIwNalP4NkFA1frlzQrX9DWUSapT6F
L+2Cgbc041ldwCV5sEl9/Nl3HB9TDybrd/CeAd9+hk/h0CiRGMUS7y/op32IP9UH
0CvYpfnlg5vs8kuROIH2/V2Mx/O10VmhXZiORdd7MGpn/jUrRWaUg2NYOXO4tIgd
7Xe4pLltLwcLIeWnlxMdKeKsl4KtpDImqE1gq9fBGgxraTziBZY0x0sWSP3m2OqK
n8Kd9yw1l4RIBIGJN1vQB3aWMMIN57ISot1hj6ppChrYFvQPSln/xbBNpTvIWAlI
JReHTr2Ikybbo810rMGogaU5UoePhYp4X2NMcLJXvkbYikloV4mMxE+/Ue7W4Gor
WcEjZXMqAHknbNY6XqXInlxiP9UQUoYtM4ydAsxvxZwzS6ebYgfc3CXJwL9zunHm
QDgQJn2wIjE4jgxugQZGEV2uhuO5H0o7gRmy5mlXGjxe0D1kymXBji53RpjDDCoX
SVU9Tb69VNSyyxm+dmWYH4Eik1yKwh/KDHmK1jIqmKwhXOWeHgrafyyH90y6JGp4
KqM6G2JxK9HrU0W8ZZUznRFaVqqZV+eccNnYCzuuyd0F+fr2DC4Bba5369aeg1gg
Da1PPoZZ3uR2VEYfNfWkeBIE4Rrw/I2dg4YvWp2pxOiW49otjHxJVicdvovmZXUO
XCIDZDlfId3TA32YqzcuG2ZS387lGkB2hpXohfApQLTA0LFylVKjJlg9Jd9+O5kH
foO/4x5VLrPud2JbYK36/0EttiW2aJZxW+/d2Y2khvIx5gs0r/robn6IR9AJwhZd
JmRJcr5QXC1YBvoekiVBc6cFJ1D84aZXx3I2sdIdLSecpQi2hdxO7oKZ4RFIuNA3
PHS20NKp2a/xes8h3PCeFTB5aamgMjEspI0PLccyQA8zyhn3tbRxDrTaSlKvEj4n
JjG8sLMMQhYm86O8jpnEKx07wdOaDbuGeWqJlOwg16aNx52QnnHAXckFfvVU7oO8
QedjCYl0BYQHkUVfE7FTO0THzdpbr0B6vQUmqbfj/8TPc8nu5jSkrmaL8iCVWwsZ
oLXt/kzOlVrGKh6UkiUpbj/1s/aFp6d0nKOKS4mxY+kL3Um740RX5qVx7En8XaBW
hkHwO+kieLTFhn/hQl99EluLCFpx9NiZVGS3Ta1CB4YaoZbaIZbh3BggMTWN2zHu
18HviWS+WAS71Ajuah8o1Aul7LB6Io3KDHQJqRIGv9xzKGROX7YxzJadeFe4InqT
Ub3AI2ZO3ChJbmdaIb0lDAhLZiv0Y80JBrlMEZoe/toriWXhZAiJBWrWjJE3Z8nz
CiCqkzOsHMRRt9meZ3OXmI7BRNu55K8I/PqvYeK5JEw2QRsShA6zdM4ITwhPOtmm
ObIp5IMPk0cbx0Uvw/f5khWtXF5HD1h7h218vspMy4vYEaCutnYz6REhYANPmxoh
vDBs/oZNPP5gCvT+gkRsZnYbvU/Qt34FYoDDCvt5poutKR+b2kklgIUhIonCZG4o
YTJfdoCiv4zkmhjm1cagd0hJymGrpLRwwnJUWrbJhBmIftyQHaGmgJe/0DwKd96r
NHsMd50SPZJlIY2+lK24yrdotvBGBpmapn7mF6kNqtvDYCAx5+BHm1oi57bX+xA4
IfmERcergtUN/9qJQiLR601DBtdPZ2NnK/GV47/kSkkSp00WSERK9DKkamJmse6Y
Af0NYZq85sbIgWh40VnBBHpjwV9DfRmxgqUcZD8dZz8dR7x0F1m1/bI2CZ1vFJ+e
eKVjS8x6DdaOHkwCutv6F+u6jJmyj/QpDK+UVPtRF2PZzpV36bvCKQ/tADi0jaJN
Tx3D46cm8QjU0zCHnond2Az4eD+DIb0zl2ljeR6AKu4g5d/iuOrDU7SMzzfsAyaJ
2r4XwQZgxXUGt0xKQmXW1ikSVhzd02HhSKBVDdQuEooPkJgt7AKDBi7yD4KQsvjG
BLy0DhmgQfGi5pIB/3jNyhGY1+OuG6KJvAHkkbuJLrvwz56S6/jQq4ZdJYnOPoSy
DF0Sa9KpTaqJaH9ZN7V71tgNlB2LyaDeBdqKjIB4Ztxd+r1kqWSSwRmoU18qpv4s
C8uO+ByXdjP4BNKKaObIH3QeRwB9hmm87sKaNNCoDxvpPiA4njoUh2S8QUnPj9aP
Li+uVVkv1SRohRzru2qQBeIbobyxpcA+iT+dN5krBtMfsIHT6B3NrP9hnUEzAOVq
WeHopVqW1kg/02ZXZJWiHaU2v8Bc0REljZobfQ32g+ImcmVLAGtqpnZaS+tARYEH
ePz2En07mCbQ7dB/LQPNVfkGBWgfJkXtRD0udybqsQaNAgTIgVP2i6ZoOkZh7AT2
wlktFbiIYVtdNX5PzRYf9pOtmT1dk22pNg63s7zI4cWB+VL0lRApD7ugkrYhq02U
TAw19dx/1sWVadCGd/l57zNA92rAjDrbVzACHNEqhbhVJ1eUtewUrCOC+1XL51Yx
Edej2VMTsS1ooho+rDWDGb030Utbl6Y5pQKeu1JEkGbAw3GYfeW4C4zTq8Y0cBR0
8kY++qwNM1GBI8u180EqGctdvDlAFFUNPFxWHo/qcn9K3edJGA5jKDhDcdZmrUlS
9y4KknYZtdI0DuxHQHYerV/L6iyU/LGjo85A2wRE2P4=
`protect END_PROTECTED
