`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZLJ1AsQPAHAQsKHVbgpGP+Tl+SD8znYFoa+91NdFmuqWRdapefi6OYNVEDjjHCdX
t9euB/7J9Hi9E2igHQS6C1ijM/igMCn6m5tOYMMtbLSOD+P6K3jS/RonhOI5EoVV
e7FxowIr9q6ZGNoaKB++lDErYRCHk/YBH/4B6iBfT6TEXSB7lzVSK5L1ogeP4WpQ
2NaLD9kp7x04oICUpnVv65wPZtFOT29799ZQVJ3Lm0HpTFiU9N39+N2Eo5lVr76X
KtdgYPwEUiwnTzrw4kpwIVdWEKro4/1Z2JQBiG+RrbO/nqjpj8wCEpfbCOM1al61
M2ajk6r9cC7+R3gO7CaAFhuyYz973RHjnSorvmRcMLrvBS4kuGIgxr1q3yTLP8zN
yhhiWMZqFHs9VlXwuUTUh+0lbD9QcpIWeEHn6RnjkD9dWO/X43FNIxu/9tO2HU4u
4qeiD71k3S1LgfOVr72riWOJCj/HbCxM7Uu2/v+S7TQU8XPScsh1IvRg59P7Xk4y
`protect END_PROTECTED
