`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6JFaw+stbKsUlr9ZFMYCMw6uz6sWmT/nU2cdfaCtePEpLAeLHSzKlVUXqt9SKuWu
47BiAiDiBhzg3FDw4EzGTj9VaIdM3HCOM8PQ+HWDgwZO/GHKkPeqZWlnAbqsrWhb
zeQs1a+AkrKuPt2SApt5QzwI+6yoi26iMXD4WwXlBjJ74+pY42AC4WjXMkNlcUPa
raD/k2YmbIiXRvFpKunkIKaxlOORx1V0yw4snWdJeOox0e2ERzNBNNctwmk4RP5u
c5thzGpvTA4LKYa/PNLr9tgPGi7lZ3ItkUoTIm2SDv8h1BTXExvojHg5SGKBHqOp
qyAFpH1b8JA1RM1kfO4UZumJV4E4IVv445ppXgj1d9ys1OxPqYU80QFgnL7M/oko
Kv3u2FRP4frkzog5jdqsYJ/x02l4XbnsAtcJ6T+1HLhakb2zZnQVE6YAZxLqi37w
`protect END_PROTECTED
