`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rgbQmbfuJTPohLclcqhzH7+SAMOwiIroglI92A3AER8lAF16TA8C1EoIyWaYyb1g
F+ZZYwp49mEv/2+u9zUx19LO1b3mVAMMInJPaqBf1u1JAnxc7MaDLKEfx+ryBUAo
Glh7W9amqp2p/SAThn1rO3bblap9+FhD2KfAN3c/T6G6vchNfS8/TPRNnOiPsxe+
CTY2696ythpVLww92K4/sjK2Kb8zqCoG3E9Seq7uUF2VG+fttAsoRSGpBCvfIY26
+h287PFGJjhz4/v0y2Zl6LPedkgdcaQShMZtn7MUkbabeE/3KqZsvrfBf4uO2L1X
n/9IGVh8jykYEZJ6T4zGLpgg0H8HCaYcCM+Rg7u7audXCSlz2SzBet2APhVF+d/h
tazbxff0o0NAQ6S+0gnRmxE7xguJNMeLiG4NpEiPy1Gq++nzXGGjOnkjoeWerU8F
hC9CE3KC/YIOMQFtgUEHf/IQ3kNtNcgs5MH6qDuIggiSY+ztWRuy04yyoVausaSB
RaMEmWudvhjj53fBNDx+bGTNIWzSwYSpTUCszFDwfbe7dnWe0aEawjEcOhSKo7Ec
egjcfz3P8dv1SpoZYtHrXK7jW0nUKi88aadOYLk14jp5MTKt8+tgJfJzXQS7fQoa
S+jwX51wgMRtxZt64oUtfK7wB0LFyDKR7f8nQMl5kLxG+uDOiQvvowiu1ZpUv2F3
JJQ/5/Y23853qEZKD8yVY2XZcTEnpvYDB11D4eYPBqo=
`protect END_PROTECTED
