`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Im0Nr3quVJWU5bfefPxJ2E5dcpokM52o6EcznF9TF2aF2SDeH/JJM/5uMzBqJ4G
vi7CSn2PJHpCWbtYh418hKTguSEVYmMzj0Fj/igFHXI8JuNyX5l1O0ktZLX5VY1a
cNK6oxM3rfT4i9y0EegKjaqrCyS0Zxm7GmEMb8p5Voauog+3lIkxWsw6NvIWzarh
7BnIVrNJyTXfW/zsogj0yn/1g53K1i8OAcSNnU63Zha8D8WtgmOZ4M6zaR45UKC5
ZSIL1NEZc2eeoHinFdCAcxt95NsrQA2lQ4bEhDBh8KguicVdBzHzRNqxEWBW486N
`protect END_PROTECTED
