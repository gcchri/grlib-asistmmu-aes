`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2SqAhLPy8otwrHQvBlPcyaLmf7j12gZzv1Btz8kObKj1JfbiGPmRlPK11fV1iGJp
2/Zw48jDogvB0tvic/S1shEAJnGvV21zxDd6FAXGayF+FI3p0vRJjwyFIyA4Asn5
M4yc0NWeCUzZNONYTWxLMgDqwvFzc0Qx+aBeSqcNIsZdNlU2HtzbGfQubSQXwJyT
F25WwdrqQriPTerIvtbIj7vM9bUPfhdMchPPh9NtqPpNHlJK6rtLYeDb0uaY6lLs
6MLGfbN7lel2ORYNg44A4VuF6iP5PrPadun84Nru93JR7pKnAw4l4SbMiCZ7+zxk
hZSFT5p0hQbokiWGtFUOyVDDRL/eaMgdB+2av5q+P7Rvdfl5XjcBM8ywr+n0qIVz
grLPvwOmyWjKFcctG0U0JCC376ST1fHtfLe7ZoBXd0Zib2hHVHMwP4D+6yukexQB
gaY+lRpPULcKokrk8O8FKd0CbQaC3zEBH74nnjSMO72UB1LYO0aGS4TkCRwl3oBJ
3/zEL6siDDGz0x5Tx5lX3nxWHOladUxUN+LzMn2vL+A4bc4BvboNGAmnCzrZD5sk
WiRhBnBEbPMzKXd0NucZI6L7GrlSW3owtrLhiIUCgXahSF9diCFtvNVBMksKczOU
`protect END_PROTECTED
