`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CIz4PVKdgIehbzqnbkGwQ4lwvlwOEMuhGoialIFMWsvZSL9fhlqTvbgn5QLcl5Wm
UkoWVLgyOYPix+3GRcVvmszAkuL08erZ4v/qoAK3UxW9xlDhIwFPcBKOA3TDwc6u
urE2Y5W8Vh6iDNXAfVrFJszci4uoGIOleJJiStK3zBapJnD17CHiodVbnOGP5Xut
EUTgKOJe/jf0LLt7dmi1RXua/qAZC2qufofsGr3yCT3BC+7Jg+vtS3Jxag93Wf14
5SkaHBfzJ7wsoLQjGTotug==
`protect END_PROTECTED
