`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7zpn4ufg/vQgndWevJM0HXy6l2uwlQ7/C23mVHb0LlbgGstqOJ2raghk9ofVpkUy
ms1r9lCHLQl/ZOc7NviR5pXo1425HbI73jyC5N9v08kXgO+AWJNtCp8htQpoUrkJ
U5OmToRzCDNtj+tC4jQSPVQ1/4HCzx3O7rJpvbg6kuEd838xh8qG3Nbkm97bJbGB
Q41IBGWmRljBzWLth9Hirc0rux065ehCyTarIEXGVUFNl4TUfAqpQpYF+8S81o5o
6ezzuiMcUyRtWQdXadlasPnnxAjYF7gE442FJd4YedMYXJhQ5HoONYYrGK+eUZ5p
sveXKAP1s167PeCLFlIzwHGGvdSLNyRY6lUdrBcXtb15VMLPipkH93XDeSdX4Kwu
EaSifVRXCLCxXrZcxvvWsmKS5bVTokaskAlhOqXW5Hp4RLFsnDJx2k6jFuPTa/Vn
oUFqCbzg620OX31PY8ujh3uaSZUTihAN2edjYwVPL9un5YthureyrQvGzGagDf9Z
VnfwWK3viYjl4TxtxbknCHG36Fqj8svV/a/r+XwqExzb0BTeUkoMulJR/cd+IyAR
hXFrAvwesj/gd2VLfSsVC9nFOpHCPsn2siIswJvX2JcrOzV3ErCQyfHGimZ1Nufi
`protect END_PROTECTED
