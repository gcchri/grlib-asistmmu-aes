`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RZIfgDfjtUVNpOf9e7u/f/a9k/qGCxkUxjK4mxddxzjFlpCmjDtxwftdB61XN+Rq
H3d1q0hNlhRgF5nG0LERD0rehL8bo6xYW4HOzD4Srb6rQPV3csWF969oCrNLdrKF
06K6tDGI1B8M3JFzIVjRc8ZsI9VoDkBvKBG6CoJC+2stzyt5VG8kxJvgLVs0yPOq
G1cj2wipWaLRSn0SfWpoG4t3iwV97Y4gbRnAKwe4ZXWXAJAwxnb6MW9nOBVfGcQF
L51o0dUc3Jzy0wv7wfq0fg==
`protect END_PROTECTED
