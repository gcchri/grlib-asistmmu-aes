`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tzGeiWIIbBfTEnaP/NtbADG2ePBn7jiEv5/Jx04527HdVYRPR5eD7d3vq24SjJnL
pXyAKdI30Reup1H7We3qcwSgjxDO9s9LhDDqxHwDo3J5DHkhgVAaXMLZMk3Re74O
EyZRVzzR6baK5F0ZLDroV8tH68N39uqtB41xpcyVh8yCfvZ/boXUvplJNhDIOjcf
CHJsgI9w0xF8NGScNW8bSDNHzh4kOHvDgGRjeF5AqqNt+Vpt8pyQLJSiic+lCfNE
yRNyZNbAVAP3OIm8M05V+M6/I6BpZWOebRd3sLVeZeiYxYHPrhvIMZmDroSn8Inl
v4qg/EyKda8Sl9vpktTMuWiMcXgj6rc6SZz8vst8CKZUSOBvioRbZ2uCwphARiem
5sIXWR1vB2R0s/7r0esoPi+T/79+RZFoPz7Ps6kIsMY0JT90EDLaS48LClQrOvQj
8rvpnMCBvsc6BCpZt3ovp7EWRXaTU/+5R6Tn6O+1DCesgzDA3x3mIRum/QciCuAv
dHE/SLmzjrAHAujTOlkoL1jpjl8MjXlkiqT+nsFtfRoHpO9osWIOwLrnecbBA7HF
RlFljj30oNaOlDdhkN+2YQ==
`protect END_PROTECTED
