`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KYZ3EcPjQpau10PrkaiO91LqRilPlcNQMKoFLJeO9RnEwkIizLBdR/bXBi3BJFGk
U/Y9FHJdJPyBHxRHHaHooiJwpZoaFtkFoUsJ3NQrVjRdXJAf1rxESNpaUYY5U+CJ
zZ/+fVvoBehbTW7tn/pCYxFGkMdW3BDvpog0fmX5ZnIdi0c5tGzmHbE2MGJ8g2Cg
vwa9t9iuAw5F1MunpqdNn680KD1BwT5/yaHjnHlgyMgSgaoDyPdjNJMv7TxtBmj6
P0Bym44tBomfg3Bz31nL2ZBUhQK8vcoZ5pbmAYZ0UNxDLzBLT04qqCV6SlrHL/DP
u9ia/YblbqM6A/LQMUZt+fyW80wv9CKqgnqjxi8wOqtrWv3l5YaEdzlN1so9k/bw
pudnc52yCvoYmp571EdbK+93TOyrw0Ruv3wSQEK9/yo=
`protect END_PROTECTED
