`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wACN9dzRX/4fnzt0RamycigtJ+Xon/ewecq6jNxA0nqRCIBhzVQ1MxDIKijCnbvS
zjpO679IkA/Me9FhoVj9/CMKBrEMr8Ux455TI4gAn2+t5zwoN6twSRVUUJtZurxF
ja4zjqMBFWpEV1Ljv2gH0aCvkoZ0FY6hB6Npr29ASZupo8ZoW6y0pwIDdoDeJSJR
EgbaiX+vSpIDyNYKeEOG44q5gFJPE07P8ynJULr3MqsZEmV5eKdvtzjImExwKxVR
gvEeWbkUYyU1XNxCfFtwQSOWUkwBUu5suOBM4pFXI1WdpG7QVIopeCywtWOY5m1B
/4U91s7xixnbXZXr1kdsLlpx8IYx1EaSn0gEFitIbSRmcRd1KB0Jn86hEw/bXTdH
njZOKd4LLktoJ0adFwmdeF/ajl6vk+iZxBD79kEy/FXHJg86DI796YCtxGuthJAT
AGkfpCo00eIGJsdNmNo4nFSljACDokoaXZN8k+Wd2uY+uE2uCBxZPaz98iVVeN3t
MVVEXBLJl5yzd2NVl5YBTsK9hyodPk6nbQYuORMSdML0t1mkdGwUX29xT2NXTwzh
VpJAddBZ8FMsVNmhVlZfGDtqt2jjZm3i+jY0hV7da6E=
`protect END_PROTECTED
