`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w2Q7DdXJPkqWnK+oiz3tEn2Fyy3b+uZy/hJQ5KOC6v2MAVDpR7mlpE2URUCoB2z1
gKKFXcnVVfHkmpfj+11LU833UGfH81KrE+oxlE8c4QvXReq44QJIKAhSjMekV5oW
9uYJS1XRs+aNzzh96W1lTqJ4kPT7vd5LqM6eoSCZvFIRjqaNtRVMymh+cvyvkBcs
A/4WstY4Bpvoyq7RVV2YV/OmprwJFBk0fdCygTAKzlKEksXqDlX/L2X/TFU3ivCu
3onU4wS1x6KScEh1hB2kIdf0+0n0ffTltqJ/TCKTFxrppK8futPPiSzW+wpS+JA4
NzWzu04FfMTYqFTqrGkd+kOShJnIlujt/ToQIn+gkcO7thM3t82R/o9zzWrMnqVe
WG2PV8dAJSEx1KWemHwjBQFMZ/ZDdDJn6C5Pj5fbU/g=
`protect END_PROTECTED
