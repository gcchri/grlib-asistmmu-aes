`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EAWBiX6BvlDV5Z+kqFyump99xkCUFObqVOZnITam09+4nsS47mvjNFvpoaye956q
tNz/g1rn/wWJH7QAqw3jzP3KkNAfsJRr1j6MFnTa16i6Po2Qsv2Hs9R3CPIjeN1c
nvgJfa/kq3OJUQwUCOvs5lE6mlz1cIvt/vzOlp+pQLFfG/Tv0em8/3k0/sh+ddDK
lTHbz9YiNp36YOSt0WU+a5PuMM2XWPwFp5mld2xIF8Vkbc5yyF3K2uEdD9ZViSyK
8uvTr5WkhpH8ZdCdgTvVx6XUR6q8Y5wVNFqGH8LIvOp9SOfptAcX6+puKYxCtMCO
G9lw1UFrUoCRg233JciZyJHA/vQijFYOM7mpSQRFdJXVgTAHE8teBvg5Jpq7h5G+
oTCceoAbGgHMDPKMvap4l4CuHFGZb6mH2XucO266A7GxPRKVAlTXNOFwikVGSDeQ
lc1+8yrTKHkeBi7IrYi55LeENLQU+3+E/tU+AMwsdiVgsAf4XEdqaXUV2+qLZovC
1JuJ+yaIdc44Lk0HnzZNuAaaK/AkJQRBVzhMInIlTqRu/TVCO7lFz9wtSXUloqho
jsBLcTnLw3u44mn5NiXGmUEgNbQBMaQE5KbkxI/9ddy2xFvlmNkCG2A8yx5+gb7F
xzFrbWr/nP0NXDynjwrJJ5QYSAW4rANsSSg9MAD/4wnfombNrCnVM2lltLpgEbNl
4HB/fQSwpAf/FLxQBbIX0hIiDUuvTVqLZH1aP/bf170dXyUeGKRGcnMpOoNsrNA9
G8RgHpL4t26KctkTYiqN9UAb02mYG6j9O+SjUCfw/FX4Q6TpWVqcAuZiy7kuxuy7
hdvyVByBDAZ40kvpVz1n7A==
`protect END_PROTECTED
