`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gCOTP0hoTR+BLtzCmhIvFkUNPHMo3pI6+d86FRDnQqSzpiKjmvPIrbpKrkIu86BY
tu3POE5x/AZf9HIGFNEu566b7LuuiHFVjVS0nblRAiGNaxy7dfo+ZBENogiccjOR
+XcfZ577KdbnYMid4EjIT2uMjUtU886Tj0zU99embQpJUlCGgj92I+aC/zYcj42/
mr1ghcqfHl4UuX722AVS0aHXP8RBrT7W+/JYl5a3j8n/xgDZfd42GWkVx07VMXzM
5HMwBbvgjb7+FISlrE/N0rtRGWruFxCKPgPr+j5WvGXzw0J9i5lUcT7eRDZNLOkh
Wc4p/Y7x7A1xJ6uDX463uetiUV1GHwuHdl6m3LOfemjHe3kg1Bpc7l/YC/ENnC/b
qyIerqgSD2Qx/DXen5SzPjPNgFnK16q5jQLml2zB2tFLzZVe+cLZ9krudagoXhia
PJhsF+baf3bFErIkANfK0pF/vUE6Q2ZgKZE5Moa0gi+QvfNly/dUggYVTfLLDV+J
FuaRnee8llZjdbUVBOXswSeycT/kCMkO9XM0sD3STM+MxyotDvOPMTI4vkby6IHD
ym2p8ps1tdbV8WvUf4+kZTmyoge7eceRyIqfFf80nmSQEvWgEAMekyl4ZU/HSm+N
c/YgVMuzCdmCb23yh7ek/Q==
`protect END_PROTECTED
