`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mEMFuyv7hMUSfgFQ6AtoRC2ba5x/Am0/FtuGv9d0yBpFmOQae4ssJlUky5gv96MC
mNubQIm8M/5exRkbBRMH0xSicBr/Qqou0aRljLIxDzDSWGikK9fRctwFcY2mU86q
3nklziNgCAUzaN0Ina94dXuezobEGr8kA2q+Cforr7EM4AQOa+DuORMWzx8NEjej
BcvSYaJxxYTv5EMDTDHNS6dLSXipvovf+/oi5/AVdPCuvex9IF3xMD3APIeIEW0Q
LPOBhXvCEIyiIl8FKCtff+nG4iQgzUPTowscsGkl4rtZ2w3Uc2GHIwEzhVsEVSkw
+8y6Ia4iiiEfWvsRATjipubaXMJLvnSIiznsXVfH9VotkkZLk8JlJ5mEicZfPAXD
8APZat2QDa59jXuwPAnJfeUKURSa6luyenvsc2njKIcnHRA6zNpfQGfUGNU/uAQm
lKqrUlCby6E9FY3DajE7s8FhuuhMyXnIFgTXarUtt/EcddFyCTykzaMYVT6YcoUa
lmmCel1SicgIbL7UOThdxFnRhkirQnqjs32V85pUbFHIEzMwO7sZ9MRdBgEqYEUt
`protect END_PROTECTED
