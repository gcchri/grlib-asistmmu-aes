`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I7Uu9vhk+h/Ze+rWsxkvIVL2TF15khgQGdOLQcK4g3O1c+qf4wQiVgtbRDuKjA3X
9gLi73Gtc1zL2OAUpt751gNj65Fo22XlUt7fXCjMJkd1yrhwkVt+I9pRjzzudgFc
LsrBh937LX/f6UaVWQgVJBFRqEAUz4sOhYDpjbM+aRgPiWHmfoPHSu0ugcner6VB
qbIus3RE5aAWnyT7yO/WsQqujRtUMRY/Ft6lxWOc0xelWc0MaYC2W4VdVqTOzLpC
tc8p1FrlRzO5+3DYWysvCayuxf/OaL0XwJ5L0JughBrbLbvqYVQUTMHrN4J8grtb
2xCD7/RMsUpu/GPTkHA7YH9DvDlFVRGHqikj477TeAWm4pLFrKiCJPMZImsdELdk
QdeK5rAZ4D5W1uAqtaoUhEt34au4jbGQ4M6C7BcqHgct1o8C+qF0x5ioQVgo5Pn6
iI4Z5b+Nxq1fPnhtvSjWI7vbvY1QEtyde1kzFQ9kTX1MeYIKD6mbEgyFR8bWxlIC
962LFE6YEMmuqiPxeK0quheGv/+5z+qpvl3D8oVaZdioPU6HkVy28HnC6UYTnq5P
eK5tVCOXXdN7j6614qOcIjOnCMcqlpP8gCX9tdfW2lv1j3FaIc7UUcnhG55zjEO3
BsDBh7onZvtd6NbpNS1zcpTH8F5Ihr1j8FpOH3E9oqZ041rFrEqHFVoTg8lFr9y8
Sn63+EbxoVASvHtpTcOcUzE6Jj6dGhl1pkkLehsnJBXZTU8UQ2suzO/sCMU9jnVG
hcd44Y/tDERv/RCTlNjmGQ==
`protect END_PROTECTED
