`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kM1L0bH+KeJm6hPxOe2IihSychPQ4Cpobojuhk3ouow8+cvTdwiav8KzPxJq5PRB
JNmODVc/QuLSgwPJJ4K3aulD0WQm2y4PqcHfQGUd/X6rQWg8vJpRHMtugH06HCHW
+K6Wr2hRy0+hZwMRZF1s8nm/t0rwZ1ImKQf53dWXONrdctTAMVzIdQIPvOSiFFSV
mgij5WH5Mnm19eHmXOs+tZC7wDZrxUj8e3/S0Ir65nqA24rltyf07Svz5BTMGNFj
9Zw02iV3cOdPLVD2RA/LkT0hvl7+PBJaOzk05Hl0JOYEwkyg2MgbGtdpTXU/xOkH
2ltR7nb1/Oe2roGMuNyWQ/QArEN2Bsb7xqhADvlpBROso/YvllxACMacZAdANrP1
EEEtbCheEDo+i9BEHBWpnhRDIwRSFdgybrm5D2BJ4feB4a7RjPFQIUya9kIX7gzk
ITh7LxshoqDOMG8boGayNDa1KD0hOvLxS3AgzvenicUyYKd13YHP8EharWEnkdLj
Y2W5GO/m3j+SwLZw6KqpT0fPT9C4tmlBYzCgP0RpD5q0hQsp0vnkfk8vBTLkAlOO
5/DDxkdzJwTskq7k3PB9pcz/Yq+97OeDYadBq/kEvBB9HgeOvOBx3skG4LyD+NW3
jE1mIUrIHFZGhh1Kd1JHeQp37A/DqXBLqd8bUH8afsIS6CtP1i0z22LW/b3tYrno
6U3uekglUoPLIa3olJd4T2dNZY5uIH2Ia5xCnvLFVnBlMWLNkm9bYWTbeByp+4sK
jTypQWMSmb4TtBrVgHhTow==
`protect END_PROTECTED
