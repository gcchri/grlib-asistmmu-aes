`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1t1BvjB35QgceAIDb3CsgOI9BJK/O2/ysS5v8VJpKgPOGlSn+aQAYWHUEo8Yu10M
wgyTJ2jhFFMIwF8K5lqAEnymOnnnqn0+ly4y3+bGrdnLzIhLLSs+xrb76vjLVpGk
bKG2YIj6NvFFdrqq/L68EphwwGq3nWK9w+wF96P57N028dJ5Q5z8OampQrfgxbRf
sF8H/DLaFrMPv5nHg5KrkenaK5m/npNGL5bnp31j9JUa5xgDcEQU4lC4MNW5Mk7W
JvXd+fLyW8Y0CFWfr3txoIBv2u/kALRmwb/P/r58HX98VYeLpusJ5dimL8MPCmi5
pK6TytM8SYsiShKdeqTvo8CPlijvjFC6BEDbnIQ+qUBslziAv0ICaXDuKVAYftoG
F9+hDw0hYXN0lAIMN5NVU5oPZaCeHkJfV7YHxvB6GlMyZd4/9e6UKc5znKEk1WuP
PgR8bjZMMEJZzCe4Qmf/LPiFIix0ROBjw9OW+7owSB0SKFb3y3T9CQufD9KnGzxx
Cg1gE17h8FvlpoIZR1usOE2BwDUKzik2ZAF0FlBmpGkdgByLxglwxj7ISf9Iok7Y
9ka+AnR6FncDpGuBPO0nt3hIkgPLV+NgA1KI/xMJPw/SN87F6u8Zl5zNIT2dm+MG
FdaU3dBFDWmeT9QcsoxbPsHNTPqKqaZF4QcERDtxqv1JgIuRZ6j2vHiV9VDQOcTQ
fm1W2p8/25pfeqJRnPULCHXeipSyflow62lfqjMTN/N3XWoyCgzcO/42ejAVpRYm
KIRGTXYwlawOdb0qE9M+vv1x5WfBTz8Uf483++keBdLbxgvSPISN0ble5tIvZVha
OB4p0CjX9oZpI88lkzohih/Kc18CyNYKIu/ibGPhNuMWvYGdZtcT0NVukR87EEp1
`protect END_PROTECTED
