`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FPPaggnD+uv+fOEvdXySAsHCgmx0f+Fk7V67az31v+PjcMHDCFKrxKZ1GU9yWelA
K1Zf16snphnWderED9yKckj3H+h9e3J7vLug7TGspcRMLir1PEbRmyYIs9DlCSZH
jeEWXiqQni/4TtI0oAbO7nsfo360PM15pp5C/iYqWRbV7IRQG88yGPwsw4CFPUct
x5mjYuL4hzG8a+4XPkF5qjNinJva0qhLbHoY0hNc3xh7a/BMfXIi8cDw5l335SuH
eJ8DVHrFWAtyPUcUK+gfXeEtVj+BjmhxwO0pdIDxPGpF59/cBzYp+gxlmYqdFM0C
Bhb7E/kw9/4Km5oEKGIABciJEozY79uXeXEMl/vWYYgwavk075T/eGfWEfL6f+hm
TVstjgyN88WLia2uaVJ4KlJCmRmfs2wSIwFNOpLkeMY=
`protect END_PROTECTED
