`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H07hKhA/gZ/RG8ZHwJco/tdFpAvS5+8nJOCD98T2fLp/F1FLYQG0zDN2Hk31fJjW
WnfFCXfC6boBeQWvyJgTrnc62VTUIitZl3AgcLOZ3c6zXJq+fZzoIT80TWFfxygN
cFL6Ckyd0GmqWRlF7LjZj1tv/mBUhAJo+j/HWoOBVzjb1YE09YcWPwW5FQbjkthO
dHioYXZIA83xUkVCOZryk5bEWoQ4vB6IAHPiHiZhzg7wj8wsOsCUh9ckgPT/bUx7
q0sro11/83pXCf7qI60U8RbVyFG/eO2zuNwKCwOhzQz0lE7woB9vzalwPY8fhmEY
yiQq5Sf8OqGISV6lmT814lSOQr5zBmzAPGCnvgyQqHh+FaIs3NQIkVEHezODJv2Y
oNXZ+Z67cs4UmJhp3bVd/AXu5u706LBaAEzHSUT7Ldt3HJ0npuPervT+YmuCiXns
iCG5KszsiqvoL67X+axAhNskN2ofbsHFHPHhp1aVdAGmKbPyZ8CzvjQLx+j7mZUD
BB5P1I8AMH33dBK6WfUHLiBb4KWzYB+tl+FZBn620uEBJyWSz5VxwWkzhEpbB2Fq
4+YQQfBnFBIg875qUueZdCHlPSXXvGmtODX14vDji8xFyeijwu6Gc9ataeeXGAxn
HKPsFPgQy0qeaJkGqqmvWYcebeHoEac6cyQ9iapDFA7X+s1ZbjF88L535A7CMta1
kpRLSc3E5/S0+VjENY+NIIqpGlzDDGTJ2t5t8GGHzZnOCrdH4KQE5CySRk2muyrw
LKQku7mkJbNhnvq02L4iODFvpTe8NeKSL/KeWgBqqMbPyBFjD41NrezP681LLNj6
UbWZzCruUlKmhdAhls03jy5xVAFK8N/+c7+ZMi35mhtDFmcP9LP4YmLqDK9FuRrd
9cRvt5UFnm6v+zt9tw9uL2gGlXKMnHHDYqnu+uXpJj9jUIyZU4OtvxfNmjU38+4e
HV8KbGe+U3PfT28eUCF2QjwokJB3jD6Zb2QMfANVo657Z7ve5miwMHeVfwAcQU0Z
wiZnUn0BUgekx0VdmoSywNs5dG1pXBKv0eG/PedFhgatn//OLloMtXNYcvrFAKZz
eUeNxFQbL01u9EI9koi5ORth7TGwpDwPZE67N5rPKxTEWQkY3MLHXXpMS75zOTlh
onn50NV4Sog/LbfuJvscHYtLvLxi3x015y+921tfwBK8uS1pj3fn1xdO0a5Jg8xd
4aGSOhJCe6I3+zLeGNgU6zKgiIsY+uLtZQFpRR9CfRc6cZy+F2rEs0c4A4m6Blqt
iABBAaeKVf7QRwBp3+jQcbAW7pYXuoQeKL8tZeTI1v8hv4J5l7uioW1Fvb+67nMd
9ZL+N4HixY3MVKhH98a9oxePNYEYDHMTDAjEQxw92tbxzOEVSWdq7/ChLkWjNpwo
LsEMTvdEeqxIqCIFXLl/cWZ3x9x1K6LpW/2LI0ifkydOxfXjbntNVzvXerA6Log4
kP8XbItt/1tTnG0PxMmcCfCwrLV5SNLr9qiJACoqhXPRW5HpvRTDZWc0eh0beqYo
jeJ5G3K4Zme7zQnh6/ql97r0NVrvdPc2LrT3DdFEeMkV+UyDQzmuFz5vIlxKbtpD
oRUDENXIsWfTG0iNSbU8/PENAxGNg3E4Hn6AFOfFACU8WoJe0g+r+O2Mu1vNioVD
9ZN+6u9pN2xa1BekxGILLheg5mgICu+bs6FOEfjeYsgRirA8dTCa1+p9mdrglNYj
ZY3UqT4HEyIcRMhkwSrUO/iAy+Adc6H4szWYHd7jwAE+q4jsJdYRA6GNEc1t8R6A
T/44481LffIfe7S+SY5gZjY08NREWHtARJp22laVT9A7SZG2c9n8HFYJTkZnHvwR
394nVraFEdEc0QfHI8WRRNf6lq95mESdXkkIXWI7FMrTBtvpwzRnzugizx4lO3gh
RaHO5PGTXs66W8TtLy/t6WAct1+k6cY+JMIeRPo461gpffhnmOcd3HC1DKyZlM2n
G+3GARa+wDYiwb1N2dHOgOtNOZe2hBcvWkUjLRSyafLFmNqEePqGqBPYp9Uj+BVQ
6iVftWFZHaziAv0TlgaPOAyk427VHcGfxo93Ly4EmXrFHNLjaJitK9j6QzmOTPxE
+lbgtW08LVbGSlpmgoNJ1iWig/VDy7V5lNITbbpPS0wus3pc575oL0h8aZ+4QrKW
NI/5M2n/Su5TFCufW0+6zZdXje5x4GLNENtAd5BbJYsq0ShOzeOU09W+JZIkxx8i
DTUGMpiW/GFCzh2hraAEH4J+DAbH4Zy6+/Sm/+hSHLcljvHw5/WXTGgfuWMVUDnf
cgFJ9iaYnZ5jqLuWkAGbWcZkLEodUkxsUTGnGQT+YXeNLhTPxpv3pBDgaNNsJ9SJ
bhY0MR/4lIGU3RaGUKlzyh6QDbkdEWxup2DV2xBECjQzTRpz3qXPDTvohtpi1dr+
zEK66JyNlZjU3IofvhLRwp4ulIZ6KY8qYjh++b4WIJQsK4rklinT7qWZDk6drwn+
UF0CHzZhne3CCEQ9hbu4A3LcT37cT0dOA7n4mfWeGl9+inRDhETZSrgsDOQwilBM
jyZxKS6fc8fuzPW1rTj2nxU8NxZmtgkkQ9V1Ph/gW/bTv5ctGtXDZ1R3KlXLU5/F
WCR5XMOSRXQs4t5VK4rCauM8DO5xM404M/YOawp0jVVikvXiK8wHeUGAWJ3GUWYf
PrGoVQa8UBEB0vT8pXvnHQ==
`protect END_PROTECTED
