`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9JV0Ax5qmIJnpcNAwpyyN8Xha1l06tkQZWqzPNwiqY5RyUZwzlXyEChRrrdLlraX
U9eWDYP9JpSRybDBbKWAT5HoGTAtBPIfOQPRWgzpe4NH2fl8xE4JOkRuv8qztAgG
vIThqn8eJkgXTUxVe9acvi7c04HqN4l+/7533FVMx9kpS/pjoXEryaJuWvpNX+R/
TzZCUzEbzGEnJeSwDtD6PepBXrcpfLuWEWI9i9ayNClqoe08yTqXwDDI0d688I1k
JeNRtVkiulDJQibudn0zTcViS3FpiiUi/u0xIPBPub4UcZYvPt/VpJ3gWAHstaES
dCdYEt8Sq5Pq4EKYtYSoNGnaEz4CMg+nW8Nx1tLnvCs=
`protect END_PROTECTED
