`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iqZH+uwbyTeV+F3a56SIhayksvWxaefJuXEq6MygZK1AH5i2c86d90PIgZeQ1nmJ
Z82V4YFatPIkMWN/mRUrk3r4n8sgUEMLCs7QE7XsTzuUGfXE0ulMRW1+V5G3CyQw
WYfMNsvWQSkU8j5Xhd3RbuTHLElkh1kiuOdqA/ZjOggsCzlzk7oxNAll/uCJLGx8
uT1SD7o405As7J4iwFqypNcYfjX7TgyW3J+iaRbq5wgerjDCRDtSd5wOxZ1GuIXM
L6+eoMUo0zTSUEkLUuemHTeZL1qhO3LCMc9gbM/1l8T0ydbD+2O2DuYqdDv5xuFv
ZYVMRAN6+qffQM73ra1LRRo8VKHntXRPs/7WOeN8Lhk54z37VXmSpW6XD1vjTVoQ
+wkPR3RoQ+U3UgGS+PaCl9wH8MxNCziAB5lq6cfjXltrXnujZOei71prxY/QQMTK
`protect END_PROTECTED
