`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pJZaeN73m9GaamCe08IOvpmqQkS/Eg54saEXKUQirS3E9VKfu0QUtF+ZsBVReFpy
jpgOSFyzZltVUuDUOOpvKY+YiwLKFMxwyxg2BylscXlaFSpnVS8lpXEEvdHKsRjR
mCzXd78i7IztR7sPGE3su0ElUWIapo2zPF+8Vp3QBqVnOusLgg4Dga4jCB2rFjAm
la/Q2yvmJHbjY8zaEpfnQrC+uHXt1KlkZ0XaIptwRPdjxqlYJpUmZiLdv8M1XS+c
cQkTOVhO5zCroNeWeXYoWnrYagd7VrN+kiU63RCzfcAVWU/HpKgHn7jdGnLvaPx7
FlmcrOQJbwkQakYjVXYOeA==
`protect END_PROTECTED
