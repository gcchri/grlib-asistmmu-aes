`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ot6ej2uElKfsT03rWZtln3f4EHGX8kicvXE2JPb1+8NT+7C2LqCYJEm0DVY8P8ON
6HC0DBEH3HZNrpkkFXKiqgAyc8xzPZ4TAmGp4w60IZTT9SWATc+AZKrRA3fVFQKe
qodpQ/n/iFOSi44phBy3QHtpKQxokB7rDkjkDDSUE5pF9l6uZAqvpAjN04KfsYQv
xDX/5xMiv37y8sjEIHPOQndb61KobH6RYXZWdNfYGmI+c5KElZcy2g6Y2hmwK1WO
CRrT87ERR0FImu0/+C2M5ujOjEJ52FmD0clP3ny08faHxCqHs78k9AjksChDIuAH
1OKdEZkBynvz2FE1ujyTPcD1VCzyOtTW7qonuelXBnbVZ8Zbu/60M66XTwzxnm9i
`protect END_PROTECTED
