`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GSj0rSjH6vNiGym8D21gtGhk4p92I9vTI9n4TUCIRqH6iDfcJsIyN4f9vO/9j3G/
UsIuJNe663hgB+5XHWK2mTwVitu4xIWvsutFZoLHqpG028Yguz79OkYiC30O+VKz
EDOOcpPyOyUiQw/Ew+T4/5I+ftxpe67xkeMW1RlMFtY+Lm3PfLPXt5QRV79Hzert
t9gN0lVDMRCBKZqVdEsNJP2cHybP0ObN5j1fDmbNiSWBCak1/rxYmy4SDER2eM6W
`protect END_PROTECTED
