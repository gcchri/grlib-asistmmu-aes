`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lD64+VTWD8X5t4s5vw6Wn+yGz4arljHgxh7orJwDxqnDqQ8g9p7GooQu+yiQ0VUg
g4mwvPpPhMeqmxR4mN5yox5ywFKD9O7q0+U2imGNUGl4N+p5dA+XR6OWbTf9372v
ILgeOpmwroBPwrPyRGYw2vagBiR6m3nvNY0jFupORUsBw9mhzNGPOtXg71v80SWE
dPT3HxsApqgTA7OyV0JB7zVJn+prhqWz+peoVGlVybNH34kMVwTXsvSOhqTsk2Oh
axk0F+UAWh92ErVZ1r6GVNWcmCiXPNaeKDvR0yWbMKOxneDWM7y77RQOEtbKPbdy
+WoYPVAtttw2xr70+8SagBv3ODPB4yG9FuheBF6/vI4G5Q2p3nOANaCjboq6ck+P
aOnjXPBL6nqGWwXJN+ve6MFdWz4sdPHtBhCgESc0diiiIzVlxJx69no4/1OpvNRH
14YcwybWXvDCANjFT2kiNrXpiQ/Fpt+7tJyLZH9lkidgeEko/NwOjnMzyLTmsbyf
tdsWuVs5hJK8dCBKhSOmK2kEn8BBc1RARurEXJ7qTHiYlih3NPxHd3GTr+6fg6In
cZaJbnaMmAOrB9hfrnKgHscIv8ws3/rMO6pdKAcclJ684iAtQ7FzGgTm9rcPj0ZF
+279mg0JG4Zn2olpdorjXMC8xA7yJURKKGWE9xaBy9zV969FKNn1wWJgNqEAxZ5q
CiRBrRr7aUAL/6HampieO5inqIChfVRsM2Wfdr9vlomTd969CNn9SweEvElxn+Dv
Mdicw92IofIgPPvynp5nytxRf1ELjpgye5dueelq8wbLwcP7q0/bLjNQGqeh9mVX
rZbzr3aq4lkd+pSuqXcS8HgOBTi5GG3LiCEKQOCjYY2x0bPHEJ93pS/hpxkxYI6n
otttA1L01R39ekDA9ZqTgKNd7TkEDNGJu/eZeOb8jO3lQvzt/+/xAfr+UA9RJeNu
4tfM7jCVuo/4YYpW/Cf/ciukL4GomFTvoEQVwq0xZtBYWOm5CB7+9+PF+tpHn4II
TLprItr3ETcQbKhsXgkCMY+5KK4PcDrdEI/3LscaXkftEsgcbvz7FJ1xcHgkYM8U
ZIjNisofAwnUSCERJA1aJIZk0SNjpmECIIi7nYGEzDZPorPmxle4TF3RdC/iXnP4
znm39SqxaywLrAZycYEsfj5JClkIa0RdpMClqCPuR09LhVva86hGgBxGB/wQ3Lme
5Ow0QhRVl7CRUu4oehtnNAArw8GSLG7GDp+zHZa+iAapXIABScoeZPAecvvfKIj1
IbLa137i2iEKC9PbNPLPmhnuDW2Sam/9oJKALR/4c1g6MB0yhoX5lXBXwJuhu2Zp
cjOiWbXpXkenk89w+hlTdRyNQdeqyn2zfjeb3TE91CruNXanJbeut/SizoxhMHbt
1Hprnv/Zk9Zexn1ONlYG7mvplz1O6bEBFrYcOFEMpYGwgh9akjnj74LL0V5pt0rs
rMSwYclpt7FQ5R9PTO3X7r9xP8xfH2i4xHX46kYK6RM5hdRnmLggwVmFSG9omREg
eUqXn2a4Thazm9P0xuyzDhS86jnCZDjxnixuGcRH6Rqfi0VA6MiRj8zyNiS44eCO
a2/BPF4mNCP0vVy7w3ge0Gox0WBhCLbj5bkU/qrhkylxLzFMFRtsPNRwL84QO8QD
lZ7f58q4aV9cC7wvA6AqrsnS+YcCHQ3uhBFLKsubkQy6z49OTTylLAT+C/xjNa+T
9R2Ri3ry9hoc5k7ySnSRE1sKXbDHzgV8EmDjL8mrbHNFO5RU7k463QqmcJQDq1NJ
xlPY+h1oZRWAYNeRAYGe/bVIkGCWu31x4P+y3neNCNAGqPH6IptUqoRU58WPA55w
QnqdayWXGlDJFnmHjOsewrgrWgPxRtDYo7FO8d40Iwc5o54GEqD3Hc4HEmV0LHqw
ZqExuc4RF3KA2EumopFRSfTe6fMMPdnn6F6ggEwnwvpu4DNmCXqvJgFEfDzkToDY
QAJTe919TCG421f76u521gDUFQORC84Ehtm7UYUFiyTA/b+273Gjl4ova9KHv8ic
ZdN6EbflKEsOpOYg9Zcpb5/jdd8n+abPA9EdJXFE6X94GJyFq5/TnZjuSSX2E8Ys
QS6zaFx2Jz/lWiGOzhtSod0NWO+s+bhTHwLqzdt+Riw2oPoHwMGdtaKlyf4VKsCg
lD+WXcr7Z5GsWvlJp+tD4mLAornmd25gNA4Sl9CxgzeldlW9SXP9FvAGWvIvtZyU
4LtIqzp1wCGQE6aLnfhiujCLSbzsHBq24DBXBDTgEOoxwUQO5TIo+lOqugyjS6MS
Kb+7c+5PDNG/t4HjjZNKWQ2Qz49CvBqjOt9X+M1aQxuDRFqg0Yk6wb+pMk4KQp+P
YatoQGTRH5jyjl25noI1WaIDAg9G2W/aYcSgQUIV2eXDQ5v929lOI06AgN8eZ25d
2IvI76W4AuAeCSZVYnUetLstpwo4cfGYWA8N9v2dY8FCxDd7OdiVPT54w+MsSlnF
jamDd2HxsellLgEQIM1lX1Hj0WyY176eZlF/Zd2yrBhvyQBjVymb8HfEosRN7ehf
oUXX3jQ2W8QrSvj4oR85faVdB+ntXim3EIQQ9AFEeIJCKhPLr+G1AOr67zWX0uxd
u4HAmN2o9k7mFmIeOqM3g//r506cqfMN5GNWa8unAyDngUWks5aXGudttUObyIfg
9M4xq+Xv+rnx/dQwj57etQbEz5RC8/mt/wM+eOn5x7xsrBD4OChCeMop/zTXcCTR
f38cpQ5S5Whyuxr5kAanr6ZwRYn5698ir+5AwNxROO1wLsX7534tZGvQLB0pDvgE
`protect END_PROTECTED
