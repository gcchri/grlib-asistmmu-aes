`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TApedMwHsQT51zu1wEV3plsuwzn4WamYGQxRu4Lj8HDW8uBl0WjPF1clXfSSMBME
jshypOmGGFqIeY/zl4EPJVSSQI8E8ZZ11KQpHqEf6wLz7s+df+NHap8+KTp7BmjO
Ckwx2uBXEaYUBLuROGRRy2azlOdR2bUpv+e7nvZj7mKjRbYaC+D4YYnYBi+SNEJW
jrj8K2YHnB7GMggVZJbWSvcxjIjgDVIkPP6eyKRKyE6d+qDTAwHx09y1XlQJvrxz
HqqzTy1R+AcS6XTpz+IN7NvjFXB8RAR6rQ+V9JmzfqIGbzHiwLDzbB7n040I9Lgv
OMwv0lALL6nKmbSGmuycQqaKlrXKkYjCwzsxJsNxooKEkH5AdmHD3hEFJv4yBUN7
FJcNYTn17wSO6JNRUR9twg==
`protect END_PROTECTED
