`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lbx8U+xNHnrlmi1PiGCcNaSpiLxCEPxu7XQNhYtaTFNkTgmmS6qc+TpPtBOlg3YR
EQEYVeIJxUHZq6/9GIi2rbZ6R+Xe8vuZpqqEK6jyKrEdGEBCi5GkLQjbYmRwNNV1
cakkmjPBhQkTLBXUdhJdNRgDA5Z8pQE0oFSRE3Wy7+O3AlxRMm92U/OoY+jkYwBZ
hy1x6PE6w7EIdVyS00ATN7li40dAuAS7qPOK3dLVdUiaT5TKiHUWhb9nmnJsNAGg
j3kyT2il1CkxsjhTL52ZupNfFlZLKiCMbmBk88FvFaNWYnz0ECUwv90FeW7rnUtr
8TeRvKeJbusLkbQTr4EWuO3dvX2vwTDgxkl14LMVnFxkcAYydMcBthm0YoLsGSGb
sMXRZlhzLL/VmBm/4O97Jfodhz4GC/EAv9vze+N6XTXrW1Ambi6hymRCpYIwCStM
HBusjnJMlPtO6EBeK8FFP1/g4O3KBC9br2IU3o9jOdorOXQse54Iao/uFscWmR5Z
3Iyur6RlMAfFepf9GzU4/cty1SxYUbG8sx9AMiywQ6/9rxZ9cTMmaHe/RtL1Ysp+
AW5tGFZ8MTXiALOV1gVftuGS5l9eq0B1vw2t/tT7rMtkuvnvNaYxvc3EIFBIAIdE
NCAAknWJgqpyuUNnqBQls3fHh5ab/FCnrfZdO4smyuY8eVIn/OlsfIEUY3swhvJK
0+KNzdFeyPHQbAVYuCVfab6rDh7W7tYM0fZAeTcesGTjanxZHlSq9gVzdVH2wQ65
I/Z8WWyPhFPfuCT1cSkT6A==
`protect END_PROTECTED
