`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i5fFhqh9JGA+mkFbg707KstB3MPAB01VnwfIZXBoBSrIy5maVLj2Wxubsf0WR4CO
2m7ZhsPzZuzjpwxwnk11fOJ+NlaBCnvyc1ltFMF/uwqdUHTy1LpvdmL24S2giqFn
xPqvM4PjgxdIJ61+xDfIWXthamzjy3x7V+Ta/h141a06qu30aN8+KMdf49VDPXZt
IAxdW8tsCn4Qhalp2kvPspBiWSC9gwfaZdJTYqml9YO3HhFeJgFQAlo9/C61m5JF
pfGz3gtepzVewV0gHSWpRFDZnVQZ8PVSxtevNvwTWlR/or66N5VkKRax64D6uUiq
NRvXxr0FFEHtFW5vq4KQ0kWFinXrCSFcfo7sgiLYZMb9joFZGQ4HXHQUh9q4OalW
riHPLCOE8JzODkykyxTqIsS9+JR8P6R0IQNJmXcoEqS245qUrXLCMx/MiexaPjtC
OJRE/g4BzEfZWe1WczwyZW99faP2s/00wwNYK5eXdChTmftSHUQLU0pM1apNkpGW
KOqux+teRg6GIfmelEoo0iLRl5YulNxYyX2U/jDBEOyaqqoAKvKeijuSNqmdhnQo
h6bH/8xEbjbUxEY2U0Y/UisP9FfdhuICtgvwpY5i4Vj+OlYPQkOfFi5YuVtCfWac
4rHU1i/jXe7QMCM8PuWTAdvIV+42HFbvNyCD/PJdEhyZYUZQutb7YJ2qY6lgxFHg
jJEXi2TXzGb3GDkxwxEUnnlzH9yeILr2CJtzR9R9e/UjinJmNteiogzC/6TUcVx6
1jOR9kfahimdgqZz2DZll+dvwtS2mUZo2VFV2lUQCWNYzBde+IXfex4aJFdWR42J
`protect END_PROTECTED
