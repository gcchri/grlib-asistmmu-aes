`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9MUqutkQK1ofvwstcpAmbOnhrbeE6mERIT720LvptjcI+h/w7k42yR42XA4hTXBP
K2PSAECIUsxqAHLC409c/j/1KPavpu4N7bObiOQffIg4cgzO1z3/e0VkMl4Q8+GC
MdPYNpXQZarnWyQAstqSbszIRc5JVRWuZBtX32YuGdHAaS4hnyfo+2nNd8cuh9gi
mUQBszGgyXDfuCcP9t03j307S3JaSnqA7VinSYNPMLYMTQkY3go2sXInXnMpE/RI
cTOwfwmJn+zpihXUiysAQdEppPOmkIMpJ5qpGkJOGFnLDmQ1yXP2iQeLn3z9pMIH
jGPyyQZhQMwl76jpDmblB/A0w/SfbNR671HK0npk+KjINGj0YBM7ziH9fS7/+dtG
YiHVYttFpPf+xi8omQ59Lk3+dI/n/J0Q/yrvXcwdnqSH4os4G6W3ITMPzS/e2yJ/
//ZHUZFHHH8rwVou3Nrvalu2Bs2AQee2rS9Ak0IiiVA33sjf/+foTIU+Vo2TvC9P
z4OBJk1HXYfo0BAK8NmDgVuApwQMjSw6YBu3mdiy3+4BJOVqQfmFy0U+5XGZ/7Qs
+NkYfBV+ttwxm8ZDgO9cFYw/am4RFxx1oqxUy59KdEMg3zluGPhTggrsixgvuyyO
T+mMzW3T6OWPgYlbfP46JszkhvS36zYksgLZNYK9aUiBEdeqAQrEteF7QIMPcEEl
Mji6eFAMv3kLf9uG5Px0dsIeGQTSUyFpEYpVoY5KAM61ikbXnGqrkk8VYHivbR1q
rMsvEiuuS2mv5tmR7w3PFwi9+Km8pqmmq79kS8mUeY8vcNwxAf/HQSBqGLAd4OZc
5MXTMzg0ZBueG4vnW51ydO5Wzo8T+6Hr6+3b89Tjij5MimOX7tW2jgsvCT2jd8mU
zFnH6e9PM7/9Mq2YugXFFCGjFgtkpioiy/9QBtsm0eDnpiB/VfvTykbFrChyj2Z6
91jOsdl+w/sNHbrmeLSkROq7sMX5LWPq2AWs1u8MDDm22Jrs8IYLcfFeCSkFF+bl
66ZPUKdQZcfOUjaKHkinbq7DniC6GCY6cNtyjNFGf0VH2xt6ZedYVOvRK80zG3fK
Mey3wnfRk1XKVPuGiphcOh+q5AvejnAOcdto6aQF4uEDxJVnz9B2gdRT501VoI1v
+kVQicW3zgyYBvjk5CBj9MpMW6KGFy5JDGEfCIkmTw+6DJ3g9Hshr8acPlWBwwSV
wIxG1zSJJ/qrjEoPsmosvunzuGrUNjFTWYfHxrIuoKlWcEryniMTgfVqNIahZA/g
RBD6Zqh4tu5xj9vbQGX+4at0/sfPzXIsl6LCmKIvGPDxo56klY71h3rrYcmaeGEq
EBefz993k7rbsq3AABL71MjCrd79oXawMOOzNwTw4AguMtkd2/jFLCl4vUri3KpA
+RHloEDcE8ItFyzNUx6ZkPcK88vTfHqBQUhs8qeUZv97AkjxjxqWXvKuITjnYDZc
/CaRQZOaU7cOIJVr6jhesLI8wpsTLY68EKqFMVDvFCz55Vsu0NTpqbpb1VFiOfbE
dWV70nXGdwVuL/PjMTFmc73m3sSvEuSZ5EgCJZLBTOh8prIYhre8lhQa5iESW+Zp
Zgto9dhY0+4DGDMz1n2lrN3bHIL526GBGu/knejIDMoIGfjq1ju7aafrlKiYm5Pq
CX7wTK6ofK07E/5NusmAlzAVML0V4bBf67Tv5X8puxqBg0TIXTqF+tMMZ6PnMW8z
yCY8t4cGijfR90fQh3LzeCG1Ln54DSZHTrOX8uMWZSKNs2DWak4cnWxsWKIFI2Ab
OCZUH0/NFDnuNGlDwMr8M+DC5rc+oFE26OaFZs7483jf9stXlATe0ZVk09V99Rgc
p9ATGYhZ+Rfdx9LJcRJMXH5v7wfcwKCGjAkAirdpRVJR1WCtZU6RQXiDl9LA5drf
eAZG9rqLuuNg4atztHCRumZH2WGLUx/KyzHW9jGABAE2/Icz7VMcMEuhr7w6izpn
KqHQEb5yqjVk8QA+Fb6HSIwzoyGxaNjOxzc23M6lnYMFPkuzirKy6P3w91PFF75j
Hi12KE8FarIogccX+QLtmzaEBXpv+SDeK6Ze+eRIA69XbUUFOfARiql7sniOoGo1
ju+7GjLgQPaCwG7rp3ZnnYDsR8TxrpJ1bcmznEhsufC1PHIkuSrEll6PM5UR7neb
6daStUDrx/pZ7S9wDLI6xnfcP5KhGqinMV0SpKPw63pSeX+MdWEJNZCTpiMVO1O7
8LzAYiaLykwEdTPtGqG+oqe0VKwbgua1ONzc2PWUhDGzxYSF9PlqUTCjz0bGrGDT
f2bk3ZIGEOu2C2WQwhoMyT/Tx3rDiAUAN37Yj4EKEpP1N5UEFv/lY1gUUgClXBxE
RxGyhCLSgmwoDrpVAbYc7Waf/3bwxonF3cVYUSYsQ55NmpDi72E6p8Ix0K26IFEC
nAVfA7tdfa5fVqAjbiNNkTaezVgvfXEet6KP4542XR4v9IZAwUuHoYHnjPzc7rw9
O/SGfEXxvy5lI2hZD31gZpToqv4pBprYobq+5b0drgQIfvDSvD/Ilf8nTiHo4pkr
Zlr4spO3rDmLxpl/jkZq24/FdylL8ciql5RSMHevlvFWbY8RCcq9UHTCbqKzHK7Y
QVgdQRNdy7zb1dBGcnIyP5PD20cKJJCqZNY40kMONt437UNQS9iJXJhvumA4NvTU
J88R4ESTvIsto5+I6RaN5cgVjk/Jl2ckVq4tverpEuuh8e8Td1tWEsHYSiBx7z22
t4PO2cefE2IQMQRucEeZS7+8jfwmjRB1TtyHrrfD4m6YWRd04vD7VlDg1EBUZ7NW
hT41SxCbs6PGjjH0tvp+9b9AMWxBNic1xO12H2x/ixV16lcicoTuUW6LdrpYeu7N
v9RZlt4C7Q3zs6ZO1es7HkYlNsBrs5z3MjRZsoBj/r3OU5e2QsAVnOMgOgGtVGow
uxVxUPeVVmAhbNX/6glBEBe9JG5sYtkvluskvDoKSTblDlbVouQ/SrywE11RocZc
Iu2Fz/ur9c+GS69jm3N7ORb9xRZi8kCscOmocxj4WAcMkekDLUKlVY6+yRGASg5+
+L9AoV3RyJ/XTPdIKuDYgo5CYUebjDzrF8pQEULUlwZlUtWIv2QikQOzurqIzpPA
G2MjTESCsR/BI3PWQSy7P2ZW50fzFMCiy42ursn1BjCgHGWPvWxoPF+xJR3CBTT3
frdj76zKSKLMg6tQn9RBYdEUw1A+RufVXQo6+Tw9+wvvpaTRayYezN4++ZbwVtN3
B8Ddbn0yharMUJp7q2oWqMGp/oVgFVgHOkOKG3Js1MS5KBnzy0qlqvT0k0x3IcSV
LS1mjOoysrhIi2+EjpCYYmWjiP2S150J445BNI/AvYo/DNrUBn2XS5C5Qgfm5snQ
vGOv64lQwKHQdsZCx6+qIFoBtL7atOSEov43TD7ogvQqEEpJcHyP/96XFIBs8jXl
e6+OVhH43o0KvIRmh7x5ynOVczcO1fzw+tW8e4Ttc4s7ABmDhij8gSOJU33Yfyio
lmN3OhV3R+BC7/GX62vpLZFC9rqOP8UXUaGlp6QhmMfoDBNCGfyjvgYOamTrXWUW
C3G7+/sMEIzALCkea1h23nDlbF98pzZOSzhcxb/BCl6uRdAbNLHTExb3WuTCV+bP
LlRHRX65JAkj1C6SfLfWQuC2KrFXYzqn5oKsHHeZqUqHkwgFyHRP/zra+0zf/OP2
VMMKHOYNW6l8mKmpEjggF8yjxNVTb6krr1bJns/uhKeIqDD2ceyE7hWJDonuHQ1W
4smylLG9Rz+fNhfBBh39MLNyd0e+VVrakr228ACxcBiVd79woRWUXED/Clk8c49c
seSNawzP7RcgOQkfaCZgVGPmu0hleMv0NmzX6phwdyObgjdwWzOcuqalrLy4ShDI
Jvv6gzriF7doCRSQxZePUXb0jyviBZ2R/89w6aLomCeQq95UjVXzkBoWHZfo54s4
kXwycz38utfV6OFPYLMjzPJ/ojp3zsWAAgRE+cJL2afXrQZyXPKB3PcB3+tLKzws
hvtG/VnbXcVB7js52rzBo0D6ScVtjSOU2E8ueUdNMfK9es8FETnnmivsRelb53Jj
58AYhlv4vOUeoLrY/27m7DMdU5ONrifgTJg7yQG4dpyUk2d6vyIDTg/y448z7lNz
cdkqbxghb+kqQ1zjZqAkO0OvtF5lX6wtGEgXckxVYwXtf4QiZuLveg9mOfmpWbwq
BnicoeI/DJUCxRJNvJGUzySH4uTgm/RgdG6ookt1w05Im2zzUSCHQAuI1xTV/lnU
Fdm4RpG4+zMHDGym0Ps+pBwsglocK67nKDuokr0ezinRnfjRUdAqC35O+V/EwJWN
gFLPnZBtQFABhqOblgdA/4CVKgQTyMKo/Tgs31Dr7OGHQZWUE7H/0nHo7u8+MqZT
+lL16hMrhlS/A1OER2WARhI7+HsqQfDva9/QBTb9uFkiC4dWNf+R+Xta0XUAfVBE
+M/xUqiAN09VBXP2P4W3IitD680Uvoyyx9O6hSeNc+67+gmJ4Mo3qO7WRiJAEfKQ
DXOjvP6lKoxy+LbHonOwtBqlvDNzaOxREpXMAN0XgfRY9x6jlFVa3dUI+HwTcYrw
8XyuKwv8886fAg100J2eRSffU8O9gQKEPAbqHebrPGs1tjr/6nWZac4K1knoTRo5
6LjRpU0YbW7raEN8hbDYjRJ0N3UxPpzMd2uxt7eMOy2vKvGzhKFoODDIm/6OYVJ1
yIMcQhfpWsedXkf+DCwV8N/EBhD7x+D+4OqWVRSu+EWjJopTr9u9+a/fFCS+k3qp
XwKbCTCa9WZg1BBu8AbyVDoMRaYK0di3ZuwMHP0o5Krjht06CStGJ4ya4G9+L2y/
lHCA3LKKuVDgHB5S+yfb6ZGVlfGhLG8wSPMNb5ehBlbczNLCo1ajOyZMyhh9Tr+H
4YduZPA1CmsaOo7+PcqlSQ==
`protect END_PROTECTED
