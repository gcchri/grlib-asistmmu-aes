`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IRWvpcE5DiREQpgkMiL9fMYfrL9WJNRK4ht1cPMvDj3aCmloBN32io7hSGqM62+p
SxPGsJRMJFXvseeNycNBr0zqREDBSrPIxOZE0N3cDbCg7MJIygxtLr24R/3tehpD
a7ZZ1ZGFGQjnwzDxs2GGTJJm6qd54hBjnsTRlssJkOUF4/9rZI1JhoIku0RUfrqD
usy1UmdrxMr+K8L8YnGaaCtPGG1xHHpZ/FXzZVheLi8ejdryirNTBWbAPmzJIsOK
pFvlzaosJ6xKnp8pqugz7bHa9crQAGh82zOTHSCk1n0pU94f0/uN+SdoDQIsqTvV
2j9ngtMGhuuTZaXeSPNHT1vs0mIRa7SJsPo0hGM9NdapbuyIK3XC3BEhQ1cALFba
fUOTB20lThShd+m0F7guJ1/Zj1wudASCPfiz74U2YpSK4ONIfYs8tNKt43WaDu9Z
Go1k8lMPcgiRiO3F5CUz3QdSNanOMgvln+Ml7Jai64yOFgbnRt931sJ9B/PVcIwh
gmy6Yo7hHeOYQ7uoQEV6sIXHwF2+QfCWKDO56NOgCxNvOJez53PNSeW2mQPVEYbl
BUv2CMgVjVowkzRD8gaC8DlP00zo+cfzdp/jgzIEkt/mkWnWGkX8kWQj3MCuekvT
EwPSplY6i1g3lws6O39aGuAOqrOaFgR7syNOi+XpAwsaBIebl6kUQA2+kb2h8Hw1
SJgQFzuGNisUW7f8pf6yCqoftrC2bbDe5KU/N3NU54s=
`protect END_PROTECTED
