`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hTEL9ccmmhUHlCvEweDWVUqckGX7QD402HiPri+cGxQrEViQiQVXGVUENS7a4qva
plbsRnIY9XG5571Jj3tTOFF6TBA+2MN6B0lpgQsVBLB+zYkiAKvJex1+7CJonq89
2wBC8/SfR+np4gIxWL8csz6q6hmWu7bUbp/WMXf/wTtICeJGIqCki204NCdFAMfG
md8psa8EKDw8DhZbPEsyT8mPhrEXzmgqRiEIxZKGXWuDwwQRizFl01koCiLF00nC
a4ozHSu0qFvfcnnylBgaaDry7YobXiS6DVklFGDmIW/pv+Ex4grCQUe1N6RL1Eze
L9wRc5X5Dj3uN3LHMdj0zCH9t51SDF0RDQbLWthKqOTDpZliPgOZqRWJqYwyQdT1
lZQo8giRM31V1m+KS6B050twM5day4Nfx0egrqx5D559PB/zbdty8I1T/5F9Q19W
J2/Cj3tC1wsslT2tVr/qyvj2dGDb9UXkxQuGz0ES8gu4y5ZVM+jzoEJk3kbEsisU
eG2Wj8ml1ieWFnhdNCPJQVLIPAbPa8uW5R1isV3//PSfO39Mw65a2tuPZ9mjeSSh
tMdj09hyjOZ0mfJ5jKh0MNjx5AXL47yyfcVOUOylzdoDZoYBYh+JQOW+yJGKMKJ2
jvcDh/RU4ieIy1ffxsKghUVzHl6P5E6Rf5TIcm7se3rC9HjmmatwY0igIpwUemU5
HOi4sgvUHMWIScRy3aSGPLMsc3oeVBGjv9pFOxq4OmVln1Z5CG6sfW0xz/1xtn1t
8BlZZmw2o63BeoSr0UWrIHkP5b9ChZQ1B2/0DP64lAAErbK8K5gTX06V5kKycPwF
aR65AaWG9NqJw9O8GsOO6Er6XtRlqy3VssEdP6Lh4Halx74i/fRl+LHSZHP1z+Ad
vUGtZBtJ0K2T3Aa+NGt4DyUnDhyqAZSnIcQNxQAvn3k2kwXCXf7ihxUXgoHl6SIo
Kbl6i+rhXm3d8Z0jCLaAR0oN9kcMu2sfTpaNgc/0cefr/ESPO2Ys/2brN7XWQRIU
SGCTQb41vF1FPeSY/MAd0ItYGCUotVFG4bblZOaru34EdrnA4RWyv/TSkCaTefCz
Rd/29wQoFmUHN4u7ySAXAA==
`protect END_PROTECTED
