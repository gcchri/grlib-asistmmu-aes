`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R+UpP3YUfMJSkdq/1appj4pzsRY5ucDB1FkpuEF1XHPekDL/vOMvHCcm9oo0S+h9
14Jo4nBJc6ggVkYqMMPHPG31mN7zFvlWPRwz8bgIJgYgSfm3dyZbEs7D8pOMFlHH
q/1Do/KafwXyTTc1PLnwbCUEyoCF1FTgV570o4xmn1Hr3wWrSzmknfmrb/eX3TuY
bGs/74CXtEjMxiuH0fiXBFvXhJ+OfTc38CIUTPe/P650tyheh5mrU5fH5xRPSHhE
V5/7Q9x+nvanbEuHKZOTAzldqnF8exYvbAJocVcNHUBknD4sPKMcBeLTVvO/3LFO
MCxf2p7kn7Xmu1e0V62BPfcvYT1n21hFGozSLg0DDUT0uAdMArmjVYAlFuHWRWVJ
qm/J+98myAB6nmvZS0kWg+ovtKyrfrUBstrWBhIuD7M=
`protect END_PROTECTED
