`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k9owxxyQ123zTNhewgf8e4E22IXC4B1I7TcitdlOFso1IkQxAnoflYQYs2rWAcTw
eaN4UFWrBACRkEa2liR9xlqLADV/JvzA7yWTQ6zRk87juW2KubmRHTdXHkEhmGrg
lPD4SgmP8QF2WBi1KX6+8/0rfpgibk28u6dzaMBT/Xp4mmOfKY9UUEheJVgXzqB5
tHY0rySs6binhFaF9+xPQsjVfZVIQoKEvwjFOX8GpTk4ZP53ysO0ITCpG9H4dRv9
VextPI7rusEZckDIk6hBNXEtuiKtTNbkZo2DQHPl3JCsC+DZUthJA97oA0gsiDy4
Ua8rrWr5KwXJr3XGGV7h1Ps5UlFYfREoaAU4+EdsWEdV2TdybwN2o+wkzbyUfDuR
`protect END_PROTECTED
