`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BlczRJqeIc88bdCbjVTfjafg7PDltqeWslBGujLTGoYEE8lHMgbwX2z6WsIzwZI0
IiTW//eD3wfzIk9PAyyK1bqXfuKmo5DSbhFa5phGlpPIg4xhpPXe3zin2yCpTH+h
fkyLRsEebM1kcXzUJobY0SowxzziKo5CgFlW6YPK7FpxMGu5LV6jsDzeG2YLWdN9
70RvD7WKoFk0ZLfyrSp1ol8SEKOIj3+BSHjbuSXFvXtSZ8COzu2HFcX3pSd4yy29
IrzPrSMbJF4AjMw9xOfZBg==
`protect END_PROTECTED
