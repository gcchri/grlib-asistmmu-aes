`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pOPLj9IvQ93nSSThs+XskwzLcQFJlDtO3B+vFfQ5Gc0U8oCWheQMhiH2p1i8JRdz
8zDY19NQu60ICOEA/irtpMTzpXbze1JXTwJKUlumZ70ZP1ThzD9ObKa/vfqqg1lm
Ut6L0mYMwiL/w4hsofnQYyoeZKmlakepEBG02pCJInTa09wvqjNurzXs9IvpAytA
yxXdS0jn63W1xIoZbeZ4FvhKPTKne6x04mmK84kFa0j5eqXQBzy10qnTUmuiHEi3
tlbhs3G/tJZ7ezWzEW/i0ZK/v9WBHhKijLlu4jTI2UTBWLRJdoqUYKL0Yd5O9l4y
kKhmyxuRda8OVk4nzwGOmHYwED7fgeZg4yEHXqVvHFTh7/+cBzeCXe3rR27sX3QL
gJdmx4PMw6ZzTcv4vrFyz2v6npQZk8adtA48GJUsG41HuM9zXuoGFmWI938e4svc
lTsmcScU36ORdGUCU6qtmFxmd9AL9ee1pfJNpWalm9QMO6vcwtBan0nnNp+Kbl+0
MzX4oZEARRuUO6e69LXIHxu9Se7yroM94U9u5jGA6VTXIpBzfRx/De63wosLXsb1
BLZXr9SPzwCdjW2K7IoIpIOogz/5qwD7eiaxb8Cqx1BdpXm4fpZZLLJPINYpr67c
kfrtPh0fvXyzRxwzO79Ez/n/a6TUjZbmRN/auFbz9i812f2bvFrXkstPqKaJd4TF
T8vR04OSUiPL5sHPvOX+mXkUdML8Z19fWgpLROjPcxotCZ9kL9WuLH/4zIV+fA28
uBUkfo7dLXjn8rfBuPPqqDhOWi1cmBY+vECDTVWGESCpJ/RQpzqWxBYVOMPHSfe+
H8laQqN5SR0WFhW7Jh8ch9kYqeVoz1tTsK7FYXQJk0JXI8Aonx94mfzDpYK5XjAv
v6PyAnmrDjukIFD6HqqNs3QYybi39UzQ0YsHQqlj9ONZLcmLdb6NuDcCUjlUQ4zF
eQqXYRdv7WmdXhewPjxQyt9yyInrAm/Qf+hF8QfpIxvmFOQXrfJtKzOXnqiyetSu
r2xi0ljNE7UwCqwGGkURRzHHoF2h317HutZ8gWrHpD8pRhDmbBThQRQgqYRJ2Nx9
Ht/JXzzGqSA6YopFc3RiURM09p1CwX2EX5iUBKa3oIii6wrEPi0ag+GN/+6pYskD
CFV8qkppf2QrTBdL7p7cO/F0NOwP7DQnZfjHAka7xjrxw59kK1TWQnSrWZPNW3uW
ub0JMkE9gAojok5HWsA1syILZ0ZNWtYA52CoREzqwrdWcUebgHzbAYAo1Q4hAlYj
Uj51aZ2RwHRbqbgyoibqmNYWkuBJU7nl+8173nuB6CTePBr3a0jCHNOPamArEmKL
G8jIjsu5PoqDxPhNnyxFFLgFjHU7kucC4dkMTYr2jolSKs5i3dcIvwdXk0JQun7w
1Bw99REn+aPF1UeDIsIvmTZYlgsJ70waN99OrbOT6bQGbDOLryVmZ+jZa0TT031U
bwf1KexjbkCRwthkEfxlsyr9KQwf4mx2m/YeKUn1zCrVPgHSw4rn5Yh2GKbTxZDr
uLnGKysYcKYfatZ9Qg14WI7oV9EoU/zNOug0Pn+JcAHNQztKtNn2gBi5j2gmT4pM
/DOU8rgM313KIy3mOr7YvjTUgm0u414qioXHqvP+VyYyT7tLXCg3+pNpXMDv/A1Z
XMmsUCYplMohH1YkYsBh80k5ZBU4RMR8ral8IOQRXRMwJQRE9lu0VP8r4AqkcyEY
1uBxKyOIYlrnc5zZhHzq53yFUPauK1Ro+w8xQeIcAxfpCdMbGI65+RNriALYej/T
mjhKHZSXpaPEPx3/QIvLqF5xjS0Ky/poE9TiPbFFfKmd4UyTxifKzbiVhiXbtEvM
zQL8t7+ZKv8AImUC+Sj17zuMbZrRWagV8VRr453S/4JgJ5LhOGfW/mcQVYmmGVDq
OFIzf4MkLE5LYtX/GNTSGesLe6Ydtwe4KWKjGpZV8fXn7ecOj1rmWLiUIaW8C6k9
KOK1pwsUve3C5qHyjBcel3OTcrMDhG7WXnQM11zR1o2Gz4z5UyUCQyLNn9UVurVp
AWWnF0VYLWQH3IJ7O4uHAMEBP0wbEXr4kSBhQ1I72oxVfu3VSmXP53JlfHBTXGnC
Iehu6bISc+XEHnKiuGz/Aj97P8LY76kPQriJvzShewY=
`protect END_PROTECTED
