`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FqzW+IGO4by0m/YaYUC7yPw67t5lCXpsbcGMZ9A2dgvy0NUDqiWY0JEIwvss37ze
+U95WBuxkSdPLJoqat1OqMhCil1O6nL8gcJ7WmXbeupVH3mBz02JYqVkvfa67Tqz
aNrElCcMRoSnMEdTdKWV1D3q3TtuwNRrb47kl4vmzszctTSX1AsJwacSdjqnHzQH
l5o1QaDpLZ9jKT/aAK7m9BWO9iQg8akH17Iq6FbrhZolQU25iifBbygFCeY57z0Z
fHnVRfZJIJFpBWTMrB9p9uAoFjYfPwGTrs1OsapEmyy05kNQ7aDk/V2wmxWM/6sV
GtpmnLTNXaEeX+O2r1eAKkIJw7C6ZEbA27pY/Pg/BzLAIBj3tdo59ylnRWEPce2y
9pNXsTQWwXKcLg33lFZHW02EY3SySZD/F7q78xGNCv78jfOKyoEnV5tHmr5PzPrM
+W6MLcdnCNT/WFJwSK8k8YZ+HWFJUL37NjhsYAqie3jqvAIXCKWXEKK3jPm/e2q7
jly8vpzpnq4/w91Uhq49Y3uZWurINUBj+WoH3Av6iIVacx3pM3tNKcEGtKnSLEqq
h3ILyfYPHz/vZKr30xj+Ko8RtPsUu33yi9C8BUshB7np4sKNxG+d5Ge/vS0E9LdY
d5ni1SzLBLzKDsSzX+0Jgwc9r0O8TUpHj12l/3AGh0B0Y3pubqlt5KuaInHbQM/7
lxOgM3FrjWFdHzWghwz0RbqKR+4uG3VxodK5u+GIVDvb5Kp1obL0uFhMhjePTRq2
SIlgHMjwGFOfgplErSI4bSlbUTeBcUjvHr3CahA4pBoM34e1pG3x/0x+9W/CuTTf
r44GFiMgZLMnCyRpkackljacR963ho0UGRQYynkBNg7xcbWAudz1YHdjd353gaHR
V8ZKrcNEmi6I/U8RLl5oc7tGPwadf7taRkH7oPegSk+q8nAFl3LZQyVSn0BAe4w2
Zj2ZC3a9/GxRp5BNILfet3M7h9ptd6FS7P1Wz7Gc4/W9szICGk4qutSmCyZ+sVJd
9/DJi8g0/Ws50FzAu4Wd2jzNI2yqU5B3N4J8+7DoPjUGNncETKN3FWGuHwTI5KvY
K0bDMoVEodzf37L5sT/4za3Lw8Xr1rcEWzafl6L0OatTrf7lNT+eJB8JLtHxtPtZ
fTUslUWFfLf0zGTU/ju4ZQY8lBb3OOE9Ap7GCf7JCc6e2HoBd0TJXxt/ejMZeN++
HF3wzcbue+nw0C6r1JjZsMS3pOHgL7H5gj+XUWyr7ByYJpc4iTbYDkzqL0yzeh8p
8WgRiZvpzwkP/f3pxvdLLxBc5lfCX34hYeuxLyzB7n6m1GtsiQXH3jwAF4LPgjD9
Z5NAFEvNJqzOLdUSBnswqR/ojt7izcLboDnuLrzgFIynCr5R9zIuAdik0tVtYurP
hg1P2mhTgoZ4ATsasRtaWRr/NyZ/tHRepsBx3pj4KuI+EDBWbbShsY38wS8e9iQC
Z/RAFXyU5l2V4PfEPQTyuttdnJuonAy/PeWzdLDsEczyJ73Yr3Hik24ZKMRLX4zV
00B1RcidYl0E/Yr+0nH/6A2t5NbNexVNH9ZjG4UWf0Q1Fo6/8f7hoOEs+08OF1qC
Vgjd03P6YkFBBvK9WS3upu9IvtSzl6gGDMKKnppUqiTFhYTwZwIzT6xvE7mBk37b
3UGAxXN5Hcjr2QyiPRxUxXUXd53OLudjK0RIXmbQW90Of8XfkIEGkYbM3Tok4pC9
GougByagwC03GwELpYmrarJkU0tSrcgKxYjhshYtQo8mThy1NlDCQ5gJ26WsQ8yz
wznyXT4rzkL9FHEh7x7CmFXwb+ny+pn7J1mQQf+41pguL/lflOC/d2+HRGFEuhAq
2KctC/5I8M4j/8ntyUjVOub7pc6e2RKT3jqI9oTXisbQh2qRHc6XdpKLv2XuwzMe
YZUQmZv1r8k8LR+xztrin8FZJb4FJqY+PG1ywyW+R25d3pMgcSh9KNOWkYP1XtWz
uDUSNdSfY42SFfoRC8anjOp+1EzVU1AD2rSicmm6r2Q5czyEfXz4IK/VQaWDItFn
Hj0VHkjo3U2nwkMdXOwX94k9N/e7LTxdILBKblKHnc7yp7mvztFLBSlywvPHNUxv
hOmUCmr7fYVmXKOtF90mMoCKlpsM9sMIjBQz43eoSDvmo7xhWJS/wrFb+DemGXgu
qeSkBASZdQZdC+Fu623Wpv9MKyG5fQz5erv64R5sNM57Mh3u+Vj6aM8zCchsp4LH
OII2oeDxDd+wlmAzdoddRH0aZOC8cyf3HzQrs4YtWqbxowwnwnEE7lLOKaTfzo5P
UV5qu5fkrTNaY7a0a0d2OU0FXYvyoW13X6WMTBtBS+2JDWIP2pKtQoe62AENzGBM
DoBwi3B4vaSFpRTiLmY/HFgYL/tQYHMp6bRttiaBLuXklhAGMxy/5wtg/Cn3BSfX
twpg8VZ4ibGMWbe9tGm858/jodcseVFo3j7AN0Ko+vLVB++erXL4xhifqqMc49lf
30xVRNg86cjc5WXTXEWN12UITYti0a6ajVtK8dw+L11Duzvu3bwefSPd3PCj6Af6
Qt/PnhZqBPafP7inPAonuGpyTK0bgmFZ93RIT6ke7iVREMAXAsFrauF0NNLw7iQ5
`protect END_PROTECTED
