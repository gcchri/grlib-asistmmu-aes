`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TzDEXz0q6H4t8zaBrzqe/2N2FB1CO4+iEl0MUZ380DP4xY5zH3OgRbcEiicR2ncO
TNSpKpWhe9Oy22wB+TrSk10cmun6hZ7HrrwAsxVj533K/JJD94h5HfBsaOuz8I7B
rUNylAliiBu8Mpau8ElTZMS4O0PEp8FecizGbw4rsh32F6GjqDi9TRi3zXe/oR4I
+Wu0FAYykqEdDZP/wld8b4QN3emYguRo7AlNsvi6PpOWvOE9rS4KjhrCp82j5vkm
mbCSCOLu/TMLATZXlxf5ugy7OgxA84Ms5GWcml2hbqTXQcVzgF5x0HX/Y7CiBCo3
mjs9rwvkLynrYvepdQVQb4TI+9wgMTtWURysX4oTc+jnX2lpRvx/U7JxRjzooGP3
8Wt59IaTN01s9kCaIt+I/utj2HULWT0LqlIIoz/DiD0JBaDVZEs12eUcmgls086R
CEap6OwyjqnsaHFGwkRPT2fdWsPshQHVxu83RxZbpEK+ZLxIkG9XFvFz3EIntyPz
jHV/MSB7pYp9qBufhZ5C8a4o/17lGIRLwiP5lyqqj1KjxwbIT0EdhhYA638gMm9U
5UKtaiuUBz7mf7fUKakJEwhTsXAHyDtCjZ6aKypXqMqMVSkp3HL73XJqczwWWAdX
KIBO2Qh6gubFXz9S4pnVF3pZESTfoQBnjvttGEIz+pWm/tak4JJFOnXCxb+CItOk
OlXKEw1q/8OOSEQtNeyFiegLGRHmcCoZo1BrVZdX08IsElpsdcx6vtPvypVA84aA
J1HiriLqp6xbY4vzzvPjkvLzlwor7O1fKI8S/qRBDEmArjwQwywrYASp3Bhv58gG
xDrK4PGdKpi7iUVHXjQo7JUbJ+8xR4EErnxl0gNe+Bd+PvkjrWO/1CPWVyu0MywQ
Z7lnTmAWTxhFKPXDQLL2rC27IvJxTQeAc5HSe7YM4Jggf0eMjMCdn0eDPV0PjRWi
B46d+ISUYtn2wond0QI4/nfOyZKpN1SpwxK+Piqmprknq9IJ7xUUw/0duIIXDpmx
4iRtAMMtdD0lcuOtcS7BwMrrCzqxZ8O5Iw4/HmenohijjhrVOePrXTjK0WCqIS7J
3vhq25nr9EsoWhJD3QwdEbALZk2JKXg7hAA/1xIJvfVZf72w3m0oIKtWEqB6kix7
2gWTY0UygfRbJB2Rr9+G/fBHuZB7xK/noLVxfi5P+HVsy1GGk7wDC9bQYHSVMc+h
2mQf7rtJvyPj+BxSShqsFz2Ch+T9O0qDPsJa4com6p9XkAxW4NC/m0uOfsoh8ZuD
6Bf9sCpBvvwkRFkU95oqqv3niqKt4MHnZJK4E0/Je+tzLbvqCRm0CEkOXLW1vv0B
eTJdV+a8jiRT8UcskNZ9ECDE3BJAp651Ud8HMXiiqfmf6F7HL5Uv5YSoNT0vSkl+
31t3/GhVBSSwwRIvJLqro/P9Yb0G+jEgNIAtLIpuwVv6hNg83ZD9IiukJ3N61rM9
S6SAkagzitgmm3KYsbfkVWUboFu8ISs8hhKHWA71Xw87ms5g7yZYCTKXffoYps2b
XvA2PEjeNM6AmgrCOnpEliblucByz9Pd43pMarl4TnpucRJ69dqgHcVx12duHFKA
wfZsGofN7t2EdcvTV0Ty2WtUyxDZEex3g7uNpV4aifES/yWMZDMtoj3TtjoI4VY4
BOdwO6lxVz35oBHlKiRdEJ6QU7cAaXrKV/aUHFaSaJ6StWJE0Rpwx8ZMVWNZwaLq
Ca0sEAu7EfZJ5fMJgUh5ZdO2EUPT/1OhqrbcQwYCDsl5hLwPp5yj8ia4dpTlguNe
BYN/Blgwv90dYzy+ogVCPZIladNg+E0CDDyg6vqqKU+8aDQDUIdVp0MoAH/eNUtZ
pOgRe3VPkELcfcigQeJ63fAeGpINkzVSVtMYAyycHJWkqEzZkKIGjM10MR+NH4Nz
qBt/4aL1Pq5DXneY6HAt9yv/0nQ3717JCdFW8apsSBpVvffYQJgYY9YocGFfns6g
72Xq+1GgtK2XPM0MIZOxX+IgwfkgadismUjKR/enbbNnE4/BxHP8IKHWbPX7mGhw
z696dqp3aDmde7ggmvKzUQrPqBtJG4Xpzr6U8k99y/Faw2BSWvAoC4UeiZLfIwmB
4DjrTcEdpfcas9zPe5Gpe6T3a1pnY6cgSRihGV8khkUHaj2uPKDB48k5duAgnH64
IALDan8XZluuaHVAOXUItUT65AYO5qZZawOWPH8VodjK48HymkxbM8zOIlTG2YGW
0icPFjOfL5yuOj0oPsQqszwx/h+5HUcQsImf0dBNyFBb5Q+CDQ8jNC0OAqVO3eUl
W0s/C+8DNDdCOsuzmj9ftFUoo6kNkhu4vGFVr/BgwM1cjCcmMw6h6lJHsaJ2Hs3q
KOUNSFziUnhMJW1xRCAN6C4zATIOUpbgKbbKKzamd7ec/uxIrq4w7hdDBh4tZfId
oPLsMRgB5Ttw3HavwqdBVs3WKftrB+sENAYlZJhUgx2mjLl0J7vRHOCdMPv5rPnp
g+V/x89YvMmVYOO3Nkeh6ViEQ1iObEmVkFvusYJtcJspuHJg6WarQTDBBbmHYWdA
RuoJeJ0zaLn07oSjfTKsBT8zhJ5ZgjtvCPuJUcoqcyBPkpkagNMQQNLYl01m2U2k
iI3222W0iHeHJDSzL/qwFEMyRqTTfhBmHOm0iEsUPc43JChADLizGxUHCj37gjd9
zFDvTd08Txk9TzDiilT6uW85rlGlSJJXqria+RMsVp3FHMUEW7Rp68hJ0qLRGE/j
4djqDv1w/K7R/gyU25ZSddZu5mGEQ5hO8glQDReGyxc/bNFOVQhvaJLlp5U+w9kr
g1y4Yth60f5PjpkEJZvYLE5y01547X5+0GonzTGLwKpFQaEUgTVEhHgKZ+RzVDxA
Aoi5w5D5L1cCfUh3d1MPH6+M7ZhV2InZEGEebNxhTxqlmt49i/goQ5wzuHIAQTOe
yCyVUD/2n59QlDQRBvtg3kQuYWXhwemGQrqb5yyDOeSASKWUOTJO8t4DsgsxtlZI
i9pi9RG613kGrHKKEh7Gea12lEULUCRqiQRKd3MCHI0uITjZGimvSdQeioyszAcq
DYrhfrahVH0/Y2skYr5k0Fna9UToq+s1VqTROYpXTIuSeg6h6QMmA2B6HtC/bnvW
8gfrnvCwrcViYJS67rZi+euB8bYGxO6oRpGCegwKtMgLQoTXV3QTrTfUZ6l28G26
lpTbpVH6y006Fo5J75gULdwnN6LFWJcWHqWcPp+71mofCPh2ZTxkuK1YkhRh2SVS
LX0pT7SCLqXO24BHQBMqARppsiazTngzRkrOtIgY7xj13hBS2j6QDaMP0CMXVMG5
mR6LHq7KrX2MsWXO0kbs8rHYBe6Ewls++9SbbrI2VCju3GTntKKHT3GNJewOQ3LR
WD2vaVdZKAZ+ResJUW3XhrQPFqeo6h25m+gu3jxJ7PGpTYy9aKKnDQ50rG5jr8Nn
tbQNDf6BmdGyK5Imca0bw22ZreUy9b3es7LtMOPIafIk7MPOUIccfKG9XaoC8BlC
7nNlJLagLOk+elSn0EY/PgZuTfqsaWv6F7E6DbNORUg=
`protect END_PROTECTED
