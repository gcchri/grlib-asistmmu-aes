`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E0x6sHCdvTXY9gQ8FFdIS8J/gmPq/fsTvUQCnn95TfK1ViBgvhbn5lN9GFPiJbKE
9fn+k5nxkZBXRwZqWKSnfF2Aqp7nHJuvMZ0g6ezHNzsqJaKaQZoSTEVnEQGbJ/Ui
OCJdNxnG7fj7sMg5WUArHeIlsiRpzx3gIKPa2CpaOxInrerGwsr+4pSAoxv1rpk1
jh6vPeobM0QX3ovm0f64OTG0M9bosk0W1qmXOcCjxF64DIMx3bcR9aqBKw8TIjYG
5A60IWCLMAcFgTdXIpYZd7L04zFttJeNbNw6mQeATN14cYS72Xl5kAgmhqKFCu9T
`protect END_PROTECTED
