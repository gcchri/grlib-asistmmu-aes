`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BUWf2ht3ndTmcKS4eEPqPowov2aKcdtS/hWSXG5tnCPDtD9BANIm3lvWexqOD0mo
oP7hBXOl95Ak5czVi8mcuSOc+9tD3xslBRDqxNHcGoiTESiefCttrTBdG5yADkwT
IaPyhtEdVLoZOuLhUVhwDnPTkQc8cV5m/d1K+6nYTwDAUYDambeFD/vj+a5W40mk
h7GHrcUx0F0qdC6UmOwW2Ce8BCeScq7QaY6319Ep21xqofOrJRlZS5orc0V+GyTN
YA3UUagCsGZrte0OAOTG8ZoImokF/IPWQpTAxkQNpYNnS0POYkaqfvStDJ631hqj
MsQp+7AF/47wTEHjH9hRUg==
`protect END_PROTECTED
