`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fw5QGTK4bQrs8pRjXytB1j0/Tzq4jG2MSFvPnJPpxMANPGlTae9MLPvKp51KHoQo
xM2z7SWcAVSkzh8+4qZccT+8mPo0XdCa37U29J/EU+qSsAXX9Y0j+O6WGuIzREGt
HF7xwubzTJ113AGkJ9VTiGZRqiRcNpQ0fLuTrV3N0IQxSKBxVAC8tH7VBkgcRh8h
Z1WLa7IxtLpwcBUY3VuekEKLMNvSh26phialbaKmCO22vRrYx5j9AKl1GbvQEBo5
D8hbaBCyxAW5QLLQra8zrB2sxZgJAIxBtHwtD3b7ji25clBEYYG5CdW8ZaAAPBuU
IQaCICrxRv64ETM0YtnAXJrg9j6j2Uh5SdVNQSPxnPPCZmoXyk9w6lH1XKnc34yX
ntqXfPpDU6M74CkUP3nh6S3TjQF8aIlKvFkOOqNY4U1WbFoo7ejqAAT8PumK9hAc
PVzOIvl11hJvXdNuz3xVPDnyzGaWGUq5bxpxGCAPvz9Nfoxclh9RFqV/NhFarlJG
LMHLorE2rDaZI8YjB4g4h/bzV4v3m50m1+Apvm2p0uVj/rspwQz351Tp6S1qEJFs
RQiwO77oycPCVFz1sBjfBvkK8KPgLmchPZJRIEjOTVXcyOXCbDXwXmD6UGTZvSzx
9wgsN45J3so7gnJMVYXxbslVFmlZBtnFGNP6PFQ8i2dstcBn3J7vD04aFgPDCDdq
w8vgH9GRU1mEyjFdNaMgkbapyaVq4Wm5QNrQJ4HZFuuq/iJKo3IUoDiIAOKFSBl2
a5WMnx9hXe3d47oBKPvkr1C93OUic37tef+LMc6reaWfJ2+jzD8XqR7rRW3QgnuN
8HrJqUksKyQLSxtnw2eooVtnhZUzP8Lzo20Qt6b011OGqLMKSIqxnvbG+Jr2fIes
H09AdmJwcrFgxFHkkZ/rCUha1mYzhk5oddYwFnE2uCQs6/0j6893RsNE+fPE6yOn
tc/cCC3ieFXSv7jwSF09fBt6S6aWYCo9rdVeoFbKn2cOAvOpoMk6Rrt7GjEFZ2Nn
2yBsaKcAhEN+6ZeVjAJShrxHh1kZMe0a/4XhPajybEEjBnP/JtMFODarhs0OT1cL
3qm01Jvr119MWhXx11yM4ekTuse18sz6jSFJQshsOxVgxwvCVpg+INGqOgERp+Ud
GRUymSba7TuhyMua9Ew+xg==
`protect END_PROTECTED
