`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h6R/MShBKiUynvjEsOpn8adPqmpZj2KgMhvklKau+XlvAIWxcgcGdAgE3wtL2WBb
IFCueVsGGWGbrdh1/Ra3/f2YQdtq1IebgPJ25RLr/bPpovJrDHwrosx4G1OQULse
CoBXZ+6/r9SuyBHYC9nVvEO9qgwhlyuVi+bIDRXN1dJo03xZx0al99TLxSsu+it9
5wGI8SY20CZoGWMWBB9MvQCY7yAPhM5DJ82twIQT40hEtcznUX7IsPS6FrSGtIeY
sMbLbzrylAsOzrXwiasrSFdaDQPApBnIv3KUW6s0CPKHUN3VOwTxoEegB0ur/rZv
3A6kjNu7pNPzrcjn0zgW1Lagxp5hoQK3idZlCbnbONJ+OwNG6t8OdQ/r71bkjUk/
1b72vkpVWwm3yUv4pLrI+baaowVdWWZh3ZcmnWrQreVvHw3PySaZkWjapaaNTGOw
I+D0waQmj6FMLuPXtYPoVqYPIoMze2j7G3zvr5hO4sYqAEOk3kim6uE2VFiyo+7w
V+ezBuGEu1fmsFY7Lt362TayYDJN5KaHpGE7td36s3P8euX97o+L+MuRI7MuR2jG
Vao8a1JuUrgdL//XnwcDahwuQXskMb8gb2nIjAmsT8GMhOo+5v5bg5TsA92mSGvY
eCOc0+5fe717N72FNJQwvdHNBVqatXPS7FmJLeT2iIzbKxj1yIRDGLRwVApATVYL
YhWamZHzNDvEc6ZjKcnQoWIxdN6PEh5kZWSWmLP3D7krDBpRCECCH4cpvirRNNvc
wEYDB+0qILd65VN08fAwCTZ4TbaPtHJ6ItKzhskFdSc9Kxjr1ZQG5SLnRxQtJl5v
9v/oRdA19gyAYhU9F/clZAWOb7rPLPWkWahOziIr9FStzINqdZCeaLt+zyypSViT
ufh8KHj6cpVaVilObR/lMiomBGF+hONTyKXfMj9xBwdChciW7P9tN/u4u4FD/SBX
OI1XyjEtZhjqTRCcjJ4wCIcv+DbRg3zKO9WEt9Wt6jDE5ho1tAL1euwXMd0tw1cv
JUpd4Kve93RkA04F71l6CpbU+gLGSO3qH1HTB2zvHj1PGyne5HtqPlG7GH+uvd7B
q/pOnCv0vNo+dtwvYMPlwhOnKWS3Ccsjemjjz+JFmwueb5ZQ0j3p2eTPM7BG4bTm
ZkfDZg6IJOgGkZFdh8Pr1CJP7QPJVcFKmd28s7XVbM9ldYHAG4F2N15hqZsLchLt
sWMPxIsDC0c6Xi+INM4Vd6hMHTk/5lbEEe1r8wvTxRP6TcVOA2avqEjDrjY2KGih
vTv2/PAejRAwjquxVfWw0JDEpaLbGdFEsZ2xgVw5Vu34h5Cf5BxXj6cN5kCnCv37
JYY26XYOGKfBa0/4dpc8goInyGfZ4s/Euhmg020mIaYSdCI2dm0MiliCUz1Lg5PS
Hj4KcRCTj0qRtAp/f5aHVDMef6EOFfwRd8iRWIZC8daeKNYZwd6YE/H1+xaSwDOO
4lEWgej1zXZTl7kC+vdDxsQ6LYirNPyhLXIWkvrpnfpXvZF/B1m89PIam2knyfBE
saW4TgNnprWqYJdD4YA8KJmOVgpggJSo/BGBQr3E/uDGFNCYfNA1Rzme/IC13XHL
lv3QK8U+WwR1QVI5USYdukI6q/h4VZqK9bB1Ahtp2dbh2fUZ7RpAozKoa8d01194
izXnAIoIY5XfEqmzy+oIaHRB1DlkMqUYxGtP7wT0jyBps7GwY6DcDT1vunPHSLBw
TfONv0OXPXwXiYCgEyu3P9iqrYI3RpYMSTeIeqom/lKov22dfdifGkOkDTzY/IcN
Ikpu6cNOmYdTmP4cB6VoOIKzYto2JyXcmjOp8Cr1IP3Kk0UNZk+VRoEPNycvpmaR
fjn+etP+euDF193jsQ2pVIBztyUHvGluSAZT5C7S0NTVWMJMZNSPl+xD3cjdhkD0
WfJbCjlBp4RfnI6c+dC2GV5ewyzjYGujcJ0Mm4UVRaV7vf3YC45wlBjTM9LVxN5r
GbazBdVS/ZP3b3y3PZ4TU9UZKKdghAM7jnHCTe3i2fQ3YTt1cchRkSnj7O6hdWfZ
wi+oKNlwYz6SPM3bIiVEtGpf7BO6SG9IK+u543TVnyzfwv4BBWXq+wXtevljGE/Q
hpFtpwcbqdVbyTZNqL4GjPfjO9nxbgdxIL4p3eRBEAKCZGSHV2tCEUrp/BvJekfi
yT9D8RPYa4OfLp/GofbQE9qEDUJ2qmDrNaFjTT6MaYIcRu5AoLsZPr46EE+mPP1j
Bx/7/c+ImmfnsBBbXZ3iH9ZtUOl1qKiXjFHWEeWULkamZro1FFyE7EvU8ETuEmqU
pA9CCxKSX3WTzc/l5YgbmH9XBFuNlIIZ1T+ykMFkd085gfk7W51F1XXS/jW/2xla
9d9L7ZGYu/1zl1jdrj+aVyjVXRoD2dLH8DRT5Dl2M2XcjMLflih184kxJ0cxHH1i
6GtSV725BgZgEQt7Qxjm5vd5Ty9TTr10jnnwnmfBQCd5jHJS10vIfmPZpMCemaNh
gOSNak6D8lSh8D1K5z5UcwuU6icsGCFcykfELtTm5gORLZ5fGc7vHO9KuTFT1dO0
TuK3BvhC9IF84hbRv/4rYqN911pB6yiykZjT1LgNwraX7+iJu9qv+vsctX+664CT
GbQ7dN9yuuqJX79iRKg/PZ+1xFQQ74n7TdVYtzTW9Ea0YX+WfA9Du7ZS5cueEPYg
FRQjqccaODgySxbEWYG2eum0QQ2ZVWxFDRWHdx2y+rn8P6uHABLfcFLjdfj/rnsx
zmGwkVlpXvGBnIexYmrfmcwPZpURGDEpoABSKq2Bxh2vZ5SJfypXZtMmHrHVeFO0
5l3wHR73Gh5C6Vu+spGgEnWXE7lAEi2wghgVgLR5JVAwGJKpH9uyqxlAThx1JYhg
lYNoMZSrLgBv2Bg57t+JHX3GQzFZpE28OEBLw3UNgQzHZPJ5HxQ4pf1LYERnd4n9
w1eejM49NMdOZvlKaBJiq/TxZ5TENLvI+T/vs99WO6DRTIV4Z0MmRJB42PCGxW0r
ZiONklb9aStJEErJcgSzz+O2RnAxTBhnPjD2+qf7QaxXt0uPUrrYQHDkS/HxPOSj
NWAhqn36qzX8OBLjtpeLy52CCuLND8A5jr/CL2Pyv6xfwBVQ1MzedooIqI3rRcIv
2xOHxtCiT3uNpjmsjcKlxdeS0r4uqtkqRMxK2P6vrmntnxSP7fVg//IHkn7+XSKE
4FFPlhoPFU9FZUKxqegR0YWGGMB4h7YWxoovyNifZ8jZvoM/WLuHiZKpNNQ9O0Gs
xQOzzxEoUc2g5qL/sc/ACutCTE8csUn2lBBvkwGJITKne2SXLxRUkOB+OnTzcsAX
ZeCME2Nrwsq6LhZTuzHxdiJFFWVG+Q/1puN3eoUr9ecpws+F0EC3DiynW+oPlDfO
DIRH8iFrNMx0o/l6mMLS7bFiWnozqXayPfmNJMf7z5Dl82fRJdPob6lMex8Ah6dT
8q00W7APRvJUqtxj/ag59fALAHxpS5NqcPRadFDgZmkrfqv8YTtlH95yQTsiL+ln
l5UpE9oTBHF41uwFVPijMIxfw0TLWKvAUXXkN1iURWq7QURi3KJuuuvXj+6ZEynw
ztZqNdj+JWz6F/eLlDE6cxMkUi64+YBnBiJHvfT61OfbDjCNwod3F0NGgQGZ8KbK
DaLWMh06uJcm+nO1FygqaZtf/aTCS3cLvNSIVvzuiof7RJkdLoTXuke06GRqLOXm
oaxzayPrJV8reylAea5xpjOLEzPywTVHZmiEMFhSMV7rOBMywdIaJpvc0+v+uVoL
87axu5J8fQyns3fsjkdgaaLYVazUnVKAMEB8v/zABR9yEbBOsZdPCnHWv+kPEy2X
elQNUxMe40QxScNLhmRh21g8+XoNGM1aUqpnFGFoAiTdOagbzyEO80Xn+t3vPPuL
lXz9IYfmj6APhA7ZzXJRdOJ6+rG4EDziRxOPY5OgDp3FzCUUNwo/c0aUB1jIlfjv
ROJtmbi7XlWDw46YA4wjTvGVHIl6F/B3dO22uQanBR1tso1rxMHq3hYVS92zXoA4
EU2AAomYOKMB//200zdZ0idpLZO/OZmp7jr/8ubmKYq308OINMSzGXin4otvQWik
BNVdsEQ00z9M0yOAvHUQNo2rqnjdZW/9a+D646mff3NzMBVCQJgTCN4uYhEj1bWM
QvFC3rkuW6+KWUwfbNLVs2s711Gs6VS+8wpdkr1KokUq9k3mYsH5H64ZxMJCyCa+
84925qs9h5ZW/rQLzeXs7FnTWoTuIG5u6Iv2+ngdkNb3j64Y4yaMXtQR9n0WVQDJ
7L81M834MWMGAt2JDwMW/A==
`protect END_PROTECTED
