`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MvY5lgmx94A7IlXKRzbpGFRz+CiM5vbT/OKKrjRHcqbJsQqGKtjgztFG7Xiychj+
VAcC7ssW9flhDGG1do3E5g5HslUCpAo0IIfZtLGU5nMOxkz4UVV4Yqm2fUO1a2Rs
ZynqF4UnboKEwKKzZ+Rp8qK4USoTUcjdxyYTQq0YeZzs4dcdlQkrjeN029KA+OOj
xOwSAU8yq/miV4JWnov1KVD43sCIVogmShw1b8JyP4jwcexTy8t0u4BA08Ot/X/R
v8UyfkPJpNs3Vv4kqsXhkTsY9gRWGNKogukA0DB3Zy0593zpO5/TQ4oNTk8rH5lw
2uUpfc+vEpOFTaVEiQ+QaN8xPZk+lh8FXrSLjMO0mpBmSDTQBxglmLXCV2sTJp3v
c5itpVtNRk6Za44uu/d0dp7NqRkX4BYhNCq8+1MSYUN4HVeYUrNqghuyWIdlAWeo
Z/ais4g6w0NecRttNpmoFTz+P45Yr1A+lvtc2QA2w00JZxaibrGO5AjiRxEeZSmL
Tda4gr5kzi8roiAQYIbKLlkXBEGZfFRfqeJ++t3p3cmWI0wVQnhlw04XuosOQ4SN
QlI9dXnzX7e7Ac8fzxXRJt2uP0E8fPqPG+aGlGvKJ7NdkpNERHIwG7gvmJR+7cC8
q871SwBzt4OdYmCseqskWcJywCKtubtPj+8wjutgl4JZ/cRYAcF/EsLuyvrTBsvE
t2LbfCrI31Ej5oeVjir8/JRucJQNw3gjnr5+UOpB03adhnF8EMF37qV5bTG/9i2G
c5HHO4wqb3Z2utEpAYHcMQ==
`protect END_PROTECTED
