`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m7Ntb8w6smBNpzX51YF86HRq5unSIXoNoj7h6Cidc48UYSASLW9VZIbiWlm4+89/
5BUnCC40dtHDwpk8CuLBK7HTVNeSgMjpGhlN1HcMeY1BPp04XA2TkbUGEZ8oKT0Q
1dYyhTq8mR/J2EGLjGydyflsNIff9gyfPRSO9183pewSo6stze3RDiUBoSRR0GPu
iSUm/BzYZ9H91zXtZvL6qk19VqT3iGp0++ePUM6xqpZtIodWJ2Hv7un57YiaQjCK
G/Og05nhUirtK9mm088MyeNpC+8Cvn6KML2i/GfBgDEOG73pSxX0yTh3KqyGX33w
hzZRL3YBDMo2xq0owx5GOWdrFMPRLuxPzxMJD7oZH7tix39R00EZfvlQI9WrmueB
1IIK7RwNDhIYCcW/uvRHXdTbpo+3dFOSGV9g3I5N3WwrhtUsp/Pl9wpDU4DhAn6c
lJUCjs+ixUaNaqAWkIo6u/WF/PuwvSbs4tTqAizj+IrqRSiq/6flDEglpx+lRo4B
nAsAIbZLDkKmACva1ZyA86XpzndtECfx0+iZjiGcsfwC1gOKJ1TLfEXuRlTPPgJT
4UPr15SCDnO3zK5vUwKKPjnuftqKnQ0iSLmGYXJebMf5gZ6jl22CnSyG5RXOuhaN
vgfYsIpkO3kTN+5POhZ05TZkTzIIjtl9NfaTQsE8MxY5azkCasOQfSW9dE/DhGaZ
wHnWkM8g9U57qQf7D5/hMmkZbQzoncD1KfSOyOC8YQOZoIQnFFuobx6tqQDbfcAw
kUptAyWCSkbnPiVDzmMxFbs37XHHEd1z/dIbBHKXw6AIlrSHCAuSYpu/w1w9SpxO
2t1KVhlRDLjq/mB1uvVzPTKf7mGAkEmQrb6jIM57D7Mt/2y5HVXSCsVZoxMIwFWF
BWjC9ArYAdQoe8cjp7ViAXXV6G4bdOWhFNp8bvIvHoy47AR/O+HKxvF9q8oeH8Do
3YvZK5v8FG32EXF88i/f+3rm7UNpgOMbvyt5v/2JV8iyahsUwx349lka376dOvbM
TiPoqg4tCCw0Ippoa6YpIMJD0g+ujzqxwgRoKjU15PqRy5qSNKcwY1COuLIHeQOB
F1/3Gjpcd1h/b1zxDrh/n85hrFNIq0Q11P1AxC+IoXPf6raA04H7kwVizeDM86dk
GZ1kYvdl1dEaDUeI2zFFLW/eq3gmsV9s7qarhNNgrzfnn0OCQ/UJJwhNYE2RF/y8
LDccFVa3kFWDVZTmvEN7t3cLbzIx/KOumSLQaNSRHPlEPLr4U3NaYHoz07obblJ5
5xiHX5LKfKojs0Bhzx9ZV1hfOQdT9AeTNd58o18MV1PXOPKq7U1PqHlzYTOpDu5e
ufUX3St9Ci6ZhFhTtFuDg2KlvmudiJfgGzfcyDhC1oPfAalsbat4vGn9wR0AAKO1
QLFx3QgUpTsMod9wXBLCZO4raQ6b1YJTsCKk1t8C/PERrDJNw6NA8fLTZyxCkmkg
+vPq1O+pIZvv/U/9TAYG+9HeYJGL2CUxUguQFkVPcWKFO0mqgzASgzsWeQJVE1dX
eN00jeCdhStfq6pYZsSp6Oen2N/wC5i+BUG/3lpTfeJg/ip/ybng571PCDbAFrGG
Jt5DvuBe9dcVUX0ftbhQXY7UbSZ4RAavTKoJo5kVrxRVRIHlAL74T7gVnMURufeQ
SM3m6sS92wWRTO9iQC9jTdDPKvB0S6aEHf20/UZifWuLGNt6XQ3jZKCYoldOCwuF
48DdTqnIXpj3CT6QQOES7bEj5Ten71M4oRF7N9UD2zXYCqK3BCf6VL5VR1X0iOor
VKsU0EDNGi9reNIPURZTpfWw8JccZYla011T9snv8sz7Zaaj/Kz/TuCasAtn19yV
zCt3tohelacnItKifhqs58mbAkSjRCP8bGjR3huqLMr9yeGwAbQzXU5jucqcMytn
yiOYUcdob/f7OY3GEoPTvH+HTCewHnQTiRamAJrW7RADe+PHyGJLbDZRL0vLA0X+
3YiU63wa8pO1VWbqiqIYMY/mRmivGJxVBlKgbl3cqvfCT2q28ZFwk/zpRk/26TWx
/M9kEf/ZzpQxgua9RLvxD7wu1MKcze6B/l9m8hE7a7Y0NjK7FEBIEqp+CG/MNypb
T91RQfyhEEqo9BMyNBhMFI03SIK7XKomWxiWNVPABmq37WgJ0qtntG7HhuVR7buQ
uJaGxEFSPglBqyz3M/uGP0QrHZyUpYfhOU1YM4RITLWiOZW6/gxINA4yl6YzTNPo
37JH2MXg466AFZpR84kMLzqj6EHHDT5Pe2Dv7eO5sEwdKU12SlH1swx78Y2mhFUF
fINzvWr+mSbX075hzIWjPmWzIH4ycMxrjbLCchMEWnVdeamUbTOApoofA+pV5ayx
Z3CWHvIKeG9dG33xkZ52esO6MXXh1COqwLOlqZ+/fKpvdfuapERGtBUCOcgD+Y4u
BElOPtz5Qt/iCjcg3Cu1KACZauKhgYwzQd3OfjmSBwWoXmiieiNaSDB/fJ1z7feG
y4gGOQHII4LWKXuB/Y9Nxyiei57no0WkNaJPZfv4rMpuEYjKzIobrs3pR2PVV5wz
/r3jX5R/AXHjinqkFmMXGNZFo+rZAP8MVwQeNk7i0g6xRSvRZR4jo7Su4LyzMvhP
mVy8woOn6JH4c8zoPNiv37oS+mBo0Jy5y6TZjcS/rs7lmRqDp3GRUvVK2CO5ma4Y
0N7+MCy1qJIQMphpZDgskrr5KY1ohumt5DDGkqvT4tkXJB7bukbKF8iwxE9+VYtR
54z2fSWyeiNOuBWvQYKt3DMHQGk2L9jnUxqg7T/49yy3wocSNMH02+oOX1KkDEVq
ydncTe2zKGgem+Jd+GnPTAAwn6Pwxh+QR27AVdph2h9Lsyw20ICNJXIFYwR2OrnT
dAX+hvFm56qFKgc2DGXXDctez6b+Vmgwf57VXKdlfLLBrnx/fiqbqMIeWkFQrItW
O0fVUW03hJIcqpxOtO/RN2Xcv6XdJ0VjV97T8hAvH0CqeMGd6EzU4tfZfiKKnTNN
KKTnux4gZJolxz2DRuVVapKBLtqOSqbRaPoddL7QKjcshq0AVuTQ1iES5pVNXj7b
UY+2Mkyz8SzjKxvoqn8FZ6iVRrtV2q4nUdKb2z5qi9neHUxM8GOQ3xk948m02Bgz
baexIuMym9bjyQyTMievcPnjtPgFrUEy0V2gkTY5Fa00GRTEUEMpsKe+6VMVUQUQ
SUhFbZcd6I/0FxmlDuqQkI9asdQSpu2EToMv/dmrSfdq8r3loBX+EtxsJAfWBiNi
F5pRqSBMgWxAjUVyYs8S3dlIFOk7094mADiOoABqMGiIcKKjQwGeTMeRW//iU6ae
6A2B7WsN1qQPt18pAhhBGYegpTY5XMUrpXqV9nFDWx2AafMKHtRJy0gA6URYLaUU
Iyh+gdsfRrrbQVkwfMlZb3e6pHo4i1NS2F2YGUlTYP9ZEpPSoQRDUFQQMDv9FnWY
T+rKgNSbe0y6jenAfAJasIES1C7GIqkvKsR+phcRfDiWyrNWB57zXgAn1AXW9LYF
UpwdhfLjRRgbaG/32FkjzUfZNaw4jynn85++pFiIFqA/+1HkfMsRFBov+eYaklpQ
n+7xoluuKY+RlKVDKE6exAXFsZpx0KEleJWFgtl8c1sSJu5lSDU+J2Jauk6aY3ax
UjVX1grDbvPdZbWhIl+BqruEpNKiOi6H57tmc0AH6kuowud5dqwFioF+agPZUg5W
CwvIx/ZLDXXl3ZEXiwCBBDPzVXprs2CwDc9xOEItIo96GeayIPuziY63ul7h2QcR
Kg9oczF0cq+SY6jY72nifSPecQiCfvHbo2PTEh6iEnv7QAO8pnCbSz0tO88icLhU
Wov8KJvsytlc56vTF9pZ0s8Uk6IHSTXIeTcGc6SWaionPPHBFy93Lxlj4dIxC/qG
vRkRpMESFkC8pd87kyLaRm1cDCoeuL8zSS9flzIQCUjjyQRsqMG/IuHIwmvN9+CR
zJPBwehIX8G5kJoEcjZgWqOQp1hjFsVUnI0+YwenjMgxJgu5DNhqoYo0IneWplb1
VPw7EgAp5g4RpM+0aO1haJ8TKyxh80jUnoiMW7GLj7ca1mQxa28WNBEFxlfzP8U8
MfVRVs4CgqTGryRMMUFYOMqrJdH2FFwamTNN1qKZrJ4w69jnx4fdqCh0DafsByDc
XDduVH4BKfxq+8dJPO3zdcotaomByRRsn43NHOcBifbRYdGAOitcATYmxPs6VYCW
I4dQ3EgkoqNP4SC94djSKGKDzHuAI8yuaXxVvLQVbyjBuxuLLFi9Ys4LgP+kmkax
ggCqojKOim1yzItL+g5wvH4105ooy3n4awxj0YcFisoumZOkevQdlkIMolk8WkpC
ak9re+kVrbOQSAguIVWwtPgPWYRBaH6/cn3R1pj/wJYFydgmSUAHDHcCKDnCzp9B
Nu5MZRZVSYmccfoJcRCFq3cLRFI6QDi+wDpjjAYHdJYY34cDqp9hLqjy6LZ1lJBk
DGAqNV4kJOWcmjd7iFn5JI3kLn4/RWxETsfDVz8oeNmaEeVEy4sj/HMoRUJnbQuh
HdtfMP+gBBtcfMpZDr63nHwQ/HbIvVBUngz5EFaNRLQZ5I1wOX+8ZGEv8E9Ia3QC
5A/Ljv9rEcjoZWyyP9k7nhlew/MmYMgmTB6Y1XLXllkgrYz09vOvar4VGA7GGBG/
JLHUj7tlOuFMjVBperXJuN/FqK9cUcijPU0YAogZLiOFIPg5kt8huURDdLI4hhCp
bGIp6JH6OyQvDMGa/FXbU+ztdyyGx+5QjrJjLLQDJxKaBPKN493yEuI9fXHesbgw
xrHeLYO7B8EdRCA/T867r9okyLBTpdakiNx2hK5HbedWfwo7P8Y9NO9gC61q0u1q
+XkXrOuvHiU0XKVcITzLsTSVtf1qvuLuZBs/FpquIdGnfsSQruk2SIgxqbeTzrdi
7iEf/yqlqS9dSxPxHez4DsKfanzGt742bmI4kyhjxNZbDOUjWhU9K8PUteCOIBTD
t7uhQiiHz4+T5zsPMxtkl/8fQ2OchVCZ5ohyPzPp0J0rc1AFUerK9D86Ldq5wOqW
VaZOaiN8FRI5bHKxDrVUjIqYtMI1Q8XiceAEFq0USWtXXLJg3tcXuQGlL89t2oRu
uCMG+H7hazT+ICkpzn6082gljor+KatuyLmjBGA7K5Q4QR/kUqsNiGjtHWlovVpf
m1bYWSzsEWXABbjCHAksvIeM4ljkArX2kCXxtVaadA0QMCE7mztMI406mY9KDDDj
zDXVujfmpUjgjUdhAJFTWinFDpCT80z36gVdnzx9CPZi02Ah4CKjA8p61eWH1pjD
4wowsX/Dh+6HTuT7SnKG8EKZMnihoPzNifSi9FEJf/zaYFlcy8I51E53FY51dkmC
qGr5AbTvoOz9fk4r8zq2U0p0zVRaYJJCuPA1CbZUUmo1TGeHdNvdYcjVCiQOJCeD
FO6PnLsocFVJkMAo1UpTZcCQXhk1EI9XOC3eibw1H4jLk5+vtrxCpdOoyCWGqZ3C
C9ymkn6WD9Qv6o0M0UsMkzskCf3cT6ncO/GIGY9QFuoaWU7MMSrJlmiEEBI4BUqO
gSApe186Iy8BLxgVKONCukrHqO3KmPQrYK9tImbzv99nKHnwIABzKaW47rG2BUBJ
9dEFIaPJoqhbWKsZmg/H5X+N50hpSdhWt2LVXqFgKWtJIuaPSp416EPII9XR1f/S
vfnzLzmUEvQgQtx4tu/I1gfooJ1FgMLdH2gxFpUtmEM8gWO7yZJsQmhAFPUiKvwB
w+/lTG6e4heVZeqKNbrWfuPWjI3+1vMD86zyPWICkenSvslOl5jc+z1CcxlQ7yAb
zmS7GmvhHrfdzl47of2o8yAJgzCBRSpVM2/yxYL8rPTbUSC8eP/LCPn09EFBExvN
5zvDlMXp40Y+abXN/058sbvdpn9GYZno7nUIQU0B2Id/J/R5F8l7Y1IhuIzUa0hl
N3nUAMl8WuDPkWHOvlKM1vLmDA/8QouZXfn/XPq+DHzIPmtO7m89RU5p/F2TiJHq
5WwICvxwbz1APQ0HGmKfXtUzo0SrqfUtSRVsV3eGKgEN+Gh8ZEKTEKLAnUeBYv5u
R5gEP2+Kv7OnMw6icdnuYAoSRCIMAQvjBFnPOCk2m3VFJQilNPtUyi0mHN/IJ0IE
Vq8nqJAdZ4nGeG9UpSZ/Uo3pcu3JthMklOozXPwNF3m4p/gogq1GWP7GEVbJXpjc
HBKPrLEzf/X22CkIeTKyQhF4LH+J3ODdNuWL+XbniNwAU+f9IOWOxjL1F/q43ImZ
NaDDvlwOAh//QUGEQr403Zh6oJQudc7/KSWFPO+k2I98ag9HFBEER5aq45vxGFUT
6KhkWMeQhcvgqUo+a4edbVZJwPNiMmjfuerU5t4eKP4WtYm7yKGn36cBMutH9IPG
70P/VFqqfM+luZjn681WDlcJTAu6n0ZScms+1LBPxQ324AC4kxgsl7zUVROEi9h5
7RWFGLcgTpI+V6AeOj9U4p/5B68TLA9yDQCyFeee1euAQ/Zvn/KC8sEHPwbK0tgs
LdecFTrs2qw3QWRhycDRXRC9EwxDQhZID295WPISOU59hWo8bhXCEZ4I1vmVPhkh
ewxcHk4RMv9vG3+hIlPHDw8u5g6uIKDEtpQP+QdY86h8ePVgo3T381SUqj7G27V0
XMxFHs0VvqwtyjSfPaOPe7o/z6l+iPbeDLYIATe8D4yjoELVZFBwD3/rh8ttIDUp
zxW+jxFTWGlFy8o2s4Jh2dh/BLk7lYuoA7xmK7DeWlGik34mJY5EbXOkJQLBAee/
dRxQHGtKlF/Hlo1F2Pss900rD8FM9DSdsbKiJkRtK/wis+7rIKP8Yp7ScaNoOG3U
7MgcdG3fYHIi6F3pEniIBt49sCzWT93Nq4rCGkpBg7zUlpQJpFCGhkS8hlBATA6A
LdGcAwBgj50SQHSZ/J8BH7FQ8NhdzwiCwv8znArguyVTxM8mxs9Z9yV3lirmPLgj
munyI9dlLePpyU/KznLe7aeIKogInkbX0SU9P8K8n50AnsHa1879OdF3oL3Znl3a
7gVvdGDhKRuOy4L/Xbi88T3LLwIrTBT8QHjMGIQxHtL0ZqT87qsyHBuGVx79wYOS
gCY4pWwZmq/JtOGXUCivbrE+h2XT2j1KDoNdNQeeaRMV40xIppz05Zg4PzJClQ1n
Yi5R6Zn9LF2c9MWKJxjeCHGd92sZOEPkmu3BTtGYXAe5J9UxIHIzjbkkq2v1ZWBk
XYKO7t16O61EtyZthWdnqJGQaaEUwfPC+mDNWo3g8ZqwrC1tjGI/JTNry1B7p+6u
09fPn+tBBstwhXVAHoO+xo3zPYLHCc27RTm704XUCrbrib3PDZCsbDgK3INmHh2x
vx11keGoKsb9logGpf1nQjoiYpWIn/sRDGl9aa4844T5kZGzhNqs/h7t2ihxKxO2
4yqNOq8lfML7fKEwN2E//peTVyu3xNLxWv7TdAhMGSjvDuenDT6NbP1zVByHsClH
Guw9OzVt7KUAhj9PI6QvOVm2I7t/X1Gb8npdIXoqCSwJlU8eyqejGiaYUILIhlJD
eWqZEEaXdzY/kem1zUwrxNaFQ1hNPLFt/Wd7HNZebYfFuF/hBubwFMreRQ/f2BxR
s4V6Gyt5o6rIseRGHELRzFZ+FWlHunPfEELSBnv2+xqXcTE9OPwZ7+qCVU09Ecm0
STvfwFoYW6gXP3on5gYxxxMys+qFyQ4OUpouXVwVh07kpWdr+YXgzy2ExWLi8a8i
BYB4Kn/8LTxI+MdnkbER2/7X0SRRDrvcHWvg59vadrbQ8RYOuD0OLOqahR/IcpnZ
iInEAdCfpFeTBoLsglG6r7nEWqohlrkYCVMpgN6apeYlV/yDdqTKf8p0U9tGolwT
wfywuYkwLzoZejUtnSyngfIv0GXxVETyx3hj48zPObvgqpu8Mjl3aa5BRp0eYJ+r
61u0ZASNrxcUqs4Zq8iGUr4c3+bncNhAF/f41VntkLBrX9zOWYd09+t5qHEFRX7T
P4KVQSjZQK6oj9XxbtgP+a9me34+vNQogmrcGOtelGKOg1b83n1FeSpGAgc69i/T
JZ3uNu7yimywc5nSCGtbPnxx3I9COaO5tKQuTJnLKBQUWqsIdlyui64/FJW8DDD4
Ci+L5R5v28KHLOL3xanfHCa2gBIgZ+8BMo7NDY1oK4J2EZ0qz/V2JjbguFSZ35BW
JRQBftykITVJmAYa7h1pl2uCVpXcV8Uc2musNiLFmp+w4dOC6/wQIfw9LrdGxH4E
YC28xZ7TBqeetRR4O+uioR/9mGaPYnStoYj2mY2GR7zWzanbiZS9zqGjbE4lSocn
v7fKfbWsLq4LmuPteGzZn9W9JQ1L1Fih3xxYYmLp7r2VW1mFKIs3/7RPGEcZryXe
kJ1vJd1olHAz8A96f5iPu55Kn/fX1bOi4FJmRQar3HozV5cjAVDCrnordp3uAA9R
mM2f99+vY7PsPjdlABR04QM2BWCA3shSnzu4XdkI0Qt9WFeeETnA0H+on8GHN+56
NNu+ANgbxKmyHzZUs0WKwqWoLkTfMpEE5uYqitvR+gxf/EBU1+glbYChRLPELyKR
SIRDnWq46Y5iAGkuEunbCURVgU6x/EJSR9v4+EKUHM7lYZRSae1JunGSTSAqikZj
vYYFwmyWY+0vQUt+df8yO1lKnm5syHothqo6ymcNUndo2vIM0+oIjg1IBJJMQupQ
o3VssNyrX7yJJlZgTdDSrSIyvQRIaUZNFJ+5nXFPiw+elg9Tv/6xg+CCKtCpsWXE
TUijk/mcci0feIB7TU2TeUqlA1uRa+XyNZo8WJMRmE3aDe62cwkWtUMmvuFx17Gz
ZPgpSIX1c7RaIdk0q7nh8hKqwHu5/CXsigqvV4JmkizQ0msW0U03VB7/1I0qSE1x
2Z9RvFHJfVOK1sIi87wJ1NisRWK0DhjYG9vLMgGZD6RC3eX0RmkX1OjI3VBn3Km/
fsL91EVKGTFdenZeGJMnxHTJqAXmUGMXDQlMTXPp5O17VUukR9Iv6v9qRmDqxcjo
Kd2Js/BKSbDeqcNrDXdhXgcs63w/2M6jW8KVxZbq1V0Ntqwf61gWsUgF/UjJTtwV
26LLBEM7gP1F8zXFchQHlV9spyN/cUfMJENqqPQ0fsh8zXeR+9B+xrT7ZMGTkSYp
fSaPuy4ylz1rUTIAYliJiFaDmaHIvkCCb0mRYY5hp0Ed8zEnQwJmSQ74E+yPsqWg
+7QNc+FSPrNcFle7+Y5mZG+ISSvbeEiHveUQgM0uivYWQigaNqP4eTZV4yP8J5cX
Td4By0O+DMU2zd0py9EtJQ0ENmp7RirP5P2kYgnvq6iiZVph9iVyzJBkciwtW5Mx
qeryT+htEKOxkl6mkYDMNAUoRHId7XUYwPPse/kLF6KqRPvhT3EB6sk3Z7E4xr2G
TcVkAfJJduqqYFodLB0K61/55RlRaPF2Dw15v3tlLyVVVwrwuTYAjZ+Q4qcRB4/8
7OGjYwM2SthDtXhX9oczpE5uRWBkNbXPva7+L00Feq/qbqjgbId4phWquwOicnHl
ul0+cJDJeNzESULlsVQ7+ylBjxkdx6Rxau5YDokHpEs9RC/wsdG8mn4eJmDDhcnG
eqI0UYG21nm6O7BQIsInC9Ol18Y8XKcMWTF26uAFVgMeursPee8OVWeuZsu0Pu58
Rl9Nu6XC5GQe5/Kg5yHlSrQhzeheoyYwUwcRbPzEGeN0LeHf42ajxbJ2kLJE+rqF
DyI84mVQRAPXRyWdLnQz4W82UIn6+lFGcHGEmUzdbQlCvHreSvupDId65Wq2Bejm
sKYGpwtuJ0Fd+iCn4QgCJ8ecDeVhaUQ+cEaJ2lctnPrgck/hHV5nN9ZvkVJxWOBp
R5x0ajfW2mDxG0YafRJSWlRJMa3GhC2QhZJQ9ip/SPukQwlnT8GUoySHnEL20udJ
aslqhAhcZ2xCBqQwhVvf5gu3SwGJfXqXHzM1ozS81eUE0M3Kbnva/wUzz2E08VrH
g6gcViULtfoTBtk7vuodTdRbdaVY+fRHMtV5gNrlb77/BxmirtO6Pubatc/xSMT3
xfa86GdAj+xzbkLR2hSTtWh6ptLq4jMwpu0LEvO/NUSsdNfxfCG5f6er8IzS/ZhM
iHnOBwkfDaCAW8VP0f61R7xusYZ9N30Dv5lcdANx3uqtF0L94p0tWVQdcndPwgkY
x36iobNlry8HzkeoEKdWlD+P/Ou9gj+SZy085/O8sJ7qh6yy3rLb9cw/T9abIaMZ
4AyDFjuDEmNQ/tK6NNLlKZXqMH+M1OrnplQG7pdT8kjmzA4oB5NKlj+6/pRo5meZ
8VVBzb65W7gqIWjvPBDdreev1qwoJyxKOesQiSUN1aIES1ntSqOZQe/rDjABhoPs
fK7rvHnAg0m7YAejVteom6p8UAD+Bjjt1u/XCouNMbfxXXyTXHREjg+UFzREpCfx
NB48W9+zwlsiSHp2ur7p85ucAkAKHhqlA3geVstoiydtbrTLhJjuas3t2k+Y/E+3
UHz8fiRHaQP0xbhOgbLAtgZiSDM51VGO8s6G1AeiTLKGgHt51QXPj8bL/BnA8hFs
40B3lJ+jk5bT1z09y1ztkuPqZnaHCjheoSGobjhqQZtXcvA32NUO9MG2UAsPbN9z
c5OvAkt529jqfIQZEf9wEKPDWKxUr3ZXUsTvTGtvFghvyTjMd96xaMY/HYE/K8Y0
LcLHINxK7Tg7ZVyztxuxCEhge1AAgOxmdCEWG9KXSJAcKw+d+Zp6Fcmau8D48tXn
GzkpZgo34+2Gx8boCUo66UjYmwutwLYDvPAyH3fPKmWbX5x9EQ5x6d+m7HuQgbrj
Yb4xgAw+VhD0Z4shYkFmxv+EQ78fthjnawyWVO/ins+YElq1SpiValHMOE0s7zMB
LLMLD74VahcuenkOc64Yw47IPFb3dR+UGd3EiExM3+B/QU5111LFuHmVhk1me/zY
v8SbhhjlG5Fdf0vItouxVAkbW673q7FO1vo6Aa6V5GhXxINhmyB/aI0r059slfAJ
C/+ZIQFAmvfuh0MoEhIGI3a3g7jVNseZZvB6SfStPGHvzDAnvWf3bRacFq37MpN9
H/cEXWdIf3O6VqgwyfkQoQcHFVD3nt8DQk3jZ5KsBbp1UXU0H/dYbecvFQbamelu
DuHw7HzVS7R8sglMs1ijtRI8ai7TidzeqfeS6RiH8UN9MeJ1y+RhlIR1DUAXszGX
sdMS77vlV96tqrKFH2O6e+9LVh4yzrqLQFbiYrZfvxsoHcmlwM9y+1I8A2zWL3OH
jTPa614zAnig53f6eAWrZOTGyPaKsG6FQlThmk35jeOUeUq1yfj65AkX7nJCbEff
mVO1OCQ6GTvR8yE0vrqFG1G83zG7xKuLBPfQIdwZxAoagQeU2y2HQ2PEVxsYEcPS
9mPgqQ04Er1XgxB8AgtjwSwAfY3U2WDRZUeQdnTHdPCVCIeyiEOuoWYW8ECN0u+S
PR2dgKpqh7/J8Cm1Oo4tlkDZ8EBkCxMYz5pLkn8aHnUPLB5leUR3ehja6mOcO1Fj
D8jjKvDMqZofL4K2lVSL+KtJlx8A0pnQ8LFQDTjGWKxYyNi+msaL383mhu2ZqFcX
TBhzRLrgw07tLeztVWPFeuo7kEqq4d8ilfu0kczMHuKjBleNdP6BcJ1AB6NZjwnI
18r1zlT1rezlW/+PciO/O7eF75UBSUGDNrjh/nIVvRvAMyhR0CU+9NdTj4eA2mcv
0YIwWLp59uzDSf57q+YBhFZIp81L9SN674CEMIbZYVr2PrznTgnyqzi2dMgzPTvH
7chl1vtDwYBpW3Ncav+KIZ06RcZHDXhKEar0SZHeTgd1nf+1jaVo904XsiPZr1SF
3hP9sdrgb6PSvs98Bi3Uq8lEAY7AE2L2edmwf+hAOwFNobHgiVa2G9WNVB46LwtR
+QPEz9jxzGB39e2M+mTIqMpxDokG3OwkcPc1hTuD8PLdzeT8Nd6zsWOYQ0WiWlBy
msqLh8VLJrd2I1kRK+0+PL8qP3t/bcUsYNwHHGK8sIGTkOf1V3gfw83GqW9OZSA7
MrgEUCczP7Fjo/jFszdOFWzBOPMymViYspv8nxk3br6vjRBz63yXvm1HaLHAW8VA
RYnAI3y/EYoSQtov2aIuJRdoJ6KwaJ1aSF0J/B7rz+DLpiSEF2trPQMxhY+KcWN4
9kPirb6cPK4qLN2EhMamaQsFl5BRaNEipUlYXEFV0T4rRSVFPtJB/nF76G5ZtgTR
`protect END_PROTECTED
