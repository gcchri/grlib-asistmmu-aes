`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pX7g9FXcMMWq5MWwctJVgLU9vnjEpX+s8o2p6QJXtBblLPOj9SE/ysH69uf/pxgQ
HQJ8Yk8/KiBIExrw5VqVX2mDEWc++tne3JjSsRmMW6UyCGvJcZhZvwdBD0y6w84w
pgVRKRj6Elu2QQGCSm+5KvAcD7if8GQoAN5O9t0JDN4hn9xqNtOw2XT41G+axBNy
R+hxqr9aB1n4fkcz++EyU1X053ccJxiZAoWMPWUMtthxwcqsobDyuFHxf9WI6JTl
G+3ZCtwnTFLmT34SoLKo4vwhwuWfXdS7y3vtL3s93aklyHtu4vqQelBlBzgMiGws
MbHNlqbowc15i+Hf01eN/Xo05n9yFX8zF0EjGmVstIgmjBg6bAXnbi/kBZlBDPiV
l6d7qR7dfmUF5v6Ie7L4afANGc0WKE+5nAk/HQAUONGNW1PwfcrMxqXClqzBFB1v
R7rtPv9k8iH9n1i7CJySI1hgquqKWGxaYIaLA/k3aXQ=
`protect END_PROTECTED
