`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y1AByTu2xMjN/d8NgLRTHKsqBBGE1VqW6rAvW8ITUKrX5IA7KYz67sHLrnksmf7c
xUbYY5g082nQfY5ENRheVrZgrxxhZYvnHGjg07Tww5LuEevP2tK4h3xwC5lEZMx0
+qxYJkmvgbKgrscLpnJMaG5b50GNsS7d0xFJcvvWtwrd/QGKiOoAWEi9a2+Ego2F
Bs8kVYf9IhpisejX0O0WJVZ1JUGYFqCai9pFjYrSRv6OzOPcKGFNrevS0okgQhXE
vojwDXke3YLHAn7OiDsI5sEyDiY/maHdqE4Lpu8yH3+PlSBWuzp/IImsA6wTVcOo
W1d8jbjHyB2aKVdSxCOtBlPzLix0dDGs3+nL+QiYrs+LDZxt9FtriPfvOI8+ExAN
bQNAn1l+JG/Vi6586PP5/QF8eIKfZX+SEHF6LeT9kO8dj1Vhh+riozczZMyEM/tU
E5yM1qnS2LJsTmvzyT+h4jC/qXl8KgVyrIukv7HHDrBYwYWwOd61d/6HL07G5nJ7
4TVEVVf/0BaQrIwrx6xTjgye34ILdfXxI5GDSjYPZuxkYoqNZ33M2Us3ugcB5FJN
/BNyQAjkXv0gFZe1wR+qV+nqB3ZHOdn7hwbPzouEE2GABHHZns7Zxt/oM65eCgwK
+vPn649StlcuEuvu1m6RnHqlliAlNC+aYqH2wqPkfEfvOK2aC7YAdlXhx85eXcJN
CT7BwK5pm3gRZC+upLgev4khcx/IbmChLunfwq83hMPKxJpzTYtU0HYb6dp6RXi+
hWS612fFGUsezLx3FFEDDscbG6lmEeSp96xt5XkD+dEy2NjRvEENCNiVUb9iuYx3
rwggt+KaOQ+dz64WY2dc3O+Yee8DcmNOse5WCaJpPa9101JsD03mt2FtH3fbn9K6
rqnfEu3kw0QkfNzWwzhqjtfFnX9mcQIxZ8LvW9+sMt+7LxfOt/N4i2y1JGIxTKhO
UbgNAgrjyfKBaR6xvJEdvO9mjTqFPrIJ+GW3LIjT4CK+EoUH82gRIuyRzTyljy4T
SwMDPIimodhIU4Tzd/3xingMreP51imGXizN8taE0t2zlw2b2t9c56Bnr3RjO//v
DrZl4bOJag3Jtc94kE2+aqHpmfatbeGrOv8EUDtrHjSSNLnb2egIaLACgR60FLy/
MT/6vJyh3j/PgVHnf7DZmoC8Jkwr5E4yDQawK4y4kh3PGKBXMDuu3TnIOiPmOKW4
AwZz8fcWxsRMCs+u4qEDocBblBvncFAX6owca1m75zhPPIIJ1Du1G45+0G/5p4tc
u7OaqhjMhYS9NyfibBuZvIjFMiJltRVA3R4Fa0myXjAd/WlNAKoFms9nZpaTLvRL
jh4INQjTpjf99AaroRQaKffMeithOG9pyKbEBpgFCQQG+sANvrY4Ufj4VzdiO+At
`protect END_PROTECTED
