`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JRRbiaxUaFQU2q2swWbJqL9iR71s6FiziDMb4vvI7QVfOSqk5dx7cXepuao3NQAE
elA32KgZG8DXlh6FEW1cXqI2NkIdOBhkItchUmt3hWnsed1EywFbFDyvj67m89WL
ZlkVAqgIziujE+fW33Psr1++NvFL9FktonB55t7IucdoPTaxxXXhEs6WyMMCa7DE
aCFuhR+aV0jUKOp+HcE2GUExAfDLMNEmvGzh9+7T71ye8tSUTJNEKZbsKKRqYFCv
4WIPty8VjeA/xQ4vIpnpnToWRHJXyRqaAWOagM3SH3kNL8cwgi7ahMmXsPACe+bw
apdVHDC1uzg96M1eLQoppA==
`protect END_PROTECTED
