`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V8HvR2MjDlTvro8JIS4oHuxq4myNa9GXpWR6m+jIAx23uQZqvsddB1a7EKkoKOAA
5Gtc86ust4ym4TWwZeQ25YdouOIeIynU0E+uM8Q8XkxAE89F2afGTwo26G6+zKtY
IPLqegJC5XPFIxeGnnpKuTtkkzA6PaZtaTPzcxnNcHW3qxXDmhiGipimP0I9gh56
PvzOI0fvJoUlXMxAktH2XHqvOm2uKb2ig10J9yf7+/3CLKeG7mJeKvfndX+dswbT
G15X5L95nopq2q2V6f40Hss/qOKPCqGf6gzH6ZJ4/ZH5oPcGTdQf3PjXsaFY3Od4
6FN4E1UJj7SF2EExg8/gI3wecam13U1GnkOpwxpKFVXRjkv+6dAWWuKG0Phjvl2/
ZIH66BTCHzldLYe39Iki0Q==
`protect END_PROTECTED
