`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
scbrnessicGfs9fve/pTaTU9nigwNlg4kCX/A5vTJD7FvKbrrj+djwBVcDeiao2c
K/KFcx9GQ57HUF0HDmU8+NARu84ZYEH/D2To1hbNDw8ta9fw1WLU++bjN0C3oybM
IpAQ/0wOlmAN2muVAuK6ycPGsa8h/wOl19/gUuoZNmOFTg9Af3qowrXVhxTeYm+U
P2zchN5YHMnWYqymZdnx4rOSuCvRw6lerXtjxKAxAFEeVtf1ARjT+uRgyptvYb6e
KeAb/nR7JBoJKLUvcGp+9A==
`protect END_PROTECTED
