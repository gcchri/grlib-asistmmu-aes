`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uG+MMiX/9z90WEVe0FBwmtSTAAs0cL2RqK4guJl9xWwlhdYVmmqz7+6m8r34Qsum
BxgHs/9wflXzIp2RH9IRJBSVxf37NsuA7PpMD8INcx/JghhXBmCaGlVbRg2BmcEz
Ey5zVogjBZHAqPkTSEC4SyZkoF0HMWPcxutok597wAzpSESx6FDR6LgSt+TV/8kp
DAUHQcmMVitFxG+Nn37A6QKpSeTM5EenUDbppFT68Gvy75NESnzN9GSCqRII+WZ4
l6IvISl9E54tsd+XQ90n6Q==
`protect END_PROTECTED
