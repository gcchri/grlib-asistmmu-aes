`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m8kIN7WWede/Q035xCWG7aNaMpakx11PpeI8sxDBj4NFRv0Z+ULvXu/wmuA7jMjA
ZEG+IwSgk9I6GmB+Exx9Uovk9xLCH2Ea6jPGlEta1G7C8rkTvPeo5Va/W+xkNW1V
pCaGkhSVv1nSR70AmBWoqbrxOm0dWrg2jSbiAEqvuDZGe4klmx9Ig9vZQtA1gBug
rsl4VpZM+B/pNIMnERxXRsVATcKcQ5iCiruPKoRDNqO3atRjiqlpdZ09cl7I9fLe
U7WsQyJeCCGNmu1wU4uL0V5irQhco21JEaubbkK6u7Zfs2Z15qpgAPLXOMGrfPSv
AvM+5jnCOo5pqtYxO2v4ms32FDLiPK5xMMaiduh3jf0VSGXsZGsv43EK0UjBSAs4
Gw356DeHNhFkH5dhy6JriFD/R+rWlR8cPFkjFS3+QctjRnQHuCeqsHZG52ei5by5
QFO8/36IjkbasF79t8NJlO9uAdDJNW1WX1rvjudgoa/G2MYmfA6Gg1G7l+tUEQf/
Dq0TUlHVNuuFb9RgeeX3YO5mtelcArt4IuUCK+rbokjb21nINRDelyBnUkAjqL0B
SKk5b3olypp/xqcnFIfLYABFBWSd30Cpj9DFY1Gk8TDv5iS6MfYRapzQxAw3HIiL
66AP/fVjtQZOjylSa4dEO05PCaBM3CsNhXBTfJa9swq00a2V5K77FB13o2qkg30O
n5YjU36yRmwyL00+mYMYE5l4dTnfEqDCrKso8NDRHLqMY6My7u1mHnp6e+GiwDG/
yjC89HDgWx/GHz5i6FAxTLKqJrgUYS05ZQ64HaIkNDitt22C9mxk5nA/ljMa4rxk
/kR1fo9I8Yrcaj5Z/mgXOHZhtJblz5eFtV/1Y8PGP5hNud13R7Hjf+SmSHYqIQlO
34t2RP6gozNO+weikm9gfrQ+IK7nsjg7EATCrOWJoOK5fhmURXRi7W0EBxv2546Y
6o7E414McyizjkHtyjCbzRAjJKOSzTio2W/EGFADboh4YKteVzcigP+4uM1wh063
CFj/VOts+opcapE3JR0zYGBxmCOg9NpP9J9faUE6tUwKmRLw8HUNvwr5j8QMfqNB
ruDBxGMQgCUmex7bqMZ1LUinSE/WSr/yvVTKH6n33SbOSKaQN4ZM17iPskVx2bKL
HyBBGMdwj3vWp8jDNVUevypuD3d7v1m8Eu2IdYyL1GzqSYadLAfqF8OxuKko9P8z
PIjeshjQHsajUSHfJDTfEx0OqkVf/ZOu5IevRlwB3L0e/BmprlRM6sa+1FF+gHdX
SvAjyA40P8sExrJQx98xpTWQz3GQCKbDra1pa5npRw1yuJKyQKN/VXzkfGa0C/wm
Bi/5U4cX/bOX/uiE4B1XnBpvuLxBuK5LIj0Lt6kK1qglTzO4hzP7Jg2rI0BkBU2r
70JqF6Y9vVUhNGeD2grSLaUqZarUR9xJ+LLe3TIfxW89i4bJKJXGLyGppVKaBG2C
hlTXRvo1u0aK7rRuyKm0XKzRCjtG5NRrLUfIbwP/AZror2SP88IICiwXiYtj02Ru
hD7Cefb0RXyCKE0bfwZAm8VyZ86knSQXKC+DbEyyfS9DU4IEQ99iT23ly253ZYUD
0KEfvwtTmLUwCCLITmndfRCTApcdzT2VkBM0YuZyQWyw3cI0yyNjHNgIrESgOz3A
m8TCI4SjcS87CEMOD0BK24uAjE7gns4btECTULUMpMmHcqgeQVWdVDojvnIGNX1I
4splwBKwt+zvSbhXw8+l59XadwHFL2ZsZS54RuEc0tPCMlCUYhgfnWSlg1ya1E5P
ZIRtoTFxnhZs7gG9REFIZdDbBkk9QzkW2tjct7r/4eIAx1ikmdIMCW4WZR+TJcHe
6WU1yrC+CJ8J3xiLbUSofHraic+FAWyzR+EDi2PDjKkpHCPjIY7XGwW3ZvLIch13
u1lzV6jVmCOlOeM7W45Af4BFLVxtCpO2C/9nyghdtEilwtj4dMITEet/VORDQ0I2
NF25a6bYr8scVkVb6P1DRV8EDge8nxXR9Qb1383ffuA3yvWl1+/7x0KUzz2lEOhP
i6W1OPsoAVug+m0lbVIc72ttG8eZ7BL+l8su8S0/zAhGuRFIJKTD0VEm2Yc6ChCu
3Qv31kwqj9eNsSp3BOPZBqy/hFpOC97cm/dZa+jpXb1oFPkkXiygz/i7CejYejwY
n9deBdkYNVZ6Rv/yhQsUFe7Hx6WdG7xsV1d8VB1LL+xtGRp+ZJo1oDO5weWmVAqS
98dzqmWRL/GLH1ONFj8vhWIE8jPA6o8PmowpkY9R+RzVpra5l7ulwxYCsyvJiN+L
klJ77MGx/to2S5qXOORNGL14wuBFIxBQ7eger325ELZHp7vlCPmDGGHOPXflQwsM
RZiOrDqzKHax9uAmL/FkSr/gF57OiMRg8iI5/6gFYrrF0Sn+Tn8rVvVr1YFm9Dc+
MGPRoljakUtP9Ra1khIM6f/YVEHdsy8IYoWhTRzbjhk8XFcLFxR3IQ0/T/RI5UI4
PsmLGyMOnHzizDs0ao7dUtn/O+3e2OCxj504wREve+PK9M6IhfTgPy223WFxprsN
hKS8iRz5Cop9hUMx8mGTvfGaWzyzL9o/g5TWOfKGQq2dElRpX/R12WvHKVJ9bOmd
pZ5tBHH/kTGFwe9tRx1DlDl7XI0ihsOYni3jFT4gJu3X2RYglbZL98LCpc3oZCyc
Sx5x3IXgtHNz9fSr+usZK/0CMmt8YRy9SbQAmveaZyQOWKBwC0SqS6mDxPvHX5vd
znFrEIRv6M7mQj0MpuaixLNTUvp0nbrdWbwvTDGOuQU1uL1ciFopZ81DPd8/qUOO
Fdv9nZHWGOQG0Pc6cToJbPVyb9mN+XzGDlHTUTLfC0AMURY79d0EQ/x1f+tOkDH3
EWjHWH9PkNfexXlnOUugfcACoKK/k6out/EhXZ68FFpMV3w5idpHU5GLuqGPfPr0
C4gklnj0wrah1vnA67QgrWawdibWFVud8TBd3esw99LUNlAlm/s01AvehBDm6wuf
8MHyqlhY8DQ6PdTuTGpEAescv/tnYSG7aGbCr1mU5/89ZfY5viGGHCRyk2n2hClm
XZb7d2PwQoz4yRRU0TLfDx979Sfa23aSauEoRqmaZDfxWpFbtT2B5/+Zt6kOzx2c
gBtOKGiGuWtl526tQyfSLJy1Z0+Gq5ETFxG8V4MprBY3HVAcnG5rxMcBVXb3HxJY
3vT0SuHDv9TztwiB4jQUXKpfcdj76oGPa1NIxJMbGjb2ErjH21Ic5fO8UzZK17yA
YLFht2rYPu2ykkK/7/KLHEb/FAwQ6EqQJeHH0G24T23WaD2UoDuoDtdBt5ADMUAg
1SBZ83DNRE7Et83Y+V9HH6wTBguY+IGHlBkozXiz/vww2qNTcmWw6QJlel9kUG3d
LMKPJblDRz8rG0udGpn34JaJF3r0Okh/35J9dkbnnCZ0u8nWMVCTtFaZXi+IHTAt
10N2mH5M0j3dJF0yxLt8sNGsCVVZ3XcISthciU4PjmOeDhaZ2msVDRxomCx8uUG0
Mum9LRyxZ4Pfn7QbbeUkn30R0PCQvV62yu7UQIQx1+dYImckiQlJpdCMER2h4aFp
DD35kV5Yp53BASOHIO9ASkWaMLVHn5DKvcTUPPzb5GOJtuf+VnTNxtPwtOMZtklf
IUtsRVZrbHfz2GfxMzNgTwIQvnCZfnD2DcHYJqeXnydgoNO5TiwkdFfpOeHeIZXJ
umkhIcxFLZBZdL7njJ9GNcu3zG+/F2VTDDNd/N+WJcINaJ3vHZKwFQTr/n2WVTTb
DC1WGYjvdaiYC7RjOyykSz0dqob2N1sU8ff2dzKi631Mwo+UXCNE/TbMeUPk2qLu
iFUJrg4knX+xNPaSIuGJvajCCxRoSabjHA4/sW0od7udj6TJOLZkm+GHAYWe7B3A
GXcyCKFi6YZcgcJuEjPbULezxQfA8GKv2idRqRPZrJwGPJiVKVD6Zf5tFPR/X26T
rJuqxSAFBHeXCxJbbBKMeg8ZERy6rSZnfh3nW21s3h2xHG7Nmkxst2UrlipaY+MY
h8hgN22ZXrPHiSPu3tAzrUdCfLW36Jnr92aoVlcwOeh2oFkGK4VTuTXBfHq8qgZo
l937lTvTVhhv0ky9Qv1bvhage0rR9i6ypSmNbvkVwD00AElOR6+D3dflKXuDTBMp
ZMKaWzWshU+qlfwLQ9zifgEHMyV6aoD/8PUfWhPDz+3j4XyghfwFx1h/myEN5Ilp
eieZ+FdnZ2FArUSlsGC5VNJ/V7cqZX1LuH4xjlUxb6udkdajBCw6YmFHyWMKhJvw
SFIn/4JJUuJTZVYLUMENSwx8NwTJb3YHUSUtN75XUY2qtflFIj3t505e9ed6Ni0r
imvZ3r6VvFWAySZTD3bSnRpd/L6FdwbCylhIWyEYGyEUVWGccQ/LDw378dTLWLcN
`protect END_PROTECTED
