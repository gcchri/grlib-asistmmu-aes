`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xq2kiiEghORof+BBC68WJPXeEW85XyVEHCoV0ZE2QCDUpF8o0Zfiz9Rm7JcGUhFN
rvXKVnnQkEoskT4rHVC8MeCBwG2IcVdLyqNPR6DeEB4unFB9ZrHRcoEHj57dxFEp
kybRzbTDiGaftACgeySP37GzhkgN5XJ2TpCdqNx3wVwWJGGTVxt39gp5CvHB8nHl
NUVwchr1mZ8a3DkECWWvLGwTmDcD7cEUr7/GT1HYGP6l86kLVcmPBijAtb1oDspt
knWO2jEQySZauwazRDYeo7LANTxBlV2ebw+JkvLeK0qtqY7VCXGynpz+pmMZWtKc
w4I4udw///nqXodP8M1ipsFMqZZ88Voaz/OJS0k9loU9/s56noBnvZeAeGvTjTo3
bqZgIHibjzyO3ZR/rRlsO3cbjyFoxZ6cjvR8/j9GPBRKZoBZ1JjlsaVRJOSg0CJh
wNa4cZPCXTvL6bEZdP5ybu4NNoLgo9kMUPn+U6+Ue0DFVjn4OiGT9FqQo7+1K8zV
`protect END_PROTECTED
