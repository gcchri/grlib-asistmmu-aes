`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tL2chg1qYhQUwCPPkpcrT8iAlhngbCqXJ+1PuPPxtHMbGRIOyF7/pbWy3S2mUjr+
tec7sLKtUP/yYFJ4LIzo8PPmn7cNseOIgOrnOFa+cM9EpV8gZXQY3VFxxyrgj5bU
vDCfH89yCPAJtxZMw3aG+wrZ2+f8BC/fRlZcUOJFqjDeVdQ/ANAcZ0u7dtePKXf4
1AERsrzgs4aEW8NBt+VYTcmohX+2abUHKigDMuAaBLJz3oBqX1LvS9uYU8asvDit
BpVH9TWdxhUZWBknFWeZiHL5ZE4N0VzJlNh+JzbIt6NAqgGQi/INXCgkbZL/LivV
4OnMLxxpr1auGiyZz+qgMRuJTRVo5DgoeUCpbwrY3Y1Rjbn9+W5m72mv/zGGZavQ
Y0uSW0PbpQSCrucD2UlBCWT6+vob4A83oJsnx5PV5Qu6AIPBYhyya+HBl9Hz/FyW
fAvS4xtGNvQlI8k8UQGuxtsPXiiFnbky0W03wLNPOXGWAHC4TqVLCRlTDuKQ5iFc
sTBe7jydTYz/qoq05djNw+kQfjVLUsKWABSxEWvHNV6rguXArzWDcchBVB5AQ2RX
oFGUJahbzTpm88XuGLJcR1M4vJCfsqaOpGjI7UbX9vuRu9kd1BehTP4xKMqTukGC
TtYC05CPpvnWs5fB1RAjT9euX8Gke27SPOsak7FPN3zbPJFPs29bv7r0hmABN+PI
95+5I7RGJutRsJ48I5yT1RTdmPGfING77At8cvrs1HJnUeWh/9+mE0ibIPqajmsk
E8qAc6uJ35Jfq2abMp6zhvpr6PAkNtjAEmxv0VRdqHUdq0dqdeyHVGc56IPKCPHu
GBpXddGE56LXynwQKvgP0vDSfqzcfSDAKZrGUj8HcHjGQ9j84lKCmCYUIRroIqQ5
+mjqyykIRdx6EO62fPbml7fhqbTiAAElFZcuetReKZ07Uhd7pG3t8G8fKK/RaMta
`protect END_PROTECTED
