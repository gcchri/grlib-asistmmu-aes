`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0jWc2xfeOB1LTZqyYVrcSXyGADB8nK4Dd0+mAwaV95sONYLsUd8ITjFS2hiIWE6l
7VwQkEdneqYqCl5gRICAF90S69sxzNjsqAe0q+5mhhfQU+feC0tHXXosqx25r7Yg
EWdpik5ogO6VBBd+BooegJRJmXUxIHPSYqY22WHKblKS+GOmUmELU1n+QAYid1sZ
l/mlYKp+eO+B0c4+Z+K8bRGFKKVDbAvYpKo/XcDyj7KZD9IkVa3sOuOnM5PqTx5l
YBi2cZBMKCEFwQ9KK/aaz6bY1eCO0qtM8HNvv9A5geKbDpubcBIhqKXAR+zPkCq7
r2wAuq2KbHTwr44NFghsW6Y6AmfgeSpDb/POHlai2trD6nLwcmz9zrm3DQeSVItO
MFD0lKrXuLi5I+IEKRmiJD1x4p7ZyA9N7VPPRwlS42c7GWPHDWPCu1hcngLsHnlv
OUE189J3KWzy/LGaYGrRQOSzr2YDXXBWnGvV+9mpi2U8+FULGE+BX710jX41IRD+
mSJf9FCcnyOpVOtBJETmGuwDpo/EnwCRg7p7Pqm54ufbEA/VglEwjj0gyW73aMUB
5wjLKt6OH1qiEO4DhAX2wLt3FWEOa8qmkKO1/M1nMEqczOLydV5t59n0lhrotsTZ
lR0ud60zJGVXs2Pj/8BKomywDl7If7YhsvE2MFThjPbGVzUa3RsQPBlqqN+v8HhG
6aZKo70K6VPIEI8Qr3MtORPBrTlZUUDOIRWaEWdOBnwsWbK9iVViPfbMRvFX+qA5
`protect END_PROTECTED
