`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
58igmE0AnnOCqkfiiNXYa/R962iVSaAns9CID0kN7yzvWUPxpAsqJAJiemTBUVD3
IxZQ6oDwTGWjPppdfTHNC/jPVTLAbY/e3iUmdx5JyQrt1JL3kb8hhgY71kk/IeUn
B9jZXHTrsI7x6WiZ6CgvGR+nwZWv2k1xkZef5z1jrafjUHVj9K8reCawpVLJ/nkL
KQsUjpzyEklKzOkoXC5lc89CSNTRzVS/ukljQFJv5gW0dTgasMnt9jnvrD5D0POT
/CkmN3l+CIjknZ7z2Bg6z+sWugs9k/GuiW5N4+J4SK7wOWC/pRnQt0pp+awytZLz
72UCLy716rlMwGjGvzi08BHL9jR9567iurCf/rYh3Illr/z5MViAdZmK+5KjP9DW
h6BHZ0jYenSUCW/zhKTRpVL75/35JBfD3yF7gvjucLZCOlBJt91HYZMmJUKya/so
ogArc3pA8sbEwN7zBwCfhpgWIl59F3+wToKcxWM61bHMy5OW4Qz+eXI5tbJ27HnI
aUm38bsI3V0Q4nQ/PtDd8VXHeX7xQpHCC1AOzo0v37fo01GCBC0gyo6WhD7wPU/g
HP/Tm7MyiBRGxhxYJA+l1lhTh8MbxG3Bs47PoP85gMXU98W5B38O1/Dc/9kc9Hgu
d8LVVHAXNjEv5TgzqlN2gQ==
`protect END_PROTECTED
