`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zjEbVtAoKSwsbxMAM8Wp3tORsICrpZBNrmbsgz0OVI/JTNFVKgcH2lCdbCI+Pnpj
t6d2H5v34izW4RU9c4xnWcd52eiBRx2NCrKRvwPO+hm/gqk3mKMYr7B5M2o/DCoJ
W19vw7yJDdeyvY+BxYA0b3uh8UMedsX8Mvf/zlyXo3p1LIbpJffGnSCRwASRjoCZ
CX9L0dNBK8+iX89nAliBXRZEFzk+yipgyrNL3pynteQMVzRpKx1JzM9Su/k2+O1h
KX043RO4IwvmRHJBG3qUvlyQ3k4pb3kpnovEE03pQyYymKwm+OseFEUfEF3iDdtp
m+6ADxLjW6xJeFhWBvXJDgAVxF4Ne3X+3oOWZef61cFHggPe41mooHb5luUTGTIH
K+TDh58Yv+FOjrdPLFmUJMXNhwrjvhyzLxklreBX17gxbSVRySACYae56ocOmlKc
iOtF0izDBu+84xjomEwKc7RuYQSw++iHUVh4W5XEL+QB0IFbbVbP1/LYRrTaUGSz
S0JhenUkBlMH5cTUO265q/YpBJ06j0WRMBFPzJ43dT4fibr5ogvhavguH+OXHYd6
bvHXde4uX791n4lS6q4MmPWMKDfVR3CPKHGSIctul8sJv9b5Gker8xxWGr0A6f9r
+pUQg9O9KBuuQjlSCuocCh76pGl9m7k9zG5zjGaW8jIVgsZVW/gv3wG1DwM2YekG
/1G9s7TCxPJJmjkMkdzMXKQ98jpGchjmyOjk3Y+SjuO1Z9o0nqSUJboKmbZyOxus
BOvMZjkAaInkuDTXB1K6HKcpJHgCivcAOpNDoanrQLRjMtSEYrhZQde66jH0E8es
mz/N9C0AYwCe6LWzXJG5U4yKiyzuRzn8dAvz/JMROuYrhzoIZRFTlX42kV1M48eL
fuv6FZR3fUJb6Uo5PMBwk6+aiQ7n4lIaNGdyEL8lzPK6Io+2mcrp6SoPvPKkSQjr
Zs+8fCIaxqyLnx7YbY0mqT2LngRXMHCMaDMEqddgltVrP5bBGNPQENATCMQ4/S10
XOGwOt7wTq+yiFw8SD+APehShtoyl9hDzTJ3jSa4CiD/BroV2lOsh5W8+zW9f+dz
EN66SzetIhZLE3zhBB7O308uu5Z7Gd815EIsMdoXZvfrWsiyi9exogN+iJVgt+7n
DLBA+vQbDlXnBHfEir0gCWZVQ0Ke3QmAI7OqDVLfnIQmA2Wk6WATdDLflnQsEGnx
g9HBtOtiVkXag7psQTT95xtT9+p46+lv3EJCvc2dJcCANraFJSIJMD3lSAR1xhwl
WVjpWjkcQwiUn4TYKIbPI42hOwyMh76XkMrmXJgyA7xCSmRuisnlQBRUZjhz5r1S
ys+cTFaPaMntjO1ss7L1DcsPkwWbDxXDkLHNoKaUvOXhT+zkDBx1Oz4b0JZVJ0si
PjIFDRnJYYQ+2NajWYT+WcCSMqTpX/ht69I881TyF1mcxmYlithrdA/6+kY02spP
sWX3SgWL5yuKVHaGVmL3ICBgRfIirZTvXYcEP1g9yb1ImfMihaRAuQXaFQCEoXE3
Px+OIlHp6foCR+5ptZMYEEZEJYHvrnSqg/r5MXBqOIYnRRLE6XqeTBz1JIURI+HE
Bh9fEcAQFh32ealBMOvAUCHEdBjcp9+B/Sb6upIpdEz3CsNF7nfxwxbfWTJS2jf4
6nHz8vv3DGCkno0sUz+tHqw6jY+xkVUw7ALoO6sL1SMBX84Xj/SvfmQ9Mpu8TlZT
P3ERI15AuDqqctQibM42BBtdRo/TfBfKtKowKpSl5O8hlTxUb8nfx+FqVPtbuwan
lL7hI62e8NuZPm4BG9LZef3+UIcrVp2eZyu7kE1+T+EwLV13u8m9QdbhVMMWWCKi
m9c1arYLbo2PSgDSlWoyd4SN1iqyfFyxnaPJYIzmN4H2/UApNOGj1kFXtwnYowFF
ADzLVaI29iaC8pDlGsCw/gcSztt0FgG3DE04AI1mQ9Yu7Cm4QwxQhU3iLvMucM0t
P08FsOAij6EUlASJAtrtodBxEt0jzECzFAna9t0GOa6qJ6nZg89HW7ZZisQfJR1u
gPZlA5GbjOKlOQAC2YRHIzOGZY9d1YbhFBVAI+ovSyOxjUZDDp29CsKlOQVdf5er
zncMZdDIkzyhyi3b9FcZJS91XaarXohcMYw0vdB16hrUzptos1PZvTvHM59i7X6e
MDkQjNmiS4KRuPIZoWre6jchamJbgo8/BcHexxo7pGHSuWYhH9adshqfdoAoNYu7
JugiVU2ZElIPXsf04MVKZF7IAs2u0zCz5OykIVVwqVbLhDBLcbz7zgTcQkHbrMN5
7QaA6QqJ9OcAv5rpnZ69Z8F/ufJfEb3FWpBfXpxpzS0EE+SYrq2V/EvTRvfTRcbA
T0NzESLF/x0NpRSUTFP2VmM4lUeS/dDw6qBIXp42c8BNnhzxMr2Spe0k/Z17iFgH
kyz0zOYpBFilzBgbsm5VaCOC1UxOoML9qompUuTc3HOlIHsFG6/GneZJnhfztO35
8biJgA7JpLz4gX5H5PsqVQwlJCsyTHQ0vIY5FYei5I7iHnwTdRGIDGJUg84WBLql
vC4BXIXsPteBk0xn1QjDtzipSXss8gNKDAG0FOjDDFAIh6RWQGfgACMKLqsr334E
PsMzo1ZUJdXABWJ6QUO4UAiJ/GWSJgrLjMlGQXPcvqH2hVeHK3VfiW4OXCg3Jt1j
qzvJjoZFg6N/Gqf3dOAIF1MhIMwXygA/rAOBIwsZp+3mmIYndVhI1tZXlewXkUDu
iYXOC0KiEnaPMh0b/5+GziHAqy2SIpmsXs8uNw92f0s5UlcJC8+AswGS2Ykf8Ft/
5QVR70VfF5rM8aBOSYu5/dG0+WvL6Vm5J2De7u8oHG2OrZpqOktIULwwK9AUc04r
om61Pq7hKAM83/jkkTKFvFyvZFTgV+5f5cT4WeZyPraYcrCFko9knLJlBHHq3fH0
KbYsgkdL0igQFOp+t+Wmf4gdCD2YNHCdNbcyG1DjEb0hvCwBT3zVVzuy2CHrfZQi
9q3rHK+LyojH34CDWfFK/A+Iuls+weS59C1987H/GsZwdVyaTWlxIBIIiAQtPgLF
eP8oUJF7WWVdOuutMN9AGkRzZQAGwdzrFXiW7/FebbNoE57w7WoJf91K7pXGA3tt
HRJDEA61CCgoZR+ZhOj+MdjzU4shMeM/uNuTvTXnRwXpyIcEOMW/8yC75jRhGC0b
EqX7B3ZvnvaxpJjJlEWXBlL27TS+sH9ihu0AJYJ2F2WTKtumr53RmyNYeWa3F64q
u9Qgp8DOifnEEN+TY8PxrDuvLvCZx1zmy0dWpaGnl9FiwVGPyGEcbXQX59Wjtiw+
R10gEdBmPvv9Nz8ufUm9T23QU/TeUsdTefswpzS8vCOx+F22uYXg5koE4zmEaNFZ
axZpKZwPd0zWTCDyDFXvHFxQfWv8IwSs6OxiZb/mdR65deMyXp1ZrkikyWaFZ7kz
9cl+wC+vAO3JLZ/qhA3ksgfJy+3gGnk8C+nolmyTuARWGBngl79fuGBD8ytUY5m8
Zx3gexBl5VaivQiygFUthHM7OgEOgnDWTHeEWV0cQCfWkPovfinuSM4uxJxHy/eL
ja0RHv7Q63nkFOCdwOMJjnSQzm4WUR5G32a7zMTEwhbGNBmSP+kcLL+ds5l5Ak4P
BgmS5PCdvOaR0vgYaQL3GmY1XXEAy/9aclsQokRRSpsu1z/zZhg/yCUASlZbXWkT
cXflsd6KGF0nh4cVbbKEcATvRjBMouxRrILWiQe5DFVarcuvVSXuiXdCmEDRqgoo
+OjTctAb0li+eDoMUPjuIeRRcUKv/r25icXzkEpx36ZH3jxGVQV9oqIlUSRSIWfJ
lSP/imnTUFMxxxAsnWniZ6rurpelEfiUc4YEG8Upw1cOCXAbrh3YDJHOHObXJ2WK
Gy8GF7pNP3Az3LKKhUsS7zwoe88ItNB7NVBM3d5sVrU2mvu9HsyYZvY1MGdtaNm1
byy+YH6UQA7FQRhs+7XSjHiBnq/F4znDVaWv26p2vWBT69aY2QIao2Bkbd7rpoYA
nfoO7krSLEQzvFGgn7h8urLGvTt4j/PZ1GmYIsRJXqsoFh44Evph5IA4BDUOySnH
CwsooKDba6cIi+/Pdajt6hvz6F9/NPFgrXeXfpxsXqodlzXCZZ+5zkFqUdJYLTw6
z9s3qCn0lph1UzNbrG1V12J4g7Ve8ws3uRCiBsy/Dy0c/KcmiczL88nTW4Bn+65I
H22/Bi5kE6WbP9I0kyeUSnX2P3l+HxJ2MB5pNJkB6Rx+XToTUwMahtu3S+Ge7kn1
rzMxDyLHhjk3LMPqdbLxKpBeQ8rmnI24t0F7xyTHfN5nmacuvJmYvXmUMHFrNHvv
Js/2uznDdvoMZ0Eh3+dFgHWR8uPwZ60dyLNAeU5UZieG8bfVqBHSJNfSpDtukn/1
ZGb9sRRe89rO8M0LkLy2IXayMsavK7vbdxdQRchbe9+bs/fv0DpKVSWuRuUXn3QN
3jZ1LiuN17P9reo0Uixu3RRKx9dOAEQ2lPi6XhuqwK9LjXA+GNAW3W5l/s3JqLDM
Er+g5MnmYVMwFl7FEg21QTf9e2H7YIe732D3Dip5AHxJMZt4XUWlJMBJ7VsjOzDU
cuLU3Gs62rHE6bIGcsp7bC3pPDHY2le99CoaYHC6mtjcUgw/By1DmKRWjg8cc9XK
1oe5n9iGEvbnjhmVJOS+hzQxTIe3LH9FqRf8PV8r3o9j/Ih/3qOePPIdjrgUByip
zw/VaulBLweSRBmpsRlAEeZGcyjqgsy+MxGuCvXO7Dpw7X2YkQ3j9k0YaaJCp61S
GUIkPitHzyWnY4ZTnTCOeeM16jhAyaS+xzGDbiq6nUz2n/POYE5PbToDdeUhnjJt
AVauaITQa3ICf/qsddUgw5YVPM/wAoZyazst1v1d4qoRuLFx3YULUaIPETw978sl
JTx86zytCSTyKrMw1jjgqOqbbMKrotozHOf7RT/Mn+naeB9tPwaqjZiUHOKLdfBo
WdGLoDESCQOC2S4ST8Cw/A2PqOmiMqEDN7A0ZUfB4MnwwvdDH4uB/5liUDv7LmO6
a7rm/L2nM9p6sMga/RlOpXwbn7u30tTHfJ/3ZC9jJ4zP9b1MF550eWT4apmmOP/f
Ou+R/7Me8F3pWEqaCAIkjlLSfu78ZKn9ek4JvYVJExu3/9p5AySDL5r85QfEmxus
QiwJTbiqY/UzkfwFmYInRl39mMt8YMXVI+w3pDMm7hHk+m14wdm55SL5j8rtS5FQ
Y/4cCr7tr4stAemur3BWPANtu1tvm5JX0VSIZ3NfyTvETUSuY59/7K7CF0ZB3S/f
/Fyot83f3dbx9fASwE7QID8ptfI5nma8551z27pk3fXRVsU7Qcrwke9xLPaL81Mv
/A6HxxRY/yc+oDz+KYuCjx+TUG3Km22Ut+wTQ8C4+ovcfK/m2p4bIM/Rbb+7lyad
B5DO68tVDKnxPsop5X1kxSwFiEfdMk+J2E6zIhCYgzbcN/9i/G2ObyrN5xRoK711
2mTL/ipHMyZrAQsCFaL6kHquVMfykhVvD9Krj0a5heDT8c9KuTM9fPt5RrRT0BrB
X8CoGYzqUYcxlaH85d8vKuMDIx0IdpFfH0T4wioVgl77V+eIojUmRrw+STK65/9W
hg/fNllgl3aaErArZX/aEX2ruIvvmBwk60+G/PdgDGKkEhii7MwaSIRJ3ni8Rykj
f6idGMYjG5PpbTVYCsr3yr8ZDVpKY0p9WBgQDG51mpMYxecX1jz7mwxfVJtleRdc
OHuG4DmqOOCcPaAGPIr/BmjH4QTq2wXNPCF4BG0X8BOWV7nLT1UszVVHuAX0cSBU
SML08MtISZQkVwzMVF44L2lGGEmpbYPTWnAdlkRUoJq0JE/AQyF5nb37LWoFUiUB
5W9+byk5+XU3aHSN60hmCrV91cWnJ+WV44RtpqfHtJvu1Q1AMkEm0iDA/ciYMbZU
AtFeCOV5eNH8LCJBbYnp0nYYWdLzjeNeXCirlnYY5BMX+XRAVJZwcsI3NadVbK+P
TeAVvQx3Cmz32rgknlGez0yO6dsnz8Dpo0noMDVZsuHcPecDJ5HFuRiU46CatE0l
MBc58BuLx8SW6S4SCoCBvaX6Ay0ucjePMSLhHtYolMpYA/ToADlx0LWwa0Mm7byi
YPXmPv1d3LUzbJikGafVggX4OmVobFxy+gA2toAQC2gxI5nzPqCSnMwW2UeQ3Y1D
8Ko4XLCyHojMwLLjIAdHZVlioWJ0R3mzMeg7EkEfe1Yo3hvsOIiZixWOUbvRSmoT
O8rB+hH9b1HzAKTjW2ChyUrgtLI8VINm6a9Dt/lgB/y17F5Dmex2MKqXQT/x2z3y
RSUms54JXQoZlqB7i2MEXH38rCaur4AUKf0y/Ye8qlBqSkwH/ERTk2rydW+DXGOI
riDdXVC04GD23tnlkTVHV5x6Qox0mvuYoYSYiZD4O/jN8/BUQ39vdeoeM+avitU8
MIrI6oS0JQyHHs6NleXUJC0yzdnm+bzzVhVZxgNgpU+WaARNdp7lid9B1avCJ/G2
fcxvCD4zQnV59ewShzsLnMfp0uGcXPZRY204bZ4DHT6sSJpm7QNZQ73IjvQEp/BH
8LWXLqsEiwuepxDkmKaHm9CuiCQwyQ46iTLhQweRKSwZsTQkg+yoAj4HshLim3Kk
fsN3SgAk3zmLQCWnLnvYnq0JYfOXNM80rYy+bhmzJyoxes7qEG5Dr0AgCuI7r8Iy
EfiGS0dynn1NHlzw4jashoceXDi+Igvo2kWg+qvj4+Be1VskB1CmZ3Rxu2Kr3Ekv
tZro/0mwj/6TN+gjjcebzHHYFF04k20xHM2T+Rg4m2S7ulFwQAXIjmKBOkpUTeh9
dp3TI47BfJi4Y42PWUj7V+Ckn6sfv/og97pYquQ8PYyVWSk0xQsZsf5lU7J+yGRa
do5O9rPbrKTZvmiPu7yLBipsBxzp4XSZ8cMq5qipDypUXO5I9NeVcTj23xpTNgBN
s3pYIedQ4cz6bhennMqy9XYX0w1Cc+Agz570Wq9YiSyLpAsm9lMdhaoDRhVtWJ6J
e8ldoNz47lMoOBZl+lUHSHzCNshB5t1sV1SeC6MOixrsNUOSWArpW0ADOK/OLlzQ
vajrCH1+p3KcP1sKAXr5buwOluNFeMc/TG9dkuWTr34x+3CRByrBTcWeRY3t8Yed
+taTT0mj/Uer7JrIIlW1v629O61FLzPcmw5oau0b33O71FjTtAm3OPCGorjcofoe
+KgeoJdyqiBvO3WRqFRsGKQ3/4a1lAb5egbFjGOheydIW0VXgyc+3trqAR71NvV8
HLLlW3LX5L7xfelj7fQG8jzQfMsCsQeAQ6FSdetUHw5D2nAH2YMjZ79zKrFsRj2F
BlXI+bxPPAMKCD3AFhhGUAq36l+rnh5zDj/rHIstmUntaqjHTsjgRJiexGKp6Spr
2bEH31cvW4RytWjXI5BB/XY7yWyAcIdN1UDF4XyxxMoC7C5inkqU+KYMStCq1exi
S08pf3PmnJZWViLyyk96jbzL2iFtNWyeZSMcWEwa0+2/Dm7l+F1Mrd3g0CCPvjVg
TJdvSmXNqQoJdq0dxUDPbNA/k2JOglmDi5cp9yRZxVWIRmAvtg2zTN6+ui5r+QNa
Cbb68l+H84DMP9N1pDP8yFyd7KAnSBhGatQ3LbpEjbTM8x7xqoDjb12JvD5U3McM
x+1aunextauCuaH2JFwZhzukPkon9YYY4Z9OOqCt7a/D+3Kg0DVKDFcRYxzMIO71
9lDJGxTJ54BsePFhqvoXVv58IxbK/woVxhZEjMgujWIx3BoKmCVzHm9f7Pvp+djx
x3CHIuWaQ4LfXY0obl0XYC50Nku5/d2OuRxwYfj1zE3Ay1bZPfT65HDOA6ocEtQ7
/OCacvjDfVn+DXhO8afthc4vDn0pDNpdqXco+obQcvAqq8iMtozCN+QGZI7bwtIV
bQbtl2RbCbJfWIoidlDi37P3tZzM+qTo1TZXAn9oRWqk8lu6qs29o3ru96vrGlLO
Fa6EWpNCzbQiOSL6CFZVZVD+WS9ONiO/zhjuQplftCxIyCW1LGPz5PBh9y/M0vmV
kkfsWJ4lu7QTpONhLLabQnfv4A1noyuDk23txpoTVHRMh4fLMPxifLMCLHniBiG4
BrVs5coMh+CmKNKDy/JmUvlpk5+8gmztI05lophb/ZSV2AlY+GWAuF5thHp8x88U
h1fYSWJU7bA5Lcnyl2t8PAHRylbvu48AZKHlofmjcobnglWHl5CRFG6FIGoULn/M
yakl4sfKZf3ETOaw0l3RSVBqTM0+ToTuDJPy2EK1m9hSgmZCejIYjNagyDuA2e5w
3wRI3LRjC5/y9dF3ApeQFRHYQCXgRiF1aGnB5kI0aQVb3DWztybbY2+uzUdupmAO
60mZgbaZmDW4qGSmrxOA+kz1wdN1q84+d4c/jpNh96Rro7scIWDq4VZbcdSbNidr
S/GwPlydP5m17vwoyDKNgXH6qDlWgD8cmAoXgeqkTuoWkgyyEY1mKTRfkNhk8koW
mraXdG3N2daWj+Uxm4WM0RKfWM2QPLc3qnqpIH3SSn89vs7gPghFUED7bjt3yIUX
cDayCnqqoBtgVAedFcqVHwgwfJBBh9B9Jtl8c9dJrkMbyb/xTOIrN3RN/t3TE3Xn
jl6TxfEVCEMoeZFmxHfMN6/mAdLp8soO7tFQhrTJtDp0/XA50Huu+lOtruXWRUWc
EWIbxusWluBj9vR/kLP+bi/54tmcUsqBlZIHe8nXxAAeX7rg2T5AzUjgdwJ3U1lL
IzAIzRb4Z1vOFhCaMusszK81FHixSHy9Ad7ljgj1XU2djcBWAPPOwTwe21DcdRMb
1I9dBAaVCR8HKvPPfY3QqZF79cjcvQ0HDjr29cyRyBSI0dRExPXcoONtyp8YMkNo
fNcEeZtK7MkVTq+jRurIHDnfVA08HG1elMKWW/o0RTeN/jWudWisvUEmzDrImkrR
1cI5LCDxXhmNO2Qy0/mOKtqg9yImELKMMGIeJKWSM5gUUfgWa71oakj4Fse4t7Ec
3RICFBWG3rDNp9Pl32mKOe0mYSVxpDRqJlEUbE2F6DxdIsN4XTLGj1dacGbAsXBF
p/CDjON56H5FUSqBEhHOq7M0v1fpPJrF85AEizK0zVEAt2CueptAE7n50q5l34d3
dJ3mnaJrDdXPIKyHNcNDE5k65j4U24rHmJ3mmxDWpJWEwWrhC/UIvtWkAZRo0BU/
NPkUfUNIkPGWhixFXWUZvIXTHxAYVlaiIs1jR+sJ4yOqAP8rOvkqgOQB2pnbC1Ab
rkjTtK+VcBeFG1BFDYQdkDui1ldrEpGiaV4bm03/K74JXcBpvmeN9ZWBSiToqra2
UwVUC22LuLqGnKEOjCVQYHJCEIRyR4JPZzBrkWBwEPCaGcLKHQQ2lA/TAShs6GdF
5GlfihKzJPX3yTu0Qt3jI7MlHT2obX0zMYO2t9lfD9Us3InsPaIQNTJu6ElzB8Wi
2Q79oT5y3b+BtXoH6TXqQFccFlOMMsGfUM/SBIEC0DMdtycRN6VaQmsszpUZB2kX
DmLS7BgIFXU4weESxIFCNxQC0VqogcHlsQprAK5ps5MDd/Fs6UvKtT4nzMgvKyYE
L+qtTjeM6UlwRrmSczou4OkPI20gKcKRy/tLVn2kuRVLjaU57UEjXdB0zO0H4j11
arhBMbNx8I5X+B73Fuxg/pDhCQUNiNWgbNbZf9elKuoI6eRQnQLUkU+xhQPczNrI
APujWQKeBn4w1Oottb//7OGxDSjtgAXJnDOGoA/d3rT70BFKfjT8PD4umFPFbL6T
+0XHfEm9h9F/H7OLQL0ugiMhT8h6H1+E9ZlTQmCeEpdd7XEVY0f7DTaUYw85Ltrh
1wSWpqhwDnNbedaWgVQ09KzKc/BSBDwClNHwVUiYe7rp7wZ7xC0v9625jjglVya5
1XtQtkDVW9LZYgeeb6Fwy9nV/23J7M1HIPZeWBp1yBtuqUwLmwu0P1lZrCTJiSOx
HRbJGij+gdrla7CPOkmttdPsSg/VKs0NdZ4OjHPalfqkStFDocB0+MXAwmknQVIG
pL5KMEtXthIAX5lwaVAXH9j8shEiwD7hPvTTst6ocwmnzMA4pAtI3BHoPTOXQD8P
CzeKVq0OgcQH9gJZ8BHGBjrRcrz7ILYHJaIWReDIF7LT6Iwfn5LiOa6zit3g45LK
BFkohU4LDWOOmTVqWNRGL2TJPb+jkvAWcBUvU9wtFURq5BcqBXuz8k3qAvlunslS
O0FPZqp95FpceTQra10hcRcOtwX7Cp2xlDwFlsPVDzfB6b1EkX9Ga2yQOi5OZi4l
gxAD1RYaYGxMCsAaA4skpwKrRJhgOIk5dg/K7O7ZwTmtEJtMjRhLLnSXMwxC8pmQ
B/UPZJrbTTHmzqajvUihlrLkeBrHwGPYr7bPzcTJdDjeAEtMs7uHKODKyOsPdo/a
3OhWIWDyBppTUegmmC1g9pbqjZdjKNUGookzGZK7+GLHohz4k9lb0weh7+cfu7ei
zr9bTdypJrqernJZtHDjPzB/jt5VdI1fy/FoaOVlgW8SNs/J+zf1f6WSAWwhB2bD
+D1WnyhJNc5oTKLi1C+cFIdzKe2YoadvzuVhKUES9G5R4l3+hlGTMPMktBMDwsvX
y1v+W2EvJhxf168DNPmmtiEDAy9TZyD3hvgRhcTWQQ0AeXd+BvZb6QQGNMxTzbVk
pyFQWwri/nlLsM3d+siDXxaV/jxY2jrtsAau8XrCIXRZnZLoQmDRX5yajvEFzY7g
sCYA7lhejsUcuuypq8ugbd9i/uW+lTSQ40dSEEIHqzTCCR/U9J/9wUsqq3r9hh7R
n7lAdY3ywhZa+Dh/WA9p8qf7y/FV+WLPBUNh6mgNfOadtbIuh+TEUfw+Z28WJRh2
B6D6wyDrROoSpFRxWcDSVuYW80x/WNxXYNIC5IwiSZ02aW5/PyeZsz+E/STGmZx2
1CD1i4tXeyz4wfqC1erjz0YyhVL1DSIUuC5AnCWgk6VCvuz1+fsgvo7WujFDUezV
hVev/+kegkNZHnioXnbDXyYTzqoWn1bAKMINYWuDy9gvYU+fGp0FZ/wrY62H8GxI
B/BbJ+DMBJiJarHEQto+nG5MA/y76JrpN6uUzPfe8HJtN4PozNssbTg6R3vzGJcs
eh/tWpaw4nqg9wmDDFwBO7ai4ot5XPmLAsw9BqbglbiE7KVbIfHX1fBqYj2SDKIn
WYBJ34SEgGW4D9F+Sr2PAKhr/niv/F76M+rSKjo7PyZuCm3a1CDrp2au0Yqr9qRP
edUA/IyPcLE/cGGXg8vdazfUGnkAqLoJvq6z4KOnoyCs1y+VgGsIFBKxfKS6WZ1+
F6klw2k3mPI7HiDcK4Eu81yvRRaI0D5kGE8xVxUjkPm99vlyzePCyJFV+tEHo38K
qqLrKRJAjqmMXLuX2ndS7JAoys7hmYSu5c9e7amfJO8ErsGcvB90+ePlJvMwnFPV
Ral4I4DRiHilO13uYrZkES6aVTV7ykvnYoR5KNUcb2g8jVUZHF4iM3Of0ho+HTSV
NplhFaOudLNGTDbFhf1JXqjWteHUe2Ooo6brCOCtxwTml9zmQldyDBi+MYbn0N06
MFChPfp6s4Pa4EMOtudScqv3qKwCwfzRiCrFrcrfOoS0/lgjpj/cDU49Q4EB871n
uZyvm30L0FMAfWen3n1D1dTLRGjd5FiG1Q2GdnL2BkfeHPK/aCLTDkgvEZSNqtO+
7Mq5xiHn8eQrgDz59G/t8wp3s2dcSpouhNOaWpsGdsaPxkpOLN/N7d2suA39+uP+
bu6zmRiRpfe0ygFKGmgvUxyvCwhFyyAOUM0eMEqMyWKwVY45bg5sks77od+Xy+VZ
bfjae8QHSneN/+x6yNbfZfDRAdIDbQ+2xCUT0TBMwgnX7AQMVyIQkKu9gC/eJlsw
D5fukZC+NU0lCuqMH6VNHtoGp73+Q4H0A7Gbqe+x16fmO8oaG467VGBqtDpB9XHe
D16ldgkRqMJVSntCg7QKZoUTA/S2nlKY4VE7n/4QmWl65gpGYeeXInqzYCljvDBZ
Om5JcPQDBcgFGT6cAVrX/X+juvqHAT8IXfau5IStK7OWvIunBhljCbTypNjdFexr
+tVd66GxtxPibIXhe6xtx/KsrKPGzsqvR9YkBn6J4c4z29SFm12MuAGDsa7ILAKx
cYww2CDdKq96Tl2wJoRikD0SGGmM6TlQXHDyyzqUl0NIJYILKKHhTwLqRb/bW3xS
QrR++eUzYbamzWnvCWqtD4I4lIzCU9+yHCmaaWZpAWUTdYb3Z6MvWhRku+F659R7
sIbxEDobyTZmin0uLrnC9xbKKBnb+BbdOQMOc8TScD2SxmBg9Bl3VwIagtXew2oC
t/G86fbPoIBxFtE/ALZDOUXxVN5yUhWMZrjL+5LtYB/s/e9bz1ABddWXZxRy/u73
xfUS5BdqqI/lHIKnfHHD7VSvB9bDGdCHgQ2WUNPD2Il9rWckIA6wUo4o2pLBjtDz
8L2xzU73oqhXjguAIJLLGt+rXFVf6E4jgXBtLFiQ/C7LBACdR5aghR3AG0eEhzBf
qq4KeDQJv1A1iQBlZkft1pT6oxMu/KUVNFK43OxIgiFRlw0IcsmxlyjpNF5tyi5u
jYzMdYkmXNHZYfHVZKjZpXFT2LKnMe7dzWvfCHG4RtwnCzL3gTMJq9Pk31uSAex/
McMdLHA+dNsfpSb6eHWQ74pjILqO0O0HR2OEWJ1LMmyHhoDLIQm+ZqJKoenU7Yws
8qHLs/FsALMUrMgzTUZx/2LiOJHIrGIdZdxEuly/QwA+K+w+zypgBjhHL3QOSdIn
ZnQIFwp6R4ADk411UZ+tFdZB3ssY11Gm6qa1BkacmIl+cIqb4n/7ohQ/MVmnmHSc
jszwY2K/EZG0osNV1BHn6wvcfjnG7fayPZQidtNWXPIofkZCO6JKqHJeF0Rb4IVr
HTErISWLC/fdGsK3tw0cjqMEwFE1JgWv3L1Zo/UdAxyoGoaQOaR88pUi4MUTRMT6
mcTLjZ1vs984q10TuIq2nkOHG4T8kE7UkH4piuCrQsMzWvoUPaBfjsyOwLftylLj
byTskjPROC5vXiiInpTB8tu1S39XIDUSBcUftp+GXbYQM2DELGXqbrwMKMiT9pT6
gFVNgpLgf0fQoSHJhF3G46syZid71AQlOMJSZ37ckDBjDNJL0U1AhrvVaTx8/n5S
N+jpanQKcmBsAfVTuG31zr3h9oz0GbV9bRzDx1pGyt/EH/r2gddSV5106fpra/gG
JGpdSyZ+fY1gEmt0NNxbrHDLOENaSshhxJzg+81kLa30yeQWXe5+z8kpHfQaZbR5
uQocp+FTulF7Mn7kj9SlPn5kDbjbjJFfnjbZtEDAyZo/ZihFb/49qyxzcE2cJfsl
HOSJxY6gOYaG5120LV8HxAIb3+GPa8oKXu6haMK777FK7/EnDPleJX+RNvDyIi4g
11peVQrwlygnOniRp+EbuJuDXCEtYbBb7ESN0KP06td+A1j5l/uceqlPrgP2/IZT
gsyr4Y2ZJBwD958DbMMCJOC9kU/7tUb1pkOI9BjZHucHcZBMOwP9351YaUJOBNIc
qYtn/ScOdvDnB2qHSAGQqQbsm3t574ejws1Cqnwk18BVtn/oW0dzH4d9X7QRYtQl
tpTmb+0PDVIhh4QnoEI00HcVieQT1XnaIEhBhNFU6UqGtdDQMLb8ewjxjlI87VY3
efdKk6wU5tX97PSTviMUb4hBFBzxt8xnEl2bMmea1QvrJpJZWDJx+w643XnjIV30
WJ7bLUe9joh2561tQUpSAe5RpQGkleEIny2LhKWV7YLFzrqKH2+6pnqHkCTRRkcW
MROGxddC0AzaXDzXloyLTG7KwLKCESod9vwYeHnoHQ60ItRqTZ8os/1sdrH+VKkD
tY2yxOV9yjhJam86ipaoAyx2ut4QPupgUcvcV9VziwetS6VasD4rrCZSXe/Cjs94
uvKuCiyhbjnYRIW9I1Ze8l55PaOgo1dT5lFabWNL7dfFI5p+68qUoLzK67MD+tPZ
avqvXExTzsoHiAhqLCwdh4vXgfIDQ1Fjn5NbrMLdl3N6WeJij13IEK4E9skZxL6K
q1SxsYZ9GE/I1CXQcfRjCIuXXGdfIjbkYWRXYuhLTv7+/WChdLSU5knjyYtu4VTm
gQ9sl2JXuyXctBXeVuMcBQXKMd1mKs82cM0jLuBT3Qt0DXPiL9r05AWoJhzG/0bq
lJoLABrp1YcHxM7YrryYNU15eTlPl4b7+x9K5Da/pmOt2pZalA0Xaf55wMm6BRQc
kM5iJugNcTtCem5vseHonwnpY/D4VAJv56LKd69Z2CnC2mowrEp2ltss81hK9mI6
L+gPVDb75W5RqDFb8HstPRJNj4DEfyN1em+0PB3Y0B+SF3E25HrE83sWAfU5k6c7
nY+pCFPl3NXNHeZNmmOTS0gOlqAWPccj60VZ38aniQkqlQrTR4fMHgLIFy5zaQa+
piMb9NmgaBfY30rQIZ7NgLboJycpucaSzhufwY/EA+1aCllGqLUvI2MiYlYlwGrf
y+cv8357w+AhHDzDpnV+tr/PCtJH9rMiv+rDXAAfjqoUQs7mr7LWMD4SADw882qj
n2AP8AMdeaAH92X3L2wGsVwERXrSKg2hosQLnkXi8X+XGmbLXj7Ir8ifkxBgASfd
RBiR/DiXNQNYlkcS+jRRylRWoNvDh5i6YojCptqoxGkA3Daje2dcN6bpcfurbStF
ac4iIZNw4XoWvKctQbjC63OvDkD4h53aeDLlj0Gema01YhRWHUMFYK48XvvqsPKN
yNvwpwdQ3TL2twzFGKt91OmdZ9uKFEgX1faD7uO+7lo7MR7VRGtnJd1Fe1EmkURa
P4gMtavi6QIaUF/K5pSbSPnjWgLlxSRTrmoJDGqjhSPC7lLZFwT5Jgpv8aeyRaK7
ldXptVh/THd04xivpDV4FMXd5UwXnEZLCei2KQH/H2QujSLZY2FiEOUwME22G3+C
ddAwWpfg4Bncw9jkrD6oHRwKCWvOK1CudOI+1I9kYqvLs5gwtEAwbDSPko2tT5yP
Uy9KFCSw2gm7yGY8SeLSaMCNAj+ubyiqUHnqCH1umEU0faU29tvavuSSaDk6oaWf
JdWtWeOeHokH/Mc2gUmo/jkWaCWiybF+G0Fc6QQapXVNvyN/TQbmaeQLRU1WNhvS
Pmt+7iHR65e4sqZuxqAhU024z/9FN8AS5NNdZ5oWQ2JLcbpCkCwVBAe9iGDNA92E
4guuL+/Rc2xXvbsBqMTaKqeJm7IpUI9gzEPKNmprWDlk383UMBDA31zUNbFEfpbz
UgNxzM78doZznCz7czY86Sz4YlShIyWGmtV0ocdBR/8keWV2t46B+GeTUVH54K7U
MjrSbqMDXxnoTyoB8CippWV+Sm+CdBNIKyMID8Oe+59rOKAQacrda/Vk1pE5vW3H
p6bE0d0zc6raW7HV68OyhyuJL0PMK2bZ+xoM3fKh000WCmjZK4UbWPN26TWMIrFj
pHLQfkn37NM84H/jJ2lYhEmNgr9ZGaIhjfRE8StknrSqnbGhJx+TlQ0aDeJ1qkmt
7bS3tOFkK3phqPJMV/GpvSLLWw5dF9xigaQU1sV2oJYCOu+bF3zpjhdiisK/vKEP
Hhgv1rLXFjy1xjY2cFYy42aRHv5KeDa/WC9g1NTilDc0aYOO3gYdDu6bDnXZ1SIq
ntaveDTkfbBTfob1e10bnCF36p51Pl6FOIUyEhU7R0OETR2ZVPqY1k4wrQO9XqJ0
HmxVbI/HxQQylTvZupPs/B4T3EK9J5qHwNrtvf6oh7QtZFlizqLpjn/9/rb5PS8i
VaBWjLdpRS9pEgwQUDTleE70HYHW2cIPveRVaMWcaM9XKHVQrUTLzc50C9uIlti0
PRu5yj8w1zR8QyuhKwvTyRlyPSvS8+EuOM/H4ry0N/eYW6rxDs9v3nGIZn1lf0/s
EjyHmQhpXPSGiK+y6togBBAusetguotcrUKFOkbJ8fJ5BAd0uCx3+0DKsRJ9Mqvt
93wvfvmNgaDOyfQYeLgZ5ljqpSig5O2Wnc07DLGvML7JbwqRw+KeDF6zDRSO93rR
5+KaGctCYPmMPPx59o3rVB+Oo9c8u4Yg/pennugAt9ovLvRBwQPI6TFu7EeLzZtg
lCigiRcIkQXeG4YQyIKT9ROtgIAt/Z/m+OGm66W0iebHL8Qopw8+tl51h0Si+Rw1
kRBixLxLHNFci+28nc33JTo1M7mQhZgtuAwV1JfrB7MrWbI2lpKFQzbQe+kjW5u9
zLA4vEYw6uP55Hdt7w6aIgVrMWYC0eXuKQvCZTfOENLAnsCoi1SOO9ugUaaBUOHg
/AjWRTIpi6niRrN08ORi9w7fI8v0VpuMwCJ436FJ+b1A/Bs64mbOSVp8QcCJrIKO
Noc8o59KpsMQ/k8fO+wsuOuGsNOu5VOtg+Pk9MRxDZ52xXS6QcXHrZlpp/1CXNNy
ebjwdJOHzlm7guJJCkKPzjWJjAt6RDimvlqZf/ZMmV4pYZ0k5hkMnvowjAUE2d9M
wD4P8Oldj2oELP0m5e1ZruTYpuTsXl7/wz+2Yio6fRbX8K+D0UspVKK4+2S6EANQ
ZnTpI26QXaxgT3nz/UjFTc7axKsrGq5CPyPyy5jctZjkxZ35GLPPKYDEbwWvn4JW
0T0X2D0pVEpqUukz0v1gWg==
`protect END_PROTECTED
