`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+4tRry9HLZziJT7vv+QAJK+8uvVe0w7oJI85pIulxbaxw+Tj0oQj10iy6KoHNnyb
U/Fbh8u6WgaIsbp2q4+CzCW7mkCMcNHjdVTRN2zj9YstFb8IxY/AEHxELqrW3Vp3
YhARvWAiAO19gfWNxek6e1wUWhCRvDIoF6bQYosE5S5WwD8OXmYgs6L/b8jMEzmW
Wz/sjM7xz7WlhhXM37otLIMaVwXbj+p1OoNIU+VKI1lGF4+t7SPRgjsBvXwagMy0
cqlGjOljbKhckU2KnYVaombcyU4oHOa79lcEezsRHjr3XbpvsAsOcDJ2qFvNiSDl
dnquG0dL8u8tWkWtu964p44jbKZvyS2pQUA0dGqGx/g2s2K97JFE7tRLDqHnOJop
`protect END_PROTECTED
