`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2e0PAnZDDmcIjRNxCSWWds3lE5syxsv5Ur+pQjhrQSFGfFkGPbMnZVQHH5NjZ6t+
uVUSslA2QBOaX0/UO7N+tHvuewuKiOBPHp2xLQi5okeK4X3LCG2rUOZRhII8Yf//
UtN3Xz+wkdqVmxLPG2BqYErN065hqPbwljzTwzXHrdmR1cbeOEJulW4PdwX1JYMO
C9UpPgMP5Jzx5+7g/cmEn8BjxW0gHFkMxLFGqe3ZXPoO8VJHnm0n4AqD2LOrS4jD
2q1igXwEf99mskvoRTfvhEAWzNazTP4nY064Di06xUxf8Er6uGRunZZHEV5PYJTw
kAgb1nY6Cro07AZxZHeaT2CqSMRs7D60x1c25RzslNafqYSSP1geY2UA2N38eLgS
9uOD0eiN5sptWZ6THfwTKb3fVA9fQD16jO1BJ9HKobPpCM9FMMV0TqNSJj3IdRdK
/AY6gwT2ASoGffBE9gANCNDFHNZt7RH21pWf/xVUaZmtu5ILNPu+9m2LuVMMdG3J
LOsGrVx4GyE5pYGQSGKbH9Q59KVOnU4efXyoLMa0HiBlFTLQV7tO/ORvq0jj5U9C
e5v45cQchgsllLtG0qfeDd+sDCGK8rm4RYCMbG0zKx7dvzYvk8wsyrezv4NGylt/
m64ee/9ae+23Hgjo3cfzfEP16x5tA5pIeKogGMYWcuzrOKEf36vnFMn/a5k1FUS+
JtBPfVdJOfWBa/aadsxehjZYembHU3HVdAPH0270JH9MvfiHyNoqpMAEo/J/2Blf
y0uHzoVDRlIDXjRKdU81igBF3EGCs9m/poA0oB64XP97vmDQ+a/vbxcD5eQhYEM9
SQH7NtotdgwVyRjYngb325z3AfUcW1TNeAgk87YcpMCkhLWNmQLgiin0yp0tumMK
K+QWNkYRfh2d359S6OMqloSo90tAXEtUPxzUmQEF8T7jo2YndXL4JBKKqb6zRIfb
Dyt5SXQigNio6Z7v44pKrhPWhC8B1LLslJZuCTCOvplIGdH5sUiAeqhh0AfMQ+HA
CA/fekBjb9yhg95xUAq1GXKEpRtcDqZ6+CC2seP74HfcCNMNzAgqw7eRuvGtSAIn
v04q47Bdy7J3wmrT4sskl2QzHP+REXTAKGD6DjKGDeZSjHH8T8+55QW55bWBsjlR
ZPpwSa0Ykf0jsAIRq4daFEn7NQq8EGwozbun5A8wydO5qTHN4ShiTjFyc7ht856a
gOJfr/npBLlEJ2Ncy0PIlPMzZjyO3GMMZ0MQy2P8axUF4/qieogH8Azdjr/FJTGf
srej54gHWS/+9nR5IEu0bVHRDTDV8xiAm4aLnwdNGnE0m8hGL9sWKjfbGqbH63Fq
P5i34IF9mgpxD8FOeO/Fb/mDBqiig7hqTyU9FXw73zBDl7nT+PB4eacFnoKYyjsd
d3s8KSadTmCIo0/SoHDdJhoj+N7iXnquOPYmlDw93P8wvlg+inBBzu+G51P7dtZU
bhyaehr1l81IO3QnUG1c279k2SdKKQdra0Jo9jfzQlaINAHt4xk1CRy2kCrmG9Io
RhVRZJLMUZ2Ec2bBJYYydz4dRGL4pd/GRTT8zn1t4jC5Yh9opG3f5UksNqv4xFOu
yh72LwQIQL+QgaA956Q+qHGjsxSG5WqCL6jitGwRWKHGsDN5G0DTR1QTZYKo0cHW
cQOWKWBu0UNRH0VDOitAkyFaxNqbJ5b0Ahq/Nrrns+K6aGY4PWFhd/WxPFqa8+uc
3/dtuH3Nc1f941RVP7vGHYkYDz0L8o6KKUPNdKHJPpUo/b4Ssr2qQFJ4SpFmrPwq
YVT6uDmL28H8YQ5sXcQqEPMJt7dFuogoUaMSQgrtJEnj8cY4noBOpLal6/UarDxx
gKnPfe9Z+BZLp7hSRugfVxwkZl71HNUcV+x9Y7SX4Ipbcsk5Oj3ez4Py5nwNsKMm
4Sb/R+/TxjPJd0hdTa4dEg8ag35bHga+wwwlxrIp7KuYO58QIz/yRTQK6YuB7Ez7
8hLhIkeonPLn/8/WVe6Zow==
`protect END_PROTECTED
