`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m89tOGnXpfX8bN2ZuDNiSQESv2nk00CY8DLo4CTtrx9NLS3sJl6IBDxabYjevy1L
BrHKLwFwVn7jR8RXUaIt2uKlU9bGTxRfiszp8hS26iEnzBSJIbt6LLAbsKlpqQv8
GamCim9IHU8pkA62wRTwf/iKl9yk2ukJeNctZnYvqksfsQhsllWsjBHYXz6/DFBf
0xIqdNBH1JCCcwSp+egcqVI0e9Z8y2dnedmLChYnPMa4W4yEDRFRqg6hdkvVV0AW
lD4jgu35qq3jdW5YZBSVRbr2IMFzpQG7f1Bp2i1yCZ+WgfRvGyf0X4lYLf8zOSMx
ymUtQIpcpiAgvjASVFIAM/p8V0tjdHB1MaYKMLM/6t/1tt1bjp0w5wHCee7QHmS7
Rj34ETbg48rzwgVR1ZPTVTqzHvB/dWyEUbTBdyEYqCe4pcRpLaskX5h7ve4y2DP1
iAGXGBEEW04PyY7eQCaujDY+UhwwbcCznR7TGzwXPsXbLWUAv5F4deQBiW+FxXQn
H5oam6hvEUkGDbKBvqwILTXA4JcI1q5kCJKxnXWietkTJhaURx77XC0DxQ/KaJ+j
ETraX76GAHJiPNLGbIojm4eKAMldAsfoZ5CG6JcPMCM/H622/rbKgY7wycYSK2HM
jKCmPnZtoaZw9V/yCXgr7wq/o71caucHCZv1I4ZDKQNieK8O3divVQETW01eJSzN
B4Y3fCryaP71Ng7gEAyNstp3GnolT/KeDaAY+Dvy++Ujeskg80pld3Fyhq2zh5k+
r7B2IaoCuvbuReQnvQ2ZLFH3O9ukOQ2BUNJwFR98fMxbAvIEetblZvkTr7IuBNX8
QWL1ry24UbMd6nncK6tG0O3QnduP6ur57GOKtmPkR7TK0CkPI/pE7QuWV8MZd7n9
IgNRwdGdrFzeflMTGl+fh8zCZrJ6ckopVZ4Bi4k8e0EpMSZLnyBbh6lkJlCBsrjJ
OM7v2bjQh5HdWWvJTOWzrxKBWJMAkXyP5IZq+sqsA/y7g+ci0RdRzeFM/ILUzjeK
4lElPOJlUHfVILiHkfhF5+dpz4CAyR7RvJFUvep8nJr8W68tiOh0t1A5BHJ8DmqB
WwswYgQwQbb7I9LNeMk3l7YPn3mNMIWQGvoSEeZjDLjmUeKvEB6LDPXvF3HZFJDP
WSuGdkKBfJ2qA+OVcmpO51xcNg9N14/WXuunVSo0+U7PFx5n6dU6s1pM+mwXEk5J
d6F9UO6s6m3jBXqr/GXCgehUkD+so3/L2kTCjIh9CuDqpDH1TLrEj2KV8KA5LOd6
j+3yj4exdgQ7yDiiYOSQw55RkFJsUJDLhVJG6O1RhFsDr0rtfhMslhrvMdgFfwCu
LmbDm7zR3M3y89AX/UyqGHii1u+3FpfYZRpJ2Jiy2M5veN5oGVCtgMr3r2deQnxl
NGF1VuOC0dCi6LMu0srdGfjksI/ooyLIY0p5zirEpZPIEtGSCDGJclknEFfjEPS8
aiD12owHL3+HkwhnjJNQeWDIwc4vAp2amv8jic+0rVdulpKJaJK5SAoBY87qC9yN
YEQViufEIPGe8Nps7/inBDchOuYrZ1hqE/URKHNnStGsv2LWNA+RSqVN3BehP2FZ
mgaXat8dm+Dkh5ZQc+jWnHfhP+UMCDQE0N/3cxI4m0VPitRseT72D9ZL7JRSOC9M
MUSDAwvtHxtwAu4ewvuMj7ZY+HE8/QiJw41gRSwAC8M+F8U1XchMeyTWYmP0HvOk
RYEyc0fgZfu5Rn/4c6o2fK/w+dN+5XEn+u1+SE2iJLXa0wQOmEr/GG7mN+14CjtU
X0xZUy1gYpGxkV50fdVTfheu54ozfpe1mfwpT766NEg0f3mAj2p1vCJY42Gf3cfj
b0aq04UnT784RI1P1pBJ2epQvFU3bWz6NtzFE+llJsSzm/Kh3FYYUI3IK7Eizv8Q
5pgggShDEq+LfkzwrOleEM++cPmwEkksE+Kdpwsg0yzgLuUv5lxoWYqnp4la2bUj
`protect END_PROTECTED
