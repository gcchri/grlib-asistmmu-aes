`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q8nrZABvZTgxiXc7wdrLnV/lLfVzaIDs+8tT68y6LxwngFRnES3ICc6RCkG/P+qo
A67u1Czg3Bx8Zrc+oGcWE39O+SjGOzSCQG1i4062IoUz4XIGNzwFxxg/c0FsGT9P
oMq1BNDtDK5IZ+e/IGbNOPOKVWADYD7uhrKNOnbe51zWjoRLIJdJ5ujK6eX53utD
HaJ6lJ5GfuZohyNz3cQGiLP2K5OWxxaApwicOFFvzVRLqZ/AnhARn4JKYryaxCEg
wjSMLEmjFehuNSCQTPddcJAaPzE1cVGpWPjqjA9SpCZpNd+aP7da2e0Ki9ME0Ti6
`protect END_PROTECTED
