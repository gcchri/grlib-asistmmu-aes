`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tkvJYPXQUiOQwmYxEap3Lt7OoZ+UGK2x/U4WKGkIaW8lJCvDBlfUmaLPxGyQu1Ab
DIHos/omxOmZsHac2hWyzTEgqi5RNcIx8DsMmHd1+HzYsTHt+H7Bl9eeXMLwo+ar
g6vXQsqRLKJk8Bs9CAPXfUd/fOGIO6uk2I02sUXdYw+WYnFhyfusT1pDj4Suof83
8oZeUVYoreSEg7CYsc6/VWW48QR6V9z7i94q8t5fbdfagiPXge1MRztFExcgT7kC
7IBOCucJ+CpngLOXRLYL/Zxhfkb5J16yWFvmYWVBn9U=
`protect END_PROTECTED
