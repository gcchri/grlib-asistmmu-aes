`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LaYIGFsr95AJ4jkp7sp7NdKZDfwuvbmwV/dbs6mzMyFLhJPWS2pLmHMaviRVmptM
ay4YDgdB+bnJFJAcBTDOFdrm2YUgpDUy2U7iJDwmiQikadKk3TOoa4HgmD6K+3bq
hq37J0N6Lf6ZeFc+4TEqbSS40uFc34ERkd2ssfyNr/YT3YSatE31XI7tGpP1MiiP
OedH4XN6easKoPXO6kQQHZ0aQ+xhfBPPmujnBJ6n1U95TPsCvV5wQMTNXGJMX9h4
2G5rJy4hLOHf2c9TmrqcrO4ci5MHVgX4leZ7zQUIYTXckQbfC9a0FBVkbi4vfGQr
EBTYElAFtOVkdOGjbY93QJ7Oda8k8Ua6JqG8YEPZ+VPUq67ovL3BRQ7Zu4pCJnkL
FZqlcqd2SR86SfkW+Oi5vkUXP4K0nTXUzuN5ZJsz35kS58ON/sQN7TXCvy/oG8HV
XkzQTWjastM/lV2BeP8yXZZil2okk7H0P5qlhkjCcozWYOR11Czzi8QaVhLUa5EE
vxxS9OweagTpJ7et1ckrZco/5iq2YAEPHz3XC6a8W4c1jE5NtPPaAYmm5CHrMnzM
bjXDZC7sAN3evG2ONSkcyCNpqBamYMtyEdyRrjQFAm5aCsgSENg1UVhCn7bS3PBh
zssoRlip0jYprFXpsXBMjp7jSd/ro6R2Q3N0W6QcAveBn1pxrzHX69En2WyTeZyN
wbInOKLnUjAeih03lheuPhOx/TcGTlwzJPrxL3t9enOGtqDQxzfzsFJqubY2lLvx
pYnggQqLSbT4wdAvl69KWYvmw5M6jfmvqDaZ3QiLNJtpJymTxkuJ/0aBmxxISVMC
G5SqulV0gkwka2o16ofG/e5EupJKeJtXEXShm76AjUuhZUwg7PLQupU1Xr1/OUeM
Wo5WGzwrDgOk5+pwJv01FID3QvyEokTULUMh8tozfAEddxugEo/mIk+LD5b6SaBW
GUUPaBpN8m7Oe57+KJ+7oUxEjF81Aqdkic1+ixLuzvOF3+vFUfdlTR+ZqaTAaFMQ
0GSaZEMPVSV/Y2gTYMw9egovgIpwCgp+0pZsgM52h5ka8M28B6yoVuI1VYPx0Xos
EWRtMRDDCvssv5gkohU6EML9Z3AvQlNWwM7B+8znXkjf9QsuElP+YcI6/DiXBi4V
`protect END_PROTECTED
