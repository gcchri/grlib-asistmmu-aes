`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9v1HZXUqw+VhITmEfYuNDTGw513l1GVxZsANPPMprWDmXu2IdfBudc2bckIwXJq1
rq31+UjwmCiR9mFkDAzUx66sPMfWTyOqpz8wvwoccB2eQGrhwgEQVAIvo4DqFZJn
S7IkwlCxcQrjuzkMepPg32e9aMCZMJ+gm3BDv4ehhJquOf57HY2HT/Yx20Qy3XW9
vabVeQ6MG5O5RIY0zqvKP9dtYw37406o3MtkcP39du0dYsGrvmzF9efmcBbSEu3w
/QEtMKafKI12j0mMNrD1NA==
`protect END_PROTECTED
