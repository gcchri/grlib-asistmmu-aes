`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AJ+a7jCfYO5EkcOz4+fkrRmH1Jr322Mo1i6ZkFnME27+sKgZxVvixu1Y3pEtr0B1
BzowFEMI3I+ecihtfUVaRDdlAQEVcor9eAJTK74OOu5EqSI7rVOC4iLTfbfutN23
V3yp9CtEUA1hBj/Cqd/LxCILhW/HxVTI5S883KvbHAwJGn2i+HdArjokHfuY/57o
1+SQKjrkRxDMkQUtxO8AW4sZ49pZgud7G5RYzCORuqv+GutSEOAZ/51xVlwbCq7o
fQk9tFneImP2Nw1EJz/HEsePIh9Kei4egFQK0GLr6NMMenwHdb3BllRYiZVa7hC1
K+dvEf3IMl9dCaET6SXCEt8243M8yAQBsJk3VHW9r5SbzA3B9pNyGCj/ZYi8aThV
blOvcSMeUY9QqWhGAQ0aabZfKE/7wqpT4dJ5Bxztvj19GGnah51MCu7zHEYXyeY0
w+TkZZIYy5+Oe5r48w7XT2rXtwJRRykU07JuBnXOG98lbZr62SKe0VMykZxt+hYp
WcPrO84ywiAYLFG6u2uxiwCzEaBxEL6y4Z8O0Ovb5hg=
`protect END_PROTECTED
