`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2znl5sYyeSrcLlUEAeAyO60cgHWxEWZyW4kvcDKR6oqr3Jb8U+XgmY3HKURC0LgH
sXPHkB53A+Jaj5mqpWCG2l38u2yK6pernMSb0pnHdmmoWS/4J4R/VMrAKvY4Nwrx
NLZgVIKBp9kg4+JsWPHphnerlM+33CmIuktjT1ta4eGH6uesuxkqg2OEuugEjD94
f7DTS+3g5vruQxB8beYr1dhpqMN9cF595wWTjIatDpjd2kTMBNOLZjX6a+sJHYAJ
smdUiePA0OxzOIXDDe4BlUDPj/rK3mpi1sVR/hSyMda371lcI5caajrv9/sod5Km
gXGze2bpFkHUp5EcE68wb1MGqPFJfUr5zcxcx9/WbwyiGABLO8X4x/GVb01jwoF9
e9YZHiSI74UXmYqlMMjRAw==
`protect END_PROTECTED
