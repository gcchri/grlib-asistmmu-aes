`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K+mNIJbs0K/nfO8amt/KUL2/YS7Nvb1nYTwfiCebxkqaVD/R/0k4qOA8n0JqzkSY
5VjZT5sKjc9YO9UPL8nBEcySy1eEWDKfeW7vOff70FkGIxmjWGlXZKyc+TI169zJ
tEt6OZeTrcr7zEzH8KFB4x6DP0uNbOnWv/cqAk1rG8XT6zPjicQ+vbwEB5oaH6WB
RCMeWsW9gejJVfoBk13hrso1nJXHe1lAk48nN51J0qSdEmuqDju87OMwCa0l2Rke
WzXDD3UaHT+XdoD98Ul5Fj1q7/rjCvE3ZRiK36d7yJmhlgA1RfUmgW2T930i9vEN
T/gfP7pNN4lF/80XO0PmBC6TCsYiKwKS5x2jEwJboVsWzzXj9EgaVniFtHCwQYWb
tdpWZxOcLcdEjWGbOno9L+f+wFGPqaIGZpUG6oImAnxYSQTfCpfJbuVYBPTMtbyI
y+Sxd8pzir9zJpJBdqr81MNY5+cX+YLdVxwD0XABZjbdj2YkVz/ex8KIQkZEDuF5
hyb2aw+oOxxVbxMsyA+MLhlFkN7aFM2mw+CvWUmozTgcCZIxtuaEtqepuJLfMLOD
RfqI5pGZ2Tmiuy6lddPqFnxZ//USZzfQbvY4AzJw+GJgItqlb9hH+ymUBZQ5kKFF
04de495nEv1ahiXbHBZnvszTPr8ke7AvT6RINiyWzoZKWSYC0l0+K9xCLoxXda9Y
05V7s9jifzHY3k6ptZsYiIpMzvjDtNiT3A/ytKw3/Vt8N8eSKs35pWsbrms22JHn
/V8ifukMYgEwBW9Kt+rLmlsjN5XqI580nUPgkBsY9+UjCbvBJs1UUxs4vOMQ2k3e
wAd59KdtahP0B4bMjoyRSW/Rdb1TT/qvhdqmjBQMoKpX5LTupJiHxYnkSTehcHNt
tg+PETQlRzgcqv3n35kDLN0qGyv81AAbSxRsl5e5FdLt52TqKhqyb8raRqO0eXAd
WR+MVh2R2mZOtRmxbymvVQ==
`protect END_PROTECTED
