`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qlbyYksfEuEMNfxheFDQDycBglrmUnAi746MqSR6Ul8x8g7Wx/ogQT6I62qbVPoj
em8wbGXG5gClXBm7GQi3qTcz9qID4aly6M/8iYn+wf4R0TKjQz0xgFdPuFRzTFh+
dpGLx5bToZ06fTOQET76aST4lfgY0WosXPCJpsThhe9uID5v7ViFNAvQ4HTYQWEF
KFi+U1GcE00pxURX5vWtbdlKDh25kt4C8C6e54IGMeucm90oD7MTdDIQaFhVQlbv
zGNtjYMTeusbIWvtZ9KLsXC8V+w65nLITucR70s6roumsxvbtVZyg6aC2TbywYKF
VJRLPlbbSFkTqTbyXaC5SSs+iQSNs/TltZJl2nSauCQi/fXiI10Nad4Hz35zLwUr
JULDK73TSrdH1gVvPj1vfQ==
`protect END_PROTECTED
