`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pXYIqh2EF2uv6/lBPTN/2mgUcsxFQVnNbwYr1h1TvAdP45Ur1ugBbJ72UcPQhkZY
YWtZnG9ESgj9KrJPtW1ZeUHlTNvV41B2vshrkI1ZazDZhkM8hHc2HfKfWg1BRYSE
C7uNh9L+hT1bzRGuJBaValXw9h6fRYhBJcE1PXRq87vMVuJTt+SDHGvFQsr/ltjM
YT5Yw2XVb17JXoWO8/hu8Fheo3cIjsxb1iGr4ZyXrMMzpN0hQp0i9dETiBWb72ZA
z9rYRZnFXdlguv4iAkQ6cgGAGuVtKRVYAUOkbnWmZXE=
`protect END_PROTECTED
