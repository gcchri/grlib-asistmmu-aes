`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+QuNVTAfmKzZUdV6WNAnsH3Fc4Tfx0Hz0izNavr0RkLuYAbFNqAiooyg/o8RWfgA
sDC6mnlbSvglHVOYB/JLqQNyuFZVbkmjXVR9dmoROT0WEnKk0gwKCCSiV6CuZcIB
Je9yLAvW4/98Ewhhm88lhYf9yI6yPTDdj8Gzlycbu2gOzoSnI45fgH04iyuLekwy
ctXJDMpH2n+6RpbRjes0mbB0NAQm/HrVMkM3MHjhP6owK63FGwfK36ImvDweatxO
PPX4VUxDUw5CrZk/izo6Yo1gCVTNPhuc0i1DdzCAebCP2zjr/sQgLZF7B5AxFYZy
arHEs+zKWutjQbRXNqGZcfOPYEneacl2C71tRUAoJxEyyQHPcqxhPftoTGN6aQwO
SrgsRbrpQitHEisWkhDEluJt7IV1mAOydEbEWMFgfxw=
`protect END_PROTECTED
