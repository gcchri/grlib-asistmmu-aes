`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7qcb8DKe5kNklNf7z9KeMZWGLShgcnmgIve+acXJzEttqumcSFUYS/pDHMY9dsYF
d5QlRRezR5a8T8GpH1VfUa/8Q6V4Lw8uypByuQb68+aiijfJvlPQWGM9Qtp3qcos
1U5Z4mK7mk+gD3BEoOqwqXrbO6TYVcc5OcSk6dXOXW7kStfuwDtjghR7Qe/NHGML
iA951iKOMTsb47Ty9tYq2hSe7cOSpomIPWqy7BEkcxRV3Qe2HgaefkwM/UWNymOa
SKABzUwUNk1r5IICrZJCy9ta2QkZcPYy7TpNK9uZOqDVEGw7E4O+C6JwvtwPrJiW
yan3aLoqsYW5fIirzbPDXBXB1BTKGHctHvSyAt6G4eROhocmxpoifhsbcu9rvMY/
6pmc1sEm0eaEwIBikHRFPDwa10vibi0bXuf2KUkXkcPpkvjAyPUZ05mbillB7U3s
UILtxquV/+s46F1rtXTer8g0XcD+/6O3KwSK17GeDm1SdXN1vAMvb1FN0CVl021t
U0Q8YrcsRJhDC+m42Q+ghy/5yziU5GTr5gmhalopA3+QCFFl6n1PMOi7Fj8P5Xqs
fhMVlkQ/alS8+Rhk5FldwcP95+ccQVAoayuDoB9cQibYyjqGURBtfXLgRyL0BZ5m
aBO150EGPIcG5CnK4SmqEDMhMKhpQ7VzCyXKwV0hKAMHAGulAPUfKMV96Yw3lx+Z
vX0qW0qqHCjKNEq3kJ2REo8VA3ikQMORcEGWxGJpsFZwPkytloeWpRL1THFhZa6u
WtEMJtMweegMuYnZpC7XbG0fXtyxNkgZ7BNvSOvFmTgM/KHYAxO5077Ii91snnYe
LgoC0GpQM5E1j/I6zmsoXdn3D+5i7ZseVv73dN5esiCMt4MGWfhuIVvdN6yr1RSC
cGnfaAmM/3KsZJ+o0dTOGzp/rlTtOwqgJ1y0S+BCBsDlSMnIvY0deP0qirqU+pGE
Ht/d4e4LWj1Kmez9MKdmUTp2UXnZi6LfTCHJ8pNLs0FdgGpCjeauylWBAF77pHeG
zCguK1eXPszl6l6y5cOQXg8cZDMgbK7+o1zPgPzMVhoLoua4APu6u/B1ysSn3qy/
yUZKMVh+jSI/3T1F6+IFxrGWqiZIv/+TVoKexdci+nm2qeCp0lykKHOzIy/5xG/1
1BbHKagO8AJ71dohW/LRmHJpfnAIdC+F9c9j11KnBq5pMVaaSPqNQjJGRKZ5+q9y
3jCjbzVD4eCVCfdfwiyU6fJNqi9Do+V1Aqkv5RP+nMdT7VgkLQr2hqsOX119wGeA
Nf1zjTg4kauQ7fVBfuwB+1xSZpoTfoj8ayGYxEStESzHO2GzK018I/yyLsHJ9Zbt
1GOJxg/VNH9ORJXGal8nvGcB/YOzdiy+wMouNzj+j0imbP2eoLvTe0YMawOgZIQK
8wcfHpo3RhZcgFIbyLaInWAp3TeIvRGN19rEeppnvVmtvP2sg5UQ6r8AvNtJU7iU
iH70FYbagqFT6t4rLRX4Hm1rhDl9v1XLktyKMbwzKyujZXE36WWx3+PnW6bkM/24
V2AlSd1aQdDUZ95FZg0x00LZJ3sao0RQIX5AiRAt/Ww6B3NcW5y+QPYJ7ngVVa/y
crXCDeOyGoU14jxKy9iFz0Wy5Gx0EkN3l+EVNM/pgUYSYxbPcF7vhESkeR5GEoX8
iCi+3P8HD6PM4nA9daSeCsFXCC4aOi8oohTr6i/r4xWiE5eI+E3SW+O9dt2w8Z1V
HkOueIGsp+od2bcAkRNbsm0xwVYrKK3gESyYyU42VX3TT4KS/J5YkHwx8HE1n9VP
TTUjXGNXV3lfmpaBVMQpDK5AzYyjt5ZnyQQBpVMKWci0yHa/qc7BgqZFbFqWug49
6oGqv8gIDon6FYBgw8Isut40QbJNXDsVdpMfIBKbN8W88PV/RV9YKGJozj+7E+fO
5xh/3Q/X3aITDXnsFCpi4Fn2RRzAWuzL8EdmP+TT7JcEkzZjDcMiut6ysSMGiQED
r8Vb9WxX72v1R8oVD0vqjJK6gseRS6EnyVPt05+ktguQUghK9aXZGq6qVibMv5n2
YQnvH8jiMNUY9eI5HpmNrl5Ympd0kkY35c6/5LSfogg1FWQVlNDAwqac7orF0miv
b5uTE/LkAoW6ihf8K2NsmS/snK6c1+yOQ5JlcsU1sug6wGCHa+pLmetumDGkJZDi
RT6bplHcW/AAhr0Iptwl4xMFjsIBHWEQd0NuCA8nfnjNaiJvdGZIDknNDCfff2pS
qrmQCXdBXVPt6uIolvROnhD2q0ZaM5zCb2x1XgdzVN1mtMHMUKIppvwftx11FLDi
2f2gOLC7iYcC3VgaleXgO47BfEsCxOFu+OS/gAQOqz0w+e72COl2lUAE9BOyRRY9
1yZ74qLPaXxDiyTE9/hj0EgzUU66D9ffGC1ftZHqFjQ1pNGdhWL4oHPsJBXTzw2P
dTsmAhed8bxslV1Ih11ZL5JzqwBsMiFNDhK63i4vV82k5dQilvhOigINUCKmyHMy
i8nRdNc1Sx6hpE9/DSr4OhuBwKYSmmVwNgXN+3wp1ogUyoYTYnVm0xtWXINzGi7W
EIRpvt7W0GD1SciIJQdJgeLhEHh7Zf5gW2TiUPH3FZ0Agu5ogIBaQJd+XhaTOq/H
AuQzFGNGD6MT4CmQDJN7PuX79/okq1h9wir8wYaE4DBtCwH/6yVebnw7wO8zc0AI
gEBiMOMmqCdx81u5jx6VLiNGWWJPlD+L8p1/R0hzR8pQIyl8OKcl+2miC1YYAYEC
DXdBspZpJ5EVoBRGX9V+V3EiPLyH1eAgiCssAFt5O0VUgVM6eCtFr0IQ73J6ouAO
54onKhW4F7Y0uWbeEseesYKqYcy1LRvlOzsapN6V8k+e8ninuMHPoQK+7GPK4Wot
rPPKQ7i9kaGZOwqV6MTNXCpD9gWBm/BYJdoA+lQcuHqqVQZcE/AZ/9e5oswRNDc1
08KVnBeuam2niLXfi31mOlHwjkQklBZNBQKfuphJYRRMlGexxjxWt1Fgl3nnMfI2
+iJvPm52dTnMQ7sa3H/wZFpMXqsl/uUHQi9S2jSwB+WGhdCwu3UTGy/dtv5r8KNR
8sdY9KYDfZFYFtrzJ0KihwY2gTFfITjMX8fpwLebzFoCxRa4s/C8U5Ei3kOTChuQ
e3gYAada1xfPrFH2W3NZHJNcnN3P5Cy9IMpeucJL2l32sx7wYUBKx8LcXeHoc2ji
ZItYPi8fOO6GxqiYrl5lCsN98aVkcC+eUuV0RzP2nCG3Mew+ebmHHAejt+G85eRQ
eb4oeGmkkMfHeyutTZxe8Ko2qkBhbfEuT5rRf8JT4MwH3fc7X76D8GDneXofyGiF
jB+nnqRmn2p7Po16E12Y0+niSRrdgsMCF4nxSGyT/IRZ/7YkO1/H1U16/NkHyuK4
P0LAAZJgQR5/0J6W9RmF2uJyJIntcq2EAuaG41BS4qoUsphLMXEBgQAE71s9HneO
Aqm5cdB4+TIpe3ieRLkbcOISsH1qm7ETR+5XGUMvNwuEFSpzX2ewGy3yDtm5DbU8
P/QtVodTNqiiaSiLc0E6nQkmAYcU1mDg9jzZ90JxM3rcXkKqObyJzFOw8C7jfKPV
ULBk2ny4IlT9t0Fa76uoFtYEbZkfsOHzmqSsFda8cLWvh/2OPOGj1lyzdoShxqUn
6rAHGLZIn6AFmxfCeEXb4jms3kLhzSGyRhgleuNzJLM4e4enVRZKmUFbQyiYpKoC
zK4PY06c2M6NAL7GuHRxZi++V9KdQXuOEHNt2LCd72AP+bCnGcr7ZUdFJTfwgZj2
VU8zh9I7ao9p5l8h0JeZsbJTgPL5Mmf0Z2BmgX2GcL++cxQxdxyUzWhl9lpQlkHH
QMAUZoL5tv3faYRjBYXGe2BsEpexp1U56W7to1MyKZHPurAKn9xC0f2gZKG60vmf
+zcJjUb4tJw016fJXEme1E/LtrDT1QeXGtKYIBI9+un3tSPv5/93JoiHtnkQCqjb
K+h179c2K0MgudUsW+HhUP6Mo/1UqQryTXkOXKEBKZk3YkxOkPh30xuipQfaJnQe
hwywHyQXm9VXi50WA75d/Foy3P4HjGg71WPbNuSw5y8yVxKUDX2o3zbd3iKns/oU
xAM7LVFqRu58Pppk++z9sqy7vfm/6zoN/7NJhCODy9rSoTzlAgx5Ptv+CakcdVFR
QbL6eWVXDGZrICCJqO7vKEoBbbk1CuArJuR/zuOpwqI7N979Vvv/kf5WsN1GA0Cu
uFON0ECs+z3+5LPkCVXVePGbutFOsoF/3JVu744ycPBTBjmwd9pi2m8Sh0vrzZfW
kTfTFsFL9X8IOPJC0ABoJWQoQEiyz76IL6UhhgWY4RJn/u59jGKT+M78xO4HQHBh
dh22ZjzbDIAuF8S00gL/uRtJPDMirpqh2sGe5W73SpvTovhNJlCLDiGZ+cxMK91e
VUsgxH4IjpBBA0XOG6N0pooSg+nnOMu6Ggq91++rRj65bHVEWMSPhOxnUlW7KLwY
FhNTSp6wk/QKzhrpwboNrs718ksTH8ZRmSV1DhQLGpkUhvBPKCyObSZRfkmZxxZC
hQmE2wd3AP4iWegjsB4G/x66hk4I1P01j8HImTVQyfpUWOwBqpNZkal/kHbAaZY/
82V2ZCp8LHTvheuvFXa56Az4XL8lJzudAGTWeaG1zkAcnUKqD4JQYYWGoiM4Orv6
Fm8XGJt6plyXDZDXldx9dGW1VyJi5WtQG3w0reQ38c+1vlvKgspOSixXXjTzDHYG
yS0j8MXGspRu0bojNPybuMki2lqI57rPltO8+yJuAXj1mUV/DA2GD6B5bpLUcFql
3M3UP5pS8z3mSEbRtZORjAD7+k5PDZnggwTFVUebmTvuSOjp1s0h/W1YfSsJGXwd
nBCHZ+K6gZA1GXo5vZjWdohbcViP+5FjMNQynWHlC3cl94xT5oVGL5pv9HxRAyMn
GrHNm2T2HjU2pO/nvQP2YrPGitVMtR3mq+2LB/YyLrFKrKrBwkXXmiim50/Bw3ZM
YtxJwAbohTvab+lUNxZafJt0okoFuluMJAulWYhsg6/S2OGNXsjPso3cZHwk34zb
PVjsh5v+tiw9Fdyx+a1ZVsejXKrkSLAqIZa2vdu6Nh92O0Og/wK4GHCKtLzihKnu
l13NIBPWnLV2eVxKxVJrM1t8a+mEZwnUINBr4wDX0cj3mWO/By70Aqvlj3wRj/pN
STMHxoyr7BC2otSorQJ+dhPv7l51uuSTgmBOxYlHWLYYFmqs+dsmget/m45QoM07
iaHIfpMe7bVkBpfQOw77tApBhyh/XAgQiTq36qgu4fouPU2a4t6QH101Yh00W4HO
q09wScJNYHvMkXlW05C8DB2MZdSjV5bbbjy3R3LLsoLIY7DMF9jJf0Hg6D1QAVh1
y56IR804ik2vpOl1Zm+ck6CrCQ1h3xfGL/WVAR1tN9U/mSJ4qtVT6A7iflayAhKh
36ZCr9Irilaf0sCGuGPODfupIOISwIW5CqGeCbLbMZOK/QYPZZVdk+MLqjOqFG0P
GgMeoAnqlDIYj6slmhB97yX+jrz+qjgjnen67ZyWZ1K7RYLZlmFkavreDtDBmm+7
hongUtmc2rmGb6o3LF+8olVdyJQJa5p6mnuk1LTZ9kas1lFqydtDzI+Dp1Jkuty5
QG8Dl4FYZKs6oBCCcbmJ/G01w/HFxnY534mdW15b5CjBL9bzP5a776ouPMxGr6G3
1f9hUWZZpWmYXnF5EfxvFttlMheIqwgzAL7fEcXcmuWR/urvhXlWg+KQrjzFTaC4
nHo3n4smpj8cu44IJ6NLAmc5/+c75ZDPZTtybSSZrbHhDrwPDSvdyAf91WdXzuWz
z9U8Lr88nh1KmkSO4S/o6MW9XSkoxQ/IhTEcHWlHG14ieCIfG+sArHjJXBb9GwWv
3pYZpJAx6BRueCmSYLuWKS7u8Y6LTMD7kADJVquWcqSVtmJ3t6fjoF3BvsmXydbz
SPaLs0MfvzRG7rg2mrilQ7UZE9yzAEvByvDxWYVR8nBZODUmXWdNQYjJQAT/SOkp
WC1EJziWVrOBsiFzUxBo5KdDQl8isagMQlopQIdQn8k9lkJ66a2cV0sWzjfXL76X
p1ieVgYy6bvbnhesYFMn8BMEXMMwdhgDDXEdCgbb77eUZTcCUBPFRiIhB4HOCFRa
pQz0AeXXJeR8pRga4PNS+/6eD4PdO9r4r9FScvIrsXXUjA4vmnoadSQl2qica3+k
k+BHVV6mKNSLN/FGd4wO45MTOlAfAJZS6QnxkmjM3twbEP8TT8+urZvlziQ9VXfG
wFazwfFm8MR4c7eW/iCON39ToFwFNdm3DgaBUpH9IkoOj7wBWZ9jl0D4G9NDYFHF
pzc3oibI8qttFmw+8dwKzMamNU8zIV0F2kOfU6kNCiy54CrtaIKEpO3wvnT9lzUY
I6FASL6pUU1nhhS2UfM8Rp4/thNkR7c8OgT2SxU6vN+CuVQD6JS90J9Mb1+v4TGg
z3EJk0SkIXkrHW2lqKKuC2nnkhsgvDEi79XDWJXHV0o2CkPJzL0Q2Ru7b4oKlVmB
hXyqAi2NVzxtygj/6UO03DOV1WWn1MIUWQW023A1MLziQZFuF97QXEZTo9MSprDk
p2XT5h5zVBlpqrXjPcLJ7wUVY+7b/8wP0TUd4+kKPAdCsHVVLp+OoZlTg7XvDO/L
2KRWBJZV3QL5PEkuOwhDzANHWN+5T/ABaX43jQBoSMkry7HJdXVqryrMlxf3URac
uRM3ssElax57fNQxV5xuXwi8qFb6L9qPRGPAJI8U+voQ4L5zteRVVnjkajiI7Z0p
UqYkFSWulzDZIxuh4uM1UInspX5UJscIgmSImOgpai6MHP2v6j4IYKdf9MyoXeAg
xfZvrl7BYfpSfAdTeAlQ87BQPSwWSRL0dw1p88kcGmTjxWcgMO8eqUvlh0BKsgV5
SNXi+MPMwQs2anoMvQE7A13LJQfrM4KjZMZq4aaeXe7vhirY3FQpo/eWCABCbMxY
mxOEA+NZei7sy9Lvk2wWeshgCppSkOn1brCF3xYkaeGID3dfKITEmmpms8KAET4w
L9PFVrsNt57BfdMUhPBU2oYJQ9YM3NHCfdMxJoNw/qrnQjZcB5COdP5ZXeXfvGZ0
cBvPQr1BD7+SXlxe3kvJa7NHeikyroTqqPmC8J3M0gwP4CRN9GJUp0OTRjQ+e2xj
HPMkwCnSSPmiZo5hlwfr1sq+eObQSsdVv1OUnDp/HpG5q0nCm4eXkL3wIJGE90by
1rucPlgrE63OJMH03oLn1qTzJ1h7j/aNXdiEAMdBQbGH2oB6j+2s02XqmV5akTmt
spW4g3Xs1LBYWzpWhmNHnVB2cRuXddwAOyDVMahc3NnIH1l7xnl+jdKk2qIAJo1R
iLoZHFnqqzIiVDIaBR6NtIOpsvAqHzIXsFqqeNFo/7euF9sc2Ml0BT9alefUwyam
cKHWIfxFX1RxdWzZz6Es6l4pua4M0lJ79mpbgCFz95tgELui3GT+/efb3FNwqaxw
K8p1BUNGu3r3jPYSaAnJD1U6IyK5xov4npQS9HWhCneup/GEmag6iNWtf/aKW8hL
ti3cvPFFUipZ9R5zRFqG6fKC8uGoKS7BwVtalzqdShF6KcD6nqMZ8+Y3KB0w2uB5
uz0+QH8oLnT6+rpPcWKV4ajtIVeCoJorb2+50QXoU5YMI/8F4qLaUeN53S+gLb/V
atc6FEf0h4HMpcc3eYx/BnnGR0D8ogamMcv/g9tEjr74OCfvRUNR9WGCpb2+3fsn
DzDVJmQ88u9xbb8zc6D5Ia/v9K03WzeQvlriyTkY7hodnGGZN6Bn1dJMbQWb56mR
pKy3jf6ipraVNf2mB95AZ+oBTKOb6hag16Hw/TVMQdBi5B2LlG914zjdG7fx/CnD
erLNUY4ZYBzTeRHQrMvTPb1JDwoY0pZXWvNh4DSTs4eHPOFgemZXElOHo8sRqjtE
b8ocuGSf2u9pk12P34rqVhn5oEvWCVNXfYeh86xB2DbLW9mngarx5sgd5Bb5UbRo
K8isE2vj+i7c0NbITxKyGrMYmcw8csppnxgOlUa9yeenhEOsLgd8sYuR/Aoi0iT8
nddcL8CtBo/utAWivJXkKiP+oQX5wo88J36KfqgYfu5KPZayy1oY9V+RnmyFTVPa
1qcPA1IfB54iNvM1CZV8AtD3XLYU4JOZup9DLuXvm+ZrVYO1UH9wlGFZ6XFKEDl3
kDPA/d0gnRO0j+r0Krk3dD76NA5iSaAeeDznNlumAblvGu7STtLi+bhwhPhOtz0h
QurqLw9tWVm4x7t1yOjO1MHciYB60lv43dlYZFCyq4dpPyJ8/FJBpzGNkTjkazrz
mFdxguVQWQkEm/csrA3mwTAUzse7XRX+GinbjPpGMKfYaJyrDYzBvMIjPj362SIn
4issnZOytKWco9QdpUEj/AuA4+4GKg8oU91wRYgMPMK0EBXMeijqTe1XyabogRp+
4TB8AIslelrUo2HN7PRzPMORXv3AX+N7FLIPTp7TB6FXxKYJvVRf8Fayp8jIx4UW
UBJ59MxGG2eIH8t5UX+DKqK4SvazdnIqzVEtHDBvw66WoKpXb2+gFZyfcaJkAgIL
DDQvMDdIdBIdJkCWLr7mZU1FJZDkVC31pO2h9AVpqPVkdhVTctUCf3URCe3xDrCQ
H8Qe+VXLBSzPfiopJpHg4nXrnqo5bjnOHNEAp/3i4uMiNl8ZLGBUiNR1fc3Tx8Ue
9QtJb7BYuy4dMpSVqWIskpr9cFUtLF+th73rigQunwpzrayNqDD/69q1uSHR38vS
WMaJbOKwtnjS0ghgfCRJlnvIMMF6brUKYWof1QUwVwGP4/VKHaMrON/O3PM+gk8E
pbryLlzpvMovWJO+JpkTH7cZLSYhi/hnd9Fs6CylcKttwx4L/K/nZ+axBrRXhHQu
5OBc66Kw3fgr6dc90tYIeciChtR1EspV2zPmOQ/zkjBeDqy7J/0wYMDYX1EYRTQs
gofA61UfxM5wJDVaLmB7ahkdn32kM7P4xa3nFzg/fYqh/M7h71mIv1QRSVwFHYl7
ujUkg3Xhng2urGd7KcoRhFnzQbbmOT9wDl9+Ifd3LxEHy86dgSC2HGtYglvIGEtv
sw1+ftPCuk754Qph5Poar+yK3e1b8vciTL7DC4wj0iPnyMhZACEGWAoRd0r1ZY2y
I64OiBYi7b3t95H6HEqr3JaEa0rTKPELNEfDrlEPSa2mLRJGyTIazE7pnBMGTUFA
Wz53zJ6A0SGnX/R8AnVUr13n27skOsKYJpOr5Unjuao2GBq6yX0wtBahGhq7yYJU
flYPT0Prcd9FbSPIfRiQM2JP0sGb2gnoVpPCQkltzubARy3pWD7ddHNK0AXnWkTK
SYFet6t814kLlRj3yb1Hw6e8bscuUuTbvVDXg7anwG+yDCfaqgaZdctCrgcxayZ/
LQ+Ygz0cgg9F5HsUAuROyt/AS8RnKffr3SRoHNUc62XLUc9vWdwVpdNraphXl2Fs
oEQixjmLvEQQZXaSD/oLced93v1CN3XJNfMr63HX49bMzwHir65eRe7+h7nsNFrI
I5DN6TCJATkKyWGv2fE+eS7FXnfKyIk4ISuhYlhCMV4aNY+dvHdoVq1y2RZ+TNLD
AHULWYeBVAHAdDPQTt9/MqmX0Jy8M+GXKhngekfBVqzqC7PygBPdkUhCuc9rpE11
I/a4YIaGnrcmiKKNxIXpekUYkaK1wh+9r1Yr9MLu8/HhRMFYF5BtceAal8JZYqwv
8vXI4UGBbNDGMLhVrzqizHV3GmiqTMpYMcVdcvlzUSwxj1e2VR2D1KUyBAh7KE2K
jDW6OAIZz2WlDSSr4GZ7GzoeQrOwMjE6V/MF4QXraA6V04qwJ9dCFH8AFclsN5iJ
aNtL/w+PHVjHCMbOaS7ar2gy9viCqZaVjsZdTbJpM2Xg4Vw4s645waKQUqKL8VTw
ArY/5AKxUHOoXC+g9Lgn1noJdt4uVX/0VY198QTcM+e3njmtek+dIt9SnPLOo6dM
k+YDYBfAk94w4o8aZyiltmtMjg2pNDX8icv1QdmhU2veny7OlELOhRl2svoNcbKm
dzN5IGjsA24V/rJE4xL+T76jow/zJ/VJOKFwhpyHtOgSNbtdlokaIhUDfq05UKGv
K0FfsY5ZLtZLi8kfrXAMDsCGn0+bBce0Copu+bcvT89BesJx73qcti7s1Msj7147
c+rLWstgHWxKeobolP0fp5VlQgaR3QA3o5xLqgcgsRuTfQ5xKytbWRyr9Jb8XWr9
0ItcBF+5+wUUjJ+ud+jp4opVHRRBXqg6KRkGib81k8kBsfzwX2osG/2Q89gptCA5
yqja1RQHvu2b1/xdXse3Ie4S6Sl2OFYve6CpkEq0JYmeY/+q45GGmXpcGBPn6lO8
A50ZpQhzKeHmUjomzID5ABBXgCED0itjCNwlUOhHS9BqEZjH+bntXevkDgC3E6f8
zTXrfKxvtff1GvRRvk/E36E7KYiz1/5lLUuUTT47kdtspXBVSMDZ80SMLp3byJrs
MEO8sa6YS1zbBTbYxNabl85YyakN1BSiU/dDz5xQC8y0ifjcY6oWHwCv4dkaHhYb
70RPFHx9cffxSjLkEd1lRtR9EmC5uhnv8ONCCgd7ldAXUPxPZ6uOEssicCJjGHBN
bB8HB6u3jTvNSqft814mr2s8rMaV3Eq45mnGQVEkLvbakECZ4YAU/SN0hXEd5WG4
vmZkgSDvwgnJOThqkmns/XGYHAEvIM+Fy5c+NDcTeoqPjzWLdgOplwVuZzxSOw0Z
khh07281d25DB1z6dnxa90SN93OIk1Xx4w8g/Bb4IodqgedKl7H1EGOqdWduhJ7p
qaVOgU69Ewkx5AMvdnIWhQHjbI7TSqDmfRtluXKjPFLjIBtDGyi5zvKRTZHDndW5
Rpc9LO4zbHOrtUowxpK6US0xKE9SWQpnT+hw/khacuc90IoFWGzINJIbcM4iZiY6
UWryFKRSJdl+fAMZMS04+siRIx68ddydh/ZXc7ClCj7moePKGW7mN6bX0vi4NihC
p67wZr6QR4c5w/CvHFgE/jyeWFWrIRfI2ef8Uy+C/b8/ltVZKQ2sjNMX+f7cdFCc
fRH3+Vul9n3KBjlqPFBljys3CiSQ/jzYQhQnPFB4bzs7k59tQpfggL22hGKNt4LP
y0xNZnDkDsLw/4Tz88ZEtL8TxIPvG2aueHo838Tict1jRr5M48oarsyre4pGsvBn
y7jpPWKb0k6VaHMAPlm+gcuH9r5OXu43UP3YwuaFogJqQ5x2gkD+XUFdhx6NxFQU
nG03WciMPfvP8uZKSwFK3E6kJPQ/VzJCKE80vCPSAJFxQ/5QdYKIvsPLDmOEYIzi
XaW87yPmZvRy0X6logqGwjtJTudfJ9aDqIYtpatuFy2WohrQag0haUBN+SY28Z+5
Gv4817OAJNyzajWjIsp/Ov0t36YSfyyTQbmFaiU3EE/nmb9bOnims2hcYZ4cybr5
YMbrl4N9rEcVKwm7mssgTNtkG+k5KoB7oMwir5DnSLITziSqIFpY4HL8eRvS4psA
l61RzZT5r6RR8paFdXnLnUqviLcBtDfhIy/qOSe2zkiiQYIZBluqSL5V6hEBEQ8J
DrgK9ZGx+RY8OdxIvo50ypKdoOmeM1IsAi02/60lXjgnCEGYThNCpJ87fWWneABG
fRCGxSO/wr5M1q/I4G/cePN6Oxlzn++0qv4qUSrMYF5dITKC9qa4p/imJ0iKRdg9
kriluOG35EdfXLJ4xsjd0imb7s0zdM9QlX0cfcRcs6zuL9+dUSbRzrrCpeFneRPb
hJkCipgYltaPo8AtWrajZfjDXV72okm8JSffm9ZMC/tuk4QF4RVddIWMMyJzcYHt
6mlXegQ08LsoxxPWarmiT/656aP7ouMHfwk5/om00oBzUcXdmhliWExFP2WMzD2e
qBiJGcYwNNoKj+H8dtBGL8sD7q7tserpuIk8EkjMOoSw3Dm6sD7eoTHAk9y1M21Z
1flarTVmRkxjR0Fc6iPwVm5M13ebIMus2BucgyVPGIPlaaWLvGvx23gheiMzoUL8
iohFeX0Dl+fSFNth/AjrMpUU34tB9o1aZZ2tvpdkltg0xGQFvNAxGHre9AVD3Z2E
d32zKa8rSEZIUKvk22vzglpin5s7uahKfqITnGOudgnheb5+Y7nEzvJrqaAmg0u4
TYcu+U2wL/st+fDRvhAyA83Mb/erbAaNLeA+HHNz186dQFawGDG0JnrkLoSmDdoo
s3kQWynBJKwt2QG7Gbhdv4kKmbpnQ83oGZdZMMbYt7xHlMb0qehbCndwMdHS+cpp
Lv5/+UDnU+L4vg9wc4vM4sN3SCSl4NwbOwQm07QYCW4FXV7skM906NytAWt9nyvZ
3jfs5Z5utkCM+uVNI1L8KGTpmNrKax3gBHPtaYezJzRSE0UdviCOFlp2YJ76GvZO
uehnLE7Fz9PRT6IZzfvvbm2THqz+eeDTxK0guA6XceCK3S3XbaM+4h9GsAb53YIZ
6EU5xTgzo2ptYe26eJ1XoIQXhICR4hvC1CzX6P5hWQKJKTL0v93FmWGlBhXqGtbk
SjUl6U5q5CAEkfW+RSV4QLMTUtKkorra8EG/N3jZAuAsfBdGk7/oV6MuBtOj8ZM8
2MMwVgbj3+Qnoqk8WX/Mt19QKD9AXhX0D3blG5KNhb7XtR5KKW/bo9W1tIY0ZuY8
zLBCbcuhNcge9zQT9Uarw4FudhFHo1VeG2Z7rMos4wZaB64XQzSmf4uaXMLGrzMc
AoovqW98xeSVpeAoKM/1t87OVvl8lNQ01XuzrFd2eTnEhI3W30tSB7qQ8lPAI3GO
ywiyNHzoEgR5HLA5F1FGTXeCdatsY37LvmQB0jiiME8ohwaKnO4FPmyCk7fZUoc/
Ym7n1/dIuxACyvyMwqllYKD2MKzoX+VRx6r3AlqBEe5BY5ypRrj77bXi4omqL00O
zKiJqFECMzWdQtTQdOzpgG9tc107yZXj1D65pQh9dtV6rggWxRrfFRbozMTIW4gb
xhjNSJB+Z57SRw1toCReaeiANiH1Ffvj2+UCVjcNeBbZ9CO1dsNXb8COZiVUezlk
J2LY3+Gh1+eNVjoZIlGSD+A4IxYLrc4wuj9S2FiJSSieoQ/VihwvzbWljLm2ggX4
mp2kn0T7FkI1VW8bguPMNXpNUF+eJnTzi/yBr0Hzgo5rxElv9DOv/w6J8+id78C0
w1gcVsAu5rLHo8SYfuLN1nOL5N86hYSzdzL2v9oxWadOVldMmtsRQ9xlGih4LRTO
16Sjtnk94dlwQZNoGGKApj1WVcOzV90yct5dFunqGUnNIWs8mI6BHp+952gepATA
d+mKdZsl+EGZ6g+tsfTjbZkvOLUVfHJ8MDUHK6QbWjNKez+HJIXVrFxwQFYljMV/
lIHIrf4YrTweDeE47YEOBffcm3/UkrVdjNIdlq1NjfRMNAI5Vtt37DqvSGJO5NlX
+3cNX1lHHGZ8GeWWNTWVLTMbNIOR0BpV8Fwhh81LamMzr1zJvmDuczTuHwku+YJs
Tbn9VmtMFk7zg54tmiqUwJQILkdd5qHtcIDNBmaIXGSBBxD6qySrkzzMfsjo02OK
03rJZ+8dP5z9JFJop0nL6GdAUMHdEX0qMsas0NKAffKq4j37lpD527MR1Py0XIZJ
5RcZqs86RzdyFrnsCAc+s/UJ9yNWUFBNTOuyrP2ASPZr5JEwdCxUJJwpmlmOa6RP
uUKSpoirgyvLCqqA4eQOKV4wKGgfjCZbwHNKZ+cjdGpcM6Cx5ERfIdca5+pa3pFd
vkqbE41bf6+EP0twKgrgVYu8rndEGZsbcPw6oeFFNzG419Eabj2ldqnZbtxsvG9/
U1XZB03/H0KycnQAtHa4fk5IHP+ImDuhfOSkP841zJETrombtknoQV4y02dPoIDd
ZDiKNdZ1L/l+KD+90rl0/GWUnDcIEQ33Bwvk3eHc6w+lmbwvLoEbhRfvCpxgPRF2
cc44fp63mKjREWPvOXrt04dEo04UKziwl0Vgpf/6cm9Ua2vjIisbBsU5TBGa01+r
oTExfPpsrpm4oAetFvOoDnR+P6tbqI/4LrHiRnbGxFwC5OKdEqFih3tr/TA1HFPv
E1PBh8Evjan5xvmBMADD4Lozq+zxjykEg/huxl3D5Py5MyT6OA1e1ZV8bRYa7Bhp
C5CcaL4uuEzCcu7bcmz9d/GTB2nPkC2W5qJYWxuAY64FPXcgyX0VU3azb6vdJduY
+LcEoEyhAMUXx4Z/4mMsO0pW/YjjnAVA6CfztITFK2REHz8oNbFYodJSyqY/vGJ1
X0J8N0VcEZXE0NG1cJ4YIoCo97d8eDFvXpT7hp2ReyCCdvEnlrzClARVap5Qhp6g
Rn72N6SPRAr9e+2FKQH01iA4hL9rSS0p7bnFfhJVrsEljRsTwbY6Hz8hI3/PC9om
Ru7+lssQDv72GorTjyC9A4RMvYcTKQVnAFfFnENeeQ+VNB/uDesds/Dngb50hddI
PnDyrL/AoQMx8BS3mip6a7DqngvJYzwKqbysh+FRyMephnfi+8Bg2hN9TevCnZEk
76FxpSqFjmtWrXLf9IozdSiFuJslK8wsBd5RZFhYzSQETYjY+37Fh5cMiigb4hr0
426gPGa+WWfGOSbVym0PuQxB3SM94lBh2AlKBJ/XJ0If+jm4MlRnM2ahEYFkyKWu
+JVosV8XR7+cmLu5vvZHDnkiJI4SA+UNDTlECDbJZi8ee2JY4rRzU3Zpz/ttqQGV
DriS2uKdY7ixbdjz4QMIa8PkoEHvq/j2iBwcLGGIuwlYdXuEU6kiU+8H0yvWRLeu
6CyHv0KEKd6H3wQPauvVatqW6LwuipqvyeDRbwJxtk0wYeCe9ywLfZNRPqTDQncl
ZKVG881g9JJck/O32kohdCEtE+gPkuBPd3DW8PVg9VrdWpDFSF9mQToUzMD5NMu+
Vk0HQ74hht50J27MWmvnmg7+xe1V+TOrVuIF4wAf8xBBV+JeMDU+EO3EkrttG8Z/
Z/LqIHDxgxMU8UQ6jx6bmL+3IVjhkNKQN15u6TEheNT7ACHx8C+nhFOsy9LVjdjD
Jxrj3/cREkcxL8K1a3WkYV9YD61apE99q0jbSZ3wh0vDgyde+5XuQvOnWFNGeTbf
JCXY5QeQBHLKq0gzstBnlcpfOCZGPav5M5BXw1X4NxowQXCurThLq3bDKR6X8lhV
vT67jo5K+A+UJ56G7zy0NkYLpVxH72PoOTk/MDpm/zwjk2X/N/dKAsOEKeaM3pSg
dW4600HOouLkzCAgqrxnhFp7uFbK3luLzzWkJG1ujYT0KOl/80Dwo5oGhAsKndwn
PwD7WRrcfZSAoaqPPDEciBz83MLIXfqwdRubw3Fzlh3leorANPrH/Sl+TE8bic+j
ksnFpaybrGa4Qx+Y0FWSnGiIRqq7zI3vOKF28hvrEGn9Qz6RlDYP9VK+Td9SLx/v
DLMXvxyb1o+SUhPSNU/UcCprdNxVkrpEQ2DgEj5zmWmp9kjJXFh60dBW+19MuI/T
Dqx7N3ZxcNsaIX6NYJ92vuBHrJZXN0/p7AYF4QjVqktzSUReAZHuSACo6qKvCuZZ
/HLAa3uY9Clfi1QCoj3M0c1MFOIEhXtTnu5lVpYyqtLRRgK2XQFmjsg1NobBjvs6
Q4ZNrj0URYRlkJnOvIphsyTkjqAzi+2jRn6iw4BBvyutIQavosnNItNa44UtxTWk
UaVk3s/4gTsYYcQ1FJioesuy/1fRWFIwLDfdQnlFFPZzlN1SsQdqGDfKjqkjCBU8
uUeLj0tFyaMFslHW0oslxdRFfmQE9kT6AynfqrYrk7K4QhWsxFMw2q3P9fn9XRfz
FrbEd1nVZDt8iXzBqLTwg/2wLFUk0ZKByCuAaVjP4kq0RoWN2GC3boD0BH1/o5Lo
3SX/0DruXQwbg3uVSRNeLrHdSRmVa7Shf8Ce8FvXqLM+nOFKLBQUGPHbJuqnV4yu
0hyQtFG0X7iJwghj+/8RaQKdTpGJU5ZvtCzNUa6fZ8mzJsVOculEK8A9xhlgOpAj
9Jzn0RwyWmFu1YHLSANKpsdv6gjiOuENwmWJxXosEAEOj8sd9Yv9U/TjDEPsHHbH
7Jcr1n8uFNjp8cLtsJ/OPvb//0bhGaL4kCtM+JXxLVDGhXoCxmAhV/a4yPbek2+J
Cn9VN0c0rFAM35qILv++RiuLTNQJF2UBuufCoqMHNqbo/Yp0snYUr/3LicPD/TgM
7V/TOpXOuj4P6JXJBTtzMTIIw+2IdLYih8E0GvexP3SYGWHwwpTXkOA2rOHfVgoj
YWGAVZtI2qb40TwMhCUjct2eePAl4T7wMB41UhSzRk8yATcVwIVNoFmq8KkaehJf
7S8ccmSQJS2dz5Ry0k0ywX6sjcuxNQ/tMa9s7pHY2ubrh1DVz+JUrSrDZAnTPZVJ
7A3bPK7bbCoATbeFb27Fe0/Zs9lj/AadkyF/+aotjKPJdxL7c70nSMio2Jefy/m9
PKz6P6MxoP0urzRAe81FbzObnp7k1fIUMeOT91fx4xjHSjZi7OStEUZv1ihZCN1Z
Z5/uqoTTroXOfea2Y7r/85jlug1zJr1kkzlrmyK34SDAwjTPk5HedQJk0NUrogbA
8rFVO4BERUMqrj6vhkdtuYMvZGzrT9ldoUIbioOdHTBmoLpXxIkAUEzKvueIGWvl
5fD8PZcqvYSz7AbmC+uOo9NfS4UV2Bk7W9teMMM6DG1bgXamMqcJzMFSPfYVdJfZ
2RESXzh/uOBeGe23j2apSJ1+RxJHuoAqrSfFSXjRk4EuzKlcbc7e2+Hs4wTcchzt
+eZZVIJf2Rc576rcI7atnoMMT5rghNQ2wVXXA5aNN+lBFCghUociaZC2/9SYGaNm
368FQWBpdQA7xmE93TvgNoq8hu+VdFVbXF5N8wyRCkypnz1F2hf+ytfYAyZk3T/O
Iz1RpRsdIys4lk2dRiOdmDa+CQvKIHnlqLBtLlhIpQWdcjyla6Iy1spHEnSEpfcG
wBgfwbSJ4v0z413eRlw7rm/CpUgoiYEi0q659u7dmt1aWDF1BfSdxlfBLjfTCeU+
ckMdBIs8cRHLhzTMGl8sVFfFqzY6n/BxQeBZIyKdHkVsuG/KVIPMcTwlARhPdA21
yqOnPlCD75N05k81EUp3Vn5y6dND0+AbN6ndL7kcystxGHZR3DPt2wxU6gp8KfB9
cDXhbD1CFUXuRXQWqC/rUt6jYTsF8USaVz8VQFhF4R5bS1wYt1IdiI9yGtrBKdkv
DsHhJLf1mzdw8SLURJpt11NMvSQZp6GSgqGk7BuK7EjRqoPG2bWD9BqRkvI0Mkmb
e+Erwn7a8ljCsggFIFC47+3M2czcYN6OOPqNTKlgVAA50sKFFVC12FO2Gr4SNuLb
cwSBzvVrjhW4L7ZnvaeGi0qB5Sgmnu9FBiCrX/YGFeoC5Yi4p1IKAXHOLuZY6Y/j
KRE/VxWb+gZNalGnwYYDpgHwF8niITKaSK5Y612Sz6ND0vI4qY9+Pip8xcSvdcnq
++35RELnJDaEheTSl4OIWkZAbTW6vmaeZF3Ch2YdDRFM9s716g/bwwZXuJ1gazaq
G2DHrVD0RhOXy/sZ6bUEOv+dKUBJaAeKi8Z1grHpv6mUYPh7a1NCfVEM1rVkx8aH
MeIQxFMG5+K+hjCT8DWw+UK9fH62Edx+xetRtU+FpR1SdCcnDp7gP/N655Kwzymx
kXkUYFZ6V/0+EhE+DS3f21dtNzz2MOTn7N0FJ2eSIqwixk4uKsH7KGx39ty08a0w
SX/kXPxfZKHZtMpwNfEeXJhoETV+nc0uD6JpUE8wPmctxXyrwVIergw5uWFDEr0Q
zuts3yCJn2rR37zQlvwLCCcJvikreUOuaRwjd5J+fk3R1QdaxHSTdQO5di3W+Mue
/Mz2xXibSsae7Ga1XpsBChxE8gCjVlmXzQRRF26vrkOWKnF7QMG0fQLimH+qJdFS
00xvBGVTZCl96jpkPHjFQ9m+fzGCFFhYhCaD8JE+d+9Ie73UcZ4Q/CA1dJ2MqJ7h
pBSTuk++zMSd+Bu6kPEBMO4NB1EA/7QzdYzIn68PWVy+kAkHFKJTkZA90wqPrVb9
VyJfiv/lY6WTxRhwEDLSs+iP7Z3re79VZsuatT8vl8ikXZ0BZ9In+gxHbaqRTJim
aKljLMFBO/pYsasgP49/ebyEYUN5swVvr73Q4t3QDEYuq7GFmS+UbdpeHFKs4l2a
SrAosGVvtmaym93WnGxL03dHZZjD3A+56pY3/5sFKVD86RR3KZiMfQkBlfXmQepa
ayWlMQbfFldIwZ152UOkxKtF2L/29w2r8rODPckVMATXaWIp9UJcmZygB3DGphwS
SuLbqXqScjSIqmH2P7KBbgcUxLlAcLcPO63GWdR6urrATJzjvveDk9X1YUdy+nto
M3xvlDMdw5j7JSJtpV2KYu3MmwW/1oMvJl19rQCHP9IBGFGNRCC3FxhI7p8Pw89u
RxFObtw7fniEiwYkxjgsb0Q3aZVkDLiUJ22HzCY+cPPFoodC2ftAc+hu7ceg64Dj
Xj4mY04tagdpzKGdoLsYcD9BGKqHKs3rMDm+VzEQ1nkKrGSmjWioB+webVPhZssz
xfCbAdr3xlm6cSzAHX2saPK/NooSglNM0hp3HfTyvq4U8IxJUAX8dZOyHyol5Cl6
dYC5mDnYL7pSmQCq80y0rd3lgC9rD70oWsNPxKTml8XTnurhhY5ntgwsDw3gC9at
Ez4jt6SqJxKKMghzE3bHOZeupwPzJR17d7NW3rMeDavdbcxfsrUjeGdPcYHlF3gy
CVhqeAsh5wPSSyZrv5kCdwyW7kiBv0Kme2t4Y0o41bwcPxxtcFONmW43pfjQGNn2
Y889TjWZA+VYh6yfv0Ua5WS9Ck+rNaWLbzKJ5kksH2s0q7rgsaBrLRfRz+YWTWI+
0/OfC/xtMvziWxrOCBFKlxvSyGdi+9Bt8/tzV+MkRYcvr0g5t9VYMmG5DVEZBaHl
5D4hW9hzkZv6UbDMR2cYo9z53VqwQQhDICUyCNz1vqGnCnLJPl3d0d7VcaZAhT4b
XMXw4aX4flKGzrws+JwhR03JfDC2vgpSMXfsn6YKSq1ELYI9pUXaay+XYn4ELdQT
rE+4qo1s6mbDfvyAlI4IcL2EN5YH25jwAotP8UFjE+rd0Eya5Fz3R897zVAsLXbs
N5KRH4gfPA1MUE/hiWO3UCcvv5QytwXvtpsnA9Fr8m3O4/a3UnI7s+0MOcOdm5Tw
EjCwWCjiXlMEoAoPdXz8qATgrdPrHBy7gcYmSn3g7TTRoTz/AJVg9FI0kYTJ6a3Q
MI+OHlzC7pki9HwmwhqsFZYJgJzlwLXz2+PIWjXhUQzFxWAxa57dvgZ73UhUFjOc
zW9Xe1FmxltcjQ5bh4bhri1iIh4gb7MTUXtrJMbNK/u+OaiX/pMyEokyyPisdPSO
1LFM85GG0OrpJVClbL0LJsQwPXfyyFh9iENB82insCR5ZmscJC9nD4iplco41ztG
nISpvvDjv0kqS4qvAmEaCz9YHX43aRWZEskPdz8kJp7euUx4+h4j21W5GcLTB7/3
id80yztZ1BrMGd0rJYtIhf3wfpoR4Lbr/1zfuVQvqwQRtVYHl2RCNaMGMbSphH1E
oHI3ZORiHuEAkPy2NsAvypAMSdMT+EwcDL0eEjPtC09nEeGtjGdwjffSWclKUzpC
Z5nK/h4l9PigZK2shGVqnVhwow58J4nkmUKFAiSABtvpshsDSouvaDhpQA4gJQ2H
VrIGTrafcIaIQtSum2ELbmWEVId64VUAMptQ5BCWBpmBIFDU9xC/e8JHBpFa4vrJ
BVHf8PoeYPpUNvNpsXq1F3gMi8moQ/3evbIg56TNLw7RzcRAPKTQ8tnIgRVAHCGq
WZBBrmn2homlHAJSJsX339oKyHMNh8Ps5tWlzHSEXQTYGeFcEJgABdGUZwoUvn49
YzhcUz8jupywcksWPbLBThvyS3jtxNoBFI/0l0yEfGYIzEC1EmbiwIKRAbbyNEaz
iwPzApKvnYkFu7WDomumPE0P9QdmSLV7/epD0hD/bJPSBz+U9821LM0oBaSVD/Rq
dtc85uBvnojjRBg/JaDV7mKnbKx5ffl7oOFz25oxzB86JbFf85qtvxOSZKRF6++0
6sB4ziBpnnFcX9o5LbNzYRo88qpCsyCosB6WgR8PZLrCwBtP8DiyQ5TjfHaJ0Hpi
QxJhxirgFiDtbPgkczpwXwlDIKkv0CN4RSxpUXrrYt+GGmmaY9w088z1xreH3Bz5
4d807DVzOmniJpa3/4P/euJIJDlHPRs1m0e4h4YZG/eSUuFlugH4g+87EkZD5ven
tdhEoVERnRkJDnBDU4OEjImvkVRn6LbL/UqcNG77vLY7KHavWW8+cl4VyebN5JbD
gXGlHJ8LKGZnuFqNJr3zdyrln0MljIbOS9T2qfi4AnO964srHWm0z/qPzRxxYzS2
kyMcknepfoclQxPhG0s16BHQPpiRNV/K6Qe+HX1zkiYtzgvVDu0CnswTgIMYP4Sa
Xl6ZVUs0k7Uo4iFmPnHG46TfDW+elz7JGAP1TFaDGEwZeGO9Pol4lKQ+kNIScTas
5pk+bGvF9F2Ok+3rMueRiHZ53JY/KNgKkFlxwI+11nbkKHIRD2uj8OpHVe51EjNT
l5sqWdn0j04kcReiKMHMUHPY/fyAhf+3smEgsWwAuEcARIiShEExkgDTx5UZAuMR
wgtpP7dQOfFuqX2GOYQoz5WDNYEZ+vDRLEIgUKqB70cY/4cXrjUoUZneHHjX+lmy
oeHBhfcLQV88XNIl6WNJo6VhZSB/9ZSYh+xOrDjkBbxvKWYwqTDU9KXoPKHhbiB4
ceOa7qS1fubqMOabwZvZGjtx5x2WJ0gxdkjSE1E8h/jLtiZKzAbQxoLlTKOoXeyK
qokKFzZ7NCY1N7CikvwZEZWS5VgxQ1ncrk4lBt6KZ97smXqX3YZIQYM6yvJqo/+H
xGsak4gHKbfjfOCKNb0Ibd83K1HhUGLa6aSw1DKx/YD+kIjg3T1kwTTD1YRm66i1
HX/YTOj9pTAxbfDaUg3AMUzM6l1RIqH/KV/XROly9xhiFyjbqDNjhMUNdH80P8Ad
obcP8eNckkGvisgjydZrKc2QWnMm+NiJ/5RgAsvs7soEVZwSeXrAA4+e9nRCsFoI
ji6K0eQwZKFEe1n2oiCK5ZqFQm/dtaUAM5PTkQ/wzbO1iGFOcUJOUsWZNgp5Logm
eMY9F9EOSMpizFwhFUbuXU9P3Usbn6mq4cQLPRCDJPtm340kJCyaxfXq+k4806bZ
IBiUct4QkfP3QKBPp1KmcwI4ONjvnK1WrgqcMA7Y/dsQbh1MbuDkKeROneFT+rK5
n7qw3Sm15Al39B0xv7cGTtIZbpSEivckuPl85EtaaYhrMPd99x+8Kh+qYjwRAM3J
cLJSwteeaz92DYxQKVcZfl6aeX09J86TrRulSpV/jmD6aDjI5Suw6INGzepPvyFw
Lpm5FtL8C/jn8omnPJbKQNQnRsWwqj29QM4HHSb0CGI3t95lJUJQg1hL/xk2wpjU
sCHuXCy+o34R9uhN0o5E1mQ0Fw07A0EIS6Wmkcf3yT7NaDQCPcfm8s4V9HD9+/Ww
OSdJrRF7MJvTzbZoK4YLdWNAEAR4Dg/ae00+tFpDjOnoJLf4A8jWDzQBm1LNK0P/
8FvSVJh3jlgGiYcfmW8UIYRezXRtRM2KrKItq3Sw6O4QL+6E848NR59jfIaGYxWY
rlAQFKkvLpMP6JhHpUlvBtb+A9iMrNvmsVRBW28MCE7YHXlNS5NhnVUxA0tFUufN
+4GlEfruubLloDOT5twONJA06Yq14TV2xAhSRDIG9Ciili3XvlqKDmOGj8XnlxDy
2AGD2owg46v0AcMrmlpJ/MSgFPkK60AqhZIdO+XGb/heVuEZ1DbcnVd2zgV6Irns
W0gJH0U+Xg7ph48qgMk4G2ZC367V55bN9nopfX/BqoOTxbILYOpUNlMDf1q7NaC4
6vz+0JN+tRtyZmwSx9QJzJCo4vmxlXTVmlUyDFjbI3PTDHuGVG2V0x8aQ4mPwEAp
Szf4hfFUDqkDjbehVTMH9FOuXk7ajCAAmtT87OPCkX806Z5fK196c9EPcD4elcjw
S5E9wE4wj2IKtzkImL2mvE8UyVVcjzRBHdn3DXj3xsP/7djrpUxwS3Hs+3rVi9xG
Oy6uR8lJyZKCnQ55nasYB85QngCL9BTb6cPd9fkON2zA6iWwAP95IiJbZvyixiuk
K5LIX55DllcDxv3Y37Rcj0o+na3QpivFVr0JO7f7WzRAq0jMNIa7daG+GCupZRUt
H++EZy3x5NVL1+oHzUPfiagmQY/iCoQPgy6O+8b/j+Gm8ziPVKVORMZ9FBtwYDPz
KgqOv9elpSGXJUF3YsOTUC980XHEtec9XD5KZo8CZf4cibItvuJyF0veeOmHpA+s
79ZknlSs03P+AlkAui9LpPCkOSvS6fMlEIfeN4Vt0zvsLFgUpmxuKHPqjwgi5ryD
xWsD+U0sCS/tJ5BWW+VQn7bVzga7nJYLt9Lxpg2MsbkxGTG9MRRLnuQpu0NNGYzj
OjCw5PLwnT1plie+P84/5uJLrsScfjwsOnQ1Ei75J/xphrOSs0BqVon7+D/ryf6E
uBcye5gmUwEmpBIy2acUSbIWpsZTYzREy5D6KmGnuwtpF50QUzW3VEKb/dtcU2PU
7t7KDQ09fkyeQNk5Zgwte1RL8lXKsFflawYx0yk/4yAWsX/E9aeUr+Lt82l/B3X9
sKbf7fYAxzCdlbBcnsDqBpgp/DI4Uy4XVQwA/XVLNeQYgzxWs17TGe0pzq15tBsl
DLL6up+KbuadDghiOsXv5ynzmdZrWNN2CKXHTdRNXaidSjEh+NhUPtRnMzAXX2wR
iLrdW7QvXaa17rihTMFKgaj4D4CEZX4+4k78jILGmJmF9M2hA7WLKoeyEEXdW5Fx
OS9rLI2RvcoNkrxVq6pBekviSGbDluzb5qclpWzasy/IHomN/H+bWZ5eBoJu8fQZ
N7BbM6mEVvUyUQm2JFu/fHArpm/+mdrcpIKHX6t4Ch7yy4lBD2dS15WqhMb7N/Wr
mwVuxnlGSckemuJQCyppBABnbVfLe5sbBxAFnx8yXOpeFqSg9kV1NIeOETFSPUhR
2oEBbeya+ror1jZW9JG2KavNaMFoTlAuOKPcXcaJMYwC+37Ic8S+jJykCtrqdNY0
XzNHZb5/jFEOngx/K1Ofv2HkniohzyPXKutHKEXgYaBSl4dZILoSL0oSP0VGeqfg
N3B7gn6qWojoiRdA0ur3ZEROz1W+EYN0C/Gn6ZBdhTYS24voMrD9bi7FdAKGTm6L
zQpgz3vXIZ96t92at0TFwc9gwbt17SpckVlqP1ND9hgMjn/uM+W7JJsg/sWSVvEX
n+YuBqgw+srwBFjitrK2ne2yToDrNG/0Dv1RSyBhLqc7+Op/MtUoooPzM/DNBiGG
iNUJWy3C5PXTheiJlC3STS43vjWmmhnG+VCw5//RvEBUmXj9tNEKBq9zJWi6uk/x
ovNoZiwW5hE4b1mhNPU73Jdqp55ch1cPEQLDXecJZU2nngYRHYV25UtWZUa4Kkij
2deLgWiQ49ps7GAVaRQHq22fENTImXFdmdK8IFsOT5b0r+0F2XtS3bGgLvpLQPRm
qG4fckZHMskdz45Hvcl+GkiAD//nMqHj1ek+x7g2bwDf1QOAMY28GKAwdlIMk/AW
WXbV5nWozP2TTJZW7HLZNdIaZ+yILPBXTuXIAukAFwBFpQ6+aaMLyx1K7vmq6tbD
Rq4Gcir4pTjFwZyIDz1TcZfN/8oGaGNRRKiM6SOfx/YveYqsNtAUnVzTRn+qSwn6
ZlTZrvtVXcPuTrrhC+zBxVnEkHOHN2SxfAn9cq8/ZaZpimYyYOPRm08tuNs33H6/
nl0YLqB12FjbgwtrTHZzECF9H3fFWIUwBc2ue6TQ6z+vpXLA3t6COFY11B+r1y1L
acbSmuUSqiEH46K0A+TciAt4Yx+M06WCkb6UqF+8+py5crv8mtUR0UFncL7RjiLJ
6wWYFqlaPgMrWL6jRe2+iYIvJVNvP7OmNvw/OzhGRYx2Oju4YOKNKuGnMrOSVWXH
AHizt5xaxB6uBFNx0BN4yMMLmAJ1s8yPrNwgHsGewrmJujcdtcnXbSLOb6JJm5qi
2ML5uIePYO3/WSFXyGlOQ1OeLRLLhY6cFa8r9C2xPB0LqxcXO2ir8SZAYoGLxezn
COnhcbfP3uzkMEs5HcyM6AeNXL4z407hPIWItTi+LDexr07+ohOSQUxjJGXa0xno
y7tTPO2AaP4qw6/0Jw7NAZe4p+wXmiroyP46BJkdyXPA3rihXca7m3+y8d8gTNSW
59rnrnN9YRvKciVK9N5DRN6iLo9oEKDe+1LI1aAOtkTRBkyjY5z+vs/QD5S6BUo+
VBjmSiUakwWwHi9epveblbkRRll44QjprDkyt73rf98+ssJgRJsVbmg7/mDT4cFa
t+XlOnpZ6bsSGKME2yuAOw45J8gHKmQlEGmeNYmD1NZtutBoXvpxDXlhBU6IoXI4
dtJ5CMR0eDpG1XlLLNO9qvnTY7Bq0Z9I5B4MuKnHxoP8nt+OkK0y9qYavd/HM5J6
Yc1/+4I9FeLFv27KxBqfD4botho6YwVZd5xD1ltpI38ADqBQt6axwelwugoEwfn6
27dGE6JyMBHYxzVy+gYnD2I8fn51J9biSaoLm3fidZ4NYgQulmboRLxrQRZmzL98
ppLsQAkpEb34SzQ7FJ1TGvFLhTbRTL648YC3rftTEU2GaAg/ECnxGxUnnw7rGy3o
vrw1T4gfI8ZVGCm4rEHNjYqrt8fQhrJHahIrVuIojtkoOjOLLSGx1wlL09LHFVeY
gKAFHEBVoW9h/jBiw5MT+4ng8E9v+RKyyXnHKSQ+cwKgf6UUfzS+JW9I68Er4J7p
0UNbL3f/oU4TPfX3s6Gu07gTD/uqCws7pGNFDXWSKd7hiYDxXNxOOCH36nsY7tUS
E9p2ECiQbmr+gOkcaQl4AAPBWAzt2DgJHMaunHBrbPvJEefx2sa/DGyC+G+tyEcX
tsXuYG6iEtegFpJHjYNrb0zxktu8/O/4S9t+u8E76yYHWfpt1V/8PxIQH/GBfLCO
skCl3uk/amYL9Q5tw9a1D9RnwaTkiDV8Dk8S5l3jjybMUsYCtoqP22ZETwmo3e8l
FD/4P5to57iCO1F1N6mAMo2IWJ23seIYOyG0k+ZbkKM0IimaZOKLIncCUh4cngWb
7PZyCEGiVZnKxoqo6It1x42bLavAPdyq3/+z2ST3j3cSsBzp86eiNDMurSoVzqZ0
Yq3qcSemrXDgeB8QucY+ZX6V3PPTOKAzAmIok9Lc0z6/iDffEaMzmfmqkEC9aSwd
1LdZ6RrZSLeyM7J+eERehe1/HHPE70msqNFnbs8wDxXF0Xtt6X7vdGGLAJ4fMamg
kdal8MCoQ6c7M7shOy5PNYA5h3Jefv/eq5xtWsA/Cbx/uaH1txahXC+t/2O0XCeK
SlNS2TwbLVdaZs2JegSxqM+7EqchJluGMrOvzSTacMrNHkJnuoVCzwEQ9QFf8/3D
UjoduQbQdNF00KQ7yuWTiSw8J6E/9xh9G3Wlvj/69+71gzmVxckzgP4pAK+xrdjV
GR67wcTo3FtAkEjb0gD9SunC/02KRZu77fbA1+cHIg80Dvl45S9PbCY9dQGc5dIL
51NUeAUAO+0gXnOz6S7WkxKb9KUWwspUhdBGeqLauemNkQ6oXiNLDjosEutEFRXW
NKJuNVWtFKEYiUuYlCHSaXV3O5hEdY8ttG4qt4Zn9gSR3pKlzKhdhkMbCOcRqz8S
Sxs6u0Yr5BY58qV8q4jwBfS3mmwPGbPgQyhun+BI2a4mUYsi4DDs0oK8+36Li9UK
jNJp4946LgTqjIRPk/qr1si4OOF67Q3h9moK9NDK8eehYRYWjgqwm7VprqNdeD56
6RmZMUw9hro5raFLv7cOpEbHgc0cBexALStidFh9OmU9tBqM9uMpAwpgfCKCI/3R
KFue2f3vZkd536jUqxKcwS2G27l4KmN9FOcEmxv9XGHJlgU+cUgyyx9W0GVurXM7
EQ0OqcLx0mc7WHGw4xUxDS33l2eqvXwZCYA5LQJpyYXftwzl1ktAwExI8QzJAedX
V2q4CbNjaqYxEhiPkFzYFkVLXFE0J4WRNpulY6qrm2TmGudjabVvUgH6cpglNrWp
+io9htPi4LvEIFmPtsqdijLMABQ9RgWXV2+DDWzo0XIbREJxRd6KvkmDtbKBdel0
/U+kd3QpynbiA2oFtmuumb1BaBCxo5TafTGte58VEDbgjaq2CRzhcAJAjybwD97f
36oQR+GdgykapKtmf91B6P1M2YTJPVrhXF8/lA6xAldt4U0tUaCVcR1TpA4QpfPn
GdgpmCqiwWcdTlXxOWi4peFf2DbUgWBYW44MOeoHmzljrDCyBpgTXBD1NGBTUzVm
3q1w/cvU1j8q49hK/21HCr3HaCl+Ex74sl3cHGPAFwgeB+9UiWdFVS2WiU6B/3P2
xlxqU6lfA2UtGISX8yBFFMz5Sp22pdZ8yY53U7YO6MWETDSBPCtVUb5Wr11Eog+Q
RBVaQC91Us2d3A5njZtzALLJ3IjLGFbAEMgXe3/TTKl4GG2voRAexZma6GcNsQEp
ynX739GAIIebSH68SevL6po0vBCrwu1YPtGXQB3X+T6Xbkp7cB/p/aGzj0q0qEVE
FkEg36DtF46dcznphRo+SBSYUOcrmlwNsS2a3Qf3R/4zsfdmibVVFnM6aB/bSSJH
2kI5rxQhZECvwRX9cYfTJGlTOr1xAhKoFU7dkj5t9r4X5iZjphaoy9icurID35ej
fhxvrQ2nFOI/4LTtqif8rOUpBV1xPRm3j7CBy60UlViuAb1jC24OtWM9KN9oRbA/
IFS422IQLqsOpl9yhSDHDIQjEQ22VAYKj8DjFwo9EryyudPTosvIFP82GVt8YkXa
oUHul5NI94pBpyghX/zhC74uK/208ytrz8/qSygOYqsiFVj9pxRnmlEY2JITf5av
NsO5HWawR/ju4dJMbbiASZ4KjKbK9Z7aEdbd2eCWGtO7HYYxJkNGVjVDuolOodHM
6TZhsXA1BBDJSpW5vvQkkBK0GjaDhri19YO/VMTz9xeWper8Ddyysk3A5MBuirTB
nMdFZzz0iFxN+TNBlhYlMpc4PL/YfBF2rImzWIbXNbjVgK/+lSGhblqBKnuqL2RG
uLr3ywch9jFxFMkGGan0xY08ChfOObDNIHM/RAGCVhO7rm97inESl36RsHYLdLGu
m+VE+V5Wbs7RwzLIzh8fZKlpDVipj9BkDaNKotrWemiOX1iG1og8VSQrIKUHK0AN
HYyu3CVLd3QFJaxfzV89vtT3xo73Dymiwh3I2/ZxZ6XlskoFgLNaLnPQ+XCr/2A+
AMQvfyPD3jSNAHZz/YqW57IQWj9xI/JibHuvUXS11Lfe99GI51LZzD7fqzwHJZrg
LAwrUPDAlP2g60gLaDN3El3N0TlbXX3YC/zKXQD1He6KX+NCYdoAzoPQAWKkoQ0h
1u06W4ShRGaPnVV4MJ58E/sbCyYrUUy+dmDAMr5VspvXV19aC+OcqYl69JH+fdDw
ML8CoQchfKai9ZwayKzhiZw8slapU0lv0DgpN3HiawPR0XMqn4fFcKjAlzUUpEbB
xvIQ1VUcTrHvbnYBX5VHn2zQWczME54jQANeme5zRutRhTB9sfAmQgcBpr6hqYCK
7aEYyJc/l1q6o0hbsKwuvaOpenVDgZzXPa/RnVp3+08nDLswrwz4iefOiWfYLTj5
1yUeXiRbfRahMBwnhTyeFCt25xnQ3NJ4kItwDFiXZGQRTgMiMz92JOOinKYforvZ
s4zlUimoz/CHms95RHjKmFX7ff5yrhOYDM6fTefwAVLVXQZZD/jNUXhLAB4OorCh
/RvR1dsgOXtZw/vhKjilY6qaUKrPBwXGsgjpk20kxTJQYY2SwWPwQzSDhuEE0pux
LQ0HCbXZRSp2NAroP0RkyKIOe+Z5V9lSoFPdh2aLMjMp/ADPhSJeA92TQEL7Hg6K
KMUgJQ5+iRGB5Z1veRM6IHG123+SNhJvGcpChnSZTxK5G3p9odf34S/2RU+YvAZV
khUx17bb1R1x1C6Lo7FsbCPTUEu7D8SfGcJup7chcr4GRtsdSXfuBxLANiAkVwJL
tagnjlOfRAQtWWFkFxrUlcuwDGv0F0MiscbyzMOSTD7XX0k4dEnqB24IpKYG27iV
4qGQ12VpMrRXemfOsPBk8OF+WN314MzydHZ41XHnh/WhW5On2gbJoADs/j9lIA0P
zCtWeYgaHct6RN/5jD+aZcynlZhBHM91P0p2KbDo+jjwKU30ejFNlbrf4Sl1iwIk
sC8EmGl9HivrHMQwbfyj3quOpeQC6RuPA0QmyWKaZ/9psU6VQqNl+aFSVHQ+eT1D
G3Nil/xQZV32od53AklQuKVh1+J/5qc42ku53HO+VtfDdlOUP+szaXmX4fQQvRSN
YMuQ6ROs1erTrL5tcuMLtNJmEBfnpm+qGZ3orRH1xMzfWCESOqRMUdk9SHSa7vhK
sGwEJtohN+l6AJoTazVFx2f170QAb+UGzpUhU5c7DyxLgIJORIR/XnYfmmXtV6I5
A1bpMh1B+gwPKrf7/SVoiyohlE6fy1dhx/B3Uda0ml1TSMmiG89+HQwwYFKeKVOw
hf3DxCaZqcpv9q446AcyoR9a/fJW6IC0zMs1xiQNwmXI4si8QQ+BuiqoI6ex4+o0
ikfqU2QIX091pnUIO6Ya9T6u0+fNU3rHXd1Q9JbQw8bg2fDNZyDiDMm8QrYO0Y+J
VfplubAlDWjGm83JniGKdJjk/fpYA88rMxu3en5CP+hqLqfwvg6pNDJs1XmjKBx9
BqZpEqX+c4bVEo6l8fwapYEfUijujxTLniYRYMeRZ3eVwcAEnzJf4t1Val6Sdewc
FcP5+0UPBrfl+bOV5gBm0FmZAdcePLuToEaHMtD9DhXozDvP455f50cn3gLl+LPp
YB5phMSWO31/lCD6x6XUZ6SAGZgc5JkslIZeQ6D+al1WWjeEpFMJu4IQE00qbzlh
ngTtEOMbrwDymfC2cuzm6zMF3OyM3h5IoDvfgg2nMdGOFrShz3RqOKo76jWbHCHs
KylbQc5mUOegLAzsKhQ9LABgowCgDnXorKOiOSxe4wYhCFMG7Svo2TvxXHdtJj0m
6dB1mgnD2goNPNg1R4mpa9gmRuiPDbS8IZZhjIymY6nrwaCRIX75jzli0er1zuAB
LaM0Jzr+iNzZKXpIV0WzxiqsneGKqPGTNAvYZSIlSlRFfAifuwTKuiNaHGViJcje
3AZsdRusiP0GyPIh64onSXQjdUhVm8pFK1qD6zkHRY7ajZd9TlsjKrI4l92ux1+J
KzgXt4L9Ig4733lTHpRpx68XG1fJAF2F82FEOZ1lwKtWAbEv6FnM9J3iNZiumAS+
7roUGKUCT1+LH15n+9XTEp/VqjfMQv8TjnkP66eIUnag3MjyHJXTP2km4An5Kw88
3YVeLNvxAHWNSw0tbfX/GZRY+j8+XbQNhALax97queuCg3zd9Tt5YgHXpM4sya7Y
OS8Lfehp6jG2VzEvm3ZYQFnUH8I8JIqeLhLNw3nGdFXBLGxiX9gpZbH6tOqtfW4C
W+p1TzXvYYPchIQffrPrBPPvL5LnXTotwLEqELQox86D7NeU9IoliNZOA+LsBd1E
ttiiTbC3bMaBF/64UPK6rq4p4kyDpk0GzVJQAtSjX6+qvS2W5UoruxScpIEGweXP
J+BdZyrmxJgrH0CjcARS+5+yfqd1tE6NXmhno97p3JXreWXkd7FubVJgWRpcfdGI
knsD9TqjqIHdLwZ/L2YIqldsOPXqIIYeXE33JnRNUpb/Lhpq+XoiU9B3myNlN035
8CF7883ieTuARBtp3Em51hoFzCxRKEcx7Ua6UUJVMM/r60UPlWC/GCs/pq4NUm69
aYKurgV3ImQNmXl0vIiqPbN9wA1cSqUN3CDDtuWxVQ19p8Fh+X5fExaI7HcZRIpY
9orFc3DSfW0vVu8a2Bp9/xAz3YGr1KZRY8soXTmCNDPNNr0sSdl17xsqQE0SuTFY
X1UM5rVvOGkBpvtw4Z/o1CvRLrqAt+NhhG1/W4jMuyF5yJH5WcdXyzczebMjzpFv
U5FL+6IxhJAYP4uJlp+deF7YgnRZu7YeBRFQjX1N8KDjt3DeEpsPCr9xjmlA7j8P
vUmfw6VkRY8EYdxExJVbykITSUFJRvK8mk4UR6mf9tIoQGzK5EVYTZQDhkxGi9Gj
TSbL7UhAaHx4LcxWdIKraDeu4dfX0nSTCtq7anRdr2or/4pOGEdLEh68Iz3JroeC
ZKB0685LnFyl162VzlqUT/pQLycFU3AVmoxwSBAj4+EedPNS4z0LxEFQkkC0+ts6
UGj96qO0TFXSXtk9tqciTXwtSFgWzOd99qhWIckV5scw3i3NBL1WJnmSWqR3irdH
RPkDShMpu6vEufYeLFMncV5UGKHn+foOYZ2RBaUOZO3pxZMrC5KMzSo/7LqXtCSK
et4bMypXXI+ay1UFOwPnHO9HEm1w+UxS//SNpd2NCWShsZUanqW6M3XPYTjl6YET
W1x20P8CivCtxUyU63esXVV0oajWVDRIfv1MUCbC3iAhEmm11OMpyLo44Q1zK/sK
197DyaDm8meTeaF8TRCfUgQNg/3VnDkfGypojjcB4AHaxaZowJu5XNn7gIMb8zmi
zk++nzgXi1xWxOnx22wc2GhcHr6rkr9fdp6d4OQ5eqDSS/ITMUmbm80xxYCRRSMk
zW4zXJxos5wPTMbXeLt29aOn+lhODmk80GhS5wOPT+k5WifGKiZ711uAuZms1eeZ
X+XDaQsV7pZ+YcqnIfReCg0lnmgApaalVw9GF/Y4FDVF5YalWlwBn7RxLEahkEbM
nmL4DaBcEh2sFvLGMr9ShqNEbcGgrnnYOm+Hs0HKpGsTn9dJrxuGiLrZVlBXmqpF
8wBMJyXIptt2PorhcKERF2iFasE9eiKkAsfpgzY/Ro4Eup/lI1SsXPCDvH12PwZZ
kXCt4sRlOMhvPpYTpr962WxU1T3Go5y4REbPvhboRilvcSgjejM2z55M31S65iEw
SqUQsCq5sqLmZZj+7hJow3i+trG7UV3nXPuPlAn/qCcAV1WS3Zg67ajvEmV6qyIE
Wlf67IHQzuDmGb408Z6skOV7tuYfr9GOG1tFP0NEs9wLRHFApV9pM2xZc+Xjk79T
N3BHaTg8q2UTtCjiyjsTpt1H4YYfFaqXQtN3c/E3ue+Hr6uw3viCia58cGwDvH4D
dFg+BGN2B8hHDe7B0f/tSnZLK8zBUmtDrDX5zVvRaWoY+Qr6I6FYh83y4kk4hals
Tx94yyjnzBKWsWSQqJuAW8jWPzAoXjbYbjqdwocv7pt9pED57Ow27t344x1wM5Dy
rYNr+KLsUxFU2nPvhZ+6y2WqalzYL+5I2mndTOZ4tIQ2xKYkJb75xmP5eH1EzjGd
dhjweC2YcXDT888SDKIgX9levndLOcnlbpJ4LgIHffrcDiYZmH1mXlQXA0dWSs6j
sqaeu5zBQDBxQa6CbZVxyTVQEuXGsnZOgb1RPvsHNNO8K1M69mX5Kt1ouUqCcuyt
/Z23SQ1luy+L9qwCZpT2ORU5YR/wiR1M5Oj1TcGWHMM4vG+ednvlXm0kWVxqLgRe
uS/zpVz8bRQCWuFKXOI0g6FenM7Rsfos1Oc0OnJE5S//CleVILVgQhq2iY7Odrlc
9/SwRlIhu+aXYSlwwNt0rFbxmF4XvA2rgPMghlPbsDMB64SSr8Wh1vmyLBGP6rk9
4eQ61PCx1vBsxrxaZBowbbzHiRrDWBkeuPJDeSWdsDbsPQmogc+RTbDKpk6jYO62
RuERA8GBRkijHewRGYVJmV84cGplfpOOWRtNmgzrp2DmLDt/DDmJpcyh3eptwVg0
2IMM6ymRdStV7rFRr56nAbLOEN93SE3lP9Kc/gp2YOv5SdlGzo+cc8b9QZp2Rf6C
kOGlrRVx3FbDYtpx1UYJdT3TYErjOCvluiy6Fuk+dYpDnxlOP+Xw5mnmc0AyztI0
jL6WovjeJ/PkMo58aJe8Q80XRo40wd2yoZMjMVN8JF1+vC7C8aDtLzxoW/XKr28n
7WcaaFF/dS9HIjIrb9eC2m0+ZQWStLdcZD8u3Z8GnMNjBP8OTZWR4lfyPQMNiGvF
catKs/s1gKy7Ug8Hza9K0lNpEAUrkNagtP84lsAeYX0RvSink6TFIsV0P5ixLGa5
fj0FlEmkH0fOxpdgGkmxWfVxKicEO07YN0dOSBQ/guNsWDzWrHtw+AuKj3hYhTAo
VL/jD/HTfrejaGV9WMU8I8+EO+0JCELFDu+aA9Mx8axVnq4nRYhw1AN+A7KFa8ya
MeVOlkwrZpa/bAP7ClPTWHrxNPyNL+khjTrqWuxlL+pwZQAEQy5a153g+c3cjmif
lXcHVw/+d1IFxp6/qt57+JYs3z/DRWqqfxyri21+LhRIpu2U9XPSEfbcGNePXKyF
6g1FrNV2q924HNAz08t9Lc7dgklo6Ku4BZ67SSmFvrJLU+iujqgTEJ7vyJTmVKb6
GsCbOiCDFZ8RlOxTMGsHDhDxpH9L2/Zbjcq3FlX3SdQChgdWM+2YsLVdqEQmWuzQ
9PlBk/3QoNVhx3aMDj2scY30HVEV8b8KmXPV3KIxFSf08m7JLsCj2xL2RuQZO2xT
1BAvkXo+Oi11nyJmkJjv9lbAixlctBaP0AIei1dVmLs2vBYCbPIAgHg0jZCRxm1A
CiIPmcrASl5QGV3bGHqcHOYFWYaxpyT2ZTKTPDcLolnpEKOU4el84QgdHUlvZxEi
huSVU9v7AUzG6y8ZGSXZIhl55Xzd7JX0ptYQIkaBh+Hjd4ze507Q7fds4sx/8mIn
YNlbzhQXDVQPu5rK/5DkNdNnWT5YeonW05a0KCn0gtGonu0QbqK9ac4B4zS78S5d
ghlTYURzuyjfqZ6coMKSgvujVBL+QPm871RK9qAYnUj3y61xXSge+N4BaSSMeY84
0oP+LS83RRWIXxbCWIaiYsLv2TojaMy5jblWWThzTS+rzxSaLYUEXUm7JDCg8ouG
rN4mwb42+/4pxTIjIk/vOLZuNI5YPqm5qkM3kbNupBvTcaLGc7Dr3Fuhjh6gioNl
gUp3t139V6epsGGlO85+YpnUbSkKyqCtqzNqPPUhw1mZHTJyqPWEjASgvEPqPQrY
62G4fqAEAeUkwT0g16RaXgKthkcyqI+OptQmcRkMcXw6Qm+XtwrCRRkoBQ5CsJzv
EwjwA2zC2NlXYTteayGhBX2rxv74HHScqC3SoRDTpInLP5aFE/V3BPgDeYZDRk2y
Qa5uNkg7Iik3l1HMpX521SLv7lguR54d2FvoX8TaInUqQpTk1MGpD5y584k5SdIN
op44mdq4fZsbn9YUq8DL7kyZYAfmVAmHiXYYIvuw6eUtx9h1hk3Jx9I10evdmiNM
S3Q5HWvEaarXkND1pYM9VMv67TQ/EiA6FXhd54Q0F/RXHYwWIDj1ajEgpgE11CYn
bOwZSATdcQq9rstSR68ICvw6VmKyvzcZIPji1B3+w7TtDT/K7N1IIg2G53T3i3xB
FqM03gcmXMolpmxkRQITZid9sz08WaDXWqUZkjjZtdrsPURk3bnTBOB2DiElsnVv
hzUG2sIrhlUbrbAkqze3MbiMcB5zccYHJaELtram8ql1vtiiSJFD2mEWaJ7Qn7z4
oaFJE3mHqjABnahDOYB35abAN7XSTj5tFXgMN6CJVgGxOqKowSHlk9GeuJs1bV3f
UvhOy6xHn7XfCMM9KZ+auf8dPyz95SPDfYT1PQ+Lh4VKgf0vFYCaSNWR/4ifBSX5
hEdcZtTla1txGENph84ktTwltFe0cq4bl5S0mR+hwUWVJ4PQApTscvNrtEVaephU
FEF1mGbRYuka5ApOeuBNHaqqRu6d9/1FmpNgBIG72X0t+Tw5vwlJQ/XwkIVIzIXs
ogvKdZ2yw3wWOlZdWh+056kW447txJba/SnqiILNFsXTDSU0mGsUmmtBWrT6sodS
iQMGy8YdeMI84BcarM+/3/vUFR6Cc8o4YuiFopMUyRziG/GVskHizUXkgwBJrZXO
RhLZFHFcCSZznQ6qzLIZDeV0ZvLpJur3A9JirqTM/BN2/QZwonNHM9zrhdSSa8Gi
CwNRToJXeZGnpjmSIVMy0aUvOM5NH7P/EE1MKBZjRYXIdzaxRZP7vJ8a3TMQnxgM
ch+tupTc/7e9opt7AKfzm6TEVk76OQKqZ/ArXRe6KXJj3ac68B4hMOSCl5y/SZwr
xoDTVAMX/SfcUU0XIONO5W22zdGHx7hLtUiChK9n/ssgr7GuQ23ezvlfXhpuYxJF
8k+EyQVbUqcneqxSv1ao1NjMaEEA9lNJNiKqAv5yxOYzNv/LKHnGhc3vapsMiyK4
XiON6rbxE4vtNXWH25nqvcAnugvTWgQK9hxnD1IJnhn3S8j48Eb3IuPphDWSNvSx
ZLDQVLn1vVo6JF6y1X7+aNcw7zSZa1z3Q/6bRoWtANx920A+JlLH4uBMuXT7yZv6
rfg0UNuIrKVvxa1JAKgy6RzW6SC3bMZKZaARZFGukHZKyZ9t2yVtSDpXlDhcpVhp
0FuCrZs6JGklSuoopzxiQL5gsYX+xOtQiqekKe/rMr10aOWZZqWGoB7gFLunGR8w
czUW4h731ki4bmvHM26hTU0ux3awXn/FLhfad04+A+0b6ui8wHM+HQXtDfNe35Ss
j55omr/BcnthNz8QEGMO6n2B7pV+W2PXTpf+UmP7txcgYVnu0kmi+Gv+w7bngP7o
ifveTFLSmJtyteMeoCo/eHijySBM52mOT0A1jUQgGMRhOS3WMUm08WDMn75jbW3f
CnbdizQzQ7WdacR5IhYZMd+Wwl37bOVq68Z9txpxSzKbE/1emTTCSitZl+N+Ypep
2pyNS5m9HgQNz9FSGpkyDSsaQXQewpoCgi4gTsauioyPq93MMtkEX1Trw0ynyKOs
86iJsEA4Ag6zf3WfBYrcgfmHcQCce6mcTzMtrHVB5Q8A8uJ4ogs/Nbm195qjHKxT
TDU56opnleq3WapaV0zpThV1ifXzFuP5pvgWp0d3nVqxbhj3czQLmNvFohhoVLys
cg1eI/ZABU0C1AZpWbpEGqGCuxT9vzNMhuGYaEAqoAuSnpH7UbvWc/QvFtf/8t42
TEIM0Wn0ijZE6jb52KMV1+dkYOiZjm5EcusdqbktDgJpV9vqo+GcdtP2YRKMdts7
5e+W8oDZXa5S2BDaPZKTq2l3KBqLe6eBJP+WVh+GA78T30phXzc/LWe/BaeF8V+B
3r5naRJyzab1C+enQzbV6G/+bkjhzL04RWAmuRBcp2pnhJziRZq/0IWMj6O1Okc/
HkRH8TTUWtePZ2ZSPwO5kuto0Zx1LlM/3ZM8QSSKbOMq14Qp8M85JDrOhQY0NNyp
8F7Xl4LmTse+0SzO5X2ndqwY2fmKJbES23m/3aEVuj4tH9PYq/bHkDEWpu6mKWLf
sLw9QjFNeyLsBOtqZLRLdmy8ujdP+2GF328WrTHmkOJ1bvUoAHmScoUT0WWhhFAP
cRa3m2OHDA7eweXWatTDRtDeppHseUW6gaxGC4vw+foq9gNJe5wGG6gtPuHQYdRH
CNchfaaIa6h5NPLsaENoAXg7DKzLbsEwPXkeIV05cRBVD1CdyONakTu0L4wUQvhd
bKxTjlen4ya1I3+zQoSXxlMcuFIcQwMOBJlxAOD6uJwPgZoVaO+VU9BF98OoBPW1
CiN3dGz3X+Pkz/Hl60JaVzwu/pZd0q7vqchyiwPu4Vq7gwIHIs+1iqJSYHonWZyq
dUGkK+iY9vd5H8GhXJWIolNilLxhjdNSPFYJEC95107Je6lXXZa9YB2ejhjsXukD
45mksWtko98wxPgOuNAd+euz8hnbQHGSKDj7Wct7FbRde32A2jixMf8gJa3hytav
ZyUjxpVKPUBW4KrcsRmctLxJHxO8PBCfLX9qBXo4ZIDkQpsUVRHx9UleHBHAVWKz
osRPBb73z1KX6OSIez59mXoUhch/JJ2kuB7QD0Z1gQu47QdM7UAJFs0TAkbS+Vkl
LQFvd7eqOit8lJj/JFiT8dGv5FpvrVs9X4ruPVl7b2Ccg1iNd9NuRWKOt/l0jHnr
UiDFOasA/gt5RCXXJOTG/4WkN4lq+UnkwGuqwK4E/nH8YzF/6GfIyClPKErH8mo7
e86MdN2uZDVHoOMQRq4mn9bXgEDgrakXSK5d1WyzwLafxLBTvanGSkLNC+5W356v
wPbVY3Y1FxH4fW8fNciRZhbXy2D94xLzW1w2ZDCcLaT3IuY6aZLUVYVN3NITx4xn
rR/BeGIpqAKpnmbfsZ3iD0pV+DKRmDzmLn0kDUuhZC02daLM6WK5gvETXg4mLoqb
4wunBfss9gPfN43qVFxSomOzRRpXjsABd5KQ40E0FEIZgUQVWm/78609kj+gYF5L
d9OfAfu3PiSrPZvR5nDH47kRlc7WKRDQuK6uZTSmN2ROC44+YdmaD0BEkzJBygvM
jSDzpclHJvW86Bn86nzVG85O3tIX+EqsFxC/jG3q5TmVxqJuEfH9qBKYc+qyQH9n
C5z2A4woMgV6MZfw2zdeiF7ZQ2jNpTCQkktYDPqANxw8mVBdw6j2Tte4LfqlTrXW
fl8QJ8GQImXcXRKub+nN2tF1Rf2s1SuQ6XvKmiePdQuShpxBcEEhDp7v5dkp7TiB
tJKWxkN2wcT0LJjExHTZ4q+ovIp0PG6BU4qjUvkmPGpmvWBuOHwDpHBEGWD4f7B4
TSIUQFd7GUmU6A+bab9myXudhASFjLKhEv5uYIDUJOgnaKprrkNRaookrJ+6IhoM
oT8TnERsPxrqo12YX2N6Usddy1Aj/7HyMJrcer3jbwG1MWSmTzwMd6reLbl4DNm2
iJ3s6tNqPuFGtoQzVU1TNE8FFDGPJDufhrhJejmAyFAV1EEpKIbsx7LiJ7++M9PH
qNA8ZCW5h2uRqOwat4w5roW7WAmI//u79or3zJtMc5BsJZOV0Sqd0QmiRSaHwWY3
g5/dYzoA+9NDk58wfIiuHymVYRp0OjQRzzHzMkTEbA6Y0QRofLMLuuRP1X1Cs7qO
81Da3QlFHxdY1+pb9LtcMRgmJjk/zlEe1MBzq3acvJXuYCCfjWYjRf9D5XNxztjQ
3MkNMvQ3Gftj0Lj24EFnO7K4p+fmQiKgD0m9FsTB6tuHafnLoYWnC8xRD0UNMhmS
jR94TVTL7uvQLo8LD405oC4spGl5gFG+sJIsFvX/LAflw2rR+ujDoHleFBHZE3jk
93n3IXNV40opmMpOXNL6MWMygStjAQnosYP1DO0g0mOYeiatfRNoqzzC6rSgPcD3
5m7JYXK5tRcOtizPfAII2a3rnZ950xbdyLwj/X/OXGDPXmnPBRe0Bv6xJwNAi7SB
yPaitcwKngUkY/lPnXA8PI7QxPkJfs0n4YNz7NEbOq9U4hDGJkJ5ZuqxPtuvWIqX
MTbOOjG3rUBK0T1Nfq2wchucIDJmCZDrrbXORHnW+3xiYOiBB1fCDhWFXlCKN/jn
m27Z/M1nCgwocsSPEfJHGfREQB9AI50BUmZUIIdIuPtybJdDAIekuJjG7QTW3Jnt
+EEYqtmJ37BDEPrR+vtKwrB/L98FxW15tHn76tJmCV+gifwb1MeW0HTZF/lPXBBA
yvUjuSam7dMJXGAuKtmQxBNkDtH1Ez4eY6gMQ2+4z2WGKsB9b6amml2HNo95d7rK
8JGPoPe/FgkaRBGYfm1bdpP5PehAMjelPlIoIDfNJVe5rQRvzZ0317FVnepuvQ3i
7+JewhL7s5FleHqKC7dMF+LSUdRaPwcI3Q0dOs9poZWPZB/6dPiNb0DEZhRm4Bk2
bOH6D+CchtD5ctmCiEPUFcbyn3fEDh6kQ6RF1gMY/thJUJ2CX17d1mhkDswmvwvO
/6qHFTB+tLrtTtqT6mQCQN4Np4+fyy9+ADHnGOyalMAfzUcpQ0vO41cuqf7lzgym
P145dHU9HsWSQG87vX28HU676Z4lnHPwFvbj7LBggJ5TIrSEhk1aa7M2p55DXsmW
TeKIfaPsutGAh2O0fFHX41jmRA3ylKn55GoBFcWUW+MNd2KERtgGNBK9jcKz9oNW
Mxw1HtNcj4Y0ZIWHwpDx1sOw2UxCtI1ai/xK0Bdi2beytBaILrvgS6S14glykWIF
e9mP2xraxhFj+iUAosbBtmHT6Blfr5kdsdR7K5MIhu8Qe0i9KFi+GOMyLc72bXmr
m8eoKZJllLTpGUedRnD2BOXIAIUOruFK7E4x2JlywPr4ujzMBom+Fqj2wvFhavkz
Ut7rGUE4HrtryPNFUgKzQDSEocTSlTE0RAVspZU8HeGCAhz3CyYfgndPHAX9QVnJ
I0nVJjVip2cnou1uhsgwaU0fyj3AUCLza3zR6GL5qC4ET6of5kwWxCzb6JCalP0o
FWHzuRyhvgkaV/ybl3bonGq6YDEfkz4/zsWryIF4LY8RNPS5wx+k28x8sOrQ1oB9
IYVge6BPakfmCk9raMDfK+AuvqwZ20BwMlaKsu9AeyG1VzogyVJoOC+7z3F5vDui
7dibECaGwCyx49orZjd0ji+gm+KqTuhwXz2v7B7jCu0RkbTrZywmpfvOEGuhE61g
HuMM5Le28p01+YAg1A3vJHGXMlSD62ZzHm4cJhDxzqHFYQgdBMpq4yB2+IMwKRLy
nQ6OuPl79nWIP+w99JI2PVm2LTSqxSM0pIXQiOxhMIgA8rDnEYrw6t8m0DPu05Q0
O7VVFyOblck+P5qS86beRYr9nH2aOJNstGBybmQB0X4qTAIDEkGzFEFYqPxE3715
A2oXJc2Ln0tNeQCfHieEmnzfikd5EZ7ec/acsWWV2ot5GZldNaEQig5v+ZE3FKY2
ELx4Ul7QDUClO3aT8asQ21+Yq4ngW3qy1WJqUonoEocyPJ1b9YeCesQA9Srte5Jm
0oTZUiBXFb5eQDkjBYtj1qHD9T7g621A+eCEEMYVhl9wzssVQrSJ11hvx4xTCdG2
4YYLVS43CjFsm3yoN/vhO4RHT3QKbFhKZBbcQzDRFzGsJhdflD4fqyn6nIuJgUh4
DXOBUQ2s8YpxRkt6CjQdJ5I/1JXj9wvpxdAVgpaLqb1OIkQnOKHERsn4w3OBA7sr
UffIMJqIyAJf4ozY/NeNIfijvS1/za/Lm/LytrEXRqxvHwV8zQaOVBbr2AdlErc7
yDDIWam7UcIJ7QqTqF8dosf/df8aCEM2UacJxMlNurxCtLYEPo6QYO8VksyfjGDy
s4jLss7zHBnbXbLtg6y16DXsd3rCzKmlneQ07QRy4K3QRxwezdUzRYD/LzwoMz6T
pHLdNY/vIG3xdLzgwJ3y5cNXraAQE03XWRdzXdCloeUzBTkvriEr7m0iZZMMxdMC
IvaqpD7HLt5fTBSOw/RSvLzClWb1egRz/o+V3xGlu4dEAfROU8YFRWwcZhGIbONE
8elWDtnLXTpci7Wp0HZqgV+Pop+g6lzunfmNF/ClU8ugjXRrObJ7FhECV7xys7l4
qmfVKw/iN2H2dQFYYOB38MqVC3FluVzA/zWQEw+gJCK1zfD43AkWEEOQJDb8/RwW
im6QZzA7xgbVfENzNGeyIR1kos2Wg7XE0Rr41iN1X6eagdAs6EDZREeoGTQPiGeX
YLdOGOV8BTixmAf4n65ciWrKwkNZJK/IcXNlY8S0w3dJsdxcHQ6p7OGElifzC+1j
Zx3gv5P4LIQsH65PvnJncCl+qQZKh8NE1R3tNsMcWsi0vqpmOglSW/G5pdUmhv1u
uS2Z+JCltZEenz/BWq3A3rEqr9smNOciX/PZGb6WJgG1Oawua7TwpQVkEH/Z71pQ
jq5syfQteBcAtsWoqtJhqmoSOuDS/JggZM/UjCWpjtEY60J1ZpRllvyhue1yiElE
SmXaMR83u92lmOoOM2LqeuJruomR89OPdhZ0e2xQR3uEOsdEjifqUOZvOLrlKGEE
jBRlBnyRVmQUt/spdI/gKfSI3b/Lurp2/23EhwEInCOSC+O0OF3m3SL2/X2IQjPN
bErTwDwlE2lRI2oFrrn3W7IyOb6T5XoOPqxZfnYlUzaDknvLayW19s1iI9UqWYCC
3UurUNdlvvs5roAC04lhdqDw+6H+wWOo4e6noO95x7n3OB+//Pm7uvCymFtuSfXq
s30S9v/+E9IZJ+/ApEIsJRZfcUzASW2hC26dDi1SMq7poST1fG9bc3ARFNJtWoll
BMOo3RnBRUWdvQIdnIxd9bGzJPLM4E5QHVeWnAX9ytsERhkoInLEH242SmKdpzSw
78fRjVkjW1jv9j865KxKPBQyjjzzvDzTxWmKVhdP/AxyCvo25F0WWMQuOo4d2uxH
cgRgQppFm72Hqw0h1oZc7nHdgkqxgxqNe6Q+3GUQKpmTWUu09waG7OMqB9h7owib
4sggL0b4T2OIaIbQZENBAefHSTChDdWsER22p3oKHGIrVc70hVVP9tG5yz28ZhNu
J4nXB9bxbY8nzwNoKRQevpSup5wiyKs559VGiOmSWPDe3AeiJy3S80Q4VD/w4pkp
LFDti0U3FKPQ4uQRL+LRCdJ0qshdREfeVL89V/CnQAaDknTSbPSa4to86Mqxa7IX
pP1LoeSIBpPCRI7hcwsXLn9ERx7QWk4gExEwsM3RclDciq3Liq/LrkTlP648Fcvk
riFrtYafC/3ZrrdMNIdZtdMNGJanM/q6Jqg2MMKoVfk3OvVADneUMCI0tSZVSghr
1MvVYu6R9OmpmGBgqBWIfCZhsR7Q/nbBFhVE2BVpI04XA73NzRGyALTCRECxcC3K
nW2I8WUbf152XZ7Cx0xpS/uT1o5/AyXhAye20e1QtZMijB+oIM9eVG6bC35jILVu
aBhS8Vu9ajgYzob8+GKGjPva+lnK8f9F43rfaAFukC11c17aaWiCbNPSTFUWdABX
S/tLPS8ewiK4uHzyxxivHp6oRmczEDkw0OwtxNmjbJs5Nim8ewxmuW3so30AeTHH
ZZeK+kT0bE6SIkOtqu9v0IFUPIwlp6BxQPfZZf5ETQTRkRzv7hzB6c2oJkb3twMF
f++pij1rsRAwHh3qsma3eZ5LYhqbYqbn0wvaCoOv02JEB59pbbDFSLM7GmDy/ibo
NxWA1LlL6JKQHvNLyodITIyg+IhjtvpbSqebQq+9ifj3SpijeqCupqGO25lGOFqS
ECd9AEIwYnh4F2+i8wAwMVSV9Xvi7RYYedKdNlAo8U6HS3d5LGNoAd0Y3UKFVLlp
uX+pQJTEaN9LAc05GrzGl4ujNyJZtEMHKHoFUFfT9bKAgoxKGGnc3CW01gthCW3A
PMLvaIzLOCwg9su479M5ZWBFaqIMISsrEiLPznOfA23Sn4Dw0mX5SNKGkw1mRWG4
BBtBBj6fNI8mpzmcgreHC6smJFxm1Y1HIHWQChBz+iIxs5ZVK53y4/KvQSVNlTN8
0eHDX6QWJIWwqNpqSFZXP6zDYmV+gHmJWAb5RLc4LaWiomFyo9hAXgnm/Vbw8RBt
5dtiBOJM1EHJzY6e6QeVwPimBfwZ7qxH1qB1tAK2YHOAyiYaoXJzENS6c5wwIykE
0hP0DRS+i8XI+MLX1/vGY8XB2+cH+UiMPIgF9i1npZodXzjWSoe5NDKwp/VfCHrz
aYoo5OzMcgPmd0C7fUzp5F30Fbe7LmuWZw/PgYg45QtSWcjYMD+DYGMb29X1V3gX
Yz5aiqQEouVQRbVgG1k7x6jB0Et+0ANVcsCIsgNzRsL0Mq/TbtAk240oSXoBql3f
HzYs6DsJfD/XKbChtNxz+gxpgH2VtezRacbqId3YVk/W/9iDn8M4tGpnrMljwuWd
GUoTqHgtiEpX4X/RIO88VJagmGy/M2kXZITDqpTxXROmdUW7cPJPQsX0fC3FwWGN
13eLzCsFHTTIVHIO+CsR5E4BZWfDiOLAfIFVXCpQD90LOyyTxueJAZelxfgsHxFw
CgBS8cO2PAOCzHaKc7as9LbBEv8XmhJlBAEgMR9un0moz7ONA5Eb7Pgm7NVwjuDc
X3/24SOGNqyw3Oyr23DXLWV/MIS4hJQx2vvLsFAlrHgWJd2wNrjvI+OZGq0bYBaX
cabvdZBA//yq8BDRaLTtgks1YyjTEyzT6v3SRELTpgr0UBpPRqwN6MpK8mFsTywW
d3OX9qiKk9nsjL5JftiljIv5/Zs+g9fcY/YptYvmQ6yAvlxyeR0R8ZowIP0BW/1c
kww0g4syZ46scDwTT24g/t6qloBCsUAOuR8J0kCgXdXuG6sxa3b7LYHS/nNFS8Qn
Kdg7ogPiFbQ92olWdkn55kKdhl2D4FSV/AT5PR7T8IIFPlNoB4Wzf29fxzPSetI0
2W0TIjza7FpLXSovgzjnjPTqlLFpF6Q/XoWH7CKOyW2nC/XArsVaq4E5BvS9SvlS
l21/uaU7GSpTWQsJjllz0hIwnLsXZohlvyiOOMFWOf0ewuxXXAjNBr/FHCCiSZMN
IfgqxAp3SOVxHAf0AP6O4oXG4xGhoPBTvcAExcXxUNDtQwrX/O2S5TaLlYBgL/RQ
PZrUf7VLThKCB34Pska/iNKx7a8R0mFnLAyrHizC66tF+dpvYhedQNxqIq3Fb6zY
Hn1cL9YC4Md6ESbH4Suuif8PUJDwwcfRWNDSN35b1tXrbNhnfPiUAZXuioeFG/0I
C9z9H54Raz1edUj8F45QqsrExb9zHYWsimi4cOT3ytouhIdE+3Ke+nOHRL1eFZ84
LwZzl9Y16S5rwIHXl41xZphvbKwMT2kpC/TQNDd0NYwcxHK4iHBeNkuI0M4EsbVQ
G4AGxzF87K0f3AterOyyu5Zosl8ddMlHaJbYBr3rUJrfMP0qZN4S8GwMXkLGFPTE
FPADRb+wpFmw+wnJH7VpFgDoF/EUnQRN/wkWp85bcfnHnoLE2fZ5CmupytXNiHpg
GQKiFsjhnDfBMoXpUljJtpmz/kkdRjOnKIpAYcs6Qt1a/7d3DKQZt3iOj+FrRv+H
1Jy0bb/L55NwT/McQn6MWRuyL2NmabqT5khiLVocsda2NN08smU+pCfr1eisNPWf
HYBFpt674+uZABcL8ioDenVfzX1DHKlpSw2YwmVVCWqKC92VHiXoiHl9iD25wy/C
kh4+3AyRJuEyYMVXScS+CUiaq+LXGdseRBE/jCBE1WJwPeu2J95MEHYm/UZLShrb
/QuEDnhURDYKYFf+3DWdYEtumq3dHjzapFcJvK/EAR5mVwaMikvLC2eIsluemOVT
3nRbMNprl4XmdtcuDh4uLjnQKpz6mMIXXoTwXhECotwt5yksR9ohrBoeY3K6Clf9
iqQC/HdCWoLDOxyfCJ53g2YmSUFjEVI9ABvfnal1/wmfUxSpJyAFXYqIAv7NQocH
jjOZU7IxTmaOJiCg3W6DEu1XZSqzMZlMY3Dejxpq4kPhFMpVnJmhnyI75/eT6RqE
xaT7vNLAZ8y5JCAF1Ih1FeCI0gXMmX8PAwycXkaQKgLywtz7uqbT1ZnsEhtwuITu
0ud3dNCQX/0ulqYf+ypOtnFXqVAnq6naGKtiCDYOG4z2sqhH1dKKf42pE8BxY5Pq
eEVJXl/EEvK2k0WnEGbfXL+QEjlaAW0pHoAG4WpYDTL5TRr/IkxXa16nwuo+unZa
yaEkQvDAORBfx+EXb+CQeLZwvITn8qb/H2Bxr0qAUAWrqjxjbg+9R750oohFfzaS
/vGJPhUPie7Ui8Y9pYfGKl3Q3rzNoytnJP4a9jdt9/3cmtTml5YIJsEQ6nRC6J7p
Xs5cJSjAPVudCC2FUrIfMZ+e7KsUAT9shTe/I833K0MvV4vNvPUoSdnXNIYCyYpl
bVx7dzu9L4Y39EjdXmF37b/Pz8AQpLWmn9F9YjQHMxbeZTPD/aQZZbZbDlei4ByW
LtKLGtwRJPcZkylttGi/1up6HArpkr+g78Qlg/rkdyw919k362mj5S044ao56mMc
r1v6OzD8pT4vbwUqIHDOYWpS5ndQWCyHa6CsHahn+jluB8yCcreWi9zXpkgaqz9q
5QEZQxg/5myThxJ0OcV66Yc2oTCwHymbM+YISRqGUp1O4UG2VVUm/yBO3s3LO20N
v9+tC+XKgSTks5nBDMJfaOL19HUe+UJz/oF7z8gu6pOecstEapWg7FW/PYFkytxh
Yt258f83bYfVHVX2Dxt8OYn17afAYgWZVBnb3LiMdZCsqbl9Roh2JFmCuuiV+uIl
453zO8XsxjlSc6xUsu335Rk8ls8N2CYDOsdtq/TBiSwDRxrDABLUudWEG7OCQzna
7b+D7W4lmp9xfwbuz19sXOITC2nB427xyd2zLsXnlH34Kd6aeI4dFdsxXNw3rUHU
NMlvL64nrj4PPm6hYEnCT7fnCYhZSrGc95fPsZMkUuwtxJ3+Ez+B0WwFgzFZk0dW
xxIThNF0pyQserhYz5bDrhyUHf/mth5uRYfeHPjpGR54LEMY+5qFBJNRK0/usj47
MLribYTlMOr2ySkSUV5cIHJGz7DaSnunAsofkDKGLkiFpXJ6L/zr+9ZFHNoyXGVT
2FwcOZoErvTLbG7fB5LYJoeRA8Iq/kqbFT3Ef9QnHio+qYhPN2Sica+hI4vUfhbr
w2PRlzc8JNtrI+FtWVIT6IPGBuwGbVbX3hxfYddAstNUvScTPrXyCYBBXOVJ1JQz
7YtPQVjBrGwKE/CR0BEGiBo0ONp05dE4jll0n/3VZFlbrjw9xbXOa/yx6Euqamzb
Ih1RkkmbR2UlyErfsPp0CIt47/HfLu+fEUpEUa2w2c4QrAGPubH9t7E4jdU8jQ1d
kOhWNvUZHKFr+nci46yX+CYoIYKJyf2vQdo2wzFT1vG3CueiK4d0tJ4oAeqR1pGF
Mbr/n2QkigPfdQJ3XFLbXxbZrybOxk+WEiZir30Zy0TtsOQqvQ3oBY7mEZC0jHoB
Bgmt+DIZtnmVbiyXX+ICJOmV9q/RqEZKHsJnX1DUg6vqdaB1uqXncDIPb/FoXecp
ojyJnAyOsSe6FyOlEE+vOdal8JalPTfWX/LlIqjlRrLlo6dpzlugJm33AvpTFrtE
HYhO8Mf9MO1S0WP+EBl1i33xlrHDDU+OFASr6G9OpP8HO/kKMvRxiP8K246f/N17
cdG2Egx5UdtXuzUQ/LbSKsV7RXIiTl0L8F0hq/3XM8sinJNDGhT4azbslP+z1WcO
W7ILFc6TzTKXqlpCT5RuBWLAa+qnZ5CWbwyxqZfMRPzzndXD9T1w9cj+XYQKFa/z
s2FmVt3FM2wnYB2jx8FBl8FXYPwgdo0fHcBCgH/0JPsJCX7mGzWcRJO7asIibMzh
5uQ/PiFnmwnLCZZGF1OFx2qyv1yAT1tgaxK7qqhFWPbS7NoW9/8ZKM1wPDB5RwRW
g0SsWF9RtgC0xoX5S3ePsySL44Ea7DuilEkiaOF6C728Q5pPMFWHRxNcv0VnvXE3
ebNIGKb5m5vUl75xtYMHsRrkRnwB75rJIUexKAWHmBalhPlRKshmIuuNSr3tJltu
dzrTMbd3XvMdW/ZskRCP+f70+MZah1hYmeLeTsCUrV6S6ZJPKdKmwxRUzoVfBgPk
I5uS13IHF9c562oYPu2k97+eby+6CWWLKFo8Gm4IFcnxkp6tEaVv6AcpdTHib59E
G0CQ1BY3Dh6O0tKJEIsspYEsJp0dGuIRbxjoDlkm0hCieZum8/PFzgi8W0Naw2yB
JtPTVY0gczzoX6z5pSav88vOUcfQhaaXd1bdpn9GSF6kl/uTILEMUPB25h7GaZ5d
Z1GbzkcxgL8bmjyejDdUij2tCdQ5rjcTN1KOvvX/kArCk5fghau1rRVGvDIDWXT0
bnyVr3IKdHUzNpXVTA15MUzkbp4krEDYSZfAHZ+ONCt/NXgUlkJAP1O/86uCf0t8
FX5bmoTLy/r6VHCF+OPTW53LkYztbGSaIzCXbJjLoApj1eneD/YP6aoNBgtLnFey
F+Evgk4aAzjZAVgxClLn4NmR1VTT5BLN0P3Sc9kXSwJvHZSIwYZGxeik/7Z3gkHl
6k1wvZsG8acKjYSAk4pc/IWma+TxAJhrKmKGEWf09ImhVqGsowZ0Ia3dIsYodjm1
ijVOt4f2Dy4CSLCXEPtHgJBbjQsGi2sUHpSEDgBowAR3MlDjuswz8kVI/PSMxZ/F
j93eNQMOzK+aRCFXmZsv5ptLCEdGMIa6vRugfY4hEd2kMoWgeqqTV+2LHs8m1zqP
LWkHszKA81DVmW5LnQRjBgk9xryRYRMmo9sUIGm67IWnVpIseI7LDwa02akWjmPk
m2lrd1evH6U/iqOCyVsfN8m8f+GxlDbLbsHf2yITL9Szvk2zUdLyPS4BpbXykxkU
jmt6xsUIeQ2VynhSAJEzHxrtlEivmifSjr8+H35Op/wObvJZt/6XpTHwgjROM6N5
efL/QBRGw6KHq/qTxFoQYd5THDYeN7m/1OJaQZX4Mg8bKQhzTHhw4g3P+9EU8puS
vhOjy9X29aaVAItA3t1eszMvCQLHQGFlY6ecNOsUws8QRUw9AnFijYnENqxDYQn0
O+mvFV0O5mql3TCvirEliqZ72cf8oPW80Om12pXjzrPRk/FBlsk6k388D3f0qov5
cuy4CxLtDka9CVopbaIwE57YNVdoLkfY/mpS9JlrsVPn7YyT4x0SxFrYhi+JExRe
3oZxMqZ+2uGRis+E2pbTRoZKWCFL6X19FX5kBNP5Ggu8TmUcsugMap7v9wSkrzDF
2+0wd6nZjkrwVjE33Sd31YUpB3TGJ+QdXBIWu2ms2ereycziLlRvOCrcQcsBfBZn
d9OUTKGgQEZv8240kQyM/at3rq7RdAm+TfhXMipdiCWL9gI5WBGaTIx+D5zpg9O0
PcuHfITGGqEeXtt2ywf2lI1NN8UygdCwv4GuSsumeCXh9KPxmuh8x0EuHKr8ta8s
fE1/w7yVeTEquIBtxei91/ob3TCWZzLgNLeQg2bSlvm3cX4EONw4izjJFYdnNVUP
z5wk+oCxtoEwFynr9t8zoqzdmhmtoO6l3SzVEfGEjfu6HZmFC/tSHMJyOQVe+FcF
9SRXIDUzKb/RZY0Snt0XsVu4XZOB0v3vGKGYlislMEnP/pH4d5bLoVy9JdnFSZPD
or8Qu4TuFSBSLSbsGYNRZ5I38RwrcRkcmG/snCscQ4oDkyOqoG+2tdnttQeIoBTQ
lg95lPd/edNkc4zJd3H9nzZQJQzuTElrmDusX1OY6PAq2pDlqDiqpUk3/J4FL2jd
C5nTS96BrEfftIPICw2x4wZr70/yW9gko1FoAqp3IPPuelnfKeJ7GDBkrWcxJPVG
4L0+LDBwAW4U/d3nyBVODaJMDEtKC4cFAG3UGVYYynw1sVUZx1Fv8xWFOxRFkDbk
0pW7QGreXyHNx3zf0n8W0FbWrrmuVlYPGOrsT1ykfufdeTb5cht+XeLRvAW5h2Aa
/GUNQ64brgETKsFLDu4DusW31MOyZF3Hig+yVfkpXWbI1IgSDVsa4E2uB23pG6QO
0BmyMWg12xUf1ejth5ReHU1x1tx/lWuAy57VTvoxEOSrxG8WCIZFWXseEQFwoViF
Ka7Xit1XCV4HMqRF6Tqg9f/TDs4AH8+cU4Tnd6scwCNidOxphJqHeEQ3HeWdZ2lS
L615iAc+QOcRCWCDJpxbH53ZIQ9T2tCMWSYNyJ509NtqERwVf33+f+EXMSMbQOAo
Iq7/41XVCxo8CytDaJAbMkHN3O74/KXU/xjZlSwefC24ftHAL/vJLF+HyR9w4M2R
de92Yzm5Qg5ZfqR/Z7zCjoK3nw8z29GybYru9YDONEC+6VJYnFmFd2t7SrA/5rSf
/jWR8P+hMlYbFhgHzvDhKAfwJi44v0r2GHKKPHlViZY4ymqrdltUx0S8XDqxQ5+m
5KKiYRICTcJECd+WZyQNatGf+d/tBx6IiOAVYK7uA65mvPZ27IyFjzZsGPEOLfLw
z1o4ExAHQpGGznRGtacR/fXU8GwY2YHZHyIA3VkpzeaYMqRX+dORczeHbGqVO4dW
kedCj9QBviFRAWxtem9adUjiCB7ov3Ve2KQhYOJ68dUSlcAbp/Nfit5JUrJc96Yi
G38dlTB122TnQpV6LSCbx7YOnM+kWiW7lihwKQqA5GE97Qqfif/4Q+wSMDP+YWy1
vcbWArG4gNBUoC7CRVWwExUdJapjJgFifJlJx6YL50Bunk8pPUsiKVki/NZTxB3a
8qA+t8iclE4UlY/nS14jj7IqJ8CAPctnscA7b8zVXsanMbv1JkTk98sIZyKNljDk
+qq/cCzPK/i55NCEJPW9+DysgxcZG4kmCDx7mxFklmKRpVf7vvFL7tVvVnO2Mt8s
K/S253WfjIeaujB0Wtl24lUP5XXOckW23fiQaYWQYdYxl3A6CWuBRIpNb5U2Wn1/
pfO/192Tpu7ca8hDJDFTZS8dvEr/ib3WUZhVX4rfpFkLTUB4rBjtD9BiUVucv2ho
HXg4H0eKHE8rk+MD7M6jzFHl16gmVI/wNxgm06jTzfqF0urcqbsqfA20UZGXiaot
0Rw5AF9ay5lJKsDN8kgZEkwBy56tDsC99X2VMI6kOFJEaHc5htBh0Chm/2AguB6F
bKj4d2OeTyF0tSAZiaZSY83zmnDZyFU34N32nlhkQPwtqVNtnc0CwTD0HvnvOVCM
V9zdfe/9jIda5XkHTNSg9wSleznO6l/jvW+dqw961w47w4s48x8/G/aFRN8Wa1o6
5jksNDURJd4cqqnAMLF3zNkruX/amJ/9dYmuVVk5FhRNqfHuVc1whOA7FfDUBXw2
QUYd378qDqiLFRHmCOyUOhpX7IQ+Q07i7ajAvrfHmQLQ/bRcHKFYGhYNcG7IDYLp
IXJ2k+Iy79yxteobW7yxm0a7Y8Rwik9xpq1WRJfP8Lq+fp50SnMRVGFFZG+wHmfx
+ui4hHX7+5F6poTKNE6rB7gNDyMFgugyxSTSxVNiviKahvhyIgcQv9pTRZBir231
5hHccUcYdZ7uaFemOA8jovvc8bFZHloLQag02NTn1rnqTSeUfE4Ej9jWDu8kjPc7
9yoETArJ0LJ6HuEDvSgjqPadTTiMRUFzVIuneuis/0dq/0ffmuVwR5CQ9/03vNh2
3NoSYIcIVBonHXDCJ3JOdLfRIEMgl79jRIlZg4JEs3krHrqfzcR5sclnZYyIap1P
oWoqeVgIxj0JQS+1D5v6zubPoWkG2zk1L25iGw4JyP1JsoUglbU8FXndWgnr5bmU
N+m1YsVwII5rU5HMsV4KOEc6sRVuF39AQGEBy+G2Nz+PKA1tVUUIQfTgB8ZZ+kAi
jNmkszMq+4diGz5rQ45j2kZyo+Yk98FFVy7JrqPKUNuuvUHcCW5Ke7Ov6WwVV0ws
gtrStLnY0TOaL2759blfUnf5zi/RVtpYe6In0765+Mggo2YYHE9baHWLQyTruIGQ
pwCGM/Y1PVulwAwCTVL//ey7C49zKHBT17UtYe6uZOXR7pVCxHnxnOZeDlRFbaSq
9c+y/gRiL2btp8F8QNevywGoJrqKvedUGmhFblOaoTyGTIaW7gPLRNTrwBJq2up1
46Gx9kAf5Gvs0Fo64PoT1IohhmrNyCP2gW6gpwqkf+KcAQ7UTkuzYu2MAExdxgZQ
hcUam8aQmgp2tn0OWfTlnMakh1vnlYLjAqZhwpW5P99TMLrnEOomSqTHk21eZ+Gq
WYvPvJ0WXnYHluhmqEazl5tCoYNtb0JiuwESeWi0NSD6M3ue5O7OUObfStvAVURw
x58RgA09vB7gOEl/voGgaUCCtHBMIRpgxWCPJyJDLITnZKuc1AKV3qkvMTatEZAo
cVKsqF68B0xP+rRfeDi+hGMfDA9Tx2jVjH1GC7YlDr3cPKwNAQ9ZWubZFIV1zSgt
9ddgxh7e+KGx5YnRst++mWHEAT8lfNY0qyS3bMuF98trxxPn17GVEKtCbeieFw1v
sMNGkMCBkezx3wTGUo5v/10xz8gKin/2pTluaDSBQm3q1UTykQTZ7fX3XDj8JG9B
APDFQtHQKg3CYxq47jg13AbNGqgQgVQmRWX7axPLNw+tOP8F1Re4axWo+ByIRo+C
z29zhebmWZbs1CWw/vbo+9xo9zmssrxXmuXJE4tkdMCoUFwcQTECWIhgfvUD6R4t
ejhQjZeQgLdt4Ykp3BlPI6imCU+KKZ8Zv/t1IeeBdHgl36HvnQMpmy02OsKj+HAX
xTp/S9CIdwheLZBz6y53rhe8RkZafUO612dBp6YJkB3JdaV5W2VPyG7CIBVcbeYC
404hFIZZQFZaA/lxnQ/9PQfH5qcuTh/EBNNhb5ZdioGZflsR2nZr+4oGok2kbBUm
Hk/3cylG6j0Nj9I1zBnsvjmJ2M3U63/sYjfZU3jimf7+9fkp8CdiCLoCjKs4FXTl
+FGbUuBMXDFIHArSXlRApOFVAx7F6BQQgS5TsJ/efMkZ/qeDr5mB91Z8JytVEkiy
lsP5bf5dVTzPgT4NUP+aeK/hW5SWDKjYST7x0s8ZVn8Lyu0uruyJEpOz3P0qzpzS
i4yefPrpjo4LzGNMtrg4Hsj3PJnahiKDViFXKASKSbtSoz4eTOIkdJLobb4f27yI
qwn2/YZfu0h2yfaVHxWMjVyIDt/wVxC3gUabMz3aGU1HuhYy/oJFXDNWcffz2FSW
U3uTl5ZRpYP5vN1oDpDNSynyVUw0+Ggw32PnW1gh4BzU5+h+fiGmsa9uGyeQqOc6
3NJYPoOjnUPCB2ZGXIcRrP+8hPS0WKjfQtJtdzsQPYAkTZ0hkeor0B/0Cw+xf80V
sjeKIhWYK8Md6k9Qr3JH5W8PfbIAIKWCOLFK/P7pjAXdEDB3lMNzGSohX5lP1kRo
ckgpr/aXMtPrYaque6zTyxyEgvZYPCGFGEVyyq8yqIn+2sJYL5WZrl8PMX315rsl
mpT4sLunG7uA/bhyYvF2Y/iGQvlbuRqKFcGisF9Sr3RNbPWjhso0BxfnTC++1ObL
ItqT4Ex1+QGw7p3yJinXVSpmFXqqmwH3Kj8BloESku4iZAQOOMpFwExyF4kFP6YU
XXeZuv/90Ljs4ybGb3THFGOj0FSTZFuw41uV073ktdnbLSNxg9c585yhJapOuQ/K
VUa/DLITz3CvIpXL65T28jksDpgc+amT1VDM9EDq6xXaegezh5pu+0ouUz6VfTNe
cbijFZpexWVQOA4VzoNR0TE8Mn8V+c/sZVSuPk0ziP8f6x+fqXupLC7N1UNSi+U3
aa6P0FCfkcYgzAnyU7g0ckLxCz4ERlnCpwySYA+uwE/rvSS7WfiWGrWsE+uoOAvR
YMn+6fogMwTCvjV6OhXNScvdsMFd9hqDktxM83Fgg/C3zCne5V7oDxZLr6vy0ObH
HZSSP6szjDpv7GTrs4vKcO8Y60uJEHeA8t0Q9Uiur47GKPZZhoAck45kNrv+n+hT
dwDfTPJUC7dinaV9dvy0/03YGtSZyGw4RYhHpIOPkDaYvXY6WoO6Nn+cTJqdmtAX
fhJWr8TK4pexH7O6PBqm4JMwIxlVr6nNs8+CdEy1R4kxkPL3PUkBlMQn3WPkQk3K
CEY30lg401y9PlnMCLtsl7YvHyKXT+sb03oesRSzVpLNCvHStnFxxPw/ynasJXeq
2jKXijEBRojXFgC7mlUxtZb4NGMYK9ElNVxCUrkHSrwsFhxsSGCSWAdLuZ1/R4rw
151kfiuqxq7yC15B2uQCE4C4C2FlDWm1hXugEa/rpPsYfpbBUeR19z3ODvQV/9j1
uycZgTr01vLEQ6Ph56U/2IXQU21xjdbyLtWsiiMSoy3E+wbC9RClExjgFGVYCuRk
oaddVp3Xs3c8SOPnQaBa7L6KBhIoTk6Uyy7avYozoQHzJ35udlJGoLi91DZ0C8gJ
UvUjgio/g5kYGkpBJiaOaWnpiudmkv+kmrx+Txw3Xibwa1bjb6aK6I+6uC9S0SEm
noRj5mVu2UKrbw5MfYH32Qf7Bw47y9wo5edS3H0CsAtZQzpA1OcAme18/CVEH9t7
8PpaS3kVZ3ybA9J2yZNPd0qKnv4fc0Ru7TYMj9d1nBqsOZU28wqYngSYmxo6YwL/
P1P58IiMp84ob53c5FtkKnUsPBv8WjWi17F1+Rb0b00nJwu3ptU3qdmqGVaaeG23
cqAiIajp9xW9pEF6j6fHmU7FTZuX3rv1ptwk9y38kkmw9aDawIvAmzc+hdewYrDt
TQeV5jUHcl+qI+lPhtglHjFytys0mR5z/pIlnlYOo8+FZP9M/rFuPPdGVvAF3gba
24J0DZgJhqa8r/d9wwawqlufmGawWDZX7TalSbjrwYpTf+Jm5WxpGKDJN1Z3yFyq
jHUSyrw2qH4CEvIQMF57E35yWaJqHSQdqEm+eon4QL/TlASq6jEbmK4E7KrDBNdG
xIKfEULhLQBovY4UluXG+E/NEVI3s/ht3KCD+tRvydFwVzlKgpQeV1vnEagc4Mqa
arzqmSMWQpop3dYYkzCxQWgO4VwsVcoW43fJMsJROjwjOy91ULr6CBHVIEglBd0U
fJoOrgFdk1YI++2t6QK4zmmy6x/tj9haB0are0XqBIs+NuD95igbPzYaX5zUJctt
1m/EhEvnf4J1ZPcyqsI/3vKPFf6Gt7mkcaZ9VNMlsexzxFod9IfuOB/iHmqqhUaz
Nm6BjjB9QYk3wmaN0rPA7SnAczSYtI5ptR3VM8EdgnYqfoGUPADAYIlHsrmTLY6F
gznyVIGH1OlxiXri0XtlhnZztWlcQzDSdz0Drom6oAWtQ3NsG4kgtbQT1PAybv7e
R63c+cKEGLdNRYk0M2+BJV5ydY4wlerYtU5I9ccAHL25jX9RDeeQMOa8BiH6xO+b
vGGgxMHPcu+jMfM/55Q0/ZTt55Ik7FdXNpYqgblmvgyFST+SkYDeDhaAsLoFVT4A
ngmVJlfrH2gyF+V2D/p7Vc+eOhYjLr1n3ye9JGjXxxYKbNapQRs7wAbMtJFPSfgQ
Otn8gMlN/5Wu8Gt4tQjKEbRjQtcInZjo6F7MRdbKLkaGbm02vBUOi4uSBoJm0RiO
JgSwDGItMCiMOc781vWBsgy0LB39jaUsD1QwzBIPg9xeDi2+Nren6TBn8Knf53Vx
E34hyeWWpHaIF48bxa5xHJ9QQwqY7Ev0qPG1gtALl0oQrqnSiT0PMZSeOlaFRlBV
aOT58rPZzpeVGSP8VvIo7VrjSceTcWYUdba8MKZW/tEFGtWhPxsEeffY7dylQNhE
Hq52tQu0xbMF4KtF2INriOfiFKiICqUjGL6eWKtaL3idI/pqRW2urGGzFfGP9F+c
LHzTwj20Qf6M4kG2KcraNOg3jG8ODRHXJfqoccsJIG9f/5nIx8GKutu2LdSL+Zje
YT0UIOKW6RYAnROVNNKk+PIkIQcLOH5NnDlEJAr0vtLb+3Y/7PS1PyD630q5rbKc
QafdS397xS5KcuE0vOGaw0SsZ7vPpQMbuv8DbP0sdhIy/6gUCTf1XOXEuYfXPoej
Js/FoqlppqWBawrlwSPkIXXxI6QOS+Uoz4qL7dpZY5FiqJYcIps0lI2+wGXvh8TT
2pcLntmpvuZGf7zYGSMQMrL6ptaF1qMyhQW06IYl743062f87jTyJy6mVjyVhrMk
rmv6GSjkLzTMIQtcxFziaYhWdDE8Rh7b2faaO/rYcCvQdp8uFP/IwF2VcIzTaTwD
NiyP1q4l95hnUlHIRs3mibcaDliWyGvZi0A8e9GN4uYxg20GXJUyl51L70pWWoI5
KkPxghQUHF2qCJnbLIWlLIh6AsXMOth12Y/Wnvb19amMCjs2LaEGhrUyOmOtDKaF
0GQaR9L/L3Vr+STkk9c4GwUsOVM05VcXMhvsou+/9mSTtQvmmudnIda+6iBMCz9W
cy4FdZhjy49SKwwz7yVLlygwA4haKqE4fVMBbc+BnlOtvkT3GrFjyLROrwDh+Kh7
ibzxiSAuPNUREQIZV0CF1X7T2/qP2MDxnl3XHr2StoNP0LPVeBkqkHjh+64esiUk
ia3tuExuGyeHSRnziGBc7jtWipF6RogjOHdo32mCYBPjJgvmTthTIYKdWt+zYumX
DIr1wOhucpZWUC0iJ8dkAeInbeIShbtIgjRh2TrwOkSpxvHS3y8OsZ+6Cid8NoCN
QNBos6puOqQRW3hvLDhkY1BEJrL42DQpWXEpt2bOPlmmRX3KcAGcLClJfCeXeah+
oUTEJFw3JHCCgDy/h5akpDq8CePXH6EH/h+oixWfvTljgXD4VdaHFMI0f3+bov1L
vxJTTETzABkW/tGqfZ6A7mLvJCfAO8gSL9nRf79tG+zCUOCuunCU9XMLvu993xfV
WIWadV3QEQ4+bKHIVlFCets/6ONQT1rQbV4WRPGdukv5XHIAUu40/zHFixm+6lsU
pRRHhkA+6oDe8KVA6F5oXWp3wE+IWf+OM5S0oOuRdPO0Uek/n/WiCLK+rvMm0mPB
XyKCcoydijUskh39g5obwNIUvPOM3C985VQagbJT+V2oKYLtqbHlXeB3yeqjELXe
4WmS6xWdaED8w+KUpALG+1EcEFGbomAzy5qysetWbxETkp4xhIczJzkwY5u5uzfp
69dbxy0JRQJ6Tt5ikwR/X/81XFAeRg9YW5RF5l/ePZbTG+d66eSJWy/QEEWBdDzI
sX+YwD5d4b33F+bZOh+ss7JuxXQOtyZBAlsdrCl3D80D6B70pScn+N6/Jn6U5uNu
ikJ5NMHFulzCp54/SQfwgGhHAJZIxgsgBnpTu07AtBo4RnfjgTG4twcl8ZRXZWyc
2mHqamtA+teL22vAgkqchD+AZBN+tYS9BDbUtBM2SGK4A3778e3Zo8Bz/ubysopW
nhgwWe1z4OSqBJWkFBwRQHDxAwCy3VWJa9hMdXjNS6IBooxZXU2cSuPcpjowQSiX
PUbu/RMEmfov0XRMXXw9KHy951v18pPVPHtmyWVP29Mrf+/feUSnyfzyUVUF5u2k
6DTp0edIgvvTuxW6FD4aMAF34yQ9zSE+G6sO5PdY/cwKAgFNldOnjiE+n8/Yo0Qj
uPY0kenLW50Y745v2YBALq8tkbHHqiAOvdcNXIGoYu5PDyUozQIEK7FfKtLY85yh
7CzejmdslhijpgKjvNelfPaV+hOR/4Cstgq5IU6jTKOjWAylbMwGM3WSKe+Zsmdu
1Ak/nhz6nBuUY9fI6qoh0vKhOvoSJm7ZQ9TY+lfl29H6XTCDT6v7bK3FwckycvUo
4qUWXmz15XbQvaVxhjxv+JU5JGTw5CT5EMGRErenTLrumXY7xvIiWy+ZL0nr100c
9B50uV0WM7w2Lf9cofr4QXmVWrzFXAgj/Njqt/gmguEZSx3tlBcqXk1WXj4gbYwB
VPBztw1X4RoxMEDCKiQjhBaYGUvhpqO00x+HWPP5MFiOevRRL6SlpsvvyqesI3PQ
8dU6I+bPfaurWfVN1W4A6CopseflRyPscIEhyEe5f1RT4nyVsTYHIeQIGEzW2cAN
9fJ3UAOJG0u1JmKse4s4TSrSeC1PWltyNl6grWJvLWycJl6zz9BFslL/c6IDrkyQ
WK6iKILfEOGSliolx/PEPzKT6HzciUEVAvmXhP9Bhr1Odczysk9GsMuMzxunCzdo
BC+QlYJIJeZUR206STI/amUIrYKphFJgvwOzTA6ocoupicsPdw62ThFiEZSfKtIh
uNHy38kwPBWKsZftVR7vSg+d9n1do3soSo5e5Vc9QKo7NAIg29PyQoGmI/WGlPhU
BHWebxJjC9GpSVcO/sZiLx/LThGJjlYbGfq4QMYH0wNt4vBtMAVgmFYg2TgnHRIa
RjW7y++NNI1pSRgFR4BSv6HgA8TnKqc4n+Ak3PBgrbES3hRvyrzlvhluzy67jC2N
dKKTj04mMuM3rDCuDCnmPf6IzetdBqQO7L7X65xB5xmhx6hXQqmRo9e6jqG7ZW4x
2dyDsVVB4fhbBhSwiWCCnpQDtvj9fSOsbbImljr30jhAI8/sWceJo0zKm/Y0BQO/
sbjXX06bPfIZrvxeVnfSYuo0JvG1dJojfe+z3wQ/DC+fa9dGr9RFI5Yza62A1G5b
8TDDeCBp97Thz2pyNsDcVg==
`protect END_PROTECTED
