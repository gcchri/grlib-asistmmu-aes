`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MuLo4AHLC3rEZ7+ucTyzpdrvaOpz93GHjYR4OxWjfMdSMjXD2NRCV0donu2C8Gr/
cqEAP0uHglONj9PhB6r0HdFt5ZZY7RMDP0DH3z9or33ozTkTdxUPUxuJy0lG183p
dI0MfF+qYwL0ZVo7vfm4dnB6sxmU8ykppK+p9g2JymwTZbU2vzVEOfg5kHfA1OXf
bc7rnHVW0cUjBUY7qeWhwHApyU8Yz/h81TG7grf1e2zdDdVyfNh51BJVgytfKiUv
5dqBtm1Gy5JFzz371+1IAhNE2WWr0345ARixSP3hNifHIcRRsMNYm8DQcEQ/+OY6
oRP7ncYT/J//bieZvS0QuNoMPUayk/L5Ip5/3TbcDGV3l92Z1dzXbwK/K0DpYCjU
HVhlABFAU11IvQSnBYbHqw==
`protect END_PROTECTED
