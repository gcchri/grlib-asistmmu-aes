`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NxTun3I5BYnoFQxPtKfW5K3NA5q5Q3AGfAs3lZKOrLAE3iYZIzgGEMsE5ctZqifd
TL4FM92iDmtA7YEshuTd05s+QaCZqgCNfPam7pFQWCzt2BZ3qULXS6qniaoJvMdX
KW8bYBFVYn8h8sClTgpY9sXiL10T77IMYyn8DpFxWFrElPlp99hS0WGZc7q4Vli+
g0USozgQlNVtslodXKbUuykaZ77Jc4aiptMgfBNt08QRquBJlz8NQQdeWadrC1ok
gXOYOfv13hkW+7w7yJKnQcI2nwP4tC03p90nM2pFOcY2UxTuiCkTX2Kj86/cbjrF
cPwimggjz72tdP8mRNjJ0kioCVGIxYX1g1Y7hG9gqWT0ioOvk515vvsv7fZ/6JGh
B0xaNMImHA51q0VvNi6/E/7hjA80fbBx4phZi4voIw320TEARw6qk3w2xEE8kPBr
mz2MF+7bRVCdWrTbDps++RpxauQlz3kATQD8cPO+jwYIEkV+Ye71eAYKzceOVFz+
tvjPRBPXK7rsECQ8WRudz0QewVqUfxn1O04gugC27cL95OWl3GialMHsFQK4/fCg
0J/g1Xm/oYbJ8vUWGgOehRP38bJdkQeshw2sYhniDgdplDkuvmcINjeXjlQVhdv3
rHBGKM+ko1dLEsdIzVDUe6Dr1jFXsOUvcvJ3YRxl0ND8E6Ei6EK1Mz/uxgKbU0aK
VwwqxT53tBJlmsJQGd/1EYk7Gd0MBOlWFyjTdAtqnBg=
`protect END_PROTECTED
