`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sRh9+17Pls1Ym1AGM7OG5IYT5ezt+KyMVa5heS3sc019K6uqdJiM1y23L5GUgozp
5eaGBVyW2ntijSoSMt/fea966dlJCHS18t8EnmuPEse77sa+SjUVmvM8b5ygSLRK
kzkrfUUOrEa0i3Hn2nAz1B4RJt/C+GylgDE2RqpWhheYuLT3tt/XkRJHZ79+2DsO
TNi42eJTF2OvzwqoTG0YypSFZl9FT65cqG0579939SXjmrAfEOYZyjWYzXKZD5Ug
q73VZKHCpmp3fRU9dsZ+theLRuS+UxSvjJhlQmufHMaa+p1NIjIKAU2duDsWBlwZ
W+2/YDL/EM90YqBeIcWNoeHkmJtmR2K7cQl42G7HzZ6HoFijI/1of0+PxlYpfszJ
d1BTWI2ZDZig6xw+JUpHRtMs+mJANb2mmPd3OqmEl5g=
`protect END_PROTECTED
