`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ViXFgV4xGsjj8vouUZERiuQn6nhlE0MDg//gJUL/ylg3ne16+2Em+NL7XqnQCMGo
TpTD9g3PCUT/5RHD5eJIEsGVkgXATzXk6+HI7gXNU0r4YHncCEhSMkhWoEFU5t+0
LV3QAi12HEs/0yvA8kgdabsMOZhOf2DuTi82dKwlp+m/fXm10m4Qzs3YBYCGORpG
wpF3RVa/nAw+wdW7LqZT6sAFmPKdmsKnV5PeU0ONux1XCUyb5jsHMvVgv365G6jR
5xvchhWZce3LbAWP/vLEh5hAjXqhpVVrLJp3BqHv5lU=
`protect END_PROTECTED
