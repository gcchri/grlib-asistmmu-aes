`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4F/HkJa/UPDxT6wbwKSg3ka4cpoC42KO6eksjzFOA61qOby6XxLTiiMK8cdD+gDu
WR6EJtCPPT50NhySDBIsjCcwl6hIQIqtNAv4rmxiaesuEgQaJ2auuvHWr/qYtG6D
9Ge/5nlyV9XVzXrR9W+3nWbyNWG3yILvbAswVmktbTeZZI9nmJ1ujJDwYEf5KO2v
2ik9hxMVNjpxeLBCajplIItU/8cFjU0Au5Zm/dFnf2BH0OHxqQbGqEa1qubsGq1G
hDecOJW4p9+bw25mRUnZP8XDQW6bKCkF2aJpAXoi6uJ16wIzLSqkQAbi5bBpn+Ht
HGJGVkgW3ts03wP6YQMatw==
`protect END_PROTECTED
