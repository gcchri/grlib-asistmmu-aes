`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8d3gM7pMJ8bQdGv3VRgeIKr6/VzdwZY2dAzo2GbLgH/5RkyF0rImb1DjPR+e9PNH
VEb40HkcdGX6TLASpABWpfzv8BcUfp+vLJ5VEWtVKm54bWHY0uynm2vg5GwMudmZ
fRqYpiKo2RH9PScqXTdCAor8kcF4NphIMtDYq7p2PmQy+jUuhdLsjfA6no/qtQSM
sH4dsbPQgGETmzYRm77PMaR8TzGAwsjnOC310h7jnKC0qQ2enguxgyrirW8l+UVV
W2L+JvOSqH8txRW5wP8XtZMnS6fzzzIf5BSZHaGYJIed4nabc+rY0DvNcV89k2rh
u6gwpzE+0qWTelge0Zxspxo+chMah5QZLaEtT6uk1mwpcNqYmrjB3qm3QJ+Hj+G3
x9ObeqGCOheVhRjYiv5Jqzr+oSxL53h8YX8Q4RowVZ0+Hgrt+U5Z/jatKKg8tull
wMwt6HVLDJh1V/3zPokEjrRzoHAHLzLAnhluKY2LCHATMNE0tLfBe/1i+I+JTAbH
pGI0r6OXU3fGknbXaDcLD47Yg7AVnm2WbMfe+w7Tpb2fBv0IDUOt7WCPZ5jjUd7j
t/1SlpiGholdL+PSpjgjxtRuolgw+1rXMNVCczRDxiFhpl7/k2FxKYqcFzuEVJT9
o/8iDVahQAtKJdFXG2FHR+n+t1CKCh0w1DLdVERfHvrL22nB3kLB2MGW6FaJWuNO
kcCx3TJWznny31RIKEQli7qj2LycouEDo6B6SjMUdF7Z4LUOgVZR0zV2TO4VyOgQ
2XkOoWvArRsHgwCpjZnh0h6toTEgJS7CGQPTRx3wv1bfZwsQ85+51ni9vporJTjs
PGGHdA8EoF/PJD9EQMOLPh3w6grMajusRoZCwSKhR46EYi4VCw5RBO+S6bhMkF5c
UBjwGqewYWIorY9cwnnaMu9npl2K3WHe2zlXYpqtgNtGfUlf3ncqYqoQNKv7cBrJ
O33OpiJq7e0AMNKE49y+bf40VHGMzm3u4H1VUgx9/tJ2BWZjMiaDHljtMmzocDAK
QJWmCDs+J9Cx0TCriYJIvC+BTdEHQbmZB3bclNgycvvwmzOCQI5hUoCRfQvnxwEx
8EaWZblBiUaL0mnEBp9eVID5BEYO7IPTwmwhwWvC3zE3o8AcRNB679yhF366zoq+
oaIKTzPmaNeAm1AkR9QxXGiUHFd22sqCf2jSkBm2czVvIdBTINfDapxWAvABmrDz
Jtno8OJXagFWSDwUk6mxyD8mQzrGI7SLnHFmTfNniPsDZ3kSV4EJ781/c646UEmY
UqRrnzRnW2Fvo3HN/9E4+abZmYOU4IpRwcUJsUfsgg8hjb/5H3H/iVZToC9hKPwF
5/qPDHdgg2ip3YTr4TsjcXzMdeP9LN7LpDOOhhsxqc3KAP+7S5XMN6mjJ2nS6d7A
`protect END_PROTECTED
