`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
++wEREo6dTlOeJSVz5gA+fX0eHVL83DFjV+cEScIRF8hn4zJOnXsrS3QmwXjfGu7
rffhZgtIcDL5qKvL17Qzl+sYfBJDbaX03PN1umAj90a1J9dyNEnwkSLirol8PR6h
4nRLHoh8y6w/DaOeiDeDisgVcMj0qHUIu0mwCD3APekuEzDHgGAiQb75exeHKIWy
84RjE0yKIGGDkHu0v9o4PA+DfVmyMXBKp3dKaxfzf503cz3kyozxUXvkNIKtU4vc
gx2qeAX2j4JniGcDY7vcAr8dGVnE2AcYdOYyEGaBuEORwRFLpCcCmObJxoMc6nEM
gR+l33EfG5qf+vlefv4QJ7BPkQCltjV3RVG0Coly/j5x7l1XuzPDl9TSUb09dTvM
`protect END_PROTECTED
