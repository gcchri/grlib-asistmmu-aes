`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ssaiz3EBPAjGQ7ClkqHz5NTeZXByMv0SaOL/lvDs526ekY2r30O+huDl3AKIq9k/
8zBuQYg3MNwqrhF8Ic7rjTdYGUf90oxPfIUwXKD3+K9LwQUeyntRQWVnlylIUYqD
JxnIGWR78Tn1FysuRfHpddYBxK+6rZs41sRio3QK/JXUd8yiHrz9MF9uSlS9wMh7
TBOmO09eE4kGhvWDf56m4N8syCsIGthKh0TxJ+3G03SDKAHvA3trB6Gb1Nwvdttp
tfn7q7x2JB9xNrmNzTebyA==
`protect END_PROTECTED
