`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aqnN6dtXDYyzsxZ7vfW06beX2cIvFY4k4r3Y+pAEuXp/baYgjvtUROW8qKHBg6Ov
Zz86U+WYPweFBIL+Yf4B37M6Tdg6mOsH/rSEEQ7S8lYlQE/NM2ruCydbnjQ8tIBd
zDaDYY69L9clzGyJTweg0KZqRxpPPc3OiGghYI5kmSM3iVIX6Hg3RjkLz6vQCjki
vCelWEH3u5s3ZAdXXia7gI/IlEr3g6pC8fNNSerZOti4eE0DCnA3Q6h/yoBv3DDe
PX9vtuTodqitZCuW30R2H5NwxPyN+FI4sUpI/n1dkAB5xoeFkHDoTh6P3UJgs/SD
RD//jRUs/qcz/m55Hs88f9d19rPjcUqwA4PRytlkXXspO+gVk+GFUoxg2+RbKQfM
ojd4XMep5cHX9jCGtFLXrB8cMflRgVM/b1qFrpV9T4+otJW1tKZqg/qdH1ruXtqA
gf0QB+quLJXVNcT0VyfJC3v7jZZSqeMGx3FTZkYjolzj4KjOwjbePuR4OjjR2nO2
raJiNGg1YxB9E2OsPL7k2j2Ohup72lyBqa/W7Mv5f+NE16viqjwHzIhAZ+veZqb8
1+hdPHFzhGCAcXl5IDQVyzZSHFVB/S6LoBdnI9jxfgBSLcCuom970Zg6KKlnUZVD
NnJn/7frQUhGKfl3+Nrequu0PDJpYGrRsFgamnX+9WR7/72ijx/ymJSLlfGArNS5
7n0t6ZTFbFKC+mgeAoBaG2b2IOx+UW324EgKBBld0e5dwJ5dX9JJ872YvbDUUdKw
VhkW4QSGGdLbUApdoWpnQcSt346ZwSptuQrrgNAuHKLAVlduYiRRnMDWdgPvcfBZ
V40TtQ7yUrdB+VepHDduG1ZjShXTHxV17fyxMUHCFvhrbUi+t2HUlISf3ZNqUKCv
i4tgQIAddQAlB/q/KS3TaT5Q4qNo6OGaujNhI01LO6DXkoleQ6ZkZcXa3lSchqjR
Po5uZCksj2fKev9iQr4vzs+PIP2rS8V94HYJp4lzOY21ex2xhoC4doOwOIMipaP/
B0NzPn5c6TeY0JkUYFGpbV0m4APCUvg7sfNzscXxzPRFoYS6Av0Y7PsT42gI8PNh
IUEVwfZcUA72qPCRWxQzPI1Vp2dhU/dTysZBHqV0QI6Brfdg2m+xrbk2q5HDlVvA
SdVu0CeU5IJ2o4aSsar7FSxjKdO/mbQqtsAAm0pU7BA=
`protect END_PROTECTED
