`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7bfePQYGNCIMvMMDdMDBufjg8LI2tcwdetHXI9T7gjeGaMbY2pnkyJ8+ySjI+d+D
g0JkOCwognCO+D1WoyGsRBFEvknJwwmZoyBoBJxSRYDySPwtsarhp/VQ8/dvqPuR
yEC+BmCrPqNMgxz/+tQxajaWvOu0puDUUWZtPc6Bf1klGCbk5gSvGZ4qWfeHRQ2o
0XD9Z5cDAdJmJS+5cd5eRKnEsyedb94jmZpoUZlBSFpi6WBsfelM/wdPuCFqLCAk
efyhZ+BH4XaizdC0s+/g72Tp9Nd6vX2JpFQ3rfvHbsVcXlshYjv8eDCfzOnY8mzH
DERlmeyzZ57it2Le1MCVwmgCtm+u2riOiRPZgSGiMrv9ts4PMXOgOh/PrMlQ/Q4/
SOeKKRMOYQgGeYefmKtIjCzyU4m3KulhRAAdqHSCauruPtDfav9JQYT+mR47Owmj
`protect END_PROTECTED
