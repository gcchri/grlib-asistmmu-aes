`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
chtcOe9B53tS4FfylxdlezTh7kLJyjq29o4q0AJokjTOPOiX2vFhmLyWhYAXHKni
hDGgB7U7LlGfBTAPitOkkAqpksusgKHaIS1gmuB9gjNy5GwQ4xkLrepR4lFo5sc7
9c+qhmH50y5ILEbNAwrFWa6iv/AHnw7RJgqYmGyIIDYzUn+tiC/w9qsALGRrjFiU
dvblqB0yzirTBHn3hIpHmraJvgHIqhe5qX2M//8Km0LncHRcIrJ+IZ2Wjv5tpDnf
3BmMzw1sISLVLLnmGrPcMsOfb029WcfnyMNgDBXUM0MdY3cEE22VeXqokNJ1oTq8
oSXavcB+NB9eeuF8IFD9W8G5JT37WXSP1ElWS94YHV9Fcfo0/ibtnADz39qUn06s
HKzAaAMvvaLLhNMehNgj1y/ZfLjIvI43ekmniwl1phUgS/HatCsNKvBaadzJRRK4
GxY34m1fElDsoSiNK4jD4FWGhHIdNNDzLmTZ0UTFaY15LKbNLypwB76UHJl4sJXa
`protect END_PROTECTED
