`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HpderpqiKmTxVisNkw63UWgDetvsZMNApCIBWkwI5mPN23cCCAeB/wx0Azh/P65s
/3ZnQNGxhAV0XHzHiIHpJf261LP1hmmN9J8F1kkpxrd7tEvKk4F8/WjSY6KYfKro
2GW8cDFMemp5r2AGlW9VCsLE/rwXhPJZFyXDskpLpQ2G1YKol5CPaXGtUonV/lD1
ibtBsmn+qlY7WCzM0XZS8clFfdsguyVSjF174f7XtE1Ie9/QD6u+ZaX7DBsySRJE
+JBlGzgCLutTFaFwxmQWbYpBbFiK0Dr6eNHFDl2kRVEhTOMC/4zR3CThdCu5IyMg
P12DUa2IUT7y0VPlhIJAP0XAi4z2RL/cuXOL52TTnkhUGnvO1JHSoRqza54Mp+5j
+t1DUhMpFyaIm142oEfjeAjOqbMPYS1bKE23XwXV9e09sOM4Eh9/sdGR9EZ1XRnL
6brVgi07V3hlQ43J2eo5/cKEiS8Gcy86ZVSvG0wJlmwL1SUgxMuO0Bu0ikJ9Wngg
G6l9+2q1ccznEUBMJaDnccJtHSts8a9BNpqJjLJGHjo8GpnTyKkhiEzOsqkdIk+S
gzYIb72EcSbyXabsPrCF5lWKDtZ1ClcYvObK/FhLQw9YtJOMaseDG74HFrRp6puW
wsKq9JPKQCehCuHOvksCEQ==
`protect END_PROTECTED
