`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mVTx73+1VKPH7FbY1BMBBU5gzL/Z1J3r3f9sWFizjmhCvHkTueFarzCSAfVBGECu
KV1HLvQG80Hj5pqydkNAzNNb9QQtU28SnDhf1WtVoyzMlA62ktfBpQ7nT52dJEaj
CGYrNxxyV6A3gldcl4h9GJcStSrgsETGQRGmjCYaZrzo5kXNwey6gkJBKg6WkcN5
mytMmNVc3sB6ROpQt7cA5KtvjWzFNcahH0uAsMF2J20ndow2EHaVosZ/zuoimlCS
bNCc848W5p6CAe1k+KjsCcI6ubVCF/i2PYpEp4ZP0IBUOfYXHr6SN3EO4mpRKbhy
+fSS07W4unlPMrHnE3UfL7SA+9nb4lyRVcl5ww1fHe97xGZ0vQ6G+X2XB2ejxRIJ
+Qw4W8Omqx6R9DiS5xw2g/690beCCsqcCQ2xCns3rgq9QPefwI1Sc+lNb94X87ci
ZPxWen+8Ynx87Y4WRv9Y5ccf1jgs6+lBWnbpjD0yECngHUFGMHft+bdj8NGaSqyD
KnE2qbJsyYX1vBpk9+vAhHvX/5KD4n+O8zkPybzVGIrzptmMqZpFMMWZO40N4sds
/654Hjc+4qEpkqEvVNVa0HVCkSF7LJTvMKDFphdm5lHUrPU3pW5tHzgjaWK/CD3+
`protect END_PROTECTED
