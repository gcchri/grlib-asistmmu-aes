`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nv1WzVFZIa/Krjl/4/1/BdmgJP+lRBkEkOi8pugcvWSrs34I8tNupLQehiZUEk22
3kjr8YKcGBKzLhGisMZqCYp0dGvZZ0xWkj+z1Wzx4zNruEqpQjd/cgeWi1qbsgI6
XT0b+y2GPaz7gPXcldgtopyVN5mEYFOEi0R+kgLsBaUQflhhRuILnR6+EuVH23Y3
vprlYaZV3x3dS1FuesZVjit9igyZH2u82z3VdhNxY0mwlWl64YmLigiLgALAcqDJ
e0PCmcMnzU7zZ8xEljU8/VV89BnA1+e3WBqZZk8YekrVizMiLCUVNDPCGv0ggFWH
KRWuOg6VbvCu42e3t+nq8iZGD1OOEu5YUoQYa7P8ZrxgwFUDHbQq62Zle31DkkVE
o9ZJe4GEBughafEKcBvddu24kDHZ0KMTUegB587yGIAfYs2aed/BD/WnGyRKmuBh
YLFlm+eUhDxi03pCBBM+lipfCJxU+2pl+tqxzP7poYoH1A9k+YFd4ea5CRYF0cWb
`protect END_PROTECTED
