`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I3gg3JIXTOtawuQJIMJ23OxuiM97ZYyEcYQlT9lmFIHWMfB2cBRmJXTNW6g2nweD
pn/hfOaAc4ZMekubNCbgzH2df0+uFK0mxTcSuVH+QhumwaiY10TGjox2uEw64r1z
4ADF8FEUbqlIC3bettetCAGlYQSq5zyT5/Ojma1pbEp4AUgbmwoY3rMacSDe9mkf
2d5FqBopA7tfXN5JdbVi/5a/GCptOXexBBJaf3z7U0uSX/HrGaMxxznqdkpkwhXL
9Hm9aS+kE18s1N5K06PbMlXlXsOleoXIfkXahoVfWyo=
`protect END_PROTECTED
