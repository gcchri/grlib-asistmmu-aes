`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m8iWu28qDNGN2zDpHKkIIKojfxjlchGU/gTtilux6kJupNzeXCS7oKACsHrcUrhi
prxshIijBiH36zhU7txRV6HicoqQPJuRRBidLMtjDu/BG0gOqz+vVvi8cK0K55GF
quwI/4NUTYwVwtGjuVfiOIxFz/Hrcz0NjCIzc1enbKFuhjoKlD7q0dCkqTAqOC73
2wmJJfWuZys3gJwFlxGO24AWRnYbqQz8cx2BV9Dz6kHavexvpKlMEoxEjMitiCzp
mg2GK2NMr1VbQhRyzTns4LOGD486R0WujpsNZHlH4lzknMHninJmuqKkVxJBBzNw
2AIs30cnoDk6YgDD6F8ymcLAN5xcosBuSgWLUFxk7kLbKhr5WK+mGziv7iz6wovK
B6VRiDtiJH4URMB19yr5IA==
`protect END_PROTECTED
