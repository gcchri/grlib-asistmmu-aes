`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vr5PW5ZjQ3tqHg+8jChFDMnxhg8sdv9/lkv0ZX4N+YkkFRV4Z+rAHB7j3LgWhT4z
rd8WbL16PT3aSkEsy+s3I+Tvj24VP5wm+9rhjCxU2gMs4G/K0uj90gjrcMaayE3G
NRLMfe9vvzf7Cgf6fObkgRwzBo7zfu84p70pZBZUBv1tVW1wj/7vk9IwpWj2t9y+
9MECyGbvct4/lR2KDaXnFhf/bkTaV8cyaUUm7QFBjlh87CNlqw1efxSb1S58L+qn
cxNXh9ENEAcqntXbY5WBfUvINoLEq2PtEiaSnbL6WTdwz3tkM639h6ULld7DZG9B
toUf2lNVRDOl/ytcf1GRVCWDuUHgCwVh49/MKp+zh8fxIcotRFt2+Se2tfw99MMe
cuAS9zlTxDaEW9t8sqPUaQ==
`protect END_PROTECTED
