`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VvnO6ZqBtj7+RQr9DBKG8W065fPE7yqlzZ4xTxXokdngth+YzGlXRtYbr1JRIUlc
0RqFkruOnAxmBPensCMIAeII3mxT9P224shZmzpLHYq4ffvS85Dg5x1gvDoOcsI5
hByi9olCq+89y13psXTgOWg+hvrRtMW0JXsks2Rvz9N+wubisA8wv4lCR6cwPUwm
YnvWu9OrbDmbhTXZnVAegZTlIZgR6lkAxoCvY7X7cgIMftaAyPLaBasnxyTS7fpI
dFmfif+bqYihbTeGMWxQ8hz+kOOADZ3Tkl1W912cvX+xJQ5WhN0QJTTstis35IDz
bvk+XipDbpjVTSx+B9edP7KvZFTfPp5AcZxjdZvbuEOvqKjhUuOnFw9pLzOMX78u
SSigiHn7eeq2c0eqtKw/+jC1qc/5RmFuUaJIKniXRaKRosjngoefuhesmK56TLcQ
`protect END_PROTECTED
