`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q1RShh+hGg+bZeUBl7sHaZ9KQ91IjDf2tYRmjL3faWRN1+n6bZNQb5s+vNCGNF5H
L/xAxi30IWqC7PxNzbuGO89UegEuTxnekghygptDCLYoSF+BOhsWqwnNWYv6O82n
WelgEz8PN6y6E2LJs5v3few6fNOQKPoqftb1eIpKMU0zobLTtIK/7b0yDRMCDpyo
wQxJf5KzloQ7RtMgCz9QTT6loc8cMqI/CRLGMHELwXQFnqN25q2zleSifyan165M
9XsPhPxsOmbW4AlCl+7w282tK7fCJsYTuTYY7Q2zw0TijpggLaGEB+OlL5VQk9/s
4fMf5ol2O4g+xzv/lY7SjD0wjJxbCzXIwqWssqn6WA1M1WOSC+t95mkNG83niYrw
NxT/k0My1wlLQMkK87WWvHPPDF6UOmGNS3vdfa6VA/VdfAEssj09E5Ib+vDDJzMk
3WhycQzcMP7aj4CnqLjMjoCWojv4q2ISDPoPEG6V8xIxfYET4oNCealdoTf3XRJ8
gfAyChnCZvkwfD/x72IYZCAMwTUHxNMKaIDsHpJhZL4xOYuaie18foivGaFMe+e2
FKzomgihfhxw5Gu8EFHFuqe5H1tCOb2wqUe7mVg7zCeg0Wcf9x/B69k4+tZbZo7d
ncD37Osr2/k3e2cdk+346AE37fHUVdRFdcUhXz7sinkMQhfQxkkosicYIfNtG4rq
Qzr3mSYwXyrK1WoFdnTVbPvfoTNi4ok1XZJ3LxJNKj1HthooGawlDUaz3/i08oNw
Kr6A4iUNhhgqDwKwoffrZ6nrpJI0860RGAy9KqovfzryDpzfjsg/0OIh3xrnlazc
b17H5CsvRodRKtWUzxhZKIHgidvBgC8P3bTrEyOAzm+MDJCRFtOehdCex9cNFhKD
+9n0Z9Vz1otdDMjt0Pd7O+NnEpmFSppR7B+HoDQZexX4dWck+uKiuJHgB7ZuHV5m
9+4v6gkklZWpAt+fMxSi/9oVFNZqqEzOS9qSHEry1aB3VM/85N0r51gtmRR7BG2y
P6TqrvYubcfPmGPo6aDxTt+gtf984ZsH1N/r6wZlWJuxPd6g5/SzN+y1KUx/i/B+
kuJFPYu+ynb5sNiq1utIfyeDjQU1YlKrNJO/C13n56vsPg1+0FwhHO+gK03LKMbc
0/8IQ0iYWh9gU+FdZVIBT3gbeox4dZEOAC9hOicFeoIHhrN1r689wmaTd0kIfT2r
Kzc1VvITS99Dcs7gQtbj/4iw++hOYkd/M7Q08GVB3GoelQGu1xDkyW8JKUMCD6Zo
s/T+b/eLvKSTu3qzHAQ7JZaPQRy0o1u1L1x57QbO3+duGsQk60Q2KTEpGFa3PT3Q
iOM/TsfovWc3ZR71kWjILOg9DKP8goabkYywXvU9GTg=
`protect END_PROTECTED
