`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0IOSorij2FIftYPbihOcHfCGDdp0/q3/no4zAz4qBsrAhTzZzBfOS31BleR/NVJP
gY82Dxp9XRwzOHkwtKWCfe224AgU4YzlgMFxDkFvMMJFf4znhlSuV8Ad7ggd2hEo
AQw7nn2zpAp8VKSVR6by/ODSMvpHC2osya0W+ESmU3fB1UU8K3vMgKZMIP18UzId
vH2qEK0/Y51lNYbyrk6gCzo4Ij7NUdPXwHBvbmG5wfyS/qMoif7pthrYr+c7SIG4
Hrx2FW7BWC63KNoDyunLCfG0Yh59mFsmIH5wFKAAaT7Vh0yFgzpDjGq0xAUcCief
q+Lhj+29wTWgvAqLqxJvGdqLnLyKTqeFT6H75HwTUxnYai02FRNEPg+XHafYPL6A
nJLFQcY3MeqaIvDlvePyBvYhe8yFgeVE10eNpj/7wOmaVvA8aoyrqbmn3fQNBsty
5FrVPf6rIQZg3UV4wdoxlzPv5D3Sl1NQr5xMQrQNrWpj06YabK45Pwe6A/+zbiUn
vafgWI7X6bHhy3A0r1EJQvZzcuhSXurJbtReMUKf5UMCo7becN/NaArk07H5CLvp
x0wtqGtBTtp4P4ggirrzTGe/fRg1HsT018b+aYLvJYUjy/A6+Bl38SEi9wxxbuxB
I6185cIwjTTFqpPKHA5Lrktgv+54zHJ+Nt9+NnTwCIEp1xKTBAwdxx9eo6hiBtam
xm75UrdSRSWpO3w0nR6YBzxeiqRo9WHHEE6Yn078V8w2hy7ihMQiIIGugIGQ9yZE
k1GQMaYrip6lijzywoZ2TeaVPTBLErEsdLZZVVP2/+NznrC/eUdNqySTaN3LNJzU
LRDFRDtWUAYvkwsjcptqocG9mroHBMn8aCJvbvQCT0pfAhJ6xN9lz9QJDmIiSgUV
VI+ujvTh2fWOrg7XQSzHjK8FJbnraxY0KCvz8/W9dShxnwZjFdrp6fEOflT4iMTP
xtdTNmrsJlXApuDFXAdwRGGunmmdnjJQcnFQCBEx81qfUgpGPnr+Z4JpvN/luzhe
`protect END_PROTECTED
