`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HXuCYsOstdKfAV6RCpVh1qGC8kk9JxFatEs6iOHDnfmPGJt7jGVWMV+kd3u+JT71
kwCevJhtiuGniDZkW3UIfs29i531h8VKjPtBY38kUfDecz8Dz1D8j+K2TkDV2u+a
PFRvBTAHuPaHfjPLWA/0ODti7z5nr1z2sIvRsGqsl9roa8ZQJ2lt1S9AjQlLghra
3gs+P124voZbSBIplqVYxbpPL3/ui0dzkYRpRZHXto9oCe0EOTSifBazUqKUEO5N
NGlmY3LQngwt+TD0CQnqBgwpdsN1f5LVkGczW2P5gS0fXKATkR/AskX7x38rXUyZ
2b3BgKF968vkMlUFf/7og3YTTxCFPBLvQ+4K3tPAuVoUoACP+8Ic08Y7uIIZhdet
BhHpgQdvyG8Hsej3i3lR3wzqw31dduNOOnfHbwm2kq5/PycgmtE1aeen4ceZCLxm
V9J5gLeKbuKOeM+gvRlPzQ8PAXguF2c1K/CZHZ8YS8m/9YR1rYV/odVr0xWwEXdZ
eiKJMXT9D9kPCUriYH9ED6QzizvavG07iEOB8MHPC82+JAO281ps89Ke+uD+IY4c
ggtLyg3VlM1guj0UEeR9Wg==
`protect END_PROTECTED
