`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fq+gI52XVOtg+UCSXBMvOVvWdVAkCFGcb7ZW+xlqxhkEoJOI2a6OGhUZXyKYmjNK
IZEc/THYnC9sHiypkc//DMjRTqh+AueW7s+mOalv9zFaU/YuiU5G15ezveIk/zxe
Rj/xnsgLhq3c4rTElW6+4YTCt44e1LVIBfRWDsEMGK6H/kkGo4PSaM5WQteg1ft0
aIvmHNSrIKG/5NWOE0oZPtWBffDSPrjQMsR/KN9aYTyGF1bZOCZtWjWdKrdbTcWk
ASY60+/tAncYCtxgLx1Dr8C0gWQM5i+aV7WOX0QNhdGYlHSzNWnDDoiEFjaHJWTt
lsa1Z9wTVhQdsS7wrXKX2svR2pfYbziCstccdCpqYAi2yiqgQhCTejVqo7aEVGAo
nhBRqRyyr+Q/pQxFeTWceLIhkcbIIXoaGsd1GXG+K/ANMYbSAuKDTM9yr5Y8LZw4
3rRBa6NY/76INffcYKi9KCwfO6O9Th9fFTL7EFWHmi+JVR46JfLgNYRVWB60I0Vp
O9V8JSd9yIaokdGIqxpTTw==
`protect END_PROTECTED
