`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DLy54TCE5Yt+pfzPWGvRLGLufvgeMoBunpxZACm0BJpFrAr4l8TN0J9FYiBKkTsM
pqfyz1Aw2k+bE4VrAx5ViqjyhswD4efeDAmgQ0LQ+1+yyWw86d2GUvfg/aeehqqG
d91rp2/gD2gG1qyMS22lDGT7Eg2wHSpdNvpks4rjnWVE83IZ5gvXMbLQp+AZQfJa
/6d9epXTLttimuWRHzBwmYtTlaw6mC07dkWef+QdTpuJm1vK//Kqr8DXuToZDxGI
tGICEXa6Jrt3OfPq9O+OOWMD4q6id54P9Dv88yMTXcLRxLYIx0cwsUt23KpGSrMu
9O+ZF3dn3pwhEd27jzN7c00qn8fMDS1rUJnP6J6ptMrVo+if1BvT3nD4pKV3YCi7
lc8ZtQL7qIyutVX3d+p1hzaQu0SgGkD7GIRlnVytt6bkvy8Hk8sTh71xeS2l1sko
HLUnCnUvMovVsuqISMzM+4gpybut442RSTRAUuilQKRN1of2UQUe7DO3m8NUwksr
`protect END_PROTECTED
