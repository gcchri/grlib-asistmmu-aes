`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v48Qkhp2a6wyiuJO7jp//z9bavnB1oCOKqg/hNZ2wqt23xy1rROUfnQU8q/wWdUL
wW/9WqnX0R6cMCjm0VLGYEcml5o+S407scSG6co/U+qjBQuXkDx5fWtUgdRIlyPe
VcJFvrjzluO7GVUa5smq+FEmtRk2KJ9R7aG06QoMuMmuo8J2L5jA6U4k7sfs0h8v
13havbRh3gIHomKHIRptul7zXnNzyvauurUd1qCACFmpe5M1ADSg5SVsYQstOmcO
FYQpUKPDk6GEi3EyK878kUHymRVtg52PI0tLvNXvTs9514NFzWv2bZFx+bS8m5QS
QzQkA4aLzKkgfel5D6luXRAVarQlwCovXphH28EKRJhxJzNshZLso6FMq/L5dwHF
TmDFlySJGdOomeAtCgotg++5R5HqRLsDsfYoFmg3pYYhSdOxS7Oj4HXKWLWFq8sK
orl2FRoZH5q8F4J52wifnwe9+UsdeUXJTsztQW1hFsV8QsAomLWDgkVDPH9wFG9E
JE+VD7LIoCm94+NmXwiDqJBmb0xAsK3y5fQ+vWRXXcst3wsQXBe58zT38AYydXJ3
2Dp5gGvKxtmDxTqnUYNH1GgMLeQv/tEQgTqoIuZGkXfqUPY/0ObjloTuYipci8Ny
k2rll4n+qlvvQYIt5Yan55g+QR6yb0HJQ6Y8WJ0unA9KzZKYp9bcLk0/Yjprgv3l
DyFAsx+Ihaz9ozhQACVlU446Rws/JLLH0TbuLCZ4opfqnOwrpWNstFyxwR0JpgR8
xXjYVZjI6iT4XrPanwC0n0cSEv/Xwue4ZKI+QhMTQMUWByG/X/br+Y5LfzDe5S8k
Re4re0Nj2xCxdhO7CFvrSxp+f74vBZ50KX9TnEoc/FSBBxL553BYxAstDW1j/ICH
lZBONCG0gkmYSZFCLHYav7iz6axlJKROzLslZf7MYvOklB2etKdQ17mn+WzZhebA
PNKOg+J/jTXicf6ZcJ2YKngdh+tb9RUTaQvDKzwHvVmDiJAAvpBJ/Tp1izkqllfr
W/sSqgRZLwQzF4LqhD19jitfAbb6kA1WNOvF1HSnoA9hIZwncvXwo2fMPeM6KZGw
HziKUzw33oxKj2HPLXciuVIIQXGiu4rOIBBydI3cc8HQGNMOx/ohg4zdbm2XdvJx
NGnCoXNt78sTQNXKN/AqEfPBt9KQKm5HTVKqq9i6xx/knmuw01QYZE+K1aXU/mrc
fj2Ur1iVCZRTvYOOXX1G8SaHscSc7A7WJt93e0+gdwTlHfEtEjKkSsdXXPLVdvA9
mKnSwy1rIlgZbqE/OMkGg3EveAgRPMHw6QHfSqo+IpIf6fJvkMfI3F/K8VaPiaWt
b4hFQr/wD3pdHsAk3hwB+37bfX5NonPuFtHDvr7qCggTax6NlhREYAOD0iOz1hNH
SyNO6dQZR1vynffYa32V55Dt1G3TFXohSywJ+REM7GNqkPWAWckw7F3XUten9nXE
5KepbqdmocKE2U1+aTvUkqXJseFtbQG9+Pj1vsQsdovs3Tk+nsL743z4BVPOrosr
`protect END_PROTECTED
