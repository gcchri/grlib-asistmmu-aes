`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CxYIm37ibbKNA+AN0ZtxsNpsD5PT4v0/lo5zV9Qb8yDWJq2y/QAh/kE5Gsvyyz/y
drqNqgOpIwzgT850+R3hVQWZ3puXU8QITQ4NcHllwLWti0iYZeWbkkSNtHUxteYn
OfCbGlZObgnqufDJqg+A//luWd2ocKD8aHvSgcFPGL6J9ZXOxBUkwYm8/fLvsSWT
0NF4ewFdN8yViETvD8q9jqSMp04/C132s4G7zSt3PyY5YGEXZwa2MRhy8+a/ItY7
wbEh87Wh6NNilQkNC2Z7XAWGgvlcKAEOR/PRmFApHma3rfG7SzgX9Jet+CjXrF3v
/OIkMJ4sTftl2Bu7eOn4SBwhoZyda1puiUDgDYU0Sjb3yJwN//ASLAbehxRTVMHM
Gl5iEszXWbF3vJqAtWlGI8eqtjL+OLmPEm+WQCyP/DyFTVY+6xhwkl/pP7i7DSkI
e88uK9em+r6LvcB/o20liJMOWaAssqtmav3RlG608ulXi5BQUEpOpHyw2QXhIa8y
eK5vRU26LfhopTtG5zW6i1lK1SYI/MrP54e6NXKQwbptz9KvL2f6tSdBf40jUGh2
xqe901nMTJVKy1a0zF3/vDcau2hFex1tYTF75elMRp2UE4VcwAdqy5uMUawVmTFg
qMM82UbaipyLkx1HqSaCjroRaY8YKRnhSfojKVA1+PMGF2OE8OZ6gk3NIx92guy9
MtfuvSJJR19skbPSGsUQcBtzb64VPxTp/Mo8AlkP27pEkGz039Ghbs77FUXIdfw7
A4hHYMlbT965R/Iw4uTMMftlX5+DLqayaZpNe2odkPnrPhMNL2vKZyV/s71cuU/F
GDxZjFeFhBtet/zBjgS10gAsMQnLb/ZLd5qcMyo0QgTCvd6HpOJggUy72Y/IxhWI
QyTBm5sw//3ZZZs9Zi1ZGJSTFGP1iIf2bGHAI5+Lmp8B9HQll33F9W/pU3kFXW+f
Gn9IlfLCoGS8OC6XJp0wbXAaFsj2gRBS69QPfuZyqDBjceG2lneSr2Fo2MbkBRpo
uhxITbERVoazHSUofLPUt/dX2ldKGEmfRgAoIqpJga1YwjDligXEoHl/QImdoC3l
sNKks3eaWBZXin0vp1dDEdOHCVUErDnH4DxVWzM7rXwwS1zU57Qa7kmfPCv5TgVW
pSz3bEbdZit6T8Fkh4SGSpiyofXVASt0BmoaGX3nwMA5CRmxoZUJoBQa2rOo2bLM
g81rzImnT+upPtxE5UJRu8OTAb7AdUqAXWItz6mRplG7eRIeT9a5cGpak/znpiP5
XQRYOy5AZa/RgZtUPI0Dsar4YUK7VUyaMvJgs1Cmy3/mXwyXxvWc22UO003azSyt
XjP5QPvJIklak9KMlmwNjO110hGsrbPBCo2CD6Sjr+dqRMrSqr+o8Orkfk9z+Wov
LmbSAAFkKHBhmHm4Fiz5qODJtfIhhIG5mRnOi/fV59cbVOW7RtI1bAJqL1AGevJ0
l9IYn+q3dtGOMHpmmZOJ5yEtguve0WL7xfcUbJzSV2yQcjOA2YYn234V0CEx6QgZ
N8hc10E1g46c6fOqpQsWw8dJrEpEK9hZushIRQZvfn0nhsjiT7CcvTDpB7ec7Xom
hUstKiElSPNxbmMaau5KSMBHI5Qi0SZc4a0zzFrTeN2Uh5OJ2jIhGaeIwEGXAomm
cK60p6BwZugektuYWnk8OdTIE4+bTF5Gon3k3Wt0TIVMTgDA71292z8gw68O022n
RgyLr9DTK5Q7nNaI45lm5erGvvRCvk0OsUvLyDcOqkVFIplWlCgz1/Yw7NyiTFA8
D2JzI9Rx8JSzJ+vPWc9AgJgL5kuYcSKmlKa85i0bPECuw2IheImccLJ0jw/pgWXc
Al9GeICM2GMyY3EiXagwjXxkQXWHpkR9NWeek6fHretA0Njaqj3F6JG/3l4UERTK
TcVlQ3BeMQD2XBRryvJSSh9IPQaLGTlfdTMpqw2YrxpH3sW5uFY959r5wBqcqJox
rlbbvswiJbW7nQGnUnPLr1OxVkkuBX6uNskB6V4GTcXJ4dmASBu/+eR7JbO+SKaL
wUgfEyABYZxylPv0KksRx32JEjXBI56MNmYUBNIBm37cFUvbOCGV68d0P487Kj4J
ykl7s9glD5DWPJPK9btES2M9PkU7UtZj2eZMiBTBgM83i1zAxRJaya57eJ8o0jvw
IlCPhbELtolGwkokxpKX1LlaocSJo1G2HBnkIQQ5TERS0Hu/hl2dW87yg+tA+wAx
r8ufXtlW7joiZBD+ttB0dJlvqRg2ubey2TRT7EoHoGWedM6IzMWZhk6iHSXZErMU
9G6d6x0VW/FJE/uGzyJuNGTiPbnJP9/UjhPiQ9WAvgAbvYM9MaKmf6RKKuDwc0p8
tK/YD5gFcuJxQAe+P9+jz1a26FOZrsOccc7miAPPLl8TFR6lzj5OLZLuWgjtbQ+1
Im6aRomWeli22scbkJyMYuN+In12dJyFQH4a+4Oc6MmOQ8VAg8zabYhzOlfTSWGw
AAAgsp4K93OwOa0DgTDx0M8vmKtp6VX48GXwR4QEjyTTf3kv33ssaORs4XWiYdvN
FJMpotYPv6kX5Jp8eBs1fRgG1Q5gumu6CYHb2q3AQB3ioDyNCRDX2OmDrssXhTGo
oD2rceYfqUfd6jobSXvp16vfvYwji5eaaH22/uQicKfA9f7xDG8RiLh3vJEI7Dze
bMIvRSCQvpzOR7FJPcZgGP5laVqiMix2kA+gVTis+I0VxqLIcJeaCIJkardu7IzG
QNYPCsNyMLBPvUQsm4FILdtoSGr8ZS+5pl6XFFwtA7p3afPsiotCq8YrqfqxAgkc
5g9X+VBCROhKrFIghGqw1ocRXDUU2PyiMOIkWajuhe6D/BilkSyxSNM36XbA0R5k
rWGDYeskwbx/HFECJnf74pXFndqYvEMLY/7ukhENq7Bd6dn8iK5lY6FQVpvVTAiM
RKx3U4ZSd77WE8FGKHPA7jKG4VNbDX3PNzUC69IQuAMl7vbR5uvO3UvILd7TCQec
spjmlTWCcyzNMihfKgqyNIO+11EwKEuqpdKfW9LwcdOa4c6ZT0ZTrXfHeaBvvRi6
S6Tn5SLcwtLHt4l4hWhr06bIos/GKfyycDhaBz+FBoiAfl2ioagvMosxIQL8sOc2
vY/GZ2iSKzhStMKktF1x6moaxr51ihtfglIB4I7KThFztNJ9x1hFeJpO9+BTNyEt
Of9r2tjjNd1paM9iLThyg6yxViLIXXTZ/36V87pwM80n+5CQCaSgBNueDTqzCZkw
tKeAC5nXg1IpRKt3hvNJ4NMVBrvvPnFY7zteSVoNc83zdb6mIFklc3eOKliiz9fQ
M1Vok35WxVLbcjX8sN5NCqnB6pa4XMNAYxtHdO6KRr5UXhzha16v1AwqoT6N0ag6
gVabRCtrsPZrC1i3T4ORk28DUGq98HQvQSKUPMNNGsCCKB99rdBikm20fQ3vdhtb
aCY1DGwFau+lwKjqdnytQztvQH+qj2/Afo9qDc73QlMjgcwYIPn7QDHI2DGSzWIs
JwjQo8ifDbvG/0XgxFych4ww9Z8OmvJZrgzOqek2Wv5Xu8rShc3Y7yULVk9BMEoG
YRfTUrPqeE8tPkVc20t1xUGXECVE0hryxj3LN8dQ7189qcuvcYc/NkHgjs3ZLNXW
3ySAvMDxs/67RW0cs23BBBcX+UVFlXxhuZHxYpiFq0FLFr6zzoTQRDQdOAo2AYhY
+fSGxU21FWFsvoMEhqkF8IVf1k3Ai6cbzPrnQgn4cae/260Ow/AaG18f+UxEn6sR
mcSt8D36xf+DWHRkNlNt31QNSYDRdu/hDpkR1drGAmqhp80pDOlKG6af9ShK4Ql0
fF+AahKgvRngB7OngFkjaFZDRPziqjXIkD3eGIat65j0BE5fj9dOCUNL/lHOcgSc
29qX9R0Zbe42iNFBte9j0eDi/716L0WvSaJ8QABdcZPFWRehrg9jnjkh62GYQOlH
2Kd2e6op0k6hHRr8Dt0NaE7ShNgcUAqod7YYClW2VVD1jhLN+SjAk6nQpmSxRMi1
mci7R9TiUncW7ppWbuXaADlNiBCz1cN+3+VrLjW2qxuoJsoIFGs1gkhov+S3Svk2
MEb7N7YWtUYaZJYaOZfTXmiabOPnJ002XQNOO+VobXGAWbJD9N9LF49jJXziqfVK
If7JUoU1R3LAXmoSl+Mi6MWBBxJT+pZkKk8W2FeNsdz5MVgA91JSc5ITNp1UDeCq
KjhiLvEso06W2xThQThgxfX8chUhr340EuQTd4XhwBH0RbuuzlUFkNrLiVdD0Vqs
FzFACH79FgerTIv2zs8z1APnzMccvNG7nG+FxNVaKZVGAlK775JGpPsyNgShAgms
WrRJSeuX+q9zr404l2q+dqrP7dyEsARLUd9H3sX3wFYCtGESZcD8UrQd21Ml3ODU
ViweIW955L+7DPERtb+qiMCcKP/ibB/2+SlQpC3W/h652M3LFM3k9SW8aBY5gLkt
dYLb45mayTLOV5oHbgfXwVD64UjL8pwkS5lvGv1LgOLa9O+luO83VPL1B8bMzPlE
z9TKkIqbRwYVbYcEPYFtOIdKmiQA1jLELqrnoyQhtLZqRTg6b0/S3tZs/s1qA0wo
P55oxZr6ArKWCDgHzJsoDmrgVtks/ZmYdy++8ImlOKt1jtxJl5kw/x/YUbgKe/Ax
sQFpR1jN+4BpxfQr86j3ey9+iftdlSVmc6ou6XOcMu+0T7sJGOq9m3mWyRNjIOqU
vU5c5K1H4usn87d0mEA596XS2Wkl+qPxIQK827GHkUkYhQUaYS6XzLc6svIu7KKp
B0+Iu18qa7nY3ukc+3sfbKefbIli3VjBoj5XysDKjx/GCsfuIzKrWFXt1AknQYjQ
1bNXu69X7IZNt3Yt71nb7hy/ojjrxwLQwuvFRXVCOjBnBxLDwB1pcFpCsoqL9ZfX
mh4JSIpjkD17dSxLZUrFN/J+saAg5RhSrcPlqemKTXn7ksSKvCKhjV84jpCeis80
gq5GuTd5F/tfOeWGWFh6aCfwrIDUFnzVpMj0SDiuYgRxg+zZ+JpVZGOyWqh3Qcaq
CzrJyQK3rqRTXqfKGDeBjGoyQzPLGiVhtN7xzlKBzfnQlozcNwUmrVN6o0kqBCwY
L0OsdWKfV1iG9ZsCtx0WMUbmwxRd9yq8bYdNC6haLc2jB7UaxkDoOkadU/uk7gUl
5SgM4DLq5FeJjgrzRyjT9BLp1X7NXXCcsYRaiijoyVc88E3SLj5L9Ww/fj1dIZAg
pgTC3ECzDV4clWCbAMl0h399WKUVPiYZZXK6TJA5lfq1sqyvxUtSvm477cfWiXuP
4yIdw1iHGltjSb2HTE32GqVg5O8UerF+9knKv5w0k6kFZ2q0AlDlyu2l4l8l9No0
Q5GwQWQgnl0vVuPPmWQ/MwVtkbH+l2rUDOZF/k9jKW0TlJax2TNnH8SvB4az47uC
SL2knTUOFX0cu96DIH2tIercsE+LFEIsI1bVQmkq2gJnsVdfSUCMp/gwEX/s5YMm
ORz4UA8JsobMCiD+V3+r1o9GEsthwaYqcQiDPXiDuxn5Op4s9dxtNZcq3kGyjt+q
nC31zN1J8kQc3Br2fRFQi6hfCIbHZab2BSn4blJzGrkpeWIswon39+1d7WBhXPWF
H6EzOSwA6WOw+oo0Id0+olTb0TX7oJQ4fc9iggcYKSua+cwlVfxygHq0sUWTllE1
JYV6jTety4Vk8eaUWc2QLHvYqakLtRXnsBQWuXlfmriSlfq2ZjkacL0R4tjito43
aoR7bm0qW2GNZAb4Dmqho7s4O1hWl2NjaOQzFlWWlBwc38ZUETUGcI5cSMr5XZkm
DNdw9XID3J8z1UrXwn4sq/FPRG17xY/hCHRpazJPdbDltXRCdIPPKeoYSbzAKwnb
ZVl5sFwJswrDodTRasl1p7DJjTk7Lm74n6udGf2OHXzhf8ICvCmNy65ODqhXgKQg
hi9MpogHPoGSJA0GBGAruzI8w+frtt34QKLRsbbk0/nhu36aBJV6PW4YkfVVp70B
65R1NksZ0jg22RPOLHpNr5pr3m0UMv8FFbdDBw47p0FHci4HElavHUZxq5YtSDKw
kSL7J2SCUfhsh9YQnqRxJUYAGYnJjSmeDLTBXoRoCJp08lhbxOCqwf9mBqWX0fkd
OQkPRLkMQDEW6g8YZXPlCpzhkzGaTK5fWy1M/qyO5M3AfZO1qCj3nUnGz5oiMXUh
3hl5Q5XdjtGuwMvz0fly0OpERSHq8GrLKtjeXy7fkuhpZjFroVkTx9WDFFXySlXH
YGdsgTDbqrPLdhvLRphgs3z+JJT9gw3JvRdEJto8pS9jWbOqeVUYpbNZV6aRUvUn
K/ECIeoCnJHwTJViVpkfn2obrY0V0GvfAJ+QQ7TvbTdaCAwszk+TW6FjLvxZl0/6
HPH7VMyjV1WOeQFnAuN2Iq78Yb9z0XrxYL4zCflA9tvc26LYJ516BoY/6+i8ZifE
9cOsydE6WKbt52x1Ok9nJsSEAyRJgNPwG83gqbh2oqyGadFxmPhxZtM0GycUou1i
hQHICnkE74Dd4pNg1wpOHOUNHK4RRXWr3JzkRCyoApE9LgmF7eFVlBGCHDzBRvso
oefE91fwfXrIe1hhTlgQ7T9XFgExZaDRAsrWAXNzlzhjGYJQ65Lh/dQILPZFGMio
u33DqRd11JCVf3sNbiDFIcCgBmkxO2XutFBkrlFRXzp+Hi/H4wmASTSyUCIdAEpZ
B1KS/qpbzDJJaWy684qKdNIHvdY+hr/iZZlJHCzF89V4QjecIds8LnjcQr0PbqyH
hNWhkt+mR0twODhjfkfT0KCnAsJtMZf7SJwMiO2blnZs3l5EcT8OtbUh2pkFyT5n
CX6CIndxuqfHzu/lI1YkThubMXPNcBhuG2uE/ILVEQ3xPESjDK0kwBT2qz4z31q0
dGY9N0cgAXfw+3Co9qtgmWB0+9nrmjB1D8+a2i20rVndhRPIPZpqLAXtFZjO3gZb
aQrnh6peQaBg+EPf0LU1qcJ6xYe65HQ/UW2AYfMWyz37HaMT2UFI2cmCJmhw8DzE
dm56Dje8DP3nNWpRftUsUKR6DfT0nNd8TNCsZKfsgfMLY8NAOX9ti/s2BA4ryCcU
dJe2rwOc8vRBCQVbByQgdBStzgAj5dBaKddLkccy7ry3oQua43Qny0N4YWxo5nTR
aWDgel6M+wvuJDyNaGUtr9r91jPwD6eHbh4J4SnnWGl3DDQdSLGwT+ycfMW45iJR
SypMDxUMqgreroNu02WNmo7vS71u5rVeL/VJVpx86Me8RPsoNS2qpoNctoLijXIQ
W2amtxoVE8PLU9nqd8hz8t6aZ4AQkfF9CxadUqa/qxgiodoEqGlEd4Ji9L7yxJ+A
iP+1VtCDls3oeUi35fzmmv+y5NC5+DHTnmhqN5CZ+X97yhHlNx+Su0QbRxT8v9+x
pKHoGfebau9g5fu/L8di2zFToiMOPdNsCcaJzvPsLQKZze/clAchtoYXjdurnhJ1
1QIhFEgKaO3LCLGlSAFD5UrOWcqt9OijrzJYIgKBm8IdXKnujedecD3FgW+X22+W
mOfLD1YfXSmzuRMwJJDtNG/0ZUmx+/jQURIGXHEcZ1gUfUUwstouBltL+FJaBnWp
13+A8vJRtAR2leVhUTFE4hNUgUo84HJsjFvgrcXKbHE07maJOqzGr3xXhSd4Rex2
xhRajX/vDmrU1+DIE62t92O9Yv+vMd6qAehoVuqza6VuNH5pw7eI422HoH7aBlgI
ITpS5mkaOGygmdpIx4bJUZfB7XbfQt6ElZsJWeo9iWmVtk+18tajD5vonLEPY/uo
ATHFtd3zzprM6BMcyOc8uRAFRwSmemFpEP+ELlvmv2pRc7BPe1usV18Tj016RJ6H
eMIw25IBe7bX/+ILtwjFu9Iknycn4/q+dO8NkD6IAHR1nqrg1h0H0S5lOijCQ72Q
Cdf+/A2mKAupHYmizFC03N46CwHEb9NMgO1wWoVIF4ZuMygNEcjrSLEltL5vy9w+
1Fo1nDzaXIcLHhF9dhr1xX8IPU5ujHNk0MPn+sIxOO1IYEwwn4k4BN/osD45hhad
rik5aSGPFA5SoV82dznif/uV6+1GfpFpbSIi7YiCECX0afW+LtAHY1V1PkkjUSJg
gQYeR+IWWxIYvQsylGXReTGPhoyrqYnp7LF2OC0zMqJAaBai4385Euoi7ntXdcyi
HTyJMBbv1/WC8HQffHZhBZvvAr4IzZiKNH7AZsy8pFX7xiT9YmkR6zIX8KjNUgjt
YcZjphBrPMOqnHax+/KjL0EwtsSltot2lPYW/Dkd1trsgiBibF9Kj4ciG1FpORBq
Z0ujDzff+7gJYbms9PfxER97Ph/abFRKbF4xZBZ7jOaPAKja5ghWFMXuo2sas5C7
QW09tUWaYWgbhLiVGdhgx5MmlgGyvbc47ecMTrUKd/1RxGGqrAIn0t9k5vEa3k3j
4Cfid0l2F6eRH/R5sfepXqciA0QwAqGaJN0956+CPOWtxj3lHqUcLMjRxCov6Eyi
s6mhyhQSMmxk2yixNjNE1rpuuJ3juYE+Q0IBFsSGfUssdx571hvOJnjF0sAIGqTl
IIA59jPlIufwyH/FZmiHR/9dTxjQmtG7rSSoMfo0A1+aaWyef0Yd1AyyftYh5XzO
jxNHpZ9KVt2Tz4aA/4LGjqRAxb6Es6l91vogRBNGbaGYCA8nTzY7IvmWFc6fWDY9
IKIyTGvVsBcHQTbNwLOsD6/qFmvLB5EYx81SvvAj1EkAZP4/plYAECdk5SZrLCMF
m4Pxafwa6h0nzJojSZK5gGjZHuNHBkLk3//gBffoSe+3Fva/uxVJd2/VaOnMCbGE
45bLdw+dbyfqRJhdoP8AlV6c9zqNHY4Y/kLV1YSEwKk13xQfkWkaWfIFa71l/vsG
yLMdLuP4rjc3sLRT0b3aRqAJX+hLpHJzgimqsf7bXX/xHEcyef7d+eRG7syLS/H9
nCuTgS50PYhnMb/GsVHYq+tHG9NPDXQ7gaxGfFsGNyxWizxTIheMQzvj41zuxkhC
d5Dl440qbvqPUHQE0xdBwV6Hey6KBe5r8qcWUqx12fMw6kPBk4FvL2iyBqeAACOm
NtWikf4mTJQu7uWgfusA3hTiFIK/6PACaYme5uZIe8WfCgTgB1SYJvZDFFebJN5i
+m/oh8t4GccCSODHsZMnaOgB6X1LN0mPqvXpk5eZjQgtlyLX+llu5/+P1bKsE/QG
uSmhTW86tsb5fvZsM1JgDmccGo2M9FWGjW1HW0pAfXd+lBDGoJwekmdor7iiLw4V
692SCObVNhu5yevPMeidNgKv4uS9FsNFkqrmbvcfHOcxDrK0icAHECLk43GWMgZm
0D6rTlgczFTOk4EjI4L3ALAEJkHCJ8oq0PV2lmUytQ4Ds1Td3g3CH7BhOTp/6Tk+
NKqJ30S7YhlCKhcU7W/mfEweLiTTCF3hLVmwwNGLM+dNieESYznZWUuBICNjZPmT
zlrKtqC53rJqMRk35bINQiRIWZOwUR86RTIihNV43c3hfiAPF4BSf883ejvTjV/g
9k9pbc/ymj9IJLW8Np7t/oSqmESf3qcO3Dq5qgYxsoGH7z1aQPthUrfuQ266jMi/
eJ2dE4VqYBRNortzzTp7wPOUKcm4+ey8tYppMGvmMzHv7303XU9r8m918DZBoKPV
kZS+2X60o7eKQb3mZ5ndgxXDkMQI0UC2TVHyghkjRn18kgSPMCeo3OgK+NsHww4m
ufXZJFfkxIop3NJuAEuX2McEuqWlz+jc+6/D0jsi3ifpXyPEW7gVUajtIsKrku7C
4Y65K9gc7mVMLozJu8Yqx+ZvIjkhiH0Zk69vaIsT+ndMt8Bst7MQPKOP+x7KuTGq
0OAOVkFaeE3mgpd3FlwAmyVri/876G5KwJy4WPkrhxd7JUApwyU9HXPYxNNS4X+F
FUAQmKN2Osc3S+dGIaRs6oEFteCVfm2fksoXGy1ilgOX7cPLO5eNFfwsUUMDZkZ2
kLLA8KK5S/LNWmzpbpf1bfx8d/vi21MvisKY9u5LnDitrBuw90sbwyWvTNcGyJS+
sbKCT0u76o9PE+BfuDNETzujmud4ufxJbOgfBOk4sPUPKVqwEhL1xNip2yuaS59s
PWuKLNlFysUhcAn2PfEHhKF/uxqhNrYAzk6dgPt8n49s0CslG02q1NEmsrMZ4ojI
tiTMbSYgT7+5tFRxoCdlMXsm2TD06AHzs7yZ9U/6WvE99Qh6FMX6aVbhXbfzpoxU
XK0hEuPTNt3CsDahy1kKEQPt6AcZCX7Gic2jOJIQ3ZtSgNGeGew2wAIQfbWx5l22
Q5sLsOKVVC1wr1uaKQelgI8AkEFI+ttbL1eUBqOXeI9PVasKWTQGFSDI4g5vg+ro
Px914s97eq9b9D3OZtyqpPwXAlcefygY8j7/t6B/4tZDns4za8rW35LGFEhAKWQA
5J9yftQkW/fzpA5GFFPgZCTLg4F9/vs/5ngNNS2An4nJTS9mko+kl7GoZisN63Xj
5GJPxe5A0exb/7QKcjHmFodrcTPYArmdpzGyxd6sZsTzbUMwGGTzhnjgvNV0tHGU
liuBme6q6QVG6W6rAi24+pxqB2TFb5VPr4lZl9oCHgEwcwFxpbCYE0UZfMWtCzq9
QnBBC1FqpxanwxpwacIEcdJoA6V0a5tq3bZyl8uAejS9LZnNTt/XF9vXqtq4Ak+b
K8ffhm01EgBzvcFx3nh592POOkP27+kzKp2V4EJRE7qkq1Occ6C5noeto6CFiyiU
MZI83PD6FEOrkIw1r4dmh4u2uxgANdqf86432Jbmz6FcbrpBR021KHFG3roPOizF
RLOtGRwsAQu7/RCq690PFTKBgdh3rcF28gTJlv7NLOP1Iqs6p+NNZKwzs6Z+Xzs3
dw9CRsICeuyDQZB7lMKgv750Esi/ZOIe+3YLzzdbn6gxI2RxN/dmjFyAYjBbrH+U
zJ+esSIO5y4XtoLwiBBJ2DKE8zFSQmXH2DDXiRcCvNK+Us2lC7maUVc+eJceqtZW
3rqvme+5+5bnGY0pmx3G9CR4IereOyfHOjJpxZ+RxOTn7axdhq8hGAHVikw3QIbk
1YHlI4irGCTSLH2zvO+t8W8TljJbvSub7jZWUunjMWkPIx4snR9/u0tCyZHIpGwr
/z4lThKlf14KSCIjS603OKRGxdxB3juulPnOxs17Kq2aMeW/rgi8tzrUaioWlk6O
eUVe+q6vUhbgLFSihq+aa8+uFBSJv/4Cvd7nHf0BWE1mIW07mFeTDso9fZerEMxl
RV+MtD9D1DZSJhm5of7RldEXg/qBXPZingFDOnjeMkm5zKD0/NzIa4wnJrZbls7v
DMlKnRpfA/v7nl64OshDvUZ2F6QgaTh0s8UEkOjZFuCXzuHPuDaxQJLeVY+t4H9t
HeccESPG2CE6QxaS+YPEdj2ETBf6NJbaPbfzJhjNQNd2lTfjOzja8G8FjhcR2MYh
sGFWjCgpa5DhAfXXX0OMgDMzYwp8MtZYOIm6UIOFh6aL7XK6D5jegZAhIAG2VAmU
vSgCpyFA7CWLvhmgd4eIcgElzck1+CrnmZi6ezY0bHSqReTvlwxtYCDSK1aXpL9s
Dcwkh0N6tthbAfZVcVeEE3VlJ5UUJnmJe1E2CESVn6hzxuSLGZ44HB84E+fv2sJU
Fvbmnc9p0B9aRzMVp3w3S2K1cyBWZkwzLh0qoFi2H4o+HH7ThsQcThPDRGErn8vd
ViYJ0tz6XuGxFAOYo83VMFgfEf0KLJi/irPsNehqptmG8VEqU5KGWVqF1agycol1
bXQ/ai+GquGinFzJnyFVVdx1w7FlBDLdAwYkIm/hOYtAnOF0BnqYExpKVAidUCcT
J6FlBiUhSYzIZ0gNVvS7fc15/EdIpzAKA2R3PiL4rV3w4o0FSKDdGve6IBvgeNlQ
/fGwMeloIDLgJLuNA6tG19wlt0eRdvBkXAjCnhoVddini1WM8zvW6ufSRh6gaVSv
1uFP8D6rLFgpMODtx1Hs6kyy2E0xuj9SJzLNnQO/yMXIk6kEtd1kQ9NAPimgx7EG
j1iStbHQKpBWN76sOR7X04F+tkKtyYgjkO/FZB1iAFY/TPkAIBqz/ib808cUDmwg
LJ7IQBA99V9rLI/SSInPasmPy9ddy/M8kaKAAdQqlKOPH+mO1YcFrm/67gpLpaW0
8q++5gW5sFCSuOVDMTjemsPBoD3ikvr1TEhFH1ln53eG0h27miGfPtZcWMdqFlWG
FWbKh+2Uv3n+SVPf5CObFuQB+h3R5Pt5ifWxVA0L+EttS4tTw7iLWpNkar6GjXRm
mYa++E8A4Ioe5ALjF9eWG3tIume/8UbAlMDGYIzpwwROe+Mfi08vLHg31RVSgou3
ndeVxrEmVSGRvwgu7U76Gk36lAOuq0mpZ+tTq0JWsV+aHyFkeqiemRWyojK6exZX
6ZN8T41Cou+VQPFM6OYXxRRiHskgoO4KHOu+Ek4Lb4zb/ZlzJQKMeo42bWLzXfcn
Ohv+RhCAZZWy1cDMw/e3ku/g7906L/TPZAHINFi15UPJSf53q09xi0fkZvjEoUwc
Kj33Q1DUf6lKeDWs1EHsv9QhhHSKMQGcnYcnfo1/ZHXh5awnjB6q1ZWbgq0C0Vq3
UqzuCNcTd+EUHzeKPde4Jmo5hW+CM6CmqJl+i/U1HKaJCdS8/pPK5ISCzR+TDw24
ZT4wZE09oK06a7AAAmhF3rM+rB6hnIjIE1ChvYKE0FiEMN62DzjGMro+6POUb56P
w7HBnJm3SKN/R4u/T81Jr6OFRsqlIkOfkxk/FH9KrcieupqEoi0Jryt/URxICYPo
71qJBqvIbGnTxD1omzJe/iSMO3XhgNkUa2o4bySUkzGJrnadZRWI5C4SWhbiygZ/
eVW15lyeEq03KIDw4OtnIxdpu7hv1CVEGVQLerUQKeNn3q28/ncysXAros8UhaS9
ipmYrz2HcpUsl/e0VRf+/UicIfOcGRdqR0ZQQbn2KeB0pK3o5Y1L9cdAdHkoGsjk
ZE7Ug3l/3FIjxb1FsLUWOcJEVM5GTmAmnWYOdWs25pzXoytq97ZYZliOJ6vMvKn/
1RpGj2CkGJ3iMAtl9xYukidjhCeLlT0cPDacTJ0O4521pyrmCQMWj+01UGuowf1i
fXZcwWXkFSfFJl4iaZEO7kUQ+4XtCFeiw4qAD7+Ua0FST68OnuyxrrlMHGYM7ey0
8e3L/RaBuXdV1Rq6hj+ZtJeFrUvLAk5s8wTH0UF7IVQI2ImPUOP0RE3hHQiU/Hv4
12mgDLk9Rldj77fIRFSKh9uC9owoUSVAp3Xybj/i36gni/EMqhiOFtFtHhKUCJu0
Jbs/ZZNUA4421Gm3f+h81g7dkMQTv8wZyirbvLAuvZ0=
`protect END_PROTECTED
