`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nrcGYJGUTA66KM51CjteWfj14EKrdK+cmoF72P0JywuGfpaR84kAdmB9oBCuwPDx
CsGk9NPQ7Jn2K1MZV0VmN0/uEjd/qjizGegbbqkBFYxLaMk5J1k+67+DW0z9sRea
IE88d6w20S6ad+WsIPyCUyGc9fftg0sPSfQH06CP34Lp9kuyTgZm9pnMXLg5jDIB
Nq5hfJFoxps7ufXy0TJNh/vGnhHhI8w1WwfKNwMqQzrwaQUF8eCYUxhJX9VsbxH6
eYoLiZAO1VlOPgdiQbHmIGBRZ+8S/VxS15AOwU+zp8Mp53uSBlIrkIq7GM/LS9az
q8T8+O3+JGcka2Pf6/wsNRKrqnLH0TqN/nCqD0UduDefN1EBO48CdCRAP7C3X5Tc
QwGOipSzJJ2XafH4vqCHHhmcX3oO5eRXuF/Wu8CR/ogQdrCwGULXD82cNAOTqaK1
8d+ChRTuzaySsTpw+1ScUFKvYGh/wpGX8aybI4GkS+ukuMyplNI0XEcjCIyQIf6O
uOm3VyZuzFkO5iT+E1rNLiO8DiRpBa6yByvBqO2LUBEKXPQRgIxzs7D6qKGdezVp
EQ05xfZXDEKoKExKU87Seo15lVZ/6uGlMcwq4XjUVqXAs546QILsidUl9rpv8KKh
NPzuxxhF9kUIzmTDoZ+nEZtwsberKfPRDOQkqxqxUszO5TC4Ej4Nn836xvnoXckY
czXzkpv4XKYWXS7/TBsGmg==
`protect END_PROTECTED
