`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Otm4XPmVOgwT1Rtdz79DTWoc3KODOyOmNz3bqlPzXM/lYjUqSwLcEt889Kru9nkE
l172qEY7gNoFwJufjwWaEn01Z9NLZh4b8euwE6bB6F8dpw9+WZ3G79+QbVsjqfP9
1wNn8dHRgUgYhtcXaKLwQFkeZJoda4LY3ei2WqV0NyXsnQPFTAsMo/tw0Y8n/y70
5eeJ4U+IHA0x+p2VJ/bZdRJi03C0rshfZxmCSSJc2wBbEAZwJyEGlExtrhNCQO8f
hT/gLM+sKB5aUnFvSATuUg==
`protect END_PROTECTED
