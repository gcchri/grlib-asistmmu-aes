`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ZX5/IX9Wsty8bqaHGqLuLQ8OShidclZPfwv79ppPDD6JFIRxfcQUQsY8FV7UWvS
zyE3tCjKe8XZyKkniP1qpJlzhehktpLCyGt8WXMSn51OPO3q5qtIP2hYeebjlgH+
sX7IB4xG4DVYGFiHp+mNoZZKhr56deW1cmmjZiMYyDn9yhLlD3B0+HUf0LbN4WMk
pdiGBS5rjWRiWg2vrKPBHs4DNhXTsnEdVloH0AxqUXyIvyB9bMY8RUteH2KsT2G0
4RL5vZ8ZDOOHAgMkyYngdWt3HnYJyjOdPL+nYYNuF8supFw1/s2OhyGFJ7Q/NLUA
ifuhpRtJxXL6217KAzNsbrNzdgQiZkMQH2WrrwmsR9NVI6TUKW3D2pE9VUPoWAWD
NkDycadLEALpQalHULwn1Q==
`protect END_PROTECTED
