`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kEshxZNlVUOOjeDiiaE4mSrW0KO2sTWbkI/tA/+qmQokM3/U3cCNRK/K30mCJpDM
MKTadZ2qKNmYVJcSj4Wt+XY3PQcVhxwEbY4VRH1sqVKfhh/RP1JXEuXr2uNyavBD
EhCQWfyfgO2EhiWcPVmJ/EHvpZDOJlVmKY235w9ZdGEvyC+ynlIS/yGw+xC44tuU
DqNQN6sZcNwa/mFYv9EZ7XPKSIg8ax+kYTRRCb92gDhh1z5U0GvGLskC+MfHsn7o
vSmzq1DFaG9s40a5Ie5dAupBWhcaWMnQAd9ARJgFYv9/4TbbLznECdhYtrzV2eJY
VTOzR2dWoHkBVkV14HQYTyxUcuJuCeby3t3B39G2r5biVAHTcWW4K7Z8nWaQVR0W
WYi3t0L5hAFF2h2eNwkmYKlbTv7iD5kDV8n8FD5PYkI=
`protect END_PROTECTED
