`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cvpSIgHRvGGDYKkxRmQt4X/TQjz5hlVoP8wb58jCekzoJ1v2hEJXqGoPJsoJz8oL
Ixu+w34PjcIAJZsd3G7dWXF3kQacg2LYFeaghXM7HEv0lztQwKFMYHB8wJ9iOK0q
99kSIcGP3UImj2Eq4lMUgypBEjjrmxTyPchVlABPlhi9xaN+DHsWnc0dT7WIwjCO
PThzZS/khJ5ShgQ+qHLdPFTDqo0Wvj7Q6m4Lw0y6RW3u1s7yGXPZHLNeSVB3ikSP
aGQlS5Z7AGY/5jYqhxqVxobFt54sttetcDayyXY39/EPh0uV27eEbSK/ybNWPDJE
A9DoNF96V3a9I2dIAUKYyeh6QmY6z4gfwt/nbEyG+Jos0y3FyZtaFeXw3W7J4TKk
tsOBwbs5IEjm95Ywj4Gh5e1XG/SBRbWjxdpwjvm5LYAGg5DahNcoyPUDqQcf2LGx
l+6Mj5c3RlReGOMYDtxaSpVl78lZeOYp4iPtLi27mQj6EE/KuyFsIayH6/kNrGCa
mFR+B/JM6m2e/3uo6rMxABvQ4Y7Yw534ftmMnAxeu1SctDSpU4z5l+ukInUMY2uW
kzXLEwJIrDTlJhS8+3EegvXR4WhwbP1Ypu7Jsj8ZNdCzVbRbloZiwmGDgTOgMln2
3+2p5W9Cf4QjpP1EbzY00W8/1AkaeDaMnll4gkK2fE8NXC5ycSB2QqbrIkwadn54
GrG4P2lSCfmNNQ7WFmGF0MLiGUBfZsiZLXPG4zGVhePV6ZAX8W9LXlvr3cB4Vzc4
ZL1OM52n6izE8RqmA2kmNA==
`protect END_PROTECTED
