`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6VTCnVN5PFWZWnE7Tm16KDM3YqQcvrimhjjszvdULIQTf8X5VUsvxgafv5dSO9mf
bMkB9khwtbR2L7klnnccRFzGFroUYkNaPqa5HA4+rOncT+ltyNbj0X7GCQb3e5l8
idI9XCwuKLWc39druXkW1CifxtS4Dm53Ew8kIcwV5mznL8w6H3kD8Cvserb4noNb
h8a/sq0J+K3Hl5H3YYLnYPJlWmbllGLxHfgfkbuzsIgsRQ/Gjd/I1kZXAIgd4gAE
2bQ4kV7CMrkBtc3OQ9JU6n33J2B3I1EjYAqVguPvpvLG8YAWTBbTMWb3g3hriIlp
4/epfLXZohr3oFFbkmxW+b4AbCZ6GvLJKAfKRiZDMfP2v0ZrW9CHYDa1eBWYKj+6
FRFimY86c/a963+rwYADSlQ+/T2P2d5EvFsYxbYzrpsgBlSBpbFOYGSZcYyfgr+R
L9XoaQJATwAiNZ2HbqbFfnyW0EH4WEg6y+e3xFl36u3Th84Oj4S6tu7U6giWrLm3
SJdlfOuYx7UfsWfKSZHIINR5j1DErOnt4GghvjKw/+HdedXjUACgXsj6U1/gCYgd
eIejAgV6EldSC124gMmu0dN7VPyPfUlDZEMzyN/Fl4hOX3w7E7qw91r7eLYfr5/N
r2H9GM1yTKsBUBgA6UBMfQw6I8J/BFJyM8fNtXpg+TMCfXWdVr4nskFiul/Y6rzt
GxeTfLqQTtIeZrwKjKNxDDbwtO2xKUAo2IKQmJRoZL12e7NoOMZQzswSBXJ5C56L
t4qI5YnneO4Xud82gZrlGm+dkAmAIuxgQIj6AeUmubRDLf73NqDlDAmq1WunrVQ2
esoi2EfPHlcY72JVkpjsLj9vUZ0M6PEXlOdBJ0d8qYZun1uRObQtpyfu3f+bw6Lw
HMn025e8kHkNfZkuerKCoMT+cyWU2vT0fhyQvIm7gG+ClIZaovEwKlO2wtKKkyXj
e1WbAuTl2IwKx58mPyNUWQ2dWgQnfMZATblqbAxjHb3rLnOd8onnddPPudJuarI5
Svv8nLHzRUETT8L35YdWNOaDk5TlGDCT0/MgwgGUbPlejc7usLO0YOimKuE6a9q5
NwXxjtsXRoaIIbJxPs1+fYPSpkKDyOMj2PeFP8+wTKq1gb+TTxobgTIpcdKLb8vq
Gxp3FMxa2c/9ILuzEgFBxmW0/yKvirCF9nowOVVsjd3Z+MKLxSFgfv/MxGWWOELV
GBAHSXram7EasmFQtELitftCOwjAn6Kj0ukcBARuwNOQbi4qflauNGdL+uvL/E0Z
7EE92OS6Nb3uje1UdsWfQDS1hc+1fCGifEtHuQD9qCfLGAH2dZTzWJYkDdLnqKQe
2Uhd+WRHsRpPFoUUMhWGrchXQrixLTTbvEg0Iro/UjVp2xNIgOgBCppDqCtJxlJn
F+qaKCDg0onFwdbdosLv1qRPiCRaxrDM+YlPgLQHvqKoWqPTZxaR1Xv2vDetJ/aY
uivi60ZpgTqEm9vkPfYBVRAvAwffQOtVSiyifLF7Y54o88VsrOXq4692KsUzKfl9
hqNSVz/4p391pUXecgxPen9DUKjC4VL2y3f1X1ChLgSomwlyukVLZEIljlXnAXHT
yxZdGhOcrrHPL9JKcUH55Lr5QIAGBkYu2p0K0CtE86HYrL8YvH2taCSU3Lpb7bIn
UiPyOhUg7Ba8MSWFj3xkkRBwnkj7H1LQ+jU3i3MWoO/YMZ5eWs5bhRWQ7WhMPeeY
UcOnI7GlvzegI3zEznkVRdugngVZuUAHuSXpwRH+MuaMB0WEqn83+8jUXp8ZERtS
UtWBGNnrOyiTQWvQYZQh+881CTG4oCvAHqphT47FXwsvkgtfWLa6v4LXD5m4TPfj
4NRRruA/IJlA2KbWpG6MrZQi8kWYDyza9m7wlGJrUBCOhcXfplU1fYXvyXKil1nt
WzCsj5iMepWFamS9fBG8NwBjdCADIj5HO2LOWf0qYFu/crKItg2kpgpKAS9mSP2n
Gyl406Ko48gWplPsw8Pqbg2JE6jwoBosyoUrjR6H1V/5tgzh2u+zzO7R45bljXat
QrfPRuzfUJ27i5GKRgFYLfRmsLUZZ855A1fE4IHjrAf6PDoYEwk5XflR6hMlUJp/
TrdEHPAb9HuZR57La9Lp6cjwIcX+M4LXgM3iQb6hf2gd5KHtnsmM6b+ZLKjRJXFR
W7j9nNkjlZOsySN8vIeemJiHF0gwVzCuzoXnaTFgEp9LHDwFqIbB0vopB4oQZ3EL
kIMUng3DkhVsG6VnyksNq+mITsRwgyP3Wi/5JgXyU13TjuduSgnVEsYmxR8EDOFs
fKlQyHeNgZFKeAH0FwE5AOou8YsKgGK3ijymvwApPO6dPDGE2/DJm0xhXWhk7LOu
i5ebOjionrU4cU1raRruu+wKmd6vP5uYqLFpwzbIBxeS7R/QNgCXriV84KLNjMCq
MpRwI8uLrIHDQbymxZoVEc9F3WhCrJcWxaeNmXoG78P+URFLZXDMo4ADxyKO8BWL
l2oCkZEX/YzW3PVSYYdF+3BRuFslIcGuuaybnCmagg1INxIlwp3FhoF7SkBq0FwB
PfpO3MfjIvUkhFwsuQSsXcpBisyqS55dYohqvGQAVXcop9TIQkQkuro83IqZR/KL
`protect END_PROTECTED
