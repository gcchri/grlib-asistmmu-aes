`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SW6zDB0MTyVQAsaROsJOCSnYWpb6J4dYlnzsGWh6cKB0kvA3hV415oKryESA2uu3
2VRjYLGlg0gXrLL3tw4p5kT6FlhPIlCoQZlZMqJt7jDu3RnPXquXRQT77ZvzsNPo
V8+B55+sR0xoYF1hiRiWV8NwydWQ2GGZFxy65df4JuuQTybB++zUWVFYehH/jEyQ
ub1UwA2y3jMWCVZmG1K+mpUvVS1ueqZL0wmwYAy52ueEg5B/al5qgMczHAdQ0/s6
pzxSBpkGFrbSGVN+CVVbq9MYUC7W7E11tSHQc6V4ftHxnvRQB5sfqRFJwEXLuu6J
DcuYdHZRVXkxd3V1R8yPD7DDOPE/c+P9QbZuq1NSppl3EmpRpeNj+YRM4qIZTjJR
EpGw1EJVS3sj7b8cu5UsKMf35QOG/uR+H44gDuBRoygzb+VD0u+OPdAg4t44HZDz
rvh8uBuIWRRanKkJtuFUnNLEVb1vmltM/HCSMYgfyNWLQXeWuIw3f3pz82FPJFyo
F7PY9qrzVw8HZFDdh5WWsObTxyfPhYoQjd2axJW9VuFCQQc8RCVUsoqfAxcp5MRh
i/Fy5MRubBJoWJYYZooUM71G6DqUqW86jcvZgc0+aVu08aaGD76KXxqqNl/elXTX
EGcMr3G8cyJVY5Lo2x54uTM9oo9I1YyqJdYJjIy7Bqv6WgFKCyCxeIPgZw0siHvr
GiP7J7oJEa3jM2kPzOuo0M8RohuDESank+ScImnu88WllSsF7Ds2kpOb3XaqHyl4
HhYQi+AbcYCBI07w0fBrRBECPNQIARv0QexQwGckIl4z0xz5jjcMcqMOlt3K7VvV
sNRDwP6r/n6YZN4lPoILX/oAt8MCJ0zZP6KwkrWWC0E4mFwZALWqJ4Ax0JfoNUw/
XCkWOxnKSZyfa9AOq2ACYnJ6JV+d3HMP4MsjQvruxGcEf8/cjWC6Sm0tJv1bOHfF
0ePjCuatMsOmYTrEtxCUfOI9lLTLNKdEMhUpT0lEz2Dqy+T0kicoKgglGV5EQZJa
iIfQan3L8Vh7EGz4K+KLKKYbRxOWOlBO9v/TciaK8meSnJgn7J/byIXrQMYpM57i
lDIS9wDjXkGbpTJYhsjRYLFdGLJD0pMtccpHkaLexCcTeK43myoIHRZGA6qLgkP3
gmie3QE4C2CI34xoIyfBzyUZPWAs/7MPx5iIFU4LzY2V94PxpFj4ose0cPb6w4gA
DhqvX5np3REInS8TvWqmahANRL1jszmz69Oj5Q5piKJPzV36tJhZ/PYAgU0ZzzQ5
IRX27UWgbUaYh2LTdf+tDvSiLKq+2ur5WCVxRCNCHK9o7pQx1dYb/m6T+N728eni
kduzy2JyFVN9t35w8gTTmhMamg4MLnc3UwxkzJwbGOyd2wQ1cNmcFhwPjn3k1v9O
11oyM+xSjLb5w+/YVUxnquiYDxO/uiZIVNzlEFzDxRwPOLgb3x/bXyhz+h7L8/Kv
bMamr8yIUHHDjvPNv6daA0B2QkcERmlk1rmM83qVGQDHnc+mdYAmpihcOfcnW+0+
mxqnw4r/c8u0+jTZ15IKXQ4rzIW2KHZneXdTNi1bRD67m4Gq6w3f8XKxzcFHSiHR
zVxwxCYmajqN47o8upTMKsGJ42qKd8w44nyPUmBuFI8mAdBJIq6KFBBM95vhKFJZ
85Dipff/HoFjU0crznkS03odLewXV0HTTrcg0sW34Bxq/sk/ivZhahYAwy5+q7r/
stpM0O1c0oNCnhlToNaKbR+c6uTFBEF1TaPbgswTuKLldiGBGTgu+BsebtU6GfiF
OnZ6Q1EZLcHX9u7Jhydk/05S5ESPvA3ADiHQj8xrmTQk3SGVoWqyn2T5OcXzhany
OqssRi3RusNK5f5V1vCqkr7KquXSvDmgBxjCZtlSTTKYhM1BGnAZKx6YdYMFux8d
BWXJ/bTvN+Amc0fJx1rtXLf+BToalaVO0QpV6lCX5afWZ6b9BVMlTaEiod1qQ+yF
NaOINNABkEIVddG2Trk5+ZzMiunIO/q2yaeGYoITE/n4UDivZY/no48MbFRPtbAs
gPjjhbOrsfJVTl4Rc7X5qbX6FCEeM2WX2rqshVwIJI63Dvnzzx4yjsLNSZ94pt/R
D7knH69mnQ01LGEApft6RW87mOqkHQqF4WR7V7VVD1qRIMV9DonJHdGEA7mRV+mJ
AFiuab07asLKdJLgSxO+CN7k78nqkIZPolOR0/86/zD/HOZIlHBIZPkkwsrgShd7
8NrnFIaCHKz1X1pst5Ht6opc0RDaZMBHTH/Pus8U/8r8grr/xH4pSgh0Oz/rtGFZ
1UQTeTWGGYjYtFpy48qAJYva1ye3TnDWamxHZqkJQJERPoIfk3XMMCCiaZPEmXnm
ho0ngtAGk26+DZppB/mmvQpzmFn9OIS1E1BFQUsUbDRjd4um1d3urvCCv9D/vyjR
ur6ocjkPfWJyqrKEwvhqlLwK843C3fCIm5IeR9CR9pmjS4QJ8DNiraCnUcl6ChRb
zvsbQ1kDB2JOcvrZSRvcRCyHgwBdE1lSwCcPYQ4iOxk5HWMTVf5JJoCC5s3zOSBw
aqStq7VszbX7DYsI5dXt5CrrE9HGQx8sep8Ft1pgRVcT973yuUqYLzJBdGjiutAJ
uTssFWrabkb1X6EN/IPtmh9OOc0PbUqPjjlLJwOBYr/RVejXmi+KZTXsAsesakPw
BB+DIy8NmE4vw03SQ6jhet53jRWIBqVpKmHrMRACv+9R/y+YBNAJMeZ0O0iJZ2n4
XrdKMX7zqPvPZPk6/2VMgcY9VR7vfrWs1LsWF84lHx3VcrNfoYE3t4eqby0M8C6T
o+cRpeoztGPfd3U4akGr2Rgc8FhJBTUrIj4twhDrytUPRH9ivzbz6k9ZNmBaDS43
yh+MTRZT6dY/zZpfuZcx/18bmLab2ugZnk8FvMz3wX4KkI6CheF08HhQL4ne/z+s
qK+71Muj22He5EQM4tdlb7Bqv04+pOO9YlHQoR+fBVDdls8GAu/Z62MUc8vmsYoF
CTZHqEUIMJOrILtExB82jlguFSWj+ZlVpBbTccv1UxrmTlDvl1K/BmAgVTIFblUs
Y4tM6784LT12hvtD8uRQ3JxGeSSbnTFMyO4bde0JG8QcQlk+YIDHsrReFZ3l9Wiv
xHSHDpNAxxv6BRtV68HqPu2q+FkugU5ttc89p2SX0YJPQVTLHhOl9249DG7WrOgj
19wuNFaHGgtLrfiP2hH1TMzKZkwn4ie4Zb0OjbQcWY+8Z4waxdOygcRBI+71Fb3P
jnfCewZUPvJj/gpP6/9zrPlTZP+e0ug75407HlC+lk/hsFt48PF5IsAfocfqOwB1
7ga1qCohzbmFcjvzWUTOaklOSE49lMNxUVfvL1FFXLI4G5lh540D0tTSAoRV3xyu
10T/8Z7kL0Tx4lmjsLRqX/ZiirjqsUyDo0jAFBYn2HBM19LjvwZlk8NZpFXU9bjz
m41hguZa2jOee6efVXXDEhrIkqHd/BnezC3e+L27gClInd9lZKDQm4pY4TIgdt/U
D/7SIEKgdh1JlgOn81EgIfdmJM7lD5G8s8ByeVDqgV8Qac8YkmXeF4Oo9fd+JP+b
zBDcckCFHdfewntOd8QY9g+LbIwgALZICJUCBLmgixuI2o1eadmYws7VTB5bt3+y
5fBJEE4XFgpezR+0W348u3GKIyD6SFo0fPuI/01TUETT/RvMAtTpduHa7VZMrT6Y
cp6C5WO8nqW8SiaozgwllXjEp0IvLXRmcCq2xXLBLgEAVdbwJ+tUuh/Em7GF2s0Q
eIWX6YXi2SATlPMQ8PL3P3vmRAedm+uaKwChmN0GuxiwQF7PmYxI+tw6G+KsuTQA
G1EhIL6bNvOGZvfAGHYurbWc0/ou51rXZkLPvtRzeT97QCAp/cybRn1BBNXJiDfp
nlgVZriqZI7jl2X1DTp1bDvJTBG7J3FWKRftFBSa/+i7opt8lawnGZl5++fClbzj
kiMHNBx35Cndue/LN740VUyBW0oNcV7SW4sb0uX3dItE9NIQh9kjAkCuCqCBDKjI
ppQ0/k26kpppG1edOHBEyOpA++U+n7UHrz2rkvoVBY7FwQ6zo02kyyBpG97xLJKC
YFhb/nCfEUDx7Z84mivY258smVu9Rdo+cyWC2cUXQoIzppItRBYrRG0e4mJnfAm6
l5JhOIdb/qdxc8qUU+GznP5aa7iI9WjF8Q0jXNX85dJgMAKEbs6BFxTZzPW4dgUK
u2Je75T0pqp1DErBLJ1YLyKUNb/fAk65RDmskQUDDw+t8Qa/WS0p3Dl+c/Awzvge
EabcitXGcqUwzayA70aV3KKJUjWsIITlZz4QbFIP/wJs5j+L11orrb47dPVRo2yE
SMCBVz2XqMhf56CAlDYHFe+GidXt2jV7H76yyzdtcUJNe2iR14eRc2EGjqZavEHH
qFRVkNPt243HD3PNF9BTiepT9ZMktp5VEtTU1pM7DNN7U44AdUZJ1LZgWEGbHK9+
gJe3ILE0vOc1fGL/vb8tzonIKeSmVTwQQpWuN4cSAz1Tk+ZvLIVVJrB3kvUYfAoI
noy51Z0kM+4BeGrUeo89uvEQ2HyjXKbtbn+7DdrgvMwrJ5TsqCgzHUQxfwJFzbwY
8sNC6m6Xf6GIhJFhBwpyImDAzMz+pR3w1YQQH38mLrapUStXFb11Wm/BVX4R9MjE
9pUAKS6W9tbLTmP1DJjjG5UBJisl8zUoX0v19cKh7HVkp0OCP6oWDsFFbu9MKbL5
sOQ7eqfcl3d2M1oKW1oCHI2DKfhJoLd+4R61f/cuobuWo6CpN6rA70GTy9g0G2Mt
BNCLlzqdDsCpdhJdjpWpEGjmcx05bRTubyVJhypJAoB0HXW3s1RJxZn1kvSp5Z6Q
r7nFGaY1avSR0BLEHJO0/dDUK7QShHwvEe4qDj6txfY52abQPL5t0HzemKuMDi/Y
T2cYQhrtaDlf2+BtqD+3vRTeG68mOg7yE5tch3wlFH91S4XukC5Id7NuRFGB3XK/
fQlF65ZtwIxKXLE7PErFbWupghd6qWDplNl3Q9jbyeD2ueGw4H2a7f9T0E+/8vtK
KCDoqD3+gr+gTCqGiajko4Pt8waPnDWerMGNfkFjGIukTbDAPlWEnNv3pt39TW7H
pICUSsQK0HFNTk7zF0RxWwvO/HzTRTPkGZaeLkdPeX4X0yoVeD/jZf4zO6c7yeAw
4LQKMs+Gtokhph9PEUlWfqLzb2fWS7EiW9D3QoKaVyyYORlLRo4ViOfu/CBeg4yH
j4SM0MDBDI8pYiJhuk3cQeLOrzo7EaZ8/wWhNkguzGn19hj9KKsPerxyRrNuwdJO
TpcCCUUd41o78fMpPnTvDnPB6ALtGa2WbqAKvlZrodCSN6YCgsciLHYE4/M4fhJ0
T4eglmt+oqxNZIsV7t9sW1CHNvNRDtHIZnNAKfwAfbYtQXg16JyTdi49Qe/+ie9I
L7/quh10DzLJbok6HorSiXygcsMEqC7pLzFParkgT/6XB8tFhr1eI/Xa8yie8zBm
hlbMEYfath7p2xWfOEKqgZZVV8ZW9sgEhNMEnn5zypeQ+lfDmkWSRBfNHU+In4YJ
Rfb4scZ47i2KDD30FbXkPNcwHZT1yKbrYu4xVfK0rNVu/eZZbjJ5L/XFftC2jnkB
z69ArxQQ/V3mBikJ3tTqOsVKZQ2+iMaTSd0+1BCRy0HTwmmAiyq2Cy1NDZloGE6s
v6mXj6srPGp8WbD9aurY4NDqBI+LHISrt2m9eNn+82Hyz50Tjy8IH56iAlYLZHzL
n5Mq6AuFtDToPSYpb+b3zb/e9694f5Zu+n6C5aTcHdJd/HdxhHKkPR/zmc6vsDvg
wjNernkvw79jWqgO6M9morMoRQfFjbf3QCYLnrFjTwEnxEteqWfxYBJGI4fp3+AN
Fc9An8AX+NiZhf60V/x8+0EQHIVs1vGdDrDgvT+fNwSTmNtHc5IeKW/5FwXn26XA
BEpcgo5uFKs/HodLBFYvMj5VROjKaKme9XU/shFuZ89jyxfgOPwZLkCAkbKPX3Ef
j2AxYiQw8rjmXZrXG6T2aT5ntj9q8clclosBcPaAbJbWLGjCyD4TWu//vpsDrzw5
x8PY37JyVfDz2azs4M8ECnTFuZtdYhEytOpXJ9mEIdtf8L4E+L5rua2XKl6cXpP5
1/SPvmwgumSIIhTr2ATg13POiS4wqL1kifQbT6R5Ya18vDNJLh/su7MXih2WzfSa
UeumSWlT7sbf8ypPZH8bAfZcIYZBlOrQCYTe3EHXyEZNcfDe+BZoZ6kO5/pkt0sH
YC58ii+YNMJiT+ENaChoskwQ/rwPW2vMoQkq224OD7gAx7blR384pEx/+38o3Cnk
lnLWBNi9AchN9lZeNvRjgPcf5bvnxLaQRuiR7ud3ZRlZlgVD7utiXBALNV7orzoC
cop7tLOlMqu6WyZcc8j6rzjlpMzMjgw2y52XkaHEVIgUAzBXD/ghQCzjkxc5ljPO
X0Dg3PADzi86y5p0qvXdAd/2zSffnG5/6bO+1mCr0p5tfsTfV4YRzp8qmtKzNu9d
qLAtEZw5yrD1RbyCQE7D9oFE5m4Heo/U00T3b9Xmm6DD9EZGscunXNwK1Y7c8dV7
EXAxJO6eBQlAMdKNJNrlJ9iMja7kinag1wwRX7Cs7tdBEApTkz0eqikD1IyP/KrY
ZoKjMg1R+iu9O2bOGqO2Y1E5i19ZfrqTS093gICrD0aQua3bv93VhmO9GWlH1fKP
tq/XtxjZonu7EmzGevT/FGB6mNB/ZzPZi8TzF6yELNWk+Sa7ZSPXXBoNM3eoNcer
89Lp6kgtUnx6fN2RZ626LxCsPDNffR0FICPTTL05aQwrVs0hlZKZFVGyQVY52BNA
DBDI7uxLmf/QjXePFI8YnULwCoup4rqWZkbVJyknhRoHpViyoszmaD91AOmljU7g
RwiEvlh4+5YlevuDEwNagiZQYxUWyEXdazY2z19TLTrodNPO2WmjohkuMy6d705H
sJU5f2geX/T3QbjKgfYEvIdJ5UBN+Q1FkycMtKpleUGMtBV28m+NqX0OB3MH9NnI
xNAiGuJKbotVDSeWZZpzb70EPoSL/DhcSgXsyZc8oEJI0cVnQ2D5BHkkqCfgKINY
RNbk7CTATJU1vEAxswy0cqFQTJe84HHQAFEhAmvLtZi1dEjW0661r+R/IYjJRI+e
UB4Q7lKSrfTFlSCXC555kfB6+tOI/n7o677VWi0rfn6P3l/6XguMfFU6ITT183Cf
XBK66I1YaD4oTYn8zhlgDpxV6s0JYPa1U9npj44krlkXw7a5QxeXRH+OttA3PLWU
LEXgVvq5Hj1FN4FSlwk5JtAoFCoq5VudXuXKEVGANmKQ25ZebcRGkiyEc9axaiqa
D6uyNowxbrO0HMJDUmNyMxm2fxQcndtf6pZforGK6/BOFigZZJjEQETi30rTX1xQ
Deozx0fbq/zc8zrtQbp/xTyEH1/OoyncQdMP5sh/4/7g5WtCtS1X7jeQOrqVbLh+
xYkl2YHQFXudecGV8EgxqbuckQg0XsBxzbD81eqr/av/xUYL9GN14sUuzEVWjwm6
zo4sftAY7o9XbVo5V7Ou7HLSriBpxCimNJC58106TyJl13WidYLQ8ICbqQyGi7Fh
HZ7a/zfhiMDnSatCTN57g8Psqu36GD4t/0HTV8W6VCDee4RJ0+7pZs7RnsnzOzB9
mNSAOOL5SxcwTKunCEBYX4UF5A/8oOG0BGEr+LxlFHgqDvcfngU+OUFxdb4IHh/t
IbRlYVg+ghKbSNpTfnvzmfJ0hcFsUk7PzSsorj8oudbnmokR5slT4n/AGIeBIFb8
ZP3xbyyey52ox5kDtjWZSj1IPzYcExo3lnmJkJ0y29vT8W/MhKS7duwnAHsLN7QT
mSuKHVVoO8jYj2FDVtSdK8VfxjQDG1+y0WFacIsZBnO/M8/1Kih4DSmHvNcDXHc0
veoNiISscbzxYYww+2drPVRaByloQyRON48IK4D8G2hLUtEGnDu7z5h/l4k7kbV3
wdm1pNiY8etDGmrvx/sES2bYb6fMs5NLBrfTLRET0on+ItozWwMmVQRqMa9VjGWg
m8HcCYqWw1jZ3K42iJj7Lg9aYnbqlqjbgoAs25zP5qVeHdLmdpCBI2e0IuURPF4L
5CF03JmIcCnPazJ+TMa5tZs/iH1hd/8/hM/WzNYQT9J0hnJ7AfxFWOFUS2lyi4rp
YYrlbTqf0+Rz/netWmV7o48JbDNiQA/LsXedDEOBCyKriIeaul6e4vQo98Cstvoq
a5I1GSSFReJ44SZuk4B+KkNK/N1ULvSJUfGD4PqIQcKDgtRNpOBPBLf1YYuG2yDA
u3EWwCxsJUmQfxKOu2eLN2dQkZ13YrershznrdLvBXvY1ukgEFD4BjQWaoz9kkU/
SGCGEhVjCw3YHOTrT6JE/+374D1P0pBVO+du/WVdCosyBcosVLKcVwMrWCI2V6FZ
PamtsnPpT2VEn0M6IkWQ6N1WspXTWJyjN6d5E4Zmrm1Kk7Br/2MLAvnZgPPtkoRM
8HH8SZ9DD1DqqX1A61+cu1PqbZPhg2gfdIGa9aqIQafG3H/sNN6cD8GvicfpgeEn
MsYhfnCDGSI0P7Kv8PDIomQcO7ug/Ty0/bcuLesyuKJy78aH5wOBZUUSGhuf/raN
uWwQUhTwC26Xz3x+CtU8/cmxLY+xNor65fw0e0jWYaPIzuOdxCMbz0KB06GOJgq2
WJ4LWNmvg+aRD3uZnYsCcq4u34BmZsp9KKAbfwCYkZCCRZqm9t9qp+cOMP6RoGav
vHpWj1B7S+MWJD6yyYzf/bgvx6FicZKTwI24bhNwQduUIYY1qTxhUWp5sq+bMXmG
xOSEKXr/HQg2Yt0b37EXqBTl61LCDXz2oxt1l3FJyl7ktjyJFStIMa5nWA00ILTh
aJbnELv9oQ9ZnPJlDyVyERtealJTxTpaCkvdqcH9Ge61sHLJbhUmedurHTNk2tg6
JefcEGCYmVo5tt91NKS6ILVZgTrNKyhdICxeWkuXXNebOCLQysAoTauXJxYGCOuB
RYKULQ8aSEWOc/KBAHFBvdbEsi+twoEL+rLSkNDVXLRAevulpMW8t90r7H6cfvHc
P31XQ0zryucw9Y7VOMWb/vmnHDk3OLaoKWT3jDbLXcTuQTAasbCXILt5j5AdePqD
UzxIDKsrySO0YjQPJBkzV7fX84rpIWvb6k4rX8QJm6LjnEewBLgJ+GTysKtojUeJ
KxgdvkvFRAzYjsqYkNf9s9Zb66DX5NYM61V+izaaoa68ymlxNR/O35SqDaa/afhO
WMzxn7E5rN+nA6QpmrTujMAhRdVM4hammVqcCfxSOqeXKyEOR7+ncI74me97teaF
pJqpUWwj2pU4UQOcbH/GbfGupy5jq8kCZW/4sM1u2KBrUohpv2po2cNqfVX2gXm7
Nsk0515EFx0X5SHfGVUOs54EEXVycM6ZtAWSH9hJn++ZFBuLE8Lz5t1MeTgtO+je
GDYvU29pPUVbEHAq66HKuoq/BGZDGdc6RW4HTmne/I9y6ye51QBeKuSl9NzpZzuN
kk69xLbVqItIBfXyfA9/2gJNURDO+gEhVtnr/v0GT99Vp8ltTvWRACZr8j/dhfXM
bNU4E8YG4+1F4hW2lg9Kn8MwEUtVV7fsSxbzs6J/PQEgD50fN3s/BCaDvV5l8HcK
ENaD80NfzVTUPtJ1AI+Y5l/xJAemu0mEdKym7GQSOkBC9G2KtR2KRXWhR7/ViqvY
FTYholk4HAeBjGQ3TtDJaPxaFb4EaZ2LuZJQauSfRugchfR7kkAwyMBnhDe5SLQ+
h4Sg2uY2n4k4ygZLEilhL06XQptiSKwuwmyXwLUjf2yLz4wVMFjA9+BjuTlQ1Z2g
vhM4+y/aVyFvPfmOQE6YBoK74H3EKbPwUNhKB9mIId9FyI9XRHRgXDU6P2P/vl1+
bZDjsxFhLvZaW9r/NZc/qQKy+gCBJF+a2kdu7T4kNoDKw0Y+9fh7X+BjJ1xIx3Fp
1OPLwPweBr4ludcHadRNGWV5nFrqI5AxqRfO/lP2k8AVhSMBgCGrqY9PnOpuZixu
xC/Nz1YghXLxtkmVFNGSZNUa8HTShQoqxRxRnahsCgQDcoyGi6GAaKv/ehLe65Ca
Gss9XNwLE1dNBd24kfs7ff03qXRQ/HqunDMhlAXMRHh/C4RYP21Nm5Z7Q7r/HsJH
qaCnfcOiMkRcRp9+I3faewu4FXSUPCYfDe8bol62shtF6bRtVha3yc6nJ0o3PQG6
NMibLb1y16jmdQUs3CquTT5SQVJQp+B+jbkKwXi+2LaEXdlob3hfXCnd9ySEcH62
oKPuEA8MdyBfKG/HaABDmhF/cFlIOyqczVKzuCFiea7m11U/R/4HmJWbCEOjOWOk
Fwx042KBkf0ox3eFGqkPEmYA8HqrqlFqmwyMkNwoGJ6jPM8H8cjs+r4OHMmFeGPF
3ZtzF8llo3X17bMeQKxDEiOnNTIRJLbZKlTCAAaMl1Q5tyFGalJqk2QSPZ6IAPDw
A/h63dPiHc8NYNzPjYY2tJzFmMYvm6wFB2HYZrksvItMBnRqkvvJnZ8N743IUz42
lLeyjsf3+DVxNOgDvSH2GH+UVZvjnSI8ERXIJRKuS1QtVB+EJdt2BFY98Jpsibz+
L3DmLR1KrGSONE9bT0je73f09vW2sAQjE/eGMo31hAsP3242CpTFxMKI7JgdAGXq
zp2Ihdav/7ja3cr5/Dr1GfMoixXeVjk2UNvyejoHmBbZopX6N3r2dsAcT6PBCM9k
yQHZ9o2JjQRww7bFCi8LwwM3pJ60HWudinKV0OYaGFmSo70qmVbAbzNwuMD3LVsK
N8gRHyidVE2V0jJEhVPDzASUH1xi76J1mvDvf29sGDncnnWBnDMfCFHQiqXKMk0K
n/Wy67WK9nOfpqUkWon3Z/7IHsWldutozaeSf9ZsEuX4nGhpYBZZk3ZYyu/33n24
Y0nV+sEXOUjwe/jsBmNJqTTfbEUta8xyzFOZAwbKgEvsHdFFBMSwe2HgUXGCdaJx
G+6BinLov+a/L++o/R6maHa1e8R5GcLihoDEMepD4OGiehSDRiq/gtOym2fv2N3L
rmtHrpd/GvlG6vDQbiM2hYRnzwhBYi6zUpsP+ULjIhpuH9dfrxl4yeBHhq8iJfEm
6m7ImbXT+XU9wQz9B59e3H8xSoYxLdcJLJDE93RomnIPVaoCBKFV+Uat5HNP/bXY
tbF+s6W/o15vyI9E48G5wq93soHf7KKgjoQ80Lfy+xirnhZY0gHWpxG8+bn28Yjx
dmJfdSYsksumtMOgF4OSsy3+9+GcRbh2u4b7sRC3YgEEEYwxpwqLxmJOt1rS9xgs
wsgt3h8Ppt7hxWLGiAkJiNW5qCXFWzWULYJjNNp2H6ESuvgeMqa9ybobSa38AYSt
vs9GU1zQcGpeU6UcCV5eGS3VeJP3V+h0ZQcnNgxkrrXydtTK75ZjcBFOuIbTULUf
x+k7CXGzMdLF4+Apy+YUoaLAjLGoFFch+D4VgUeiaRcg54Nl4I9ysEHqaFdwg1nj
g/T/YPHkKtfiH48Fg+xDhy4PNysH5BMxAUG1WLDNNcrgANERKQs3IPBswpHxfMvt
Ext8yQfvvAaitjL3f3+n8c4V18ZTBQQ+m/5eURFUmTKvNy27l8vEDgK0Rz7dUcxA
0nH16Anu3aY0n/4s6owaGx3fz6Bud1GnPgZlVnIzz7pmshgRoZk+GM/eSX5Bspxc
oBLQ2nkMYS1BWZ4FnTCsIaWc/D9hMOQMP+6WwfeqPuUpIaruLbeQjVRldmyNS2jk
0hqEnurAwqFePDRei76kg/mb2ZFwCUJaNVXuBLaFwrYMXFqN462hrO14sX4yCqFU
31Auz/IX8mtvKTZaeb4o5Ap029EWStSNqMCtreemAVKkMpObQe6BZlawQ4siovaN
6RY2UMNaEKz0aO0l2kWlsuwWrReUnrIWIafBf5CvQgHsEwyJBSh4LYb3Yyy27qNj
2w/7MV+9i9TD1R+DqDP6aXUcbjZEzH3VlKGYeCg1Y4HQDQbLMrY1lWqnlVnfkEAk
XQsDt4Y4Jtmqn+Q+MH5CzPeUBaH9TNvsXz6aWkLtNZ5ElAlm8A6EKrH5+BY4opLG
wnR+uJzqxdM7EFm5NP6bi50LxnrBb11xmnxgG3nVuIp6XlEbIrPeQ9Q/kXZ4zfjG
oj8gE0zOFVKPxlsD+zaY97nD7NkRziSTFY2CoXozfYOtn/MxSXgZ7Bh1mj+/DMw1
BgfZmPBfmUUHVm2dnZQMe42ngyIggrgIkX8DEdBbdnbFsksprAINTIKtYz+u9txb
OvQrBH5TphxmI4CRlfcGxyOzdfrSkGXxazKu/k6Q/F+nKEbd/zRwn9fyHtWUxE3+
bV97d65ZE3fplYa3yTgiMO+j7MBOfl1VZk+DPvXb4OmO6CmyCD6pZ37VXonc8Fvr
3oOoXxg2KP1gQn5d1bY0s1WH51M0CK6FUWhDyoxs3S93FoIwFGxzDmYBwMtETPsO
QIb4m4lV12sgfGDk5q2u2OTpp/q3tL/YqKFgNv9gaFrZroT9mokJ8PCHa04oQDCW
/kTnDYaSGpYBkqwylrD04AKIIec8EPEr7GEBAri5ejYocYx1HOsqbtpIFf2vfm06
xYZMdK7XEWeNuercupjLS7lQIkFPQhzGJqxN/kvEBDUVSW4B6H8zUR+w5bFTrIwO
vrg4ZSJwynjiJOMec+W39VgoCefNyGN1yOeX0XMShi2b/2p1A2cyPMxRblvuJRLG
HEEzARH4vBEhwJNbj10S+8QLb17F0BRHH5j7YHBhucaKyEHjoC1mXXj9ZiLLvlb5
6OmGO63vfj4dfzVdEFT0G1vEyuXpw24GQagGcUF9lnzftiIN71Kh5W5sPwNoez96
bXNUELFTEaqM4OHMruEnAILoTSQH2RBrel+Wckr3TvmgnI5ZIYC4Js9Qwa+UWFdC
f2TCFAP5UtimyTL9xwJmnMwwuK7scBftZlGVH97ItqRwJGieTHdmtq9xhlVbhRfM
jxNDlUiTmuXZsHY0lTQEV0w9FPxujVhIIJYB+v/ZQ7FCZLXkqOxDk60tGqynE3IY
BPW8hd2lF/h/H8Eu55MkJsyJJQQqI2QRLo40NVb4rX60wSKYuBdaHa/iQ0VVrOfX
k57VzY9A7PGE5bgvQKWvF4x6ETlMkZoLh/ZrASbcjmylBXzjNabPQE0xMJer+BVL
Zgk5Pnb3skf4SnqXNZfi5DilePwQSGfxzKddMU1MtFN4NnL15f/EmP8z/GPYSdig
VUpQBtCeGGGyMknTnMJc098884CFG91qjPoyf/3kLJndVZmerszUj7Mi8NEuQyhL
oDNguxQonQt+Nvrk93oOQxEHxpOgzTuxWBvnGFhIeagh5h7DFpPpCPXQ0+hVV8uv
eBDH0ugzEW5m70bFlwp05R1fbN23/+F+SweL3IbkKJ3c6fvT/Fwc67SPzgYB83o1
/ug8Blv2EcAUJeujMXvdgmsWC0QHNu9nAAmDNWtGmnuf35wb0zMkwhxD8b8mw+f6
/R0I9OmuEN6+cQ2QhYV+x6bpW4psDBQNQ2SL/OpL/8r8O3u12rtLW9pzDu/kT1w4
XhHDx34FwtcA6POQArYI/8+fdxtnVwlxFccnNhvcFANA1P1viO+HXIOj2LdQtGDG
jG5KMmIXzGdN2WC0N53ff+jo6ZJF1KiHiEBGkeIFoF4VTvNQHl97mzBU1mKfPJNl
wljJ1+ABcRTcTzB8XPA6kSuh5/i9+ihei7z+jZq88dnLFVAeU6vA8Zhdp75unne6
Vx50yEd9MWq1cVuHaUZEmznj87zxepKg61MlQK9Govc1FuCo1jEckB38efpK8nO8
/xAHMWhJfqAsfO0G5J5G0+hLhTpmvHdDTxWjet58mSYfYta75TqbaL7LrifYRa/X
qrSXZXIUQp5hYv8Ja7Y98K0R1/JeuM5VMlH9S0I2nRqzdviUkSUFzaEfseObbM0f
IT19CvBbctxLujQHG/Jw61PWwnPCxwQ1RUd3eSjbGZ9Gref5PcUESn8edK20qk24
0KHM2ojMtIu6XnebQvEgLso88n3TxNt5qjDzK5NuXW9pEzp2X6XdIOcjMK9l93ra
sG1fYN84AwEeLtkg5LEcST+1prOBJzj9S3h8NMhd8uwn6aXBTIohJzBlu270GdlZ
SievBj1QLw70TZXQRoEvpwzEpYwzPrige2mJdzKbR4TUJByD3+otN2br2QnWrfQw
gHDuG56kQX56iEeUu1JPE5tdjh5ovNXK3byMa5/iN+28NlSrCNq6y31ti1wlUKfh
Qwgx+JFkhMk6xSz7umLI+/G8/442f0Yu8HUBH0KuWSrfjDaMsrwbtQlKMm950q0u
AYdzYAd+IKER0f4qAkYgvXVFqgfFTW2MeRwBE85l29BBHfwcRwTB6XVvNLVISh9M
JjDV+Uz/l2MPzAsGKX7vClf8xJg+hP5u1Gti3JawkOtx3bjeMtCUp37QNJ9hRgeQ
5TChMrUSZBLbJK5BSKEISUtXSgmlHskms6X3WHM/0HvfoQoMxYQ83DiBr1zbSEcu
XPNN1BshDTINn+n/M48SyjsnP6gBh67wL9iIVTNKJWUTNzMvc8q7JwdyBj0jlIO4
Ostbe9x0FeDg/f0pTSU3MNOZtMLaunJkQGcwQj7u2b2vwsyNOcvx2P+n5pmGFrRH
8TpKxZpdmPO7sH83ektQRMes10z0SNBgNvY6scTVvVETlYGdFrCWF+ZNe+qUAoXB
dJGYOdwIIrGelv4Nq+9WZOBWjxdb7Po6GMasykxgGyP+vXgZo5a+NPu0Nujp69av
D1t7Ge5j8AdWn7HRJECsVg5WBbmqj8Ul2UNZOTKcI8Wrj71+0OkvYTOYMOpt+drT
5xaFRPfngrnAzisagJa0UqBuccWFMCj4517o83ryCT/I8PdfzxNmdbyfXMkjbGKB
h65jhTw1med1d5VBY9lAVOwhKCGa/Zu0ZiXVA0MIfxFnxKCqFvltGV9ACEsjP6FX
TZIwML25GZO5DMpzX2hMQTvF2ykNUGF3kdMa89RlIyzBdOlYGzWfZwo5f+FkSo4b
0bU52GvD4i3zXFPqKlVEGi3r2mRU2vR/dpIz4GYu9ZzeCLnMVA5KW07vHi24TywZ
S6u+hLMxLdclIXIrKVnmT+z1jeAUFw1EHgcASydhWQsYvNmCWTzYq6Tzv3S/Bwm/
Vdn+unSawPp+ZmyKVmtEe3WrBXp4dirMP+wGq1oEgZzMijwqN/K9NHKITWoilLYg
X8amjG9vV/u1Qs6Q+GEIx1ucDnQ0isA8rXdPigwThQc+ZSl57u8UM+QlzYrszjDw
0ImY4imKXGFxk3YLX5WFFJq8fprDVuaSx4ocXYIj1wGduCgcjgfoA5ODrY65miPH
Ont93GHMb5VMhlQqIjyD9MCs64mU0uxw97T2SuKDZhvOk4NtcaeCuUrOVX82hrAH
DwJiM0L4VLnCFJFBiI2ElrNcYfbnhLPtVbd2QG+y3mHbHtNo2aO/GOg1yTxBe6hj
qHK6r7nZ1409VDF5u6DjuhVlQNETrSxoRULh2fCNMN5/063gX1eg7LrCREH3I1fn
z4ry6uGkpMwpWo5XAa3GgPZOupuFpFluB3SSu7i9oDX0kRTEJjy5vguHlxyCsz9F
lxF2dOGG74SSzUc+jdESwAwbPHC50gFUuZoLpiXfJ/rrWCsc8XdiFbYCOhAW0b5A
W1lKVWhmX/ClB+GrsISrHOFEqoZ46w2MtG8E1b9YDSC5L4UO6PSvbmwoV0ASq/E4
iHRkNn/UC5H64V/Gd4O2w9xonflj7KK1WcW7ns9KY5E2AjpgvltfVQZV9aFUvG+V
XeKydJhbXq722CAKzs99n7RLUvy/UXWj1xbeQvaaJZaZn8Fq2JJyUdYl62swBXpf
ccluHQv4IYOlX0IgYUJUW2/KW4Y8p7Kqg65dl3ZoF8+GmUSsDPXHqwS5nz/hZVeQ
it8hnew72H7INYKFjNuxWcsXEQFByVXhzI8qJ42YYkQ0LaqjkTDvYfH5KuwWi3zu
0YmdhvLDJ2RBJKJALWOQbYlOSLryAstluoVf8wn/HBCzNnA4xCGtlLP3RDV//VjQ
HZiWgvm+rya9ycJ7fSwx1J16xTtmTsmxrb2j7lzL2sud1ivYgfqaTNw4Ep0s9Qqh
8E1zd1USKEKRk1unaGr+QORglRTlMBYVRsZT+rnB9s97JWdzlQ5a5sVwKBamob9u
DaDydMvgD0b35iUIzQigw8uLkkMFY8oyz/wDFc0gsK+F0X3UR4lH9d+3bO9JR9rG
yglSYcxeALT54PNBmChzNwwgzu6KTWQw/yo1xLnx12AcS+C3j+92t41RERmbK1Ra
TOq+wE4K5htqVqiBaf1B0/7cwQDRjGdVevoEU6KzNHRzE136TtQfk3PMD8Fyxt5k
G1P+cbYfDW4R/xUESBqez+GZKVVhywh+f+LRBHADPT8JEuc4RjqtIern3Z76aI9L
mU6095VzT4vZ2Rk8c2juAuLstZ+XyOrGQaDW/g0823kyyublkl+Fs/H967wfkv62
sRlHVcjOSiOYVmL3zujg26lcB1GmR0FWRTjZY3OJpFeabjZIdCMBOCd2tlX992r7
iyZmklgRM6iOb7FqO07miyuoxtF+ldlW+rZHYkzf+0cgzWkEXMEqlnX+6213Q4fZ
DgAmKeuDCev5h/aN9XG8IHj2X1TSMdwHl8Q1WvmVSeH5Uf4O4VQH47B8qJzzup/W
1voQ8EMxkfVqT6uL8niB7AJgNP6x8gxLT5KRL6n+9B7dbLVyGNac1mtFQjYtly3y
PaDwGr6eGq1vLPjU0TXL0+ryt8Mi6Y7uGnJgK13o1YpYczhuNbCU5AaWeK+lXYkG
YM9CUqjpbhOMIKwShlpr7Ru8ynqOSOFrQnmHpDNLt9nutN9pBBxCaBsu6HMbS9h1
GWOE4Z65+xNyp3PCJW38pBWz94T7+b0QGU/PXLQrNvgZo7HG+hc5v08pgUTi3yF3
PWt0b6h2dnM1h0bAm0+PL1FzvyAnR6goiE5tDQWYrrmW1Te1Bg5+4W3gwSNmCBo/
jGj+Yl9yqzhEYOKs16AfEzlR92+zIFbwvaX9JMotxUUge9k2ap8JRW9Bc8k/xtPd
enGVcl9UTDCaBr8JX1W+By2x1iFUFMNW3ByxB1Efd/SAFxB5ft0vQ8bc6oODB0RF
aQIm5CTmzXiR1+4GJ9i3JSzOot81LeMnn2xLtIBCIp3iNkQ7Oh2Sjl3/tObG2nJ8
G/GDekLexibHJZFb64043Pn9naArMBHRlBkZhuvnW9o2h6vUS4E7ZmZvZ35ACpmo
WtRX5NCQrR/M2pAsFzKPW7TgpCMrhLVDOSDn49F8MZf41TJjhsS7nMHk3pKu3vYp
M4CoZGlI63GgSLSz/mE5rsVxP9SIBQJ5LfwMZ6EFD7ugYH5XoxVWQr6bmTSiUdgl
4V2x9oJHZrnBUmd5UHePY6T8sdW/5/y5W550vT8xOBenneXzQmp0jEQDwjvP78E9
8iph2zFKZTf113LtuO6FyMvgMvf1xa6b+Y+AHmOGLgcZVC+Qnd6/zcv5SVlFJ6jM
2GUxS3TfPr7OwAcUU+F/bp6rqEexZGBiBCRpbWxz7rFGHj0EPZvMAYUIECYCEjzX
dJWfAesf10/tqf0D5+NpiMMtdXiRYXR3BL5MUFYLpWQZSaeTJA8EjMoJkqDHxjle
RYM3m0arJqbedHkoAjfXLIdChXCG+4CjHSNf/PeMeaZN0yVWUiEYrRBqpnS1Z3mu
M1RrIJiK0AJG7zadg66Zm45qUK0TbQKYPp8sQ6nmgtpgVE9qXtdXI+WFLs7UhMyF
4XoFxJKmxW0+c3Ipw4bwWaqBDe9O4Wd4R8tXpvRfftkI9NwMSGRLq/WeFnkWGqXX
QUGrcv6N4Fc+Xmk9uvGsepBMEKednRbXItXBoVkXpuCyjxFtNn9z4U72cKRxJYTO
uNbkT80WACkBf5naLvDVbwMcDFpL63MXn00G8nQvLjjcpYvVx5/AfqTjUtkWLCW6
nT3Lj/FJ2Bh9wFattfrHe9xA2KOIdaMqB8w3Eav1IG4jjCPkyGumb1/gGkty/RIy
LrXaHoer4YxIhoLQ8qH9EVImwIQyGuem1R2pwJb/VIovZroqavj4IRD9Wl2gp/tm
Z4nTnuyotLo/X2HMDMEM6yhKpo8EVPbFmQFXZLn/F2nTvDR/eAdBx2VSxrym5Soq
34VvevjhZ1OmAkcfSjl3/TWyqksbi9MAKUhUPF8BeLXV72WIUDVTsZMgzV46Fb2O
mAyrWhQy5uTo/rueSIz5SHZpA996AphL8f1rIOZkDPY4Eu+pFU69CvDT5kkdFzNu
x0A7KkqiMj3KLukX7fBo8KxATRisraKRAuu+Q1CihGbXGeS9YwQHsnDZTqcnUxkD
vg+cZMRVcwRWxo1vXHC56ChZ+ZrWF/U5jI0D8yAM4z+PzVmzPqYdCuIy5B2czZNo
UPQbckzG1K5ZEqXmdxgJcsfQtIGtPvtBaEd+CdyGTmazFXINkGPdZZk5TFdHjzVr
feUExQuJ2fDT02iBrQkssBqi8X5tU4WoBzGUvzBgf9lts5JB9fjVt8r2OAHt1PLq
7B98D4TiSCtKKf+lAbSacFD8AeptlGwAEyCTGZvl4+CdTE6cBZO2tNAX/HkEwzlc
IhW392h6BKJdkhz7rdVRWn97us4YFO/aniFSAHv1j2ddWRDMgVwjT+YbDmqfkJGU
A5AbXeSVyaz32M8HjV+Np6XgSrJC4JhaQVc/6wYL+7BQ5lil7icuJS3RS0QJXzBW
hFCUFUevmNP5az8EnXVb8bahBOwukIWLXczCGFforkGi3WtPQjp8Ld0dSN9MOfFS
MfnUW2PDrLk6KDtCt5u584W9/nUPDTmKhwty9eI52eE+ZvUzVchZZiXmaNDOElze
MZzr/sDgAa+vLRSwQEXJlkNwM9JgLOiQ1+oyqiy7ACmhoKo2mVsTxGh07qkRvjM0
sKbBPF8rx0H5ar7AqW0gsJg11dqkXmIRqF95eeDJm93p1LwUtT4xuOddU5f+LrHP
YxzkItWpVvZLuY25DUul6u9zDaDpKVM+MUvpBoeVIi+61rIOyM68RlfEW5oS2w+n
jHzCBeNQHIrai1XfqMaSioYDfqVx3Q45yyK05hNGj0BR/BJO5PjiKIODX3NO7scd
l8VquZo8mzMVgN8DIc4qqoyVeRdhQSlN1GQrvVEmmpNgR7/ptnNvH/whvFATdps+
BxfkMWwsrFDn1VCYI8fm4PlNOEmkWs6G+/TVodTG2aIDgXLQcCg0Vav/pnfW/vJk
rVxWvuc3e6/0t+17Q9jA/YUoL+h7d2oJ2L6I9FB1YQygaQrLFt66bT2EPAZq10nY
s6PxhuXi6Yo1ViDOOj594XuvF5v3vZINEMsROZaoben8SWSdMYMuodUXjDxCs0Ck
51clK4omX3jdJxlNiuK7+X2MCnIE7BmhdIElGxQXtFfA0wI5W6h06IF/kFG06MNs
qoqOKpkZ4/JaIh0gMDdWoiQqHGbSC3PHb7i/LLqu7Sripp2jjicLrfk5SEwlrLEa
rk5ElReeBC27czjqQIbTHr4IEPaWDH4yq0v5teH92fiqvor1kha42gAEOgsTFw1u
8I3oKMvIGHyM2zBxtnsqjKHrMZaPB5mKuzyULepgI+3sP0Y30dmLtJL6vSBBM1Ko
NGsqLRXultVnl6j+PMbAv1md6HZrdKU7hLCYXIqUfUF5yC1TuvaZvo/7UcT5eIAl
f8iUufXeSeYA1i9sq+kbgbmCWvqYJBlwf5SWlTr1q8hdIvi7BiFlnwI4hwPaYMwJ
DNMDJEXen23EXT6C9opeEoHfMrykuauINdAH7Kl7Uf7vnsntX50NUmmkYAXBpctA
NpJsV9TfbVxao7+vLQ1bVYm8ov7YizCKjcwuWCwK/9UTul8ELEXKn61R1OaO0iNF
EJDqNYK/5Hpj5qOleDgWuRrBgxrYTCRhuSea6zayqq8inWQx6Ndab7o3AOhhaAjv
pDS/chhPdY/6/jjVkYJC4GCwKu/NPi5X/XsC/90tJVp4tTc1Y4vdSSkpqw0Lvfdf
AK+IKUf6i4V3TLVwU1wVuGUOVhg6GIDCj9gkgci+7+2W8wA3DZqVcu/+W12babNS
EfwjGNUDKzwRSPCa6KJK6hs/ROJ+8o4n614vY0jOyk2UxhEWRH/zY5o0ia36dZp0
Du9Kaf6pmqDacxKPQocTOyEJbttKpYKK1HeCWIcCoN7u29cvCnnzytrY2mPtd1qv
KZJYCtV/IUpxRkXHCE/8MBM5VXW3x3O0PaWmjrgqQHoE6G3Zhg4RusG4WDBep3XH
FP3nxhVnVN4TwcAqfu+F4srrtx9B3x95Xr3hfBrZxtgSR3oRnV3WPxM3SqdDJA7U
cLYyzKt8THS8MmiUGkzI2TWqSfdoctxDgA3gRAvoytV3CO2zkwP+lOYldj5fOrZd
RaGBfjkEd4PATsWoNbyjd6Gl3lEO1MFWvRv/TfQgzfRmXHnNMeZEDQSr//5qtoLv
uYmi9ZyeWYFnYON29728pC4uE9dRHjUOSuiegttllzGrAA39Mkbe+WJXkpKiEytr
HUDq7tD4HO+vSH4lJ+yqqVmXG57Gzcp5Wie3RtnnkyK0JLDerTJaS6ujyx0HUqjF
mJ6XAqi1pdef9wx+zwTRaVXLErpyVuq9JwSGLs/YYKxb0VwlLB5K9eqYXEFyjE4m
l8bsi+9cWoUi1OSkQHIwEQbzvZlusPT1s+fbzRvzrP/UJDbGBLBURq4iSXt9cKse
ZC7efCnPxA/aCFf2/cpvpF44ZNdDiCL9770ek1ZGdrhC28A9OA0oFyammkS2gTCh
SARq41QSmULqLiz8J9iYNojl4e8UjAjxvXInobG0g5YLGbCVXZP1vlYkhILEXo3S
4OObiheHCRZaDbQD3YGx33HesFN92dmwvaPBq31eUeecKJBQFtT5rGh6+82qQDuE
jfGsSQpqYccNxc5aV0qkm2Ox1PkXbuzeyMgdCcLwDr0uq6TKGjjovMjFiLkvi8WO
GvfMjwpJQpt5usiDCt3tKt61zmm2ODDbAswhJEkBzz3P3q2YJvpgw67x6fP1fTeR
BZCDElORBpr5utIgYoIB0GdOHPxasY7xqOqiR7Jr1tsHmxnSnMJa0YW+yfga6kzW
BoIx+Hc+aor3JL+htoTVfYCtd/EuC7XHUEzaeTYYR7HnOrQAR3UFLPmktNaNAKPU
WVvSsJOEr3Y22iJSq200nguCAoGh8vfkUcSfuo52CldllXYA7mdPoDE4F84okeUV
W48lhb1VMxqJouQ9hV0YvX7P9Jba5EyKH4P22/jRo3fNgqXn4JVCMq845sloCBmc
wzLJSs5LU6925Bn/Nzu3MUt+DOGxw8JS++22H2G/lhTXUgRoBGxUffiVUhukspz3
jzv6+2psiCTCLdDiVUeKQPCOACmNq0+lBDqnibS2s8eSU3/Jc9S1Lm55XZgTyiyo
auMKJrU7IoPNznVD0ULh7jpnF5v0qNLZjBHRiXlAE7US8msSC/tFdU37M4rIL0/y
e1GBGEbqdxGyhi3qA1C55hYfUCM0zPiyRe4rDZVwLG1AT1ez+810wa1n/LqWuceQ
pA6EmElQJ5rkFAxgcXxW/tPZVcYv+Ls5b7+cQzXi3bXeFAa4JQZeebL2eM1SNUg4
W9yMcv9+o+nTKHSYQ20PChNa5Jxr4AHufVpqI6wKeOs6Ljo9F3jOixrCHi6TuBS6
/T83DRlMVsQBuqcaHS8YGQ8wok7thnY4293KJPq8yfuiSGLg3Zr5RRi48kqooXWW
J+CsTzI90MGAg/zZemzN0v2ZYeaFz9HD6ojeBcduUB/Wmx+YzKer3fdp82q1o/uk
okXsMNGiv4Fyq5nbcm9WWiev2J8AHtmzSb4nXbcLgyTkF/nOwbfKp39rIeyipxAZ
1/2E6wt4SGbqk9b0Xyhxm5Cvd7y/MIaPWTL7qwlkxXmM7q0Ql62gzoK7uFla/JTg
hD/tcsJ3r6vTg9Zs3hu+8eb95nhhBOerev6u4OlPjloV3KvZa4QldV30fGpQ03Mt
JmOidk71o8r835BoTcxgQmKrEDu1LGXQMxwQ+evmdmUW02O11YF3MezIp2TmPA8I
Vg+zsRWGEj3lGRV+5Hib3nIz/cHZkBmF3m0Nvfyr3a4P7A1FFBXcTiWh703otCTq
jlB2nZVA7kS+e0+AXZJW/3FyMwVy30eH6cl+ENz12SeThHKNd2hTcj/Iz79pPy93
AtsErn8EigPLxfcEnO2MwIkAp1G57W/sBN7IvEL0X0PiiNVtm+4YPynt4HM2oWfZ
1US2f8lfLJ2NzO0S1aKANWnIt/J7A3jbJ/lalklV5baprNX+Zv/3x5dgxJ0rk64T
l7dP+NySCpPMqjCNtMlObccySgJytQilFsc/GfQuRLRLf4pHY2iAqJHe5ZM7g1bz
iVQhjAn17PvgXxYz1oq4rpaH+U58Eb3hd39sKuORX92hckybQaLqM2HNGdIlEtTo
v6T7uK6sNlLj00qc0vGrlmn02XJihbFKk/6InnTQVadM2LgaMPZSMdcuJtFbH0kG
UxNDYlZHDHVQZLzSkx4l0Lze1V8gGIvkr5XXtakl74n+TMwfe6riYSuwzZ2D36n2
nZnS8oVG0MwqdnhkKFTa3JvNQ2tGOgYLdI2GkTrnwiMz9pj7Q+HQ1AHi8rztuzcL
TOciw4FffAbb0LJ8lkKLVQz3oy44a8Beb5szoeckLkrWxJbqRFAUiOIqVHQDGAnC
tNMSDS0M0NoMbQUqfnVYmwGK609V7QCDthYOcHXZdwdkXP8xEhDVMp4iF5g2yFor
gZUCOn9QAJXStsbaoRJkaEdmCQO0srjA/2XkBn1jpIZUkSFcuBJak+xd7AL/pU+3
efAEeu7lh+emRgxQ210tzTcJ+9mOGSlMciLzV+Nroc+8+S/9R6FDIQgkalHUpMHD
M3phjnJ/KRPwE/i78cU3j4YSEHaT1MTIY+nIOYFhMliNCB0PnBSuwyfyp28X9rqu
Y4upX1/rM4Mk2qEH4pz57m8zQfIBk313PpLk2QPd3khDh6++9vgaOXl/fYBncxSV
IJ/zHurazeeAkjilrGjSlGyzgvRA62ETyjse6Cmwn1SYlgsi7sZvE0xleLDD/tuz
8cD6ui8FW3t9PUpoXVDDRxGM20WZNu7MIJhjgzQTYyRpTuZAOWCj+MaQIQV+gua2
B0EDQuRwJwtadytQdGqRSEmo3u6zdsLAWIjQqa6LrrV+Z/IZsnJwWK5rl5TGBXYT
lxzE/o9CutmlcufT5rij2uZHxeygJXDwcXMgzok3T7a0ndL1S7UvsfEl3H51Kqfb
HLUGtrW2kpvglDtcOtNMIQnG2Pmq7XQWpYmQGBp0+IUwRMvWWW+v2iqy+qthsF6K
tbR7YiMzrCTyyYLjTEX4UEOF9oH0k4996UX+HG5Iku/BoOJ6EAukfogT6IOTF6r0
Xk3EbwMKnwTXyLIbbHavtXeT3ToDA7DVbRTPD7jkSFHordm3wsZJPpL/+YkRLgnM
X/kYMl1uSp2ssViFfiPKDG/hys2AnNMkPzr8Umsy/Mo/6vpc/KXsW50rVUAYVOFs
7yExVaKZyNAHWwbIoHWYvC9ZSemQ62SPrIshPLijU76GsPCLUYfJhqTGSCOMV8HY
y+GURT+1XosCnpLNhYldkuDXKR30JNvOSTbpXxl3VKu+Iqm+9ig3+jIMgfGaW/ey
qCgIhVGVHGZwHh5NMSM2jiJAoaa4RI55V0Mb3G/fibpy6Sos1JVm3av7AmRYOoI5
ETIC+v7i80iBJkSlNzPRNIV4PFYFnzxRHoldEDeV6VTtzEoOHUTTzPZL9lLVljb/
GcwkuRxtz9NGq8gwNHEt4Lx1yVJJ+ZfjBf6JBv7wq+YJ9d2usWZdDmIlq7MbnqN6
xdDTft0pa/plLTICgwZeEPYGm/WL/feBLjFTTC42nclD3tQGV20b5s0QEgr0+pbm
oL1D3UApwMrjQ1vW6kcLZwbcAyOWMDk5DzZSE1JyE+Fm63W51kuVk/OqTKQ0YlGc
cVF7zKYCq/GKphEl6caskqR3tpOo4ivvVe/f+GV5OM527rgghM8iavRcnka+LKi0
UwwTyZ2FOhzS+ssmNGcPYCuKJ21anrRTEjGmZVPsK7BL+diYpcgT7fgXUSdUZ4D4
YH0z62KlGa73g2p3bUChTIIH8KK00GPiO8u6Fb+h1tp8jT0w26kZlWKa6NSHmkKs
vx9M7msxFIAUQkZpJBqCxy3rVIU1Ue3/UoLDP1Qkem/ei1YslzoSet04WXXZo6zM
AymSTYEpoQEunYdBodr+2McIuQIj0AyxWoGLf5SoEO7QTvbk2o27Pif+Ee2XRK1q
VbF7+2ho168imr9AziV2TbIbenYrp3sO5GXD/xyw4vBkmQ5RX7ydqJC5NKvlds41
I37oGocYpKJGNatqbOWlS6yf0zILIHlVsdJZN4UbtMKGUtg/GebSoKLkWR0Z/dXQ
pE7HOu4zPvJVS2i/NuGi168kMvXAyaMp4VX+Mz7AwunpLRduzvIQjm4RXC84jpM5
iC3NSXuxlEH6Bg816MGqXc2GXGL+I3Dk5qk/nDmB4JdLzVL7oMqIPRzfVRC/Hvi1
MTqtq3//kY4lOI/860lD3zcM61uM72eP6nJ49gMbMR1XKVdErLJYYQnjP2H1sf1Y
8/pxMLUIuFYswfZZmPruPlc0kUfnqRo0T3e5gAMnxtKwfgCRxdVqW6a5QcFnVOft
HyaeOPpSHLzvggg4SpdHyTHBg53YSDeZPRkNcVIXBHvBsMJH1RObJBO/bin38gKi
VZenxVHfTWjyEpRwb5aaVWOKqKaK984++hUixiiNEACWJlkUZQTy5P8hsUC5E0sz
aFp4IK91nw1iWcr4yi3Y+qFTXm8z4A4ds4A0BsS5cetOpHgX/BnymPCY5/yRydH9
L9hFAEXhJdZDUBvRRPQWKEe/sdPBrJiZAEUmPbUk0rMCIrZzuLKtum87mTPjicov
Rpm4N4+gpoQqU9VmHXgvDkPtL5avY50JsSzQG0Ip2U0CToIpDmFSoHfBz0gbZ2qv
gSkg2DYU+WNBJPvjrxUnv1uRjj4Mh5xsqzBKIjnF+AJ09ZOufOHA9Joaj9mGRKta
d+zJ0ZFaI8QOZ61676JbcZPCR4BLk0ylsnYbv0vVW2BiWOiWEme+ggjX/mVwVONB
aRYOxTA3OCG56ub/a6+k0n6Qta9pCBtUPAKi7EC5lDiHEXhGuh0D3anpu6xqLikF
g8FJaHlQpoTM/O4WyHT/010ciRrggGDn0TbhCONZDxaw4zXzh663vHXXBx7+F35j
Oe21wurLSB4f+tRlXGlyIkFFpanZOvXUV+sfFqa1P/HgfRktbZKumACvpfVoQSU6
C/GxRf/V6DwFRZ+HDdFtyWnexW+PDtBxiY4KgzAZOLpQu6mcMb/8NWSvzmLlqTaZ
Je+6lHikAEi1Kpxv0xbtJKNxVQBiJTAsAsfK4GanOYDojNnh87gYz6WVc/hgmkMg
FRddjexDHTNC8aFeidVT5ERHGG3CywSmJv8tNAhHWVboDvEz6d+cHTA3WfKI0LeY
SgwrZ9T8LCjkatw0PpvNyqMFjKVGlPn9wfiX3xCB345+rpV7Fe4b0rZIvV/0Mseo
UVqxcNM5ARr98dRH10eEHx8k15ViNstkt6c7AwgaI2mwM1Ky9ZagHLTOabqYSumX
h4OxcocKrT8skS8/E4iDe0vdfXUWcmykekmsH1RAPz9b2Z5e99FrtnthO1sAtJ97
9LBDOLevxMwZqvWHAmpzDzTyocOfFvOXM/F1qSATvJGnBhxM6Myon+9Pt+49vrmO
leEPcWph7uJ0TlHuVTPnUeYr39h0GXgWMy7eCtWEr7YgtU8y60qsifg49trKagY8
67OUyaxkdSKZ94CLX4U/EU41oVz8+pLlaLkEgTlS3LBkeXW0M44Biiiw+TnctVLF
gtzbVTqcbnSnk3BXe3BXv+TkEgiRHSyDt5xBQH8UKyzf8QnQ4AQXt4uYoC0yq8gP
UzMfC8IdJoQFkVnVSKx7EvJdovNBv/tAfe6uY1buNcDO6v4mNQ6GwxwpFmfkjxSl
Gt58UDRptnkqxfOx9OR6Q8EIC+QmxkvkVbxgiY+coNerv2mxKvvkEv/vxzwakE+a
pVMf8siqcWSxx3lhnxcRBYpVwcHf66HBf3gjQTcj1iKuPwA0MtmRDwkTWVmJJFE0
OwyZgaEEsXN2LIyr9yPAUIwaBGp4O2cgNLYYsWD/CsLuPv2egoImSdKF8WpCMZnM
KXDJzWEBJ6W3ppWqaS+WpsVRaStVaYiWdFtNU331ai2JI1glwSsxla3y8Xe8dZJu
cERXOMSRKL6bNyQqA30rfAY0F+mASKZEqXbhqvHolOvDNjtBTj2Fu3SRm7I4fxAJ
f8Lv1YobfBaLpQYtOvT/VAdFYeI9pajjCkFbOlg3HN7YzPyBXZXjFdScbDA3FUJp
GNa7uK78N+uAS89x4asJtwlmE6lE+YF1gQX4C48JmVtL9EvBMogs8UKF9ZUqj6rc
dgnZJ8I6PrKFvIrYIISvJAOUnW91twcIXM1iwMjst2E2kQbbi00cHskgjf+lhw2q
/89Nn2RxUgHd5Hbn3DCslGOuq3HY4RdoVGOdj3iLJOOvZlpHl+GlO2Ggvllk5mUW
mI6Y3u9kgjErO06gGYVEWznS/2xAcSQhec5hudk7YupwuKeAbCyq7AfPdmK5ASa6
c4PCaezt0/Hg6qC+xrse9fCbu5nPtoPsRLHymi/LQXxxFA3V2TtWSO3nqAxT0O7M
KixzIrQz3b4XU4U7d5Y0Q8auV9GC1EoaHHV9O+DdD6DiT69h5rvjKDHCILlhxl8h
7N/Yd3GwqNj4bGwvMiCa69BDRBEwYGQM+YrCwN/86SBkxryO1TApzGCrhYcyRKph
m0wt87R24oY21lUI4LUhuExZY9/DG4dgAFE9AVm1fX3qqRtElqjaARiJUUG/mM1U
r9Z2AHPPOdd+I68HlCs6gwYcDNhOFDQbHow7u2Dp6Q2O/Q76bVleXcv16F6GGVTQ
PmRjlakx9SKt4q5Rc141G8+UowSrGMeJrxh2SoOy8tADd+0Y272SX5m7cyydyU75
W2XrTD+KFmFfCz7Yv0Rp2SE+qHRpAcCtwndmc9Rt7kobTmOvdkE+JbvAdYWRk1S7
2gVY3lUF0ZmDBWmimXsctbDxhF6Jj9nFFjH/IbGuoRpXUFGIE95bXTW285CnGcSk
X/EQCfGdqOyrnkl2m2xyt9QjEvneR6qS1mKCLCkfWia4bQG5zXKGk9Lhpjfx6NFs
LuEVnAEZLhqYmNu+xUOFxBkFkivXUfUBpySoMig/H+2Gfy+65Uuy5oZVZZsaXxY7
iANG29bu+pD74pxBkkHdeumVgmB27cDfD6c5ZWIJRwGfAJsaOxxNWRzG8PR2y8+d
9RnNQDIUDgp2f1ypvroYSSg9wyHCn3L667OJZrQPQR/vQssKI7Pt2s7wZCgkEUH/
3NR+zO5Vi0V8A3cLF6VJxCD+38eNp2L9M2V7cYwIwVWRISFaBwmo1qPHPV7bxEwV
zkrAXwrG3hXrJ2iAkccGWOpKhyBP74JoZ8d7R/WkFOpz3cX6gfCqVqBXjgZLILK7
ZzBUg7Q9FpfmHQsgMwAvWrFZjCGYmwpV3dsdfKfXyRPZW5jcQ2b5G9PT4CH190Fz
1MRaRVPxhL8jb70KUap6VoPMXL2TdtKTrvF31DnyOgYcaNw8hmISa/gvJ1zOzsCD
jXStDWBCjtwYqTlYO6CMQ29rZ5QUDtrryPxqAWxl0IB4YHoUHsh+02gbhf++ZBik
/mLOYWTvoY4SheOMPt2tOWHL9UIKVG0NzF0+dbYkp3bvkhVE+tU6yhaBhihOe5eH
/B0gghDW00lIEk+PaE9TN73oK8CApWaybJNLp33jNwmsWViXwiAB7FfedmUuqc4K
IYqKzievggfN47gK803WjNzIyRlmDK+dpwz8RZ7gv/hnJmgANRIhPDZACB9X6xZt
GSojVsKgEi62QawEVtTmGGHY80PW9FGSi2Gb1bL30cX2yekecooW490Z9p2VMMaU
zcA+6fjNs915XCPC4yyJ3VTSHji7JF3bAEBV5rGE2seuRu2Ws3RSxfz81jReIo7J
MChmks4QDUaYY4w34TlYftU4g0gMMHauBrdEQYjkJpUyv1ZbBZdcVFkGusCU4I17
o4wtkfC70cEWtWmwi7lxqRTpJVywp/XnEmqJVUdhZab1cgoxjp/BCk+I7tCXann4
88RuWtro3LoUAQt9swxnBmQd7MO9PnLrXeZCx8ZSaTUbWx4ktaWRAGQ91Ir5sM6e
c0TnIGqDcdL1iQ/q3bGrrJ8wjio4jzahO02zdXRp5lMn2Fd0ymULtkbqmPWv5swi
I2u4YofRfsfO+ekuRhh9ETQyO/uG8LZJ6YWbedlFP/6F0jzXAbNc7IrGhOuJE01O
uz7fPhmALScWfy8Vde5jZnvkDEiWU8YSZk6PbJ1rkoiy4Gygxk0YHO4kylJGlraA
O/KU5E37td/fE2Y0pSy8A9C+K0oQlGs6gwR1KV9AXS/f4XJPIzKmL9mEx+BiGCGN
0oLRTUTNfr2ZzwOULc5Jip/nhYJmwf75woRICJLOh5DQHn1bTnCkOIdWpp7YGZ6p
SvHsmgrczp7ebNK1oHjSK5AtHCRZ8jcnwpQEzPz4nSfyAJhnT2Q1M8Cadq1U9y53
Nj8AmiS8hN6HaPNsC5D98uOq4IwjEdUmDWckCOSjQQfIom6aD1vQ1jkSIkh/BAMx
+6F3dD14FwVAbCM19WXrvV0aZCkMpuEpe3nPNq1tNuKEYGSFHMPGRMnUW7KF1Mww
eRguvvGEL1pyBwE28ECLvvAVMSN4srQr9Pnx0BWLpiwbEQYetr4uB1ITSpCR4bjn
mGY008wtflXUKCH/4oOuhCM3nE8tkubKfAtMbQMuP4cpyCAovTeK228iN/Iw/1sj
iy5tz6rHa5R+GB/RqI6DBViCmPKUIDgnR00JhuK9mlhEEafpU2JBImmZDOrlyzxY
VhnP4pFkaLAWon/w6WJUN+1qWeCrELeBSilU7jDpOqbK6ldaXUjNW2maI+2jcoSZ
4TlvjuMVsVVtoVGaXaZ4mf72BkuqiGYVsI+JdXtdBIkLvK/W2s46Ya7MlLoUenXw
KD0fpH97RAOsaIac/v/ZoTraVN+FC3i0jq7FxUr0Vv93NT16RA65pOyC7YtN/Obf
7CC+FVFPPbiYuAQqli82A1aJvyFLa9ohs+PhNelc0ix+RDKBYYdurf/xWWfuEEdY
hFq1pEN9qGK5s8EC00UTa/ukYXa5KFWzgg8um4R7irUe8qPssF8Vi2qVWDj9LwqU
3uqrG41hJdPmfIlm5ZrSg3LaR9yP44dHSX0LAsnp6grMhDroVOILKRAgIDAUaVxy
aqT8jYvY2FWU2hdBMQbOHB9lgrz+zfZal8o0TB5ycJBxiTKE/+MqtsIfNYN+0ums
coTM0tYkGXqQ/eqsMg/PaTo2wLOf7NlGgreqNB2OaOTY+HBaRHKfXkpETORoZkCp
z/GmpfQlkJa7tjVlB8LvcWJps9OV/SLoE7GnH6fbVmclSeSFuQmIyZswA0mMu1MJ
+TJobeol+iRER9xEuBYolnVglsqXDMIniU0DfXIdXd50oD5Apo0kT3ibvYjK6oVE
iAokqc30tgg1eAkLyB2/tBcQCi+VpdCUpjnkkjMCSCwQfInCz9+I85NuAxy1EW27
cWtVUYTv9VIOtBrprDPsfVBLiI1u4seJfivBtQHUSPvxfKq3KNC35FrpLEo8J99X
iDeDJigkjuYJ4SfCHHRPUGzzSAEAsnX1waYvdV5uzbVsYwnz5M0SPMRfxZpORSp8
uNxwB+yWaZ9xAeSU+psCSFoX8whqUn1PtW0fFkVUT0dviP/X7bBcWDhXQbmxx8fv
ERRTmun6kCzwI2ik5MO2G5oWDhCCWP0vXfms0KQi13cyjo922mFeLsDvxMqcGE4I
TcJP5Xql0A+yglj/lRa9u3Rf+EUPBgvtGaSY6miCsRq80qzDohZJQv2CSoNtnSr2
jV8J4TK+i1OyR135pZsNaWD7Wwg7a0kU0iMFeRcIFZpo0QPaLuqYQGRFF2kPuFX4
htrwiKMkHb0z3ueURHLgbh6aKJIfcuwhYY7cwrnnJRTj59L9A/2Y3KeUwL8kpl88
phyzF3smdffaZo/RY8Hbq978bD9m5QXH8gihb1CDDlwJB77HsEk+iOj8Ku0oseGC
XLdnXLsVnAirvoYj9PQ2s4inG/f++oMJ39IaheLJfgocrzHpinaFU/51bctFtttd
iESD35Ny4uXKLSJjU4euX5ex6843zEdZU4R7dLuCRDb8UZtXeu5fpkj8lSu/Y5wg
iARFxjun5FzFTtk2xyngKg8dCeZ2NmS/FGs5Swv1wIURJ04rZFyK3jNVWpM5/49d
6OqqegkWOaw2+kszeHwDk8XQAKqnCasLx4x9h/TirU0HIdd/wdTIOgAltSInGRtR
XgNH4IMteqqL6uDQZV9b3cwCKmOmpxJEkoh3BdIP7H+ZIPlf3F/cAVEtoYPLNS6A
odZGx+Y5J5zLlK4Iuwet54/zjyqanQktKAX/mLnCXwIXaa7v2DtyUHxDnIAeZVfB
F51SRlYBKkaJfbXydSbXTC/Ljz+2Qcx7stOldrVBz7QEyrIUTXs6bKt7z+JLdzmR
JGs9GdeL0IbYnNeEcS+OheZWsa+TyyrCCMZrKKY/Ya7TG9fgMDmuHbF5jtI/AM0b
d8s6ZfASc2XQLgJJoVGerE+bSVQM9M+KKbK1UmG888WmkdPQfpf/Pw+3yqGQzNg5
0+7nhHopt8YiilPSqMBIsmSVU8o/n+hiIpVN8JuzyTdAnjzvSWtXHw6Om43MPPKe
5Nbx7UVGvlFyisfpah7lKzS61x9RJZ+2DTijUwsPGxwx7caI2J9ni01Cr2/zIdqN
vVu+gZtu0ZCJ0FSLXHImRYn+Dt5r7zN81lW8DTP+RfDlkF2jw2itjjuZg4f/lKZE
HvlpEV74g35atjtQ3BvZSEJjhfRdYojpuFlY4wMxo6QeS6GyS/om8+mkFFkUGEIo
PIAmNfbY3qzp0Agx7xp5IL5N4rarMji+47Me35ZnTe03lguwNB8Dc55+QjLcRQB9
QgcbhuSlLNYnkZJP7cY1VsxZW4UsG3Qj0vX1WW5+5dqp7oPyyUIWz9PHdwuJ61AB
osJ1UJY4VJVfCU2zIwp88rfk0qeXAR3SgWNbiSuP15TA9JRwzLZHChZ5DTh0iCpV
EhXW6HjoVp0VVdJKPTw1bGclO1MyUm2yBUjtaW/d6bKXug1Mqx+CersFie944HcM
YBIoalG7QA4SHreoN8X+RcMjBfflubHwQEQPPHrR7wMGEvnHCK+54sIg9BowsHOR
eYzuLWkx//T+oCqUYgmhJGNbuKBOsVEM6Ci4rGqR0rYUhrNGmwgnvgfs3y/HReYD
/kn7EfwnL/vCJz0BATjxdXTxNiyYOZOR0oR7nbK5F5NFvsf3+CF8gqN13N0otPZN
NyOL3NtxqvaAS2kh+wKg+uZQqOunxKe0cemG0a1Tcr6dnSASgHkJ9JZf7Mm57HZr
3Pg4CLpRnFsZ/O3xjtSabobSoktyfWqAzWSh8q4SvwBN93UKs38KmH4U4gY5sE23
cJe3y/QtvbsVRdm07ik9IYs7Z7eWELdeW/6mefSzRqO54DzzJxO15gQ94BdJAEKs
bycpMAoxAgvuO3OO+kwsVo/wyST46knTZNzuZsjpXdjrhBcvvTbrdRtIhQ9z8hgb
3AtVLhCXOEWbmP4nUoTvOdu/HRx8RyDEGzRiNIfwVtPmd/w8MqhUxKzclvvaML/j
T+/oQEnYxn/9eKn5p8KQY49WgNdZBWfPGFtcjMsZML8sQdc7cR3Y/T1pqb89JisJ
IutdH/73e6SrGjHRFKrk/jf0FNfMEvs9mwq7/YnIf0nUHim8bx2+O8LlZxna5Vuk
zWjNkX7VXtdwej7nQzRGjDp2yWb7XfgH3KIsKQDz3iuRHtXg95B4w2fwJeXeph5M
0icBX5FjnOKQB3NOzjeeyxTYdHjVzh42swALwt1EN5fN7OoF6qyzirv+YqMXAEJp
f+0only4H897wNZsauy/9fEkzrZ34xA6JKasoo6Su0/Jne643mSS0qQcXaBD1ciX
qNWxvSfWNIyPj81WrW/rVYGQqLs6gjz50rY+jEe4wsDMeLV+VpgvqU5tPmEFHT57
3GpIIsXwYyVNTfsBMLBsFcyniOOcgjg9AxWlN6BepP+7QKTBTDB2wlq1z1I+ZivI
cH7uzXqYxbSM3whN8YbLKrkurAkZwT+kUN4jUpbgY/QCnpFyTheAH806WP6VUgWt
MAbL+FS6u0kzxnLP6QgSb4umighgjbNf4StPnovUv+BBggjmc12tuT19r2f6LaMB
tGNhPHKKmv6UuqJfgm+Ayu0JM/B895td2iR71DBfWRqNzIVPvUnpAZbVXjwfjmJ2
atXC0X84FN5XiyAXGpwIpbh8UgT0+HWphWI1u5L9PrXkYgdp69sRbrMPiBfWpZw5
7S702H4Lh0vpcwD34YgvOiwdnXNwv0RB390sHIG9+FkJyIJQqnfvY5xGfmNIkowg
sXt8fq3ypV/ROW5EnsFDb4bZXgCJ4RGEmqWsdJ1C327/3xVucXhat3sI9BET2fvj
ejEaqIAQS80nSStWtUYaGykN2mb2peIxskAVmrGIi5iFK05kx2JNo3SCUAI83KLy
wuMbfUKtzmy1lL+HIAXJuTLmfeKXOV0uRUUp1Jq0qkmgqJfub5bIffnOBbBDTcPr
zidbQXS9MN+bvKTL44fEyYniYtA/qJy9wzpc0FuignhX2tGOWlQ8UnC86/pNuB1P
i3akxeD+eGyloltGxwZi/vP+VImDJ0Ssal8Omg7VWadP38HIFQz5MEGT2iEX288U
dQcNHHT/2x9Xp55IpdCHVFI/6y1o9dHJxC61IbjdLYBA7XR44R9ugrglXk01teTB
Dq6RgNypjnPUAKL0p/zFeu34bPm6D1U9CbfLI1cqt6PFT4UADqtCl7Fz/mXrEdIL
1z6ayjP3WsQXXnnuvlTNgAs9rtB01W+Jzrj+6vSvhsHUO7BwjjMm8CMLCyySRhYJ
FaFKhDEh6wh/KGTy9iK+FqEMgk3/O7vaoxN4+5rcSZURbPC/PMMK6NNnPDorGwdG
7N+Mua89z1iLfgUomKipNU70QZkHY6PmkwtKtypV1J1eyvXY+asPU1qVJhUVFA8F
RQG4XMmWUkzO4LyxgGsyl1xtURcs9ySBK2hAM/X7Iy0yzEZpdsMosOLY4G+wcSGA
OHejO+LoAiuJdJifhkgw9R5/LbqLUuQXqWDpEgEGc243tDl8w9hvtJ0pZNsHJE2n
R6mZjYoBjXj8ezubSf+0mS6fwOn6jEdmJhiHEy+74y+/glGAZmklPlbxjzFLCaRH
nlneahm71bD4A99E2083WNI3AvtOddNWfqDXQ+zPXAYtJRRvnoc3o8gAZ8u5m0Ej
JVRusuNOHdvjnfW4kTRWJXDm5EW8nnLHfnWpyUxc6eOYGLpZVy2CwPle3BFV6ZdM
9ADQULR/oG2KMlnNOcDds1YkTSCeC4z36U5JnyqB+SNrFa9JIG++FFsMukRQvZLd
QiPvdEHb/5Y0ccY2yP9QlzOojV8cpOHfcFG4BRZPljkHooE8sYuMiDJUoZijHC6/
p3kf5u7SGIpbOb2BacG1BEuF+LRAITfVvkX4lht2M9vUEOJ6pvaNzWcuW0wJNv9+
U/TY6Hfr1uyl76DU4wqYT/f2NfzwibFqW9rWQBIr0IjNpKgqF4xBR/zIzswAvHun
gQj18eucg9XOom6s0a4iTFoh4/iMTiDNFgFSlKhfHc++AY9NPo4BNiqdz6IIIfOJ
Y38e5vqsYvU/gvbicNCePKyaIbvZXHHA9cQ782Wv/Ek5vW7UvbFEAAUe5T5Jfu3f
Ql2o6bsNTOvdVRk840J6Jb3txgcKSY5dNaZWjwgEpf4ECawWPOxmkGkQKboJRdhe
tf9gP6sEcuZkBMjm/B51PoncVX/fhCwOlXIBf9WfIb42RA4mKfGJiGJyNgKf4y3S
2nPSqm9lA8mOHv95Lawsl22QOQczNFGKGpNFJHbpMaxUQOq2NaIc0sGG+d0JgMZn
C4UdJCQgUA1vcyD7mWzncSj7FCEPwZmbCYBD4CqRiXxu17ffcQc/6QUt0Z3VGWG+
BJbzoXSBxFBLQ5a4ORj8dwR9YdbaB2zD+TnIp7tRpVft4wXdzgB8xpbHJ0ljt3Gf
XI5nf5RXQb5RtQOPZQ4KEhRaOMhU32ybnRrJYzX8uLkQ9OD8JuaUyvQd4Z5bM/Qc
bQzJMS7OmxNz+D+otpqhoBFXP5vdsfK9aZwedVD7f9PX0As6d1OSPaFLS+H2b60d
i3pAdGliSuLaf+k/JJT0m4FZ6Im/CFAaGEbgSXX87+CVvA40xp8qT6JP/9+qTJHH
4+J1Oga2O7pDg+8x5MVdVtu5BY09yufPphvfA1Hvm4kexUWIrNl8LtJ6qzH+3gvj
74iCbmDfPXJwzW4UUFaPzFvbBYAQseOWhSPCSiThYzoBBc740FBl9umn/3RT9IZc
1xr3sar7SNu3CEL1C6YKKKrg/7Vz3e5H3KnEdQE48IrqAi6Skp8H8jr6rDdTg1To
2g04PC/95JP7Gjs0hUUTet2pUnbt9PTrA6+IDVCHsjtypCu0FuJcs81/2ej7BBnf
W6oqe8mD+7c286AcOrZ6oZaR5B4HRtfHGspqLS+zpt+5eqIIydO705O93i/MIABC
5EfN6nNxeHCMg0japt8j2adwb/O937Fhd1XJHCQFbs/VndzAr23ShyzO7V8jwY8A
scQb8bskn59gdvwTZ7gXx7+G9ANoIicoNlVHnxU6tvOdJHPxgOnzcgffbQGpj/2G
Rl/jHegpu1YFa2iSnbjZYm8KpGNI4dlR0+81xWmVVeaJzJwjDqaek5CcogvDcebk
gz/Es9NuFfRlSv0uff1RbRAVe29XXgEYvUct9l6RbV2Srqdl6Yt8dqJN8JkhWkHA
anExhpWR01Szuw7DHu4bwXB8APfjgMREi+28OhKekmY2hWMckBZWaimWt7djAJS+
NHk/5SEhOYa8wQui9qR32xXtQ3N9lF0sv1SKJAYW1Dppzd1TvPTOuBsWV5mjjox2
KIyhbwZ0DhvYEomQHc0xJvH1exVo6wHAeiotPSYDmMEeE7d2OU8Hquq3nXMVI6wG
sFz5SRowNseZvD1cf1pgFx1XTWeTbqKQx7Rz9Z1waPgrGJctwKV+iqTMcZbvjuae
Rv781JJbK9sQT9ruTua8to7Xx8mA84Ebpe80QaWI9Mn94+D/D1WxYvFgo/O4b/cM
A46fuF1fEwq0uTVWSQR7GGtw57S3EUnW/R2vImY8+azETKE+ItPkm2eINUTEE+RZ
OqiuMmikcTwPT5QxE0TRS574xwe1Tc/oOJ8HL3J2Aw5aXIXuQeFFAsNlO8cbnzSi
ZaZ94TAz2jzl8Zbp3vQAeDUY29lgiPOrV5PNY1ukpWhNK4ttjKSLH7mBWWWH/L/N
zr4mqa3QIP8qcHzhe7p5yRHfandYd/nW3qr+dpYjyqjXygTJ8osHaiuiO+5NJuKO
ZBm5a/HvKnAThcPMaGA7hhHHDVxyvtvrcQ6dNKjyuKMJ2UiuVqbSij8aCoGOyQMB
wKlRjnF0JBhz5bkTNRbFQrNgcHY9SA/RV1wmBvupCNCtQXLnYnDvGdfjfGTcevYU
YjZ7oxV19TO69yLZtzIeb8xpeo4DcGBLWOma7pYVtEipwX5T2yOwte06ydKKVlB3
WqtWO5ISqGWr8QIz191ubrrdY7qgGIaYYoU7R5KmOWVMhnmQ7RyEWuf0jTwIm5kB
WoyNBBOF6y39mhSpTw7wK026eQAvdD7xIejeJL6reS7bTfXKtjRR5UzpT+LZCE+G
k9ZniESQpRyTAbONUG2MLAIn89e5CknT+39AWa5kQ9j1ozR9N0Bz3MTfM2eL8Tof
T8LU0JKtFYF887aq2KrWKU0O3zHapcU+crq+xs8ICpP0Pe4vNehv0PDyvJsavjDM
xL8tdCZAFVhBu+V/crjfcOWteOV2pfPqTniMv4ucFmZiDdWr//gr7yF249nHZktz
awecuxbnx0sAmQ5mPLtUjMhxJuhOilywzd9dpie0g7vgN7FAbhJhtQq9YN0VgtNL
/diaj7KjfHEh9TBAgEg3LCdv88va0eGYKPGWl9i0jcIy/gpVaH4xH/p3HckAu/V2
+bkKeaE4BvOM9yOnFnIYqSUS+yf2wbJ/fVLYXpot00s3gxoRuWA1NDBAdO0o4De9
vaVEtXdoC2hesEEiVTQ4/kNMlY2p54tyBBNOzfhJUpdPvjLt865qJFr+G/BnWTmo
C1syFXOGbWOwXWmumbsXAVVP9srAF9KAI05u12NUlfxXn5JtjESKRHvfNitPeJzw
vw6mUwgOUsUwa+WgRasdQPR9skkEIc+Sk+GZC1ER0Mw3Yrh66MJtuwNRDFe3NM2n
NMhKL5efxVYUYiJuhkqF+u4EXsAbSlc14xudNFw7E9OS7YdfTY19Q+11GNt4tmYx
k1ZAK2A1+JYRRbSPjXhtNF6Zs6uiQf7zpkUnRWkOpcQZynaERaMHFg8W8h1O6T7Q
zl7kDhVLCaR8L3M5Oz+PhPieKo6D71AA8h1yaCjJyG+QyOVYbx4RD3VZGE1WTYuD
gAeVrQobHzvKrBHlU/VCif6+9kta7LvLPJQeqelGR2VuxbWuyJOaQtIJkgKV9iD1
oMV9a60os9B97UYSoxXqAchCEhOBv8ohf5rC22sppNyAFf6m3LKtfA3752mTY7N5
jd0ckfeWJcpECqlmsAVizc3Wvglf+NhVxcbbM43vdLcdVrq7Gp1spnUeNXwgyRvq
UNEjqG1GeBRQDTHTylZoMLnMfNKhG1gXX+H8qvaQyrE+PAkZpJ8eSbxdtegZB93V
o1osum74XFEGyftFy+HD/Z4c54B06ZJtj7+ULt6UJXzoJ48hYJeX01Ud552oEy39
ab/lHw7h88insoS4J/lIhMO1rWk6wFBEXsmRLNjC+5OknlH23TjOQmnNWTL05aPN
uzUuQ4tfg/Ye/qofXttgK6m5N8ZJNbFAlZYHMJUnVMY88kfywSfydsTFjK06HzTN
bps0jknhI3Ov8YjRcZd1KiaxSyiZtT0tbv14Xh/P/vasS9fTAC0rsDxwXwvTqZ4Q
2oGFkpOgvT6j5KYxz6jdaUHYc7AnF01wg0OdpRZuU1MK20skisBcEGmC1h4bv6yn
v9LAdqLvtfOkaL+IdoofpmBcjSWyV3ScKGwKYj+4vim79MtFJC5rRcXxCBa+rlHc
+cO3OeatwlM0XhiMTmV/Fs8xjQJ+QtRGJab4gbal8rDSWUocAgIf8MUlyhg2JhOe
ClJw/VWrQIlVgSmlJ9BkekxcPaw740xeKoqFBVzPf6OzZ0v2DORa0cngxWDMNxuu
GCQz5/T3tjaTOjevYs9ObmrHoZVKoHA+XvrirRjnGV8YEYhPe0oym0tPHSBTqd1j
gw5mscYLxzpDRIt0lZpAzwL+j4wQCqH4WLJeIA/txZV23yBX1to6OYGQDe13c3N8
+fLMVGjiNBIpaDRN8dN8ru+hMOkRjQ9mOVNMcB0XoUPk8XyYMofYzeFEqUnipeZx
nkQQisvkj8yAOjWz2MWKrugmKr+Eys6uIhsj8fADHYpBBVyn7OM/XnKr/geVVmKm
k8RhLD7gE3nIAxQZPHa3eHl813uamTWkW76uKdnJuJcQylZaqvV48csomUN6GjtR
meQdPhrCEl+0R/q70yNW20s/yhvcisdllWUYhTE7aIrhRqkr2P0ne+hJ2MbftCpI
zH+1/qznhX+k4P8+vesXksslJiENdZ1WSx6KRco6VtWpPc8Mce5jXSG/q0DIuSdc
h2MfmbBIPp50wXRv8nCjaMUUBc7+5OOHsvEvvp4jSQVJUowACmFlZGpj4n0WFhZM
nnjFW4FVGGprnns44Ta0mXnGKEo+NiSM4/EGW4JLVN5pd/PwrhXV1zue/l2u0B4t
SAEXhFx6gOaBos6ev0I6FvX0REN0gTEkfv+9LJQbUCHeTJBdRMfc5RY5fdJ2hmkt
5Z3zEFJRwDdL4tADmIoQyw5x7vmtNXMgMQs4XXgjTDFcKKPg6iP8+T4uKf/+wJ2I
o19cGpFjPs6WN+UkBd7rsSglUHWbRjDoIR7yeU//LeV5Osa9SwumZxn/BUPo6fz+
iaFeQ9bB1FKO0iT11JaPj74LbO0v4l5aucE9CROQCzRIEd1yRYl7+fJl6CsMretB
0wk+kbsCr60KRGYLmZBBvD054WtNMY6uDeQv3kTxazRdP6PYlXa5X1NNWEGKhakC
rJnDOb1cg5P2tvJD6SlDJbMSLzKuu4bNj6v+0N+bu/+Y6AGBCFHw4xsiBUBt5Jr1
Tvs9O1rWRPi3P/YP2FMTl0nmKu+e3KrUBSyvurLiaUKwmIk6K6/oVm2FCreB37c+
xBtJNSpmrgkYMu7ggm1GTKE9hC9AQR9cE5koEAL1/67bUM318bS3O+0oPsLEltUZ
ZTpmQC9T7acRfdy64aUOTPnvi/vPWI6n89+b1gSYUUVtuPQWuivGVPJajROm/VJh
dnlH1oGchv6BhGBpq7DS7fflcE4GbQwO1U1rpG4+jReu/V9M2GouQHoOsDGTFapN
cK/8DqVqVQW49yzJ3SQTgnopXeDHZt1NEDlYtoXAFLtxZX8km6fyKr/9J1741MG7
YP2hkplJkUoTlbRTSf1n+egSC5ubcOgIP5erLfMiLZqGin5hokdW67KyWdNoxbHY
1Ual8mJUBOZqwqyOEJlayu1fgGCgkBG+APbbVUVe0H1VHJCXSvkNWBpUTXblqHmu
jOU3I1mWWL5xjU4kA5VH/twWLVgBAHOISfESL7ZlFUmFwsrR3wND7+P77jXBzyri
oaUpxkV3nUb/f1PPCLWODMZdZtS2sR1lLuGAuzSZ7MQMbF3AYPO4kZ88+sWbi0JA
wH7OM4dhxYURV1WlDZ/VW18G34FjLdkLjgTwEF6LXNLTTKbYyLIqUbhyOCZiPmSg
BYxENfFXg3eFeh649D/7t5L0RCD9DGCW0RBRWHWWXfcfBe8WajJsmoDRZMm4r7Ce
Is7tqRAhq2nD80ySgy8uoT0EtC0P9bGhnhlpO9YPto1LIUFLykq2n4eiZ030rm1I
T6FrngSLW26g4JPvRJY2AnbnljWpGpkCu7VDeznbuYoMenWI1rvS66nik2+W0Pua
jE3B9qU5UrCcTx93DsS2WsjGL30oRAcJXxLDuzYruWo72o86QirYtLilhv4lebsA
1BWR3KClo9iFJk38tRnh9Xtc6YanO+Vm1hK+yasa5Ahgfr8dOj7yt8Mtc+Vw7w/4
3tmGCN4SOrZWXEUZ1qfWTFxhFk4oLZHXml+7kXNe4rdhpvmKI6m4y4Vo6fimuUsU
S6HbV5Kw1LGNumVvDTEdIWrp1m5wKIqnWTV7KpE/sDxpE861uMmdrANrV7w8caA8
0exixxv2LQSytAwQTlLxCGrPBXtauIwwdZ0jG3gQo8i1FoqDtxMUVDsn+PweXjhz
qEkUxB1y75DGelKsrlCEl4huKtm+CFqaK39HQWDSFTlnA47gh9mRX15GuueXIpXi
o6uujfowTKq+HynzKb6lzK6igEf2ax+8YXgla06RZImt1ld2ncUGXmEhusb2r4cX
VYiqkSBtazpO2vwiEdZanyn2sMS9QO7by+CqG9OMiu7ycC0mipzGLzYXgynNB6dZ
kYrWwTo+P8RyCjSa5dRRIpG9smm+f2d8qJzxpQ08t41ccrmoL+hcDKcQe9GSbOG8
XqU1WLu2RoO6rqr4nvSg3ZLCchXWo5Nihr7StGOTEVFO/G4o/0IwQkRITXGqZ3ix
FWD4CN7eN49Z7i6KgwXlD/FPfKkYJWJ4KLtIgTtTXt8axBYow4JepuxsIEZxNVOv
bqobM7ZIUAp1Ye4zYzqX6Y1TNAjudNBS0dr+CU+skT5x4ycopHBGOBWMUQkWEdDu
//nFNrkwyn6kxQIJXVbstS6ueDoFZp2HMr2cciQgdFaAZUeNsUpTCteIU4ATTxXp
H8tO6fCMbcmmuhQL2AMwf4rYYwLONXLWUpoOm7d6FaGbR+sm/YUmb92NnklWiG03
D8xS4KsM0dRiPLFx4OkBI3cckmUaXeCxMFsPEEeW1XNGIkFBNmCKDcLJu71rlZr7
+eSBBCiOoctmjqB5CRDsESx9ERz44XW735ZSQiI5efmS6zRq/UUrcIy4ZmvSd07w
RXpUqFfESMBPIqTMW8MYQRAKJCKMpbA99kNV/HSwD/uLhNlutpkxugZAezQEBGdA
gA13AGT1PFMhRjoEzZ1ydLhL1qBe2duL5e7RfSFh6wWLkuWxyJ5WU6PPV01YFwhx
8We9jatVoR1JNNk3m+ZORgu8GwjX//4WlztwbpBlSoOZqGaPavyWdtE6FE+tT22E
khOfUwa6qwVcmmZydPwb+rT4Xnc0UD4o8R+b2BMOGj03qRI1gXy4bMvT2VoxyNfD
LOqkNQw70ptaL3+ionmEZNuFZhlk9h1IAJc2yoC5M2sg3KJb+cwQJhy/VMQy6HqL
UUZyJyEvD/QveaxJRchdKw2tvtSVxs9bxWrWLEGPgYK5Fmq+EIiXkQ9SCOZj8omM
zcIupoEUcfbb4+mFzEkWUehYIZ2xYy1xGjD+O/RgKGEIJFrAIsTTGS+L/DsITA0F
kAAdSfcajkybjGIXIR7MgLBGnDFTt+ruUYwzANv1RH0/VdqfYUyrQa6OpzjK7HDp
qkUhy6Z09zuL43cWu2b9bFYEWrdVf1cpBDoXqoWrVl4+ysgULtI9SgKdbVB0wkog
vSBBkARQGRPHgXvda7T5DYmTmX7tLo9DQJBK3+8HPE2xdTwZhZIye4p3CS8wJIb+
pNH3/6eAP+KtFiUOHWxmjT3qQ9OECR51mtinMFnlCBIXl/i3BxQ97Heu2mqYUse4
MHyeNd5p/70TS5PoeSMsQx+qAoF5hfR+dB6vy//fg3FchyDoN09QsqBL2GfIGFK1
jBILBqfyrBpd5ysMXgEuuAvk9gdrcKnUgdX3MJYZPci7NqEsoDdOru4Wv8RnXeV1
GHt6wu5PfF8ILZbBbIh9/U1ZHnixCRrym4LBpn0xENxjaB5ppwt3B3iC5+zYQ+iV
FMKNgDKNovAiS8GlEx/aqGeijy5QmVmLayiHlVs11eZ+iwbuDvLcSkMqJqh1e+Ac
iLivGU8gcG6OemYGzDQhY0bCg5l1p0a15hp74/+BvHx8jbcMMNTXkJy4OTRjGSSo
irO+06mPWFU+L436h7Es7radpXlwZ1PcnKde6NGa9ivfHjgutvr8GCyosY/Byo7P
etBeLX3A3AVWc2cVxmXDxpblPZbp6BMEhpKTrVLjI5GVEaAAhzlFh4aEG0YvIM+9
chVGdcEcfb2MFCguDQGi7oIOWnnh3xNOI7ackkYAaW7GBS0dn+c0s/nXnVW6HrU1
FElmuxJKIVS5NmigBcc2y9udqWhVTv3kCyvo8yvN/z+g0cc4XFSHPzgu4IF5mcWp
W6Z68blvVY0Uj+C0S8+QNPcdPCtspbfYhgF02xNGVDq7hXJ5FXRFD9nGPX2EzbCE
E9NZk+GTmJguxLbuBWYv8GJ3QG7isDr15GMvFgnCiGzZQylIKwJ96+zMdM5r73Jf
UR+PqRg//tKH7fb6Ghpbl2qWTajGS27/Kfz8pg8dZkLC5SChUai0QYIYGAIjoQPC
kBjaar0ovdx/BPXeLHyU+azTuEGoGSsQecSuvMVze+7+O3pUilWp/6b9yzZBoSjC
TV6mYW06GiV9XPmKU/2p0hvVnt5vSvQ4TeTmtWqVdxsj2TXw90wVRYfVo9skhJYL
re57FSn7cIxmNr84OwfRGLT8GkaXRccQ3SBy8L/r07bw2cZ3/fm94KJrTDqEeVnA
T+dGFoLOTLKSnr6ZMuW6lYm9ytTEbzFPoFN6aWOZ4ZCs2RtjSNGisB9jlL/65e9X
ln/zpFdPSqGXj7Mg6eJB8OIyvtmopCZWCHUHecxGDbJMK0kn+rDuQ4j83FBs2GSC
pO5//k3xlOcFQo67UKJiZZfJtmZHGpBwPF9slxuIiDuDbqm9p3sTJ6oX2dCsTXXP
SAN7EFJsBJ7yZQgkh3J6SXoySFWABpf7BjrmxcsyrD44iDspacvfa2novs2SK9LW
tuoZCW8Qrxe+OA0qpjNBh4q5NPUd1kmoIHmEX93dbpu/rWIvds8ybH8XAfii9xGG
aDcMSY4fobYpMBznXoLcpaAZCTES9ma/mk4ep2gJVrrrO/yCCgpB+kwYeUiXgltl
e9vvZ+gCmTDj+QYLhtSNX39jiVTsG2LjcWTmwABqNIUzANQjIrePIzhVsrNkkfr0
zzLluz+FZ+giI1ixm6uNdb0hX2HisA5tMQzsBUtM6DSjgfQMUADvlxSucoo/MlED
kRUcoV9XhhS5JL4XDat1ISP0LUBIZK3ZIwEokWRLArnogw2JxJC0IwZUJxjqLlDf
N/EzDnRCHrLOoBJM5zkB4V66QZpnxCbujxiOeF0q2iE1vNGnnpcwZUdvWTRokDml
VovPg5rHCkTAj0PRPEknaYidQSr3P2hK0lqvLeYXVvTuoOgwdP+3yOP+4tT6Rmad
xfQOt8JEG7HJjymHczeaQeINPyxDy+vxcX3deyliP9Dz3poi6BiTB753a1LzzgTl
Jkq5thn3alU5qaXn9P6q8WbdblAX2TqNkMuMpanaUsmqKWBw3ttEd+0oNivxDwnM
tJ0+aQqS2jotEsMjOSOxLrhV/TUp4cKW4Gr0qN4mAMJXUaI9ZwUut1WvnpW+b+Il
B1RpQyynSxd4s2Cnqk5Z/4xJ/eFd6Vhr7O7vk+x7WyEbyANtOuyskqjbarHP+MnB
Vk6aujGAa4iCV1vtrbRej951S3gZ82Ac7rDgEJ+59C3TGELIrs/JRh49bEHdLPIe
jke5pY8kCKKl32rjNmz1cVcIonFVutUPKlb/eYuXD4EHjvBA7XT0sT8aIBQDDiKL
0LfAhQ5JwIu2aIiFMfknaA1X9PNpZNQF119m5qLJibkNzgEmTZunHtWRsTOdwl1G
pDbaX40fiuBDiY3Ajl2FrHGD2wUSZgSqneLwprdrSml7RNQ/dJiexS4Zn01Z+j3R
LHhzh5gQw+uafmadEIwWAZ+C3FHKSF5wy9e3EWngPza2Ucy+65wYiXmwFhpVqtT1
hkf6HatWRKyC6/KmysPuCeEfDrjM53eFzoBmnXS1RYn3pVamKbMK4XCGkcpNNw5j
V5kdN9eErwAxxGw9B/57BUyeejRmFNv+EmB3lI6WlpJlr6x1TBL3BELStXkJAlYR
ksxc1wOyyeHt/aZqKBkMiJS4hwHsSZYIL7jO40YkkB4VlUZRiqXwYOSDRH6vWwK+
QKURPhgy8tumpAtjQjZtueF/C0GvUz5VQ8TNayayOaQW+icsls3ZRxEtx4uUQAAh
gf6oIHcKYs9SDgJlICh+XOUNdxt3pImvP9n5+PCAnwEPT57LXgEY8n9/0oAKD8eX
DBe/zr0endoR703h3rgEKp6K1xvfbishkBmN7w1LZt5slrnax+e8JqQQtQkR2Jyr
D+aX91Es8/r3Yr1bKDgBDr9rHNSNF1HbV+9PASpd+W+F+6x4RNvk3DdVoNRAXeJf
IJhQUE7BcIFqgCYHJXAWPLVggk4RPdAWe7ztkGfzeR3QWNbj6SO5GtAJBUg0Hqcu
TkDnbZA9VJcL5MyzbWuhsd4+RyGFFI8KQtiJwh5YgKAUmp9ZfIYQuwxW42kSUVWz
0reLc7wrf2P1Wwc3zsi5TKJuF/dSUIwg6dMLQWWgV7s3AK/Bfadl4QLtZf8eLdnI
Nu2VnZw/4MqOCaaVefUfD+ybyw21hi75c7aX+Ed2IdzF5Qc5ht58bM+Z4wV5PffP
MaEZ0vpxNy5OEBGkawF8fbIFynQjpdI+uyEzwOZRG2Aly3WYDmkc2gqJ43BCYmum
GhTR9BmdlJSFhDzA/+3bpuWmB2UhSh5FvCuQTzOLo3YPe9IAh+252wfHr4Iz+jqd
zm8ibtqhXTFRMsrpKbHdh7ACaK+S+yE0uv/6KFOgdylWzOPng0NaO9Y/MWdFeqXy
df3DM8DH/u7Q4385q0Y+KzSiMLD0mJVJ1L/olthz9t9cB3glVuMScFy6w0Ad53GO
tpXZ8SkLfK2bsbsocqvFpjphfzmxSmur9mCcwtmt0cIro2zymEl6HJHBPAa6k3oq
r3u15befU8/xb/OrRgLF2rcD7YjmgjBsFfdOo0zRv6/uLSQOljM75P8LYQVO87q4
mYrgeexSgwsNHu4vzOoxo4rD5TOPCAbV5ajtAhndcFNIpTC6mxNQXAR4gkyLjEET
i5scLCvXpHIfdE1oHnPap5Ohbp6T7ydh9wJy+l1GKYJOwdFjpzYOXkGqtuR3XwpN
/t+OK3Snlmcdl2KG68YdETt8ywyS3Ztrx0AU/T3fQtGKA0MduylzQ39ZRJU5IFlh
VFHwSdDjpAR3bcRqXFSnNkZAaGy631ozswHH/PLruGNhsMRNZvxRgFldrmrPtLXH
J3gW4vc2p0Pp9jdBnW5UHvlOtPwcpl19KwwwZWfDmpJ9lWcgjwcsK0a1vWD7JmIy
+CZTJWYAm7C1M/K3t4ODQ+0SVscjUNXbqiTeH40rds9qMA7lJB8i5n4JCSWtFypX
L71e3FX6VdxZuGs7ypNRYKJiWXS8uEM2zIjJq5mTxc6cG0YLTJkMtTFjl/MiMdDb
NKqaKl0w1Og7s0ld0sjd6cJLvuOBAzbC787ZM58oPMTwt/QNgVfd7TfMxirz8vEm
BlzJ7Dj6W8/sJVW5bat8rQo1i/OV6HM7CWWKnG9FHTFQOefRctUjohRDbJqTAeiB
3qevfgztsMd8VP/FviFz7qmLiFsukn4ggFIWShYPWksraUB8eCLTfqxh/mQfj9Nn
0p+mN+MqVEZtLqVnwUErTIxsyt3T+I/GuISX1Ix2MPWIJ2v39RV4NOry0Oe6789m
f5Lrkt4m4OZXDJVaAb9MTQLQtQCaUbB94rQxxatLSZZhzTvvBk6hs/7+/D2fNkpb
fw2uD4SZ6RqLUpHOWJIxpSaMQrv9H8Yy+zBNxGvMecomold42UGe1Srzf18E8T1q
KfZ/jhs12UrQdvproyatKZ20mKSsTwJZE6F+hHleHF9qf+u5f25LcXSigx9O7I+7
QgfvQzH4DpbzugcvplZv8vz3esk7lQnU8OkWgK3TgP31xY+McW7p729qcFbur9Ji
/vsif8ocALNvYbYBaXegla5L/DINWUkY/11cRB/ARlhjbgD8v9aPvToQ3N+ipqOu
xbHx6ILgXn6/625pe4lqiitssNraoEMpN5hwA0K4w1TRynj+rsyaQXcYV3bymhpK
w3aqeGj2L7TGb/grfYxGcHdwRvPwT/BlNhgUVclT4oAHF/Buik0+4R6I0D89C+qK
3cmDk/a8pDJFfHuZCZEadUv658wVd546LOGjT7Iw2Oe58bJlXfZ+tRLke+TFzzdX
Q08825VpWS7JfytQr538rLz0QF6WbTc1MWM4LJPxxFGk6Fd8urGT8QoP/squUa+d
b6OLA5MKW5x0P77OdUJrCBDYAEc1WsYZUx7EZjN7KyDi1agNRpmb7iA2qd2TaOVB
txLFHUVgkGUcz3s32v8PN1ynMORIQQIfkEyYhuYHfgvSeiDB6sWVSnmlwEa9mh/I
GXeun2qNoxyK2aWnItzLa6eMdH+uUhrTkzZG7PAY0TS3r9im9QEdHYYWAGiPfZdV
cT16Kx01Ip/Iaq4hN3poiFPUCYWKv3t1nkdtZnHnsjjjeYaIM0ZxLWQgW1nHfShw
AiDaTJjY5bbUxtZ4b5gABUCUhM4fBRbwTQ9m+5UbaZq6hvBg6/DMNjCEgq3JqsYP
SkNSIDmwhm6SiPTq6nvpS48SxqC3g0w9Q+R9wj46N8qq1auTA0LJPIhRhkLrpt/c
86MFlSmi3Ops2f8H5/Uh1MzpgId6viRHUIbUFdDYaZ0XilGyRyxt2CYYFPXBDWBw
C0BKVmTG3C2ZIAifnyUzKv8gT8wgdkKcGOHU8PlxfFgEcIV6nDNlkG4X5HRDHCCl
+eU3qBWv/yU56IjtcxyeoRiumsDQGQhZB5P+WzTJeZgSjQGCMQybL7aN1MJxQCVY
sTqLeF+mBYfXF4o/sOY8f0Krd8IJdPLBabL4O5lIBepQor7D+p0/DmeO9aeNJJnn
DLEi1yTOUrB0da1dA3754od/lokiaj8Ka6jVR8sdszUnzBPLsE7DVY4xqkdav3ag
2NcHJNwGwOWiAsZ+X5QXYpiQ5emuuy7B92+lyxgAsvQORa+5Z7Ah5bt+Ew8qUTgT
8E5JMVV2S135luPF1maK6CoiLSAmbR69Cg0v0y2JCtMYrc7veBuahdUwOntpVGkw
+tqZrXpjPSDvln2OtvV1abHtyG7eSXDQa02qvGD1QmShKVm/WCTHpFBKRo8GRogu
fbrifkm01DxkGHct5ez8TbxS5KXXB7+T9ecGYTH3C2VcL0QsGzbfUzdYp7Sjc1/x
dYgswinBNWHkXsvaEePwJfU8wj1PnpQvWmYgtJgsl0tec2SLCE7NxGJBG2YJRLF5
5jKz8eEY6d2sOZ94VMe/t6wr+LYcokbXNWlnxpVM+zBTm/gLYk81vSYurfxe1cUK
m/iaXxcqa09bKSTvzTEeH8WKi9NouDoZl523jbxcrbtDiAxQiUhgJTVKiYavWfyh
Yf+DjEqva+6EcZ3vPQtTLZu5quglgRiMA2YSdOg1tMCnAeUh+/TqxTMNZCGf8xub
dGJ55yEHDRiW0Lk8bhAlzwbomtDkaFzyn0uTNdou9+SQ+K9jCIhZFHXI6yp5O1TC
1vc3ZVTnR4d0n+kjEUudTbWkKXaZGfYgDqKUAX/EmyBNWzzIUGYQkgqEvO5K8BVq
s7N4wtQgqbIVqe9eW6yp1mqjP2f/iBEv0n7UID4zentc+m+1K0b5gE4gOeJceKS+
fUC5H7TeToxavrZ+bLbkqPuDX+fmQVeAEwuPcCgnE4xp070VnssejWxJzhk66tko
jK/njU/5W3c5D8EIPfV2pEX7v7Qvn91rRIZl6lCEz2IdAVtvPlR50YZuNGsh8In1
XmA6T7HJ658ao1+uVEcGXD1/cxvzBOaigMRgxsLo/ASKdmnlwlAdPmi3VJeDYbx3
ZZq0KbzvEgmXJRm8/gyrdM7HsvQomihBUdyaZczYJ1kDEyf5bWg413Xr5Qz1LhFs
slrCdifOZ/NG0p3ulK80J/6ABpkUehPGNpk6VgA2giOUQtPC7X1dZ5byiSWIgxG/
ib+4uW1xUqMinzSP0q1hRAqI0t2hDbxG/S/BqL1zcY8FlAfST/1qd7ueP4uX9h27
FCMp/x0cecuxeMV+aRqOul7ED+iBGh7Lu7pNVd7ztlFDQucFCYB8tNxGBnIZyNt2
lT4wSc/YZOdzawy+nc49NyqK6mSh8P2DiW/HzcTwHEswa+QvHuSD5Wm9ENDLKOeS
FBGpSZMvgQKWoXMULV5Wr6dgddHJZ3kcw5iAs7kceKMIq6gHoVK1GPp+zs6Rylo+
uvPV8CwOyrkU48HDiYl+noQbYO6aLP4LgHa4+LX24VpPJvqyiJNgWOTeVIyJkXZd
Nqo/OQgY3Vak3ZqgCaaM8BPiHNUbpqdPjVZq81RpoB4UqoTVQwLHgHG+S22cFIz/
oWpLlEK9pqe97egDOU6DoIb7RpiKOFe6cNSStvnEk1y/NIEfUQR9yNgBpgU0Ncld
cv9NWBxVS7a6yMRxYowHhq4J9YUCRucU73ypE0HdzYxDx4+Es4aHk0934WUlAnoF
Se+MTNff7+hj6Merd7nnXk3fqhTgeaq1gxBPnJ5Z0qNpm0BNffdn0bOReXYp9piQ
8Awq7LI/A8adMjYcG+XiSJ8ZbB7UmeMnLLI/eyuxaz590BHtq61iMTag2rDcDr+g
v3bGxVNrdjBUxx/VVxjpGff+UbL9KTBVOn1GVgoeyVIkjCvsmbKV2p6S526Kzf+z
bD6vpOF/EaqeVgIsI/+gXLxqr7LOGcA89RPsEfoLN6zRr0oaCGTXytyYOGSzms0j
J+9TIw3+//lmgNn5tiPdz9fLPpY/cfl50GqtpgUzXdj5cQFRFVOWO6DY6NCiNFq6
XPyCnZDOUzH/cGIEod2hF17dKnSyQKBpRyGKhWU5oGhw8AXq5E99cKvhEsgU61eC
n4Nps2iFqueJfS/UULvhWlWs1RvB5+grlSTAqr6oGkG2jiGid4YewDfp0Uh8xGxq
IQUQp1oOw1UZx+rTHchVqHDw7aP1Fv4z8KvQyYzX9SLS9yQkN0Qm4m0rL56tOfil
8QnJCMvkWGI98Lpf+C/loSJ7JkjduSd7NuyidQl6PXunQYxA8q4AilM2RFjnutVl
aDPEu8wlRdpNQoCTr1mw9ZZUM1sr2jNn51t7kqcc9idzObWTVWdQnLOd5n99p2/O
0tn9YUlWchfp6GZEJFDbWAgConU0d/gN78pSnA6cDwHETCr3iOIJT7s0q4JLYzmU
gF0X+dEE8s4w14XrImGfko962aDgKb29zKpu9oOOGkm4NjBPjHUxPk7Jpfj80gHn
E9Tg9U3HVGhz19LaHzjJFeOxP2k2cxHZtmyYhOHUtjHSyxndPzUcCIVEwE+/7KWg
atqIN/SCuRV6ewlDCJhUlbFTkPDaMtLoIiIfsjQlw1Qll1WnO78OAL8ATmjuqEeZ
XIvIGTzz5zS0FDTWfhcTFVGvOCdN1e4tHSHYMh7vDk+jpn21fjBRR+9hOgYbhItS
ts4fokOx8doadOUGtotjwRqhWbJgud7b8AWZcOfgrdR2rOTpHwOgsp+EHC7V1u3Q
ZN1EoKiBTNTt4Ew4ZPjmvgx2JqTuZ43UrHqKWpRLhctBwoNg0VUoSeAcQwgKMOm7
HxEY0wVOdf7KxA/B0sVI2tyUC986NBHud1wCF03nuUermdaYx/m15m/pYitIWld6
kDMLxiYjTH9BtDUiKWI1Z+BW6jtcXU0N78pyvWoNJdUz7NsDXNxcl/Lzvh7kCXTz
kZT9CCS5zYBHYuLiB57EdmJJgtQGO3lxH/+gi0LAaFoD51nW8KDzhQPuGKpqoDwN
IPTaNpwFpuf+CXKtZ30MqBhBnU47tuwiWNFCZLNj/0NGmyNY2BwLnCIP9kxhx2uE
o3Y5RREoa9slVIVP2ScPDbQxYTXzlJ5u5aIqAxawPZkt+XKfe+PXi+r2pjNMtynX
xfOa3vF9dq9840ZH4MSz8aq1MKkC0FQ4zwXu+gVSvvDXT32Or/SMrR2BkoXkOI4b
57vBTczFvgID5a+5csrxiFWVipI0hAnsOWTxotCeK70zlM7Cd4aex0hpIfIcpptf
hEPgxyKULomTWCaxH1iAldeQIAyBnlM7mmgpjTIJt4kRR6vLQzTaN0sGsrhik13L
zhO9ozXVDkijVgeTC3m8xbbXiXrBsfCw4rpnAaN34/TBEsfPtgziDNdGtsQyAPti
PTqeYF5Xiu7fyWw8wMJ49HBkybVq/vrkCPO5TtDBEqUFkexzo5Hx50VVjBzBuGCm
B5ujlTVLGFuWQQEUUfKrxVaV5PngAgXRwpGmlLIIBPmmyIyVQkagaWDvmKhP6LOQ
MqkOFwP1+BV6ZPOzO4xRvQjYUr2dyJ/og2ckMIycHfjYaPgVgB1yh2xdRBxihs8P
abU6vks6HEhtvt+zkxhVHqicFbsLAo9HyrhL+e4Vlk2Q0tQ9FWxZeet5IYmaOVvw
ZSgTPYF+TQeJMYIafRnMObdGxAnIi206p+oxqoyxrvPB85/wYH4ogpYtw0uXQ7h+
OmkrGPAkv8N5AfG7vWE+n1SpSEGpP7fvqtLUbXlx+Yfq2t/qr/K/gfo+sqr/tywV
GiO5CGTl+ar4J09mIZV8aZYos67qSwruGtEQUML6WW6LLE30r4xXhecyBK2y+G6/
WPRttFkVGV7x12XRJMStS9aP4ykagPKQlYdAITZXq/kb0MTmhWxMxRFqspt9/g7/
zyjL9Olxfb6GRGg0KSGv8AcGnTDwXNGnX9mwAvUGTZQiUprBrv7Zlhu6IGs2Ma5/
WqEfKdpj/J5gnJo08dSKOJyqEfh2MpSsCY1PxGTj99b5Fp4FmkCdg5VV4HjoN4bV
5FO84kZDEM4AHbbtSsS4TgGZNs9+8jX7cPAz0ezhzjbygjZ1ualmFkf1Knvyo5Ri
f2Pcp+bdGK1C3gJ1LVGUhpGHslfPFDgi93TcSsrNWpwD4eMi3wlLJuB/RRwneOih
/CezEYCzvNKl2VFXoeoY0rzOzb02ctss3COhZ4HQceGCHK2NK1IOHOg+aVsCogU0
qsjkjZ9Q/IsFnHdcqQtgHApjPWdWsBc4wO9v2CnMJ6fVrHVgaSXljP+ZTcCQ2hn8
ybEukIj0mvY15gE49ijdBsaWWrCxvHykT8XMXILxKtx6WK7geGbnn7JooQx9KM1i
mzGxPDiKJ2qGTIK5wnOjkszxNpGFT+3UV91GwHIjKJfVcTppzpR8XTLPvksgYYgs
cOwNvMotP4B8af0SZ30B1wJjIkbwI3EGGu+CvmGHUDgSoBg+EorCk2Ms7tnZtUrN
CgxQPXLosBnqA7ivuLpvrynFWJtnszCmzNjeygeTZTwieiWpZexJpszjP5yGsHiC
lIllZsSWTJw2DUZzme2GUYgIaeDF0BX/YAzSpYLoz44BrqubqZw5CGSbYzK/KohE
PyogMGYo3+UuPAuMh1sVi29gVxIOArqungV/s7yKs7FLJ5INigsrd5NjUGVf1LVF
3Puetm25N/QafItj1E0x1Tm/s6cxfxl2y0hGuv/nuuEbOujZXtYTGF6VyfDveRkc
Y7jlwQtMwcfPUELV5Iy0U4WaurfoLZRxuw+LXHOO03g03FPnd8ilHQiCpYMPSctb
nl0qzUfA/g0X3VDyriwFzQoVkUgaNvULInmZme4YgLsB7vrN/ROxCpmWJk3Zg1EC
a71dEe4Bh51qg7WcVVhRVI++ro9KOII1UGxv3IPqqqn9EsqDi9qxfS33BuuWhMpd
lIgDEHMNMcsTDsfm41kT9moKqeLUc+FKenAPLirLbjfG3yvrX7Ua1072lVED5ped
0BxRPyj5+QyLIP+wMrPFxrbiOKbfwV2yy2PWOEtH5paivXPaJY+8uz08Xg0q/V0T
ZGEbYvH3ANEpZL5iqhsFYLApGQaVaTo1/P/0nqscOjjUKGisTznsENSJ8lB6Dgk+
TSsvNlOSG2q/hMTfAI3FJD62kqHBDUfKxIAQ9a7P4Q4uGLVeyDnA53xlz80LD9Xf
n/tUIGEkyQizYwZR7ysFLtp7F6euoxIEhGhgJZrztZcmvMuXH1r9iDvQWTvGeoPs
IrVhiK59B0HdG0DBaiqybS4cjIBdEkvsT0B96cTeTNGjnCPNIMz80HiCw+LeVpGX
drDkQVfRLC6q7+p2x6cS6n0JiQuFPSSd8ppNpOWsEnTGDyyqkLZgDOICZ43Ot+kO
KJi8z0H9u8v5g68Zbms6pjyksw4VFzH+EtNnSEk1ltxuAkgnsYUeWH6tOlsG2jT/
I+adFHEihb1kbZ4NJSt6++2dBeOZ7mvQM+6mDCDxJGmAnDI67bSEmP0RVGLon1rT
LpHDg9NY+pf1wzpzOxvF37xcOGtl4o29BqTf7shBM9lc9C5lZ5hosDLz6cT7uky7
foh0jwM9lOEXz7gNMdAIZJWZi6dwDNknZoTJ8GoMXEAKmXYo/rJsYban9MXf1DGC
p4Y6J/qiCjnmSL9i2GMBXkf+hAnlgfBphfjiz33aGlgSV9GgqeiOAzo6JAcIX7hv
l4a4MiF9P8WNv/eOJI7ab83IbQ3oc4iC/WtbEuyjsAZ/9dPmhUJO+kl/dzVdrhfb
SA1eq7UPLBOmP1qoioFCD9yCgB2Zp9BS9r1AS3l8WeX+168b+QJZEPnMtX5qyB76
Yo9eAqV0gvBynSWW534gTpsC6lrxwwKlaR7Eq1ilshnzfQjARB4T7h3Pi5VucDr5
iJvcS/jDU9QzBCc6Zw4qxk/RJy8v5xdAgb8CdoNDWe774AB/Dgpzup0V01xAxVql
Uwac3j7v8z9FOrJkR9nxy1BY+NhtjI72e8D0FvpZyW2tg21QRdTT6yxtqi9Q+l7n
rYJQo3B3dZdqyYRPMfUMi4XfZo5vt7DYA8DhUZeliSUNcdCoZfFEOkv0evQ0dE8e
jEFqpeOrcwMklZH/P/aAqvMn9Ftb7z5zAE8aiCh7njhZI2Ms4w6VE6f2Yl0F8wnx
`protect END_PROTECTED
