`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eyVyf2co0tu27exbmCfjs2wbSsqRUuPctckC4JF5RtNHnxNG6eZeaJKB+YYvcZls
BV1r7iEMic9dKBz+ypyng2zPoC7O8WLeX25PfmyxPg9yhAyv6cONO6/qN1C34yKd
wymiAEvlvX5VbE9xJWKdTV5s+19vPZbaCm9La/+52z455fREZrtGnjSWGBVzULCX
ClYBh+3zeCEfKnMFoKStXTqYiBPKUZ8TAPbLmrZCq3zQpVQGXEiPDCoQvzjDD0Sx
Fb3c2q3XGs8edKEuqUaAA5Bh1m0kylHvY+jZaCVo0hKy5TN74NheymCz4cJh011j
F/E5RFcrWGUauNJKx3GxaUAbgnXKTxtGLcdZWBPAmMLuj7U0a823wXog7PZByu+f
47TK1isu5HpvOiCd6cMl2bPKuJO2YHyxppaEIs6fvx+3+aMPnWiY48SOL2Djl9G1
gHr1yoPJHag93XhbNyF4ArnF77atRZ1+4VPKaKhrBdWQB+LktqlT00LPETnBs4kZ
`protect END_PROTECTED
