`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RpW1KBYna8ITf0fhzFkI9pb0YGXvvHitiXeEH7JMIZ9NxnrZYjB5U/DVBKhVXzi8
WWBGFVswEucNynkJEoLO/HYiZ5ozC+l8UlO6RM8rGrWST8XnEW0zXtyL6dKwxfsu
no8BRBvPtRsH9OnHNhEV7rFkm7itR9Bh3AXffmROS9UzpLaOovIZQ1AOnbg7V0/I
e6agvWMf6Od1yMGbZ2Sb4d66/Aw7RXQk61+IkGJWAmkhRWLiUqjTvVDLiYrY6P0H
P5S63WcXWtG7QuICTry1O1Li7aWThb9nzR027OaLBcSV7i5W2hcszewI5qQng8r/
Uw925QUyTkoSGgaPHjQXe4uLc+Ik/HJqiviuXJ0reUHTMCUeh5Ycj7QASWSkvbwy
LFQGscem3DHCGuvtmJ7OcUT+Swa4+Oi4YsqARaIbjas1dAHLSa2AwqSQz4PTwBVU
IETGW5yfnf9B7EyhudkE56uSdHtxSj3jFjLbHqzyxWXv41fiMzv2B1MHyuGqF545
6QusKxlp24AZQee9MZu51aUlg5xRXO63yswoRKz/SFP7mZPVk6SK4mFjCCB0f4KN
ViqAk4brzeAH2vtZmSbhGnhcykEdo0We1ynqtXzozfpw8lPiyGt+perXAbRngaTu
xR2JGEFeMiU3aMXYhPCJjJW4joTyxtfNG9aFecaFyGM=
`protect END_PROTECTED
