`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iXjU13gm3Kaic0N7q7/tyeTkDcj/qzlayGcOPEc0wW9ID6ADjhsXmIZy4B70G8SY
fXY9IC8Qha6IW8K0nqtZ5P5dCpnIQE7brijC5PP1OsqkmQq9IXziLXrZ4Q7H0Mw5
2XnAMjqaVHoaHrJAYKN2qiGaTConH5GU66o7lUFbn1o2swO3HOAoSzj5byGJaFlg
EXgF7u56+Sl3e3klJwRUAAlVkYei3K/FamaKYaV/3BRWcHWXLueRaLyvcy6Upkes
3jsOsli4rh0fL4LRCY11oDKGy7jAoK41SCsgQChnf605koQ+UD5VKHtbyJBD/hcr
Sdub+KA1eocn40JkMXSOj2gHd0R053gPvbQYgPwB4FnMcfT17W4a8cvznODXVi3j
BhxeRziuGvEPP9GMordKNSazyZcpSnl96+8ZsujNVeU=
`protect END_PROTECTED
