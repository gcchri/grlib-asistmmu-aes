`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
avrc+WsKdvtFCF7rySmf8VJOiUZd8pWIKhdO9aIcVZJD/OYuxkX4jjn2OZlDTnSR
w+4jglq35NrVhSV8k2Y7Ph2mUuLhobFy4PYsOfDBuIdr/wPS3+kh9EPxbPyQWNdR
QDp/sgRPND9DWOiQyuXP+Vjz8R+4o+7TjXc7gqPQF+SMz3ShppNcOSrymHUx+/XM
jlD3dLUSSj9fNOnuSNF4W1OufoUgwvxtp7uppUBsvOHtLigomgdY/v2zUQN0h68U
Ozhx8oW7+YSG4OFoODcNX06J8a/k1T1tpBMU5QmZW4Bhs3fM6kE3O4a/xZ3Kb1ON
PKY8oI8WP5/y9q0LRNPzfIMgjGjqHOANfmdEPecvXBJc3grRS/gPgfHynZ2lIcZY
PtAFKQqLOlYJr/NER2b5KpkNmvjYgI+cnppAb9CZU/SN6BI22L5mD1DWLiu0EMi8
xP3GgcyEmlTlLd/r1lr/Jb0EJaxo8QFgxdvFFSjMHKpC1DV6llnL9gzCnmgmqRxD
qC9E6ZDRaeFN4L3lPwvzeIWpwHjs88wJoGrtIkitZnlaybhmPcDvC2UGUgHIQzpV
J8GG8GnaVQPJSQ5+bZCvr9AUbH+zhnifu/nwCPwic1pvD+U5unlT0BRT4NORWS4H
0Usz8apOIJCbP6KkZ2+Go00NWHYzyZtrVXmD2JRD/VVVToyC+sh2EpkHRqwl9e4W
3fGbmqAww0NT1Nwf4KNI4T4VxHFkqvp4UFPzuE7SD7qsf60MLFu0xAihQy6t6OrF
2xG1bb8f7z2oTehRp4TOioMu14JUzH3UZJRosVi3HNrrg6onzBPXx4KdpwSUjOsJ
yZmMA1CS42BALAzrZ9M67LtWzn6kdb6VZLdPkXin8hp+C4CJN80sl41gkbHR8vvm
t+CDxldv8AGiqs65pDPH91I8mx5jF2VX5ns6V108pWGKgWexBrqijYGXFQ5Ju/fM
g0u6nSoDZnfqLjNdFoUcqeypYDWDCrY4zIXQP/B3OKma3augdcppGUaBql8pSIPj
uEMcnWUiPgfwG1VHyshX3M2DwuX5MMwHGCsZNFsBP8VlcjWFfDW5Gsow6Rsl2f5n
cSZ/iJpKM67tCzuROqb8fGIC5OPIyQY9YDgVwGPT6iGKbOWGi2S48AqY5Lvryua7
QkVTA6gj1KQNB0eI7yWkcex6C25UgNHiqbYPhfsZwSBXUlH2ahz05ycT2EwA2WsC
4OVmyVwcel6lkMSLRNNefsV5K7XqtU15mrtewWt1EWEKqfNjlcBWqEbaT1+sLbgH
tt4TbDRBFNl7OJTzvYv0M64Q60R/WJFzyE/qYQWe/7KonpI9hGkECzV7dl+jCnh4
p58zFO+j7H/YIp8X+0ssTlOwRZvOVOL+Zu8S8TrM3wMw34N2LP1iJ0V9cs/DhVYq
se1tmaaTGfaixxItz2LddEGdUuaEbz0lOFVzP2Fa2NzClGId2BcsUwSdu+oLpTBU
F46Ivu9pc2o4nrLf2/PTlqB8tF4ygqySLeEyTT/i7Feu29LCY1P5l7PIDTVP5k+A
9Gi1X9TCca64x876hNUT3LhFHO0U3OQgvAHlcVmdFUltx4vnlI3vMksSoROXdJ5S
9vyO1e01jUz0Ojfs2D2SJqpr5Xq032Nm7toYZP6Aw7Zm8Atg5SwHftduGRMVZ2T7
Nq8gLN8szj8MrX2eoFjybGsCPtilyjd20WCWEZ/1dozXv/Ei1j2AVFSwNRoTxEir
5q9M9lDVnZiXk6SigWAPWl3o46uz/aWHOZDMIhgk4qfDeMMSv4yX3qljzKYD+x6h
OerLBBRnTD8bZY7yT7qHNbeyyeofXi7R+tACo5b1J+UP4HRTSv9qfAEDfPz/sSwE
5dOK0/Js/OHIjSES+yQ1bGPkUu68YWFp0Kyhyq5f7x97CCccePbN+zc2TRNg03ed
m/e7lFyvccgCuRAdWp5yErEU7qmnceayWV7eW8yxo797M5Y7/4Oz6hFEfj9PUej4
emPZNMjmG6UW4jlesJUwxjLz2+bIeRj7SpmJXYGvCJyK2AxcHvoewQAzDguqVr5Q
orevKAVP/X/XZ5qiqgsaXrApviLtB2X4g/a7qto9bz2V/Wt7idHYHdCh2tY67863
YLgnITBTccYXUObo67SUqRGV/uF5evUXypKvkQzoKpMh5hyjHcbAxmr5Ni5He/ry
FtrsTO4cZN9rrjQeLazxsMw2GPatQ1OnN762Y7ZpI3khNmYuwRkXfCgQGNCnkks3
ax+uNJaWdQxL7uR4toVM8qdCgKppa29QAApdkuGOvKV8IqN/EKUGO+Fm60H55Uxz
plNjZs0DyzSGfB+MtnyEUC8U3rmyRthrPavcaU0z3L83RyjwKT9rgvAFTHFsqsGF
T2S3TbChFwXskIJxV19IV7U3CWHmtU/wR7Iat+qY1OcIXU82LzU+/qBQTDnF5v/7
wVI1DD/77TfrGqxKqFCtsnvTlzfiHcM6YzdcDVrpXIvIG/d84XKOJhM+HdW6+KJd
odoaMSweDtsE7MPCgu3ioVJaJ2SqCI3p9moid8hirzITaSi7ffrK3EhcLCa5GHJ7
rPjjs5gNxBRT51mF05UYqjW5mB6XYlfgYM1QoljX/znKFC2PbuXPKymuFuuvrtY6
lv00lNwWcTK0nBklHj+bFXBANgiKsR3w0raSawOzaac0fjiRl5K05hpukfov+2pe
Ev0+Qphyh1yyiMX6Sya0SYooFpmJXR/jxTnjZzd1hhFVgbNbQ1cAsM+srA2+Mn3d
KvZ6/Sg9/3qXuc6zPGTokfdHKjHFEiLzIorp/7Q5KSUZP2EOEHOi7pD0XAfaeawy
sZt++zX5/O7BgPqwW+lSc1EXJVTLJ77j+u9PmT3JEZn7wSwB5WgVULI8dPPsDEuI
12LCov1DEoTHwvMULXDSyepDT4i3bfHM7QIfX22bT3bQVo1CmPShHqVRctM5+VeO
Ll6W43u3PtmFpkpZVJX89nFWkB6CA/NIzStflq7J52dMFgLqkrd5+5DoVD7wiYIx
XvMurer2EeuhZvUWyxqQy0NAP9O97fKq6qlsWLWKZCAP1cf2dDgbNxmOZGuoTMcL
F+VCHZFWgqXUMMFT0lCEU8h1WZVId71Xk/dpvOUNWExyxjY9yOPZ6HwfhtDDUc92
KA0laag0g5RVg9ZCBfcxHMs4WSgDo5jU2ZgeZts9x71BpzDXJ1TNi3egAJVWCTI5
wrfB7F9wlPPF6BzBvKmt65UB7BKIRiAtgNcfbxQTCTGWR4/aRYYdhh9bs2+ERU8s
/+jAK/hXIZoAIDx82lTMvS2ZLIyh8M5Gnm7RWPHAVpjt8XodA3fzHVt4OexpL5LE
+K31LvKh06RGSUrgLJ6aWtxu1M+cJUH4e5egfLRt3xDCYh9MJnHNosEuOMBSD/g/
QmkEvcMDGUjR7l+Q7iGiqoy+kX34Y0q587Q8au9dzFkuXVJlnwycPIF3pFPf70aQ
drUVpEphi57d1WM0ZRzSeza45SCKzFLiMmyk6xTbMd0ZCFIAXNjeqsT5eOPBKmyV
pKHmc7UXf0TjIPN8FschJkTMKYPZHErjFmX13YhaF8RCwNh219QccIte0GVJU2BA
s3ZQu1dcRWvd8b8d1JKfL1en8LI/H2WP02Ks9s+Mhr9ExcBb/VNBy9AqQ5ldsaZx
e/L4BXhpQdU1M4NS9PBeJzBrIL0XeIA9BsknrNWi23M2ZjAGVhrxlmqJKYqi5pkJ
MR+YvhNe/3/dbhKvHx1g3UUdwJ2zWn7pgZIyHtE7oiNg+x4CLYTrFYKaa2O3u4qx
I2cwgVQNP46uBEoyrHDeuDy1x1zaF7F4wmscAKt7YznDFsKRGfhtUnpgtkURdD/x
/M+HfLtktYIhu/+QWtnwRKVeplkyLIbP/WEd4UUu1saVVIHBIFVEhuWFz8Uup8eV
YKIL333f0ap7fRAy/nU7RDjuSTLTgxworBPttoasiA9t8/g79eYQ6RD3NJzDhmQU
lUv7suugi6vNukOpl/ffVJWo2J/mMurSACs3IsZCE0L3pQkqfGtCBc872MdQo39Q
NZOmC9YETKmASW5WzqoQEUJXRBvelCUeGyUWLwCqST1UKyP+c+rizQ1agEoPfw1e
wWkhYK2sHD/XONCGEROkq4vN6YvOYO3FqYSuYVDCeKfsI35BRcKYaV8JhhchuXEm
NMI2XNPQPkE39X6ocOYIVrJVvMnFeYQuKhqUnXzoNgEOSvpPmKmQ8IsDY2VsSxmk
PMZL0HkotSzAEidysKXTpfxwKKrHMM4YpVfiHdA3XmZLRueMVn7RStE1mQqOalUS
qdADMuvcED8E0a1nMqhJybq/LMNwNRzA46wTqIo44FTSViY1KI7+67HcGalal6en
HD39EbKO4uv3vVnN23f//flZfVB1oiIHSkFTHIwqXZIH3BqPX4mbXD9jwmHH0bjp
Ja+0iRMxy7rCyQcA6YNqhYN0blysKf7RR7Yx3XArmhvr6EgtLRvl400RkjtjzvNn
asLpAgLdJjoVYNDFz9JX5OhYeCf2mXOuQaGC+Lils1YiebMT+Z/aBP8GnV4R8CjS
uGj/KyavLq0iztmxqwznLIMrkpkOQzAOBxGGwiNFjdIi0SVISyXepnMt8tR4FhBG
ECwchZ5vZKbxBeT7s8hPm8RF4Mnw39/IHWGFwps2BAa2cxqoWEYu4gcdyFNTO6br
IPiR0qHAnEngYnwaSNN2B790iiPGSpJtbdRagS6x53C6jay3+pyv3MKmOzvVYFa8
F3XyxMBPWw/xrlk8z64TZFzQXmkXzSlMze84o2M4FnUK9pc1XCGgk4YvUcIHq24B
ri8+IBSpu/wQjiXyMgtUPhAylarliGo4wVcqb8D5r9xrCc/8Z7TCpw+NhCGgcR4W
Ivp+w/LXxZKPylBw5oo/R7TMB8lUL+0tj3F7viuNbGmmS3hIY+fPEvAywhRyfg+J
Uvyu6n8gx2fnPiY7Hd2q1Zcw5c1s35Kz9DJ4nI58WVrcMTwKNLxyxBjKObv1X17o
bYqtVa+8D4/7bbMiX4df55x2y+7uaACSEfen6dmTUz5n9DmE0y3tIDrcuFdvvojO
VP8g/lG2Q0qxYBpWslrNsiu09e4PDWXxRYvti3dQVZY2fxW+DeSy/XaX63osDudg
TYikSwHfAxo3hY0bWwcrgN44WbGPdbZ4SQRjkU8sZZbP5IjuZQWw/AKKnxo2kyn/
a4+bPH+MV/Oebs6QsA7ZGdYELycEPN17PMRYxELSQj3//LAsaLbC63QUVRYuhw/7
S25D6VP/UICKyC9aoD1tXy9bF29PQI6QcAXOitBsp6Wse9e41/YjGxSzWC2xUaxF
reLkPLSRo5btyYbWHwDK3JGsI4LZINc7gP6gFJPllCXZO/rbUgvVqIxFp1Soglra
LrhmUQyqiLjQPpisJrxgty2EJLnNMN9sVnpsf3SVIxr0qic8ReB3lyg1hSREuRbf
wpY4bhxsoq2p2Pn9eTj9HYzJHM2O8dKy13wLtmkC10tLiebu/GXDO1lnuRHf8V0l
bJG49Dpxpn2FHGxVQBO6pUt5E1VdzkvKkLyjPCt/4zKPSPeEBkKf7rqiuoVQSIwO
C7AgA+2KZbVWmaNtey0UNZP8hk/8jw0HMkHm5l3Y7IDbsZAV8ryhKrNYgxtA7UaD
uo+/feNjWnwKGgaOvwkdJDUQIdDJvVY2Jbec08CHFe86CclCz10Q6enMgiOQSHPi
w74pgyj+AjGvl5IX0eaLUa+l551ebvQteYyQGHTCsrEUMUlRHkHjdez1+tURUkRO
znpgLETXnlTyYOxTAi8UOfun9nei/tfKGWu7Y2KeIQem/ny3xY3G9fuF9zanj/nM
PE6cg8rVoAnzz27ZbRNWke6O+d4LaF/U86YmxXxt5LkCnN7c9dPrhiZw74aX+CMQ
cdcr6oYIL9NyTovUxB/nb/D5+cGtPZX2hkT50wPB9VBwPIlkPpOByl4LccaAEzRa
BnZj6jwiPjj0lsPCsO4JRl35ByAxGtIh2KtwtrCdzvVXZR3jdmEqMINSheAyA4tD
l/uE65n8lg1FY8vhDuGQjq0SbGSWGPGA6q5YqkBhKgJFBfX6Qc23mm/o/HLAbtpX
4kh7yqwLtsZ1pA47d8rOHY0C2BFU0LSxq63RqkxNqTU0qQgI/BPmE7hhyUhbyjfH
5rQdP6M5ald2T7UOnI435ItkUTmqNZgkEof8ZCArtjZh5lj6rsU2h5/I0Oi6qiaA
VZ4zE+PJvOwf5+ucmlVbc7289z/24uDqWpzKxZCdtJPqkCnEVdDM11DVcofDb3ui
06rCbU+eTbitI4onsBel/4wwvDLHRAzwQL7AUUPb1DJ94rPTxaDK2dD0jL4yJcKZ
VSpEaCLOu9CydFz637+ws6+YlScRB2+Xf2Xtf0Mp62rHPMWPTglWDcgh3maY37vf
p+hqE6Col3TcV3Di8pJIkCZt669qiWEg7pr4NDaCH70JzepniqvNCX1CA+uN3/TP
rDB660/+Hem2stxpWuIbCsNczEqX6QpLmrUS4u2QUlqFwcSiAPDf/WPeoORoTaUD
+6xPncukd2w06JSwuvS/Jag6bWjRzBlsQHBx18Z5xX+sJ2az+Wub1fxgpDTaxl+o
tJT1e9H/muJzK/x4Tts0kxJL5N0J+PLvgRjV3m++lZlJvYLSYg//X0iqMaKZuuMU
60lnbYhIU9RwglLh3jJtrkRd0uGk+0+zLIegDH50T14SVVfj8CEHy5u2qRUsB/7V
hh99PPJpP7yZRPbFJV/3ONHleA+n5HpMnfyR5ZL8i2ReLBJjjaIAmXGTvU0iSpNq
45IQGYNMv1MTGWW4RQ5LXeBcU81UKpAM9sf6IhrIjpp+F6LSqqYl0hhNFNulFXaU
tlEVzTwM1Uwqycw6kJAkOIMui+B4Sm+j6wrf7hAlaMWlrMhcy7TkBFVEDzFE9Iif
ZShwaE7tpsOCrysycmEHCDsKYU8YtWeo6MWgLr6qqewQHZr/Q9e/K+DOTejYvP/J
85qVj0rqNIYB5B/0e/vzH41Ij7xTAR6cs0x6aaLO8CDCHjPnRo8OP/oo94bgje0p
whgv2w9ZcsIxAvDhjZLV9cFijcLCuntkIr4h5c1BVc0mPpCL2Kycdk+vUR69apGJ
BS51GajdIFwL254AUkN1Q0AoWU/saULB0W8gZhjrZPR4p4mBx2fvZP7fy2EtM9nR
aN6bzK/nCOroFLGARLGUWrRiJB6YH2GMKn1t7+EBNb3euKkTqsr/reaEH99ZxaEG
F6dX7rtNnFLxV24TCboq2ihH3xpg6l/e5qsWw4WCGwPtyxgIGcQzzRt/wlXIgCbo
ti+WS7fJOOkZaPmjqhVTSVNRkZEpA5wg6pVYEr71irmP8UaKVwGNb8Di61xj8fe5
Mw4jeNQVeGSxFa2pksaFPcpl02Mz7riVtYkMyR+4spb0Zoq/TZg7m+SCWVr6UlEy
+fWuI/gCMwcMgvbOklgfAH6gePljliSXdOZ5rcr5gWf0Q+vMFIk5C1REDMr+6vhk
SqxYPUhEiI5ZkPKuoVpm4drFEclabEcfbig0+To0n7j9LtXd1Vocn6TS+SRWtRkO
K596+q+SYBalCUxVhouYny7ngg4/nSM423cXeGtp/BK/MeTeidCRqT7enkRuJGv+
Y3qoLdY3eUsGXjjRUsBAQGmSx2st7n7dDuPOZ862efNs906kANwZt3+ic9Nga7KH
7Bh6PDcz68GCE0WOfWh+evM1Muh7AyBliLvBuw1xG87Rjt0xtSzkAyKLDb2ggxso
o4g/LkKKeRE4uNWTliOct+zs6gWwfrNvscbMutZUcFU/838DcxdJJgunaBGF1yqm
RvWoji4GbROOPw0ZAXijmZRmrNauCOmlEXhgfH9/WPwq2z9wILJhfFq7lE3ZzDss
IIZxz1BOsH0C+31dzlsn8qMDVwJGnX5cI37PFUBzgLyFiQGxfUQWhE/vzLjcSwCJ
gy1y9upASEuY76BAbeImJTSfZXk50qM+JRsiWR8BDYdgqMRcQuzVcXMo4kBUaQQw
h0j3OK4gCQK/XDoSYg2W4VoY7w31mgs9vZdtkoK81hWZkTeP97YEoHGc0CdSRj3n
Mv5JxQSlBTe/fhYITV3llpCPa7ttQOH5N3y0hh0k+Ihc/sPgSrkULQmD6nzysfHO
8pX06kcmUol9UhARmufhSyvzNNOdAtTAch3L88KRReAL7kfwbZOc2TjVNITRl7Cy
Do/CEE23mv40fBwl4A2prSziLJl035jcoF/aAGcE5n5O6q0KT+3uBt+StEMwkvOo
z2Vl7wY1P3Kwoi1MoFlzdaAn1a+hAPRv+agoDMWuMc5O8GWUbisQnKvdSGLtEKcQ
l5haTTFM8mW2/wCf8x5w1UtqcqOr5IysShEz+pBSsJi1kVZMMLzyMIY9s0iJLQXx
SPB5W4G8G5rl8E+L7tla081b/s3Bv+YECmbHkPXLOnBMl1BMSRtpQmOpBSzIuRwd
c9sDoopcf3Ywx+clG3iblK0wlQgb7O3anw6K+ElZFhxWc9sxZ77zHj8qTGZBYV2u
OrgwhMWjP6UsKWHjuOi8DggxRlkTh9g5UaO2HplPvcJyBbhRxBamBDzTT496v1R+
EiSwWzh+kQvk5F8i+FFyEiyC2SwyRukPvDomM1/TGY5vGGt500F0JmckxGhSAmhr
DhiLMV9n2wFWZPRaVgpEtYxDZtotB06tqXduSfGAaH+K9pOJj0S0Cu8uRyHbw63u
RGKf7j5tD+22L2fixqPK56X9IlfSfhUkJt6YnDDHurxjBuYCTLacuFrHiYuxeTT7
MNINxN16AU077bxMD09l5JJ3YyZIaPZbyxmaLbstzsTm2DrY63t8rz7qem8pbrU8
R3O/Qqib9UPBnIgEATk07A8FXomsrsmOaBW8N300t/6jM0+RyURpsGtontPnDhka
2vSYZ90//VKGvZuJwBxF3UpuP9/C3bDDF+DC0ptukFCGbO0Ww3Vl24Z06CZ0sPb7
NJPb6BqOz6nCNjql7TbTYGGiK85IG4UZUbwbYKwoV6z0Z9I6OnOLZ1dTzLfARjpV
s9K4Y2eUJ57Jz2xG80mDvKV0/ygAUJ/TGS9Meh3YBdZQc/BlDbZWw09oIMzBh79j
7wQxAtU5CncpZ93kf2BFWRvlGi33LzrOBUO/L/tKOo+hVhAFiZ65Tz31PaIEu6NI
i1xZFY+bxLMtssiFcGwCPA7chCjD/E1ZHs9gQvBkPo7r+y8C3hsK8GrkcbnMDQTk
K3s0f/0uL5a02gnQrOjek5/iUO3qqlkS5ipnntg5P21zVKEjVE8hOKteDu3hqI4X
I8RnZO4cJcjOiPMmM/seLLD6FpDuQmcI60f7Ki53Yfg5DlBDL5kJ+Em/hNYka36y
4xuU4yjOQ/A1V1sgx/qLlTMhf5UGAfAK3VBJOHOkPJqi318J6ymu98EvpXWHMiPz
cG0oBSvTpHWbJvmQ2MJfgUoNsLN7p+EiMxOYnANsX811a0pKKcOgDSfY3M/LPPuc
809XsGSqbT79EiPIxRBcTdHZYIBoiCVFTZgZXOmVWZ9V885EN5JBEUJ9pgHz5iw0
vNWxBEFuHsD8zhs3D0f34T5Z+R7Avgsag13xflGyo7415aL3LfCRQ5HgGffPjENe
1sHTRfCG3865zRGdq8o4cIxDXDd/QXzy43mFZgpA9DR/wJ5D4qIfZNkveor4hAlA
aAguS3nO0ZwMsE7ta0YZS+pUvU9WGckFV8WHJ+n5QmyGPvhJ4jZf4871YuEJGdbp
7gKAqTbNJtTpV5HIOUv0Tr3Cih9LsA2lNwM4TMdlATej/dVGUeeezIB2QrJchFTx
pNUEJmpagGFko1B4uvbNm5qqZXnORDFicxEvNyr/tfRy5uD/f8+xzQ2aPIixQ0DD
yP+jE1tS86UYPg5MQTX79j1Vi9HYmD3IyMQ25JlsvFeF/C33vjlJ17eQiK4m7iz6
oh6DY7hlV19sXACDfpinPYfScCqEiy8TgSEVehJKaRsHWnJ/fhZ6OVPI6BxWLrhs
xgjJSIxLBljWTAl4HfxJZo/MWUpriFrE3e+nA/PSR7tfeXq88GueYu+FIYj70h60
OG+kizG6awe1+zprjxSx0inkkZQbqzPg9IZQ1JrdeDqcTHbttQkO6Jj/jcxHnxrd
IcQ1vEC9JEF2GJwdsD9Z5keTOnxPmHePImPxJ3Ll30KFgT6S+4DTWweuG1zYeMtf
mkwVYIiidjggPxUdk9Dy751sob22h6IKz8GJZchl7a27siUq3wNSV0qSM51R8dJ+
LPIooh1D45BZsXmistt7DcJAy6gkTqvcyk59Z5ifRBIVoD5bBUpiQHLjPMcFmWrs
obMfWYimYvueoMctA74r9SMAnq5c2UqWM8DjPKQ/sVFtb1LgkbzKpUAJyaOTzpyn
QzNv+qD2tZnzEu5+4ayfOG4BKbgkrjqh0OWV3wFcuAurFqByewDrE04IgZu+X6LG
YFkUQKX5g/bMuGUb7XKHaiYYSSaTKWzKvIKodoAS/I+5a4Gv0CkZkp1dNYdaF6+U
Jn1z7c/hhkXmb/eTXhhzCmfo024d4WDi6NyFMiybd72/XNPW8psrfPCdFF15hO5N
y8GEuMd5ITmQc0rfuYJ3JB7RuZtU0fL6A0Kk0ETXroikHYhEr8ELKmYVJK14fSkX
nGbGQ0+AQyMG0r0Cu3fRVfVIZZezLyHIHeAMPW0d+beBcVfLqOxmS3SPCSIgzgaw
8OpwliPo8OvF2a4+OhQEm2RYx7r4zvqU7uC7py5kOck9OO11BjNWRZnpRkfRa3Vq
MakRzVerNOHeKECjmvVzr0VTBxjdBCVVvFLSW1CaYDwdq1aM5ay9LWRP5jLfe/uV
VmhyVN5rO6BQ7PDiclaDU3OLf00hSqLqtw5BV3iUlqpQszDMNl4ZTnkduFI0HUar
L/E5Q+maakFY1JFiyxKxWQQQpI+S8o5jnz5zbBDXqxQvz8BVr6xQO27jRvCvLNbN
WQxRbd5RPh3Mke4A6A1tyKeYb7qL8OHi+ORnl7VVExzE0hY4/sN7Libq67X2wtMe
14rwt2uIKLGIJVcJDo5HyKgPSKBwRqZ4o7aBhInVdJKqDf7kcKabpeH+KzDHI+VX
Nt2jKb4yE7Trb3YSfxEWHsyldQrUnj1Sk6s6UM1d/2Y15qEJu2zIpTbQFGIihVKU
bBTQedAWwUUqR1cVwmKCw+5uB0tHnxPbWuh55ge4U4YiNNz/Pev8fWs89DV7iJXC
7AtW5GDDNxaorsCGHI56T8iKh/n1AnmFO7cNdUXsDmMBgnJQLKaTaFe9qVzZOdkH
/DacxbgXpa9t4PRY2LNGOsDSZEotMY0cOSqmDPZ7KVq9d+PRFTPdjMxq1E1coelo
cuJbaOcQ0TinyWB3ePYvomdpqj2lqWD5irUPMhBY0Y+Are0S2YdUicGuG0+UM6Qu
74NCgmie9Rm1HUxe7kWbqOjKqT5IieR8mbCIxi9KlXSt7JD8PYc+LB6/tUVp6igI
gl2bvY0edjhiuhwKUIjt09Z7Yr3NuxIqFZVOt2zGio7P56jOFE//1egMWV+9vJ6F
fGsRwR8lrJjJ5GAGtjZDKZfrAsR8OyKZv6sWiP/dNWLVBcK7zHDxPiJr5nhvLOhf
/S/dxDwwlaXkldxASwNqUD/o2vaP9RyFzLeFbLpDOClpMb753dlW/Rju8vGtuj6N
bvPvci54iBoAy2ru3ZFLH/gK45pWBN+oN4D3Db2B11IlBx5mzIZVTu0tGJjw1ZCH
0mLNOJOdiMESpIsHiifltd0qlPTQrAkU2R1fB3iSVeFSdt6SX3deI7nUBFr2+qHT
mADQjg3IXrG0Dddsj8KCDMk8168c/W5bpHTEX46+Zf/URl/c0/M7FiLk/DIT8MAd
o3jPwLHZAoQYN2BuXGtPRN6MSn8KWZu/vYWXtYkRn4yd+DqF9Y8IzoJqKpMM6Jzd
4nt8BGIXHCIkbwmVXGZv+cezmvjH3hkBQSI3+5s7bSDe1UPNvrdCEjso4LSFTR2P
pf+SUuGE1vP0VZSbrA0AP3jmT56NXrvouo4njN3SBFSjEFYGWxsn1rWZiIX7vACz
6ftVHtMZC0Mefo28M20P2iqXGudBU4JDwhmvUsqlIX4q2hsBWLoUYqalyrkKYgEe
k98te9rVto3TuBv3pNAYg9cAOBXE3PiV1Y35Yf3KEijDYlWvmZ+AgdWWX03PkuIS
eCTSoNRVbLOtiXAUznx5tFEuc96Vgb7f02DV9q8DMmtL9BT9PKS0qu0mGNw/vbOk
0IGujCffZ/dcZYH413jOXaKn7L45hz5BSHCArjRvQC0Ln0HgV7hlFMwIci0jTi21
yrEfi0RmUWa1yC1LwHLo6LK4QPMp1Bskf7Y91HhgTTFXIo7bLRrmV3WmwnLJYBTv
WYNusv0BH2WSAe44VMaYL0hf8U5MRSNI9pqebbI+DqNPQwNXF4EXmoHgxVnEgcL7
1Ho2vhIjBLpRjH9btCVB2iziwTsddqz1D4DAeXqg8vMu0DPgHDtFLYHvdTjrenQt
2eQpHoiwsnweYmEpXHdVBZepqUiSqrcpi80x/DlaSpkVEuyEVPoPBXOL7cRUmbP7
ecxfiiDma37M1Dlv7nrBbEbz3PjAYze9Qw+K7WRJL5IE/R+8IM4b9by583TaBsHe
bVfPPidxqo5FUibfJ5FqY2ynFqJC9Zqmb+V9/Vy1eBcjTtz1tNk8QAA8Ee+FZcCN
EYVM1f9xzQGHCPgIgAvWLvM8AdQRdfwrv/KZ0YAXm6p8l/QHf3tupHW3NTW7Njsf
jf9w8g8tckzcJY57WHvcnZ4N+ZFJkWMK3gmCC/C6tIt1VNmd+HYWxd30wt8OvzIk
LyWtEsp0ETc9Mmv+hrN/g2VWP+JuHnUdWtS8YB0owPX0eQaB1MnUC2DImi9qSyBV
88bPNNIxdVks+FMnrn54mDfmCus6XLyWub5/WUKAtQVYWw4dbVqCrugtL5u1q+wY
8rzPdcCzOAQ9Cj0cuhBioa04y5vf8qGr/wgK2u878+635/Vwd3LwJTciNNwWBjBK
TcPLCDv0tOL67+mvzoO7+EYriBRNGXDUl3M+rBP71fekXV2A6wvj4JrZqQSYeHRr
FIlhh0BgrI7ojtS9uJPjb8LBx0d5Dbskf6DSpTTVN8YJ1hA4bsi6gMT4enhgfGWb
u2zoUTlDNLmFGB/LCQ41FaNTrS70JVb4J3Yjy8QRVnos4b/1J2+g6Y8S21pxp0V2
3suW6ty/7M/CeSeoVzG5YtbKCbqs7JUrjMQE+382KUbz9YkxVf+8LwXJw6XUY2M/
M3qifJPNmdpg/CpcQJskQtOzeB2M8BxOidmHlHyv1ojHtDxfaoM967PZW0OB8nKg
iRBl8V1cfBG17c2HTQpjMQ1m4KDzSK4uxJIAEfcXHq24YDSgah82TrG7ov3k4URV
mhmn7BTnIwF7ssyBkIqP6Nexu/QF65v7MpWIqzFMchx9/Eod4dN20Ht3qScZb3lj
7RkAtjscosWhFn6g2MwMYwaY+U1aa3f9cndCGzSroOlIf12EGXrdNYZkv09vkdtO
BItkRPQIIlEcM/x2Ve0YUchUQsM+7Xu+n/3oNfdwIhiICEpz4VXRU9UWsGnZre+b
cfJLP13BzR+y/pIi75IDW06JfUngJbUiQ1hrZW1ylARuM51LONi3mEds6hScpTKa
av6zpaWV2R8hgedZvYFFiptuW4D7oapDU5SVGWgpL5VdpF9VjAh/v5R1VSFHpy6o
tFK11vSIt1dOIJh3VnwAAOoUIiEsTSI7lMl2WgFuEAtUtm7x9gOF1puLAlC6Lmjq
K1iDHpCWq8GzcPm9Rk0iqc9vaj1HTc2RoJ4jRE7RJRWZ4cIc2vdCU7TubYoZdrTS
RpEH4l/gRlJrdQhNd654Sr5EzLYR5xtmPwvsqLQI0xN4ogRsjtPOaXiKijeHSqhd
wa05W7JZf833WczJdbIL6+BU8IXQJPQ87XuKlURLdE3OEU/WdA/CdRKvUO6jI32t
ZtrnCYY992dvhiydTWSlsuE2x55PRqGo2/yUEJ4wtD8zkcQuBCnPlNCMBKWn2sLs
uY1Y/bMy0L/8vDaTEMPE03/w8Vc/JCvhLK6Rq0ad1KpUCSWH3p+iso5JcAKsKX04
osm/dEmzQq1gZdYpIEqOVX7BKeRZ5hQNJ4R0n7YdC3YJo2kCAK2qYzljlhoopuzm
UPICObXbFM1Rz9uQ7NQAmOlojR1+puBuaM7g2eYM6jRiTo7qghG+6+N5E5y9/fs5
E337jsk7SetAVzczDiweYhM4kAvboAIxaOYmFk9PakpQojl7oLdNEt4qcN45PLlc
k1VliOmvZlWdnKWihWN5U21ib+jt8+pADc+dI6IgiSaGXnd8ZMGtu4YVmtagLPdp
CVn8uwDC2EsAxA/8bcaZ/fu2dAxnZzVIeLUDxZ9EsxHajndWV2Jva2hBQw7YvtbG
XHo9BUKgVwL7G8krfS0OTLl1H8b/brid3o0Kxkh8+saJeuqRJ0/MG7irlC2w914s
a7zrMFEgxYiCDt59v4Wfy/fTZtvH8EbF724CkEPhPRNJcrz7rGRNF0kKfVddrBfn
2E3uCcFzr7pH7nEdS/x5vZKZnxTeovEWMRsqajbNK5WKnPGMaJEMlayj0Cu2KsZ/
1LiURXGy6DL68DTvSW67siNgoZXM6/ee+rQeqfqgfyRGA/EKY0L+k28a7C3OZc9t
az/XVb0vJ6yl5yfOmtbGz1ETte3XKY8VsmWmlv2KrQWXIihE2NRWscLzTWQ+PpI1
4687wZIL5rno0b5pq9UGisG1KqAcBorc+F5JdRyPkE9q00Y2o+kDxNJdea6DKpua
5B/SL5TaseVoQ4OTOKsZmIU/uSp2zzPvju/E99iX5gjY7u4hWGpQ8c4nd6awfk7v
Ka7PZjQ7V4tLbYNd2wSLm7PFVL2ajDlkxZlx3aUl24O0y63Tcikik4zsjB7JoXMw
Yw+rWvk7pdVylDgJxaDUv1r7khrzMQraupRy8p7AW7F1GNhoaroRPB1DB9McRCmk
dnoeyhj+XxvKT1Jzb9hqqHTvtv0rR71tMXBYgAlJT/UZ/WcDwgFLLmI+YuUkcpcN
5uTYaUwR87DrxSw/CEOXAIvZ06Q/kqXDcfqms5i4SorOBtwFwTwo6UbtnBCj2q3i
X2ol2E5SA19E5lTIK3AlvOsfT/33EEKrkmtUgCIbcloZlC7ax/bOd7FevHWCQGxP
1m7TfhKlW9Fl13uIrsEfQRMzXNDSup/h6a8cQc7VtOCFf/UVq+jtHBIOPePEuWjY
qWMLh6T1/6F4Vl7wJokG9KuIh8FbV33R7KTvkywvooBk9QVgYySWolQq+rP3AEvY
L/s4W4jiz99umHdNAx2Upc4yp39j8cLynzO1MKBX01fyUNnb23zb5zuOoM0ymf+/
M85F9nb+kYg6YAxxUwyuBNkq5jxOHy2cDNXrKxkGfy2Qr6c4suyGczZqmlmW/o4p
ttbYyp0p2iBWFh98mEJ61/N1a03zw8ViafEUZ+fLhNdwvpe5ZNNSvjeRew/jYMfd
vORUQWo+o+0E24WKyCszSzedZaz7mRS5GxO7thAaHipORMZVKLzLgyhUKv43NotW
/w31Nm3OcVIpgLJ9IupDCD3OhOzPkW0DIHK5nPv09rv+HQnyn/H4cF+kce3h2Lat
r6kvWL1beX/nQPpznm2SSjo93u7Q7qQOPhVOT5DG6dcudIx+15XQJaOgi4aKKzea
Nvp2zqAQhz7XXpevgN09TMYd8hwe6dp0ZojSizQ/eiuucaqhCe5ULXGcWQWBCQqT
M6wl/T3W4CeL0XJZQ0fgZk50rULQTKIG6AQ23EeLJhVvn0GWV7d5Wma1UH5cQ3ck
kQEJopYaJRjnBuYCcIvJ/YFwE+dweyXjm8W+uEW2AkplcTMv5/IXBdrjMHfm8eBm
AaxbG1DENup5c5pGsGACPVnwRy03KmaHmk6V8mkuIDmxC7OyKBJ/vbFv8q+OiJsp
9oJIh5MQ2EJB+mEamRPZO9wyWCfDHiu+EHa40Ys8R0Auxbe+9PBAdlYlsGWKUtwa
aKuRmA54hZgt5bYxCsspm/UUDRin7LMzvz9sZNgeN8LoVsH2BzNl5YN/CJjvoB6o
fY3xKEVDWr23W2221ROcQ2UNKeISKEDZGda+pkWUrExiZrOYzecq/lv910iSEvsG
CabXQniEhG7OEjknU9pVZffIFVU8B+L/Z5mcW0q1HoOvUHSBYWzBJqpl3u+exd30
IJrcNlTnhZXO5rfsy+u8mhWIhz7DkGmzhxQsLfceB+y3/+mFFrE6b/TDWiTTWJGk
XiYAA6TiZCE4MFKAMR6YtRxRShoAh4QRlhuNj4AHvliT+k9n6v6Twwh2u+tQRR0q
xFoPTA5zwp1vB6ieTnq1y/BQDnllqEMxr0uqcUcFhtBurQnLxGETzmJYMsWMx8bm
KuOT2WupwAMCSY+qmFGL6fxLLj1H/3j1xCN2rE6ShIDfixKvFwcOrLmsTQEqPP49
6SqOytCP9Dh/L35xFDOl+AHZNDfc89VQxomhPTFvJwSBdnVjIMh1/ARbC0K0WaY3
8DPb/PwgmyvoljOyTE2tHuDZkEX0Zc6ztIdaneU4vt7kd4V1kUzMRhowqFZoJ/VE
5FeI4jFQoYPm3IYDurvc8QlAUF0JCr379qUawQzvNGdZNBKRs0zMkPTNzi3dYXRN
/OtXvsSkP5ox6vCLLn1PzriHkK3JKQzCYtt3e/r25FSrFP7/TYusr51U4fHgX8az
OBkqDhGBTa/ZyrWycwVWqgdaLaD9nkLqgYy6kgQhBRtaVsnLBB7VEvrAQwjkoM0Z
tQMdWSzk/9I8IIokDTKyfwceJFXe4xfH8Ek4o/dXPwBKtd251h/7y76+z1yoAsiy
ZZPiHfSePXq90IUM6kAv0Aj9WKs3ZjzRHdINB7ImMXz5CIV2mvM6BAROwV0j6/KH
FRpV5hkGA2FZ8woQ/a4qY5nqhpPqHTTTUKMIuHrGL+QVUok/SutP9h9NMF4ldgB2
ChWShr+V/+UjDu6nec3VMiYy5QFsTilp7imIaB4lrJqR/gXY0QcYj0kCeNOkV5S0
zjCC4vNy+dkuYZuG/KwSJ1JEPph3hmmhQMf6fswT0EFNDd03mnyaiimAGzkea43K
lqmOtQnq5oYx0n4s+GR6jb7+I3RG4fR/NQZ3CPU8hQv5w1QYrxQ2xBFPUnZViu45
fvCkh7ClpMskYE/bTKbkciFIEkt06L2M08wFlpeahnYDfxA1m/9VNXBQINje5L3t
7BUGzr1MCtgao5eGA16W4jhjuKX2qauDd5XbB0bVxqM8PJArC6bxoZXdJxhtQ53T
Ozu8GExja5GX6U/Kk79oWGFZ8eArcXaEcG4k2uy2TscOT64DdqtOw/KqbgK5tGoP
WZsM3RlWQiTz0T2VAFxKloCOKxpus647YnECBOUs0BXLE50NRe6/TEPWRsmXbKpr
v7QJQve6aAtV3UH2Wi+A8xEdjrn9hGvjJpUF5K0DPJni728GzOAsxnWzdUQG8IxS
khKyAiBZZ+T9Pi3wrcT4og6ug/mN5SvDGOni0NpvN30NbUiqo4oTkRP+PPij83a/
TGTJ3268rab7qIVmgl1XRq++SxVJf3BT3y0SgCF+sJHniBqreuYYSy1QDbOwmEb5
819BXb9NxD5lc3kS1+8wI5vq+s0FB983bDfqh5Bza64GsvMGpjvwK6VEkbUvmLWy
Kjk0z1DnQb++CMav5YnohbOB4/19EecgCACONRD5OxSYr9Creq94Y+EagE5nwJ0u
ymLhv4c3VYgJkZl2WAVi2HpwzWU6N+eyIDueLak16XgvJl+SwcU9e0zUX5m5RV78
WhZbcMoQIh7fpbHzGV+2feI9J9VVH80BbwvKu6Evm48/j6tiavQFZvfUwS4wsBpI
oEx57BH6amvW3LwetEuX+cxBzEyk3yXjATMsH8VpV1jFbJQykHOcrhxYgysP63t0
+jLYsLu5FRpkOCywEJuG+YBeXshVlkOlgx73VeZVmuVAcE4DwWKHKMUZs7vXaKDA
Ma83LH4uLGMFB/uFf2b72b2axulnvAk9i0symkXLDKfwcGOV2puDrw+Yh93WJFXL
FkQC7SyWRZ2f6OkSa4j1WUOqruL34wgWVRZZF1nz0rwD4wpUZmA8QbY59LWAk/l1
IIaldCZphzvelM7raDWz1nablH0c2CbMIkytYZba1C+n2sNhxebl0G/FBIMfFVBd
d/bTJxFppffGgatHiP1lGm1m7f2gpq85sobNIM3ffdtP7S5WcqKWCcXPRxXulz2g
1AaKskWJCUTXuHFfKdiRrDJpBpYczmDexK0BFcRKwHI5LwFTdzGmw0AHOvybocNh
F0Ih7KgHkGZWVVy6PDVM0cw5tVHuP92rw1upH1AakQYW46W2aIJEAZKQKGNR3jFV
jjjSqoZBANHnia5IKp3bleu8xm40hQWq9DbV1WQSpUDVMtxmafUgqK/EEUWISyT4
S26gIOM9ZHkMQWY50OYEKyDgEL/WKjzSwseNOWlVxIofeplAh/Wtaokn5sQHzjUs
+AwGGAuBTG5sotHurf7Uz8vGtgiH6D/Vj0j19Bve3CJ/aKV4kxTllzNVPkh5Prfg
oJozqRhjfKVGNtSfWPOhI4GAtZ1T48EBX2pRvEu+hrai0g5tHRfQsKvpPnSmQSCr
pebiKeTqINK6NTRd7zzC3MTwf0o6XH5sJTG7kw2ur4nldDnvbGUgjbu0Wo1OmN8g
vXgGczYyI//hQ6+PHOlC7XGG98COYNBxiMYkFv+rD9YMpcb0Qi2M3gRCR/UZ96eB
uKh1moX2n1pL0A8H7RoA9PUfhoeGJu4BSp25UgY6pSvLkwYsPSQWFZE4HerY4/RI
8iVccrIa/q5SInLpHJUKBlsvDaHVE8GHrsDUHByRGt/oZfIyVVoMziSjsoV1DNsv
m3vg9MhfaTc1UaF7zXZ6A69BFrxMgf8vhMOqvUKlqO8zpa6ljd6JZma3g8JoJmWy
H3uFvXH7z4MwcTLZ8y6A+cKlndZuD5Dy9+J0X1O9jt3P0QyKuSxFf8+T69tl92CI
68sRSJyjY0Rv9MLvO1LlAcxhQcKQiWDg7tjc3saWftPUuphfKai9mmMbeS5G7wfX
AyFEBjV1V+/OCiIOAPJ8fUA5z+wubzhB7pbvx7PrnyAR+Qns4MaYRS2RBLrLEZvI
FhesavxFVkKKBeG+S80ohYmngLkvc4eIxYILBYo4SGrNY2J9hk+b6GHooWi5lP1N
KXM8GF2QvfRvhyi/Q2vZUqVrwSQh8Yi4bd/m8pwHDPD9LP5k7cRPLBgdBKBDXmeN
C+9EnpfTvRGaz7LwrL0TzPaf9bOLTB1iLQp3HwJ7nfHA7w0mwA5K9W6C88QNqBPp
9nnqn1ncyJjmruwIBasXqAGVRAREScQyPvN2UWJah/8VnSlHeByN/3c1tMGQz4tY
LwiElLNyrPP41Ln56sI8Y2iLmr0Ag1yYnodZNLpy3FcpSHRkJMRo5UJHOicLCMzd
9LENg3J3iRAG3lRXmd+V2cdTOUfOt9rb8yEZwkEvHm+S0+Rv7si4lazwU0oHpI2B
1BNyXF6OESSaVJjn/2Vu1wW95a5AurRx2bD7o++7abmAgNXO4KALG+ArZTCf6S61
yBsKmeLsajyDgXCGijAUs+m3jFC9bRNBwjnDyyH4gueCAc2Id79CBGEmyuMtYYUt
yk8hx7p4Q0FG/Mec9KugC2aTid+Bk5y/QHcDXc3vhQmV2NcMI6P5R9UySH5MHCw2
NndfvNGsCQmyb89iDhwY1iQnOoZBNJGfa4DldRaykktrzD/CeWVYilh/qDQgAGNC
qeko3CmeoijYYPs9hSCLQBmzSd1+YcbL4xHCEd7kG/ApxnLSztALPJUb/QhUalH9
g2IHnmw4NNcd7dH/KMH/wNTMOekBznxpboNf5MYqg+xaQn7HveIxKFNLq5Ha1cyx
1xLFV/3+4VFce2QQRaLroQ4LUwitSsC0N87FWPQvua118rceiLNjmNwFIX+qgxAi
eUgemOv6mPHWcufT9JhBUYBrSkRao38quWmBiDpF4zLTLbjOyAgt8yChSGHyg+1B
yRA8RcsipV7ZFR6YAt6bcU76kxn4FdwUX46EcKFf7yAQI4Ew78MeLwTZ/lJHrP6R
0eulZG9DaHm8Y+9PtAjUCz3bLtmDMXOj0O2pgS3Eq2SCMUpIm8ZBs+U2EQjF/5u+
haken5RMblp/RGrjEKwa829C6enzdIeOOvqi0SmVdGrsNyj/2c964xxJFFR8Ru8a
Y6PzTzLmdGNhapuTOFWvPu/QibQnHHqTM7/GSlmUUlL682v/p9wuCXGOujaChCwq
f306IpQ1T3YxHx2Cpx5wd/Y6kiSU384pmnU178vPaeLzfz4R6B/o/qCKFetu9WTI
Gnl99SgqIVp6ISjZpszxyIp5++uLSXF7gFIm2Z8mH7zVfdU4LrI5JUdtBtmIvJLT
j+BvZJMLyF0gWN/BqswTK05AkLegPtUKKWTT8oN3nTaANbiSOjmlKYboExwQwhr2
cFeVxNAWzaB4pjWq7En8aADHUhr6FhfjQpr1f8pKTh/wWO5MtB2xznA0o5KVVduI
8xmtLGpMdQ5sdMehtbcjwYkbHjN2G2nij9o2CpotXu/uX+vdlQb6/jmX98X2jViJ
aHxIO6FHPrFODp5Jjv4gMHlaau9ttT6q6U+CGmeNSY4WJqv2xA0kceqg08eVVeXU
/TDeWKeTVi55Uu+/8fDYac2jig4r+TQdpguLPJ1gTT+wTx9gM719gsEveZE2cTmT
Nxg9VtdrSTkK6Mw4GUHUCgPGQYTYSsk2ZBIe1riW5dBNlic/Kh5dsr6Q/Mh3MD1h
tXV2yLVx9MDDdJW4w/DlwSf717Ip+ipyxM/XbJwdakyKAKtJuM/xhNpau4trBx5l
Yh/+ONiOqKShb2y0S+m78m7wGJICy+HTy55iCT+g796bO4GRSqbPicFQ5NgrpdzO
q8M6zRYTZrQssbousaV3aOfkQ/YdxC5781KDkGF80vToZJkL4qWrEEdwjX1bojOW
JTbmdZCViaqCg6uINawyjlzXh7xfKF5mnWDLJFg6dT4Aiw3U75QHjZCvADlz4nZ5
8dnLDIvFhV/QfxdpPnbIvVkHAKgRUCTWI+KG0kqeEUCFzvuIgMpMn/cCDDphgF+u
YToiodrSSjGYYi8rvt5TdBheu4Gw6NXjg3gJqEFUJ1FKPu+S7MGjblnighqTaKLU
eAUsS387TIS0LqghTpoD+lAgu2hY2ubROxgTrB8rxR+U6iHSrTia/ZJH8xsRi68X
HJ5vFPF5Ar+J/8Fc1QOR3wPuVknONM01BLxWbHyEO1d5JjiAhzva3rl2JCvILmRe
VrgnVr9DBG+kCgt/lbTSptA5TclXW72B01HWdY2xTGb+D9PZanlmgKrjeT8zG/G3
jVklgD2Qjh9KgG00FIcgI9NKd6Y0x1b3wFQ6wOy6N7czmx+jcdq6izY1xCgJNQTC
jO9YrBdojOF0AaOpZ120axqBRLPjirVtvmx4QRfRs9rIUehcRv3T2IDbpEtv4ag7
Pse/UdbCcse4jNimXxSqzl5FXwd4tzjQdw2UUkj8ffRUS02gc9AE4AQVTX4YnjEp
f/FhMJwc6VcAEInoCvAUkQTQO11ww4dyRCoNLMeJQJQl91opzUYFNpsz52u82T+P
e3kIzjoop+urru52Uk3S+heTS5EjWYpuN6i/R/w7BKstv6srArMEI/yGZhxSAl3g
8U1TmZoSXgTHeNnUceHswEV2kMa7WdyGRNkbGZr3lPHbBJ71Y0IVa/fyk1d1yUMq
Be5KNlbbNHQrbrz+7VEtBBTGkdF/ztmXO8ys8i2v6sP6PAtgF6V4+Ll29MT2aPuE
jDfA1mISeN9RXYDC4Oall0SmcfaLiPE90sq7cBLyuHlhUMsxCsk+xwsqhgx0Q3na
4yk4hLirGX5E+eSgxz48zRj+Cje9zlUgMnbKjyoEDHMbIILFMHHUunP/7Iuq4gSi
heBqrKwgWHWKM+6fZoi/EwLEAN8HZg6358ZCf4fvnC5EqYCzdKEPOaRNf05pZbSm
X5vmMHnQRTnQXaou5ZgN+kp3uYT0qePDmx6hj7CqVjYoyiTFKv85kRNA65Dquxrj
trvb3LO9ajf4mkPT5e/BShawm3tSYOuhupAhabxBOpHfqx3kCY7Z/ekoXzWaviTa
JfJbGUFnBs/LB/kbAtTcpw5kIf8NNeTaWWGuPYto9wChT/FDP88kYRyepqkXJmMe
muQNIU8ptFDerejkw91Mu0c01cjsmTljOwx38hkcEkBbfVXbX9ty4rU4DC3dmilY
zU17SLAeVxFeeq1OF75ZP/+/0RZdMd62h/PxEU2bceCearzbF6CtIj/ymiVs3CNj
rZuMlEVGLJvfdGfi7bMojSSTkwZjiTh7Qc+dMlbpybMAhsGqXY7Zh1yglI0NmqBH
hvruXlCRpn6MV9ClgodFRONv07XNplYPjKUNbUeYKBsawARVJZ8YwzL+ZWrvuqRQ
iekyaQ2AoCgmM3zRakYpnFJgGEplSGMTwy/9s1run6SxDry0dCqrEKT4dNleZNra
zM7AeLpnu5d+BQJUl3ORskhkPu5BU5poQ8NhLZnJ+PTSisYfw3diW8VYceTA8rqS
+3FlOYQHHn1qGIAD6Qn8v6NKdyBD64fbka97bZ4D+v8VH2yIQYrpOk1WWFnFuJRc
DGKnJ3P8hBvmsOw4CHaekoByoiB6RwgU5HZFYISRCmB9MB3hg6nu0WSwbm2NqikO
zQMrXKKPPlML7+jLZlH9m7JLWG3YwcL8vUaIUuWjFl/8R0Ij+6KQqDuWzhqc0MnF
TEg+6OFnkIJPe1U3D+IVKGhXG3rLL5qGWBCY4S+OY16iDdp8CF7cYuZrn62aHkUw
kA1NQsl4Pwtvswvebl4JsDmnw+0bRcbVQAjY1rQfTeCXyPyrKj8AEOs7ew0tTQys
bVN8hVyiNP88SNoyfpvOTmvJr3cUj0+QXzC6JsHD8/aDfr8gyyidZ9QQGVtRJS5h
ysbI9O60JfncN8iVX0xXKgWLbnqI68cqOTh9EvDmS+PQkAx6DEz2o8n4rpecJy8B
zMCeO0YTaUxxEFDRDK1z2xs+N53iiiy/6HsO4iDP75HhpnmNem8qq4rySK+BLRKX
6qm8bFktD9CmOEQWGGWgUfG0mPcQ+iTwDe5xOvCjnXANKgYA8PoH4Zn4RO8iZ/Sn
UxlSoUssSjCLRjiviHCtnC2q52bofH5QTgB3H9fBNXkhniTmQe8cNDdpTJcoWQOo
zfMlFMO7K6DWo8Gqwhyk5rRgrGpte13KeJenqn8Og26AREqQhiEPYrHX2XYpEPTz
fgbyaOMr2hqVFvDfXzGe1cats5SMqwEHzYuhQfvMGnUj4epxtIwINGVPlbbVZwA4
mkmrDviQQkgz+ze+JIPTKIj7J2zw9uJ6J7rvC9q5w6ALNEqKteVcwtfw5+Gql+7T
7m3vVO3fnx5Z5Yw6WW4SbPfL8zDB04r/+DSF5Pbx3EfydteJN2ooB7spFM+14Hcx
SHrPu8wwDmG7y4kpuWwFBvDtUnP0UIso+XxIRXdtFAk/elLEZTLOg0TpfmIbHC3I
J76hJhIbBLT8bDtlUInrtr7jG786cRC6WEApY/Ed1mXZqHwqg3AOA8At2gGkq9qr
vFZNy/H6k3MqguwXk4BidPrbDndWmeF55M6w63uYKeo+ykGG2NCxec4xsPeivEid
uWfFphwOhg9CvRzEtbMAur3n3hMCpnVsb1/G2X1s1J9/93w3KrrINoqkbV5vEBnq
K4XV+P0qQ23iNeN69BHqMFxDbbUEV2jhiavkB72m50RnuUdOB09Pb362icMJJ2+r
BsOrQj/ECr0lZoRhuGS1qpoj6l1V6akhFGl4NEMLp9Bw7Rld2AD8y18XwykRFJ0y
QUL1E3j4AWnXJXNoreuSdUhNsrbEhz5tdCHk13fpsCUT1K13Uy2i+eyr6mNpINng
4MKV5qOJyXHkDMKlJTw9spx/eIp8rRzTRcoRFtusa0Uwk3V9iCoZA9tToV0bvA/r
fL+m3yI0MIYx+Zw3mZwj846brGZbrrfB/Gk/5V0ag4yKWS1h9WRtzMHgIWunwAVd
DdtiN+brMLrvkM/80bjmQaQoiEDOwPVnpoZHkRlNQhxWo9Nl1ynZCwUx4wa95Usz
V6884Gst8TzJro8mdjvk8z83oLN3Uk84QMPOHHWRYfPEFBfKU14vZewvtMD5YUE+
JdgHP6uij0tw3J01+eOTlj5lNwseSuznXEZ1B4ly9Js/tnk0aneFGHQG8F5+uBdo
IFH4Tqod8zE0cmAeKpojM516ifnwd60AYaooJzgRPCF3AyrWkM0a8C4+IhyhTpIW
EN2Lha33a0ZR5vCKixstZrMe3nqJe2BL6U6zWFTwmKvWpLKwPEFWlqzbi+/tGyX6
juY30VWXJ/xgEBe7vumwDXSJvAv5KNaI5TvRoNbE+KzOuP1FvpU+OR3OZ1HAfQwL
PKRimgEskhKU/g3f3bRoxSll+wfomHwbIoBYkjs8gp87z/LukU/tLN5+/7quPmzG
p61cecFa/nDT2nkP82DcDVbOhqNfkz3DU+nw7Lx/VNOkgYE3wCEm9MwCbx7FhLxG
sgwNNNC7lO6NQECHSg0NwDAi8DUVZEjNWpRmPWNJ7XFHwRyEMPRer4qXnBQyA8Aw
OikIZlpnTX++o0ZWF6m5BgmZkasbHlKuzvdEwjkCuoRYuJUZJcsKlqISAnLy8TWX
T7cWIbAWJ9zDszeNIGMHsz/Ptdk7+WZ6A+aBNcAJG0mEQjAL8KhTd7JaTUoIWJ6P
8IxeTWT4ZydhKEovT5q0k5BC0FLlmQ2po+5ieeDyjczJOBM92HER4P+dF8M3n2JA
lmhqGCUSYpRAcBRW6SS565NuRepQiW9sL5yAkz6i48E5W8cSqW+zPQUksL6kB9sK
6Tl8uEpVmjJhcMwqpc6SMGfpom/X0oNu6mGY5DeNUaBZh19oZ7LD6w2i1nXM9ann
1EW6zyhEsyDDZpk9BzbUO5l11Lh/F3rQGO/IhfN11kil3E/IswFjAgBBGSVCQrv/
yolgCdM0hfakQ7/2ev04WhG4byC522BjappyTPbzDuDcFuaHKhe2wTT/UKbzftLo
jVXGqYTGer1nfG8IpQJR2A/v0hQNKiNbqunDu/MFpa5YWHWraCoHSByI7amfDSPM
tiQnJoIe27l8pX0hV7NT2PIy0WILRKbl7rSjANnzlo5GikwkICmV1dgsi7KR8NcA
S5irgQZZQmf0qIyt3nZTGMMNWyTlmrzwiQOBjQvc9iLlLicUWLCw35KCEUc5qhil
DNarmMy2koUlgR5s+DCVh93D7N/bHUZUhJWSwaoWJ1YpdBYv21RIqVmrw+hB7rsm
RQnP//jolt5lH7/1seQfdR/nN/SS5iPLoFQWiXkVxTE+xNzxFz9BXQWP50OBpQZi
VirRj/QUdTbq08LccKmYQwB2FqKsAawzCVi4RL3osnMbkzqM9GbVPqnrJAAq3kx+
+2PhjEtE5H5DLDuNj9gGI3V8d7X8XiIFF0AwxD1BtnN0slC/vwabhEEqCTieb5RA
8GzJpYCCyIRwCKUfytGeiRndVNFSND0toZrpNEcT0HQ5QlmdzCetnKAYOfDcTL4x
AF7GS8jjDWotm5j5nmtBhgqQAo0I+aDnWyXYJbriswFFBUsPFotq4f8XlYu0eQcu
jAs8KIAwf+Uc3v0n9QUoVGtXLNkFGrMdH9OeJTk6Xt2tIy42slSq5rSYPzGIaL8e
7X1b8Qh2/qxuWq/HUQlsM8cHJUcfor22lmyKXKmF7TXWTmoUFIzPl+XDvJeK4MuJ
Ntqh3wMcfqWmRdFr+a5U0MmnTFu6dYKXw3oAuguxCTwF2qk9P4gPs4P8Iz0LtSMh
Hxk2bNEkNhhflV2XACgJAynZL3VNY7aisHVYOspUVeB+2R5Y/b2uvbwy6rs1urxN
ePb30JzAWOpQ6v/xeFNau6KD8NoCTgrmpAefZmkl5yiMi9Zx2TtWTxqvxnP06IZs
QkkU8bLd2q5HLQGsNRjFVeVStzccOFLHmrUUgg7MiqNZc/U/8zhm7yL8b+2IAGKC
avlpF5u+b8yg5PFRVcgMT/6ii6CO6YmMYmN1P19oBmpEp98BHpXS/Cr5iiyyAZUk
0ztwYdSNW05UGLSGh/upmgS+vCbIDuIim4hnsmog+GcJBgsvtiswt3U9wH1PnWO1
h3GNXr8S5+1ctc/ENURm59JeRW6JoJxYwbyZgE6VCm0/jdO4cx3r3h5lFfDn3X0Y
vyw8I5DyACqs6+h/y0UaAgLdqm+uwYb0reJ3vYT1w1UM+aaKLIvWGO4h4ZxuRE6O
3ntaMovuXmt92jVTEypKMWDInmmXIUlmrMLXqQbCSHbTcvcBjYK605sKMN9OgqnA
kpZEdNdEpK95geMqZlP9ro6tFFPjkRJ2wXEt1PsWeIjoRUzunxS4aFSwglTrROk4
8dH5wQrLwK8i/6KJVcGjbUU/mbzPboyNjceC6xX6GI3qiiEX/SIBGixS2SDP317I
80nyLHle9nvtWDIu/cqrP4BHfdtAACmfBsScBGr3C4NsqV3VtXBC5smFLAC43/Ym
U1H5Ogg3XeVi/L7wmfvfw7B3XEgQsZy67AYJuyA5kSmz7WZPdPbkNhFECJGOkLCj
JnsrwCqLxRVX+9iChtVopShIiV+/6qvydRDy4+56bgJUGIUcC5wwR8et+cKZzRes
hHlMwvlBHMzf2D1S+OZM06CkZzVT2v1HtTQJfY5mrqY2DuHGpiHYZdOZZ00zTKgq
L3cIfYwsQt0xAzCSePQIzaa7biGY1nWEhhQeIiM+muKbRo+3oitTMBPJKgldJ5Df
EKhegyMQh3fRhNJg31BwVINZ0ChsX3b9IBBJIeqqxyAs4C1y6dWa3Xyv9k6dPfF2
i8vED3pS2rvv7CQgbfAt00yBGLx14SxkgpbYC109CweAKCSm6B+OP39uBQ4Tx20S
ySru6utfkYE1/qlUHfx7fVlj9k697mBQuuk0uqspCBG4l1gJr2jERTzu6TCr28UH
N61k/zAfcz4jzL82Bwww6XZslwP5LTcZz7DWuPXsHhiWjzwMtv1Yy/IMkWfGwOh5
5Y2viV7IyUc+9gaK/g+lGvCrX9H2Yu/tb0xcg0OgYgGlOk6E/Ka2bShripUUFEE9
v0xbeXHT+49aO4xemxrQ9xiPr688wzbhPBkYWZywgEhC2GAl64vpZgDHIx6o2Ok4
53nfF0CiKq3yqoaAxdiJcuq4dYdh1eZnrky5ib2ppvaPOKBvqqxjUcggZlz1eNuj
BBo6/rqQ2ZahMu52udM6AyfsQwcytHdpoRilmRWVmO5wMWI4nIUadek8Yk+OiQw/
ndery+3sunZZAHzaI6ZvhOqtC5icUmeyoP46D+RTzfdNNQR5M5IiKdw6Cj1JM3tf
u258oYq8lMBJttT5b/vsCOC/V3xsPii8JSsKW3C1e6BYWYyDWQ1TT/rPq2D0YhEJ
HXXxOLCcce5G3jHQG/m2WJIxFVguK9Vu+O5Xw+m07AvdPHuemoDs1/OyGk+e0mVd
xZ7m76YVNin78hGb6G6ltYcyUGKq0YcQdKmvE1qNsq0LcR5LkePioh5MMq8A5EMI
q/IlvbCc0IpyUdGs3hZ8DoKdBw6et5rr0v+xWdAl2W0wf2fF7o82KCaAcsotYkdy
s2sbpnhN1PjJxfozqRhv31hgXaeU56aJD/oUItTYXe++apRMNtrlpSYBIcWbh+Va
t2kVamyRcs5iklX/zsCpCevleU4jjuDldN3HwLZTwDtXFU+PlGHRkQrcgcsCspfR
bSjndmovqiaIb6pJSE8gStDp2OowEOgQIndaF0zdDXN7N5sbbeTAfnB9PQtowpfF
N8zL1dz+ardlZb+PaZGEkgmBU5uif2tVjojzSz+BH8v5V8g5aDA61zOSr9NmyJkz
tv47SkNjHKPYlSsbDQ3W/OIokj+VnINY4+qXJBOxBdzEKTU3ZvgXgKQA96r0QWkl
XgzWkmUmsHc60tU7jsf2ReHczXFMBE+RGPQnNyUAgByK/eezLlb62vNcY7iQbhRN
M1luvceU2rvHEH9p8a9+1GHmMQf64SsRgd39BFTwPtrakKhciLKUimZ7kr9DnQZk
Gd19P/vKH8HnxsEPoXY/sh6HbvMne9jIMnCMdbfWNlutb+/tm6EaY1Zb+iqs2ahb
pmcnnojtAduolQF0DhfQaijjMA7Qa6LrQOykOyY5cFLgW1WGkzK7dAFS71VRUa1n
ZKqV+W4hbgLVtLJ1MoEha7vqGXCNyRwHM9hJD8mWwSnKni8+7ilg2gamsZA7XKwY
eWraEzDtFEZTGVPmu2aw7MkoN1eUd7dqMT9C2lRhT+uWkdT3U73Bhatrc6sA71Wu
3Hl2wvgJGnHfTkaGNeu2H6A9nzLv3uZiZHKIZmcMrj+I3bjFiiMrgxlJr9SJGl7m
GTc+p7S90VqT27YEaGEdl8B1CAJ4KKN+JWak2q/sjObxVhgWvApUSd1yD2bQkunS
peam0PhDv9Tzih9UylQs79PhyJVGwdJXJI7Cv2UE079DqpLuayx6dhUrqB+lISa2
PEtfJzqYBGzy/VO9cqXzxoU3RZyARJaF/XyCpHgudBRR6U8X/+eHvw4unZQJVMK2
UteOiiGzvrsa68QoakIRN2MyWp/QBvcfWFYw5aR+BjIRHzp63ueqczor5nLvh0yI
R2mfJ9XW5kkdwVSR8C3DfPnTukUzd6Ll0vXNG2s95tQKsQKMWNq413dU0bLbbvpE
X99e8KkH2K9rLUyL2H5SD4DERZWOX6XmfpcjjQq4+ZIZIYNO5895DJm1lFJKGY3v
b/nLfCkbLriDMMRbK19juMx9w+CVvgsX4TJwbUZplxk3Iox18sEdO0/1jSS3odfC
8iPuVk2PEBrJoJm/z/VgHfNLdkj/mc2MmGJZQPeodnFmtY1UBvXEfaDG0CJ3ef6P
N8Hf4FqbLTMbRciFTGU417CBMYW55u5CoEdX9zepOKcD7ybmnyqZAntZm5ix9+P7
8cG8dOdHZsRLk7ya1dQ1ihK4CMlyi31iltm0r/hyXKXL36muNtngYNtp1D9XGqPo
nMVmLFpY7wPhsxQHkS0Bb+hq4Oo5sHGDudGnkVPdtfMFhqytBXJXAGM0Lv5IqpT+
k0NOSA6OzlQ6cb0WFdTOQHd2z4NkHOxtzTvfbBqAQdoP4+r/8ogx0NkculiO498W
ErDASLzWUQYjFEyMNp5BdzvC26WGuYlLENsU+EJ8otA3F53DEQqp3/zmbGxbic/+
CFd7MUb5caGk2//VQ1epQgAYf5FY8U63veohYM1bGxDPRXGZAgdqU9zu2C6Wce2n
WGHkJcZ8Xl8Gc+yCkuZ4/2/7okS8Tl6Gr6+h19zP5r955wywbB/J6tUIG4rP55Y8
S4awqgionalP1sREQui7hxXhw43/zhjYPxAUo/W3fVmpUXfvhie/C0nTSWargALW
ni4ZGF6I7MLCNGVKmy4RdcsGgRMA//FRyZMt5O/AC6GqlMsEPTP41jqZ1AmhJ2gI
UglsC1moT6lWwkgOVGLVUOayloBnk7OeQ2kZpjipD9HDzlgK6irS7Rcvk6G3Sj7N
bwJd1s6nJnmtdj3yyAz1TDY9wW7S5aV2woq+ETqh1XHx0/WV+izv03f64+7ENALS
8PswPXNjW5Ov6oKcnpJkK0NAWylaPgN13ldb1syaxjhs6eT+3OFg1nw8xk7oT2A4
nZNkRhbdUpsMsyFbjUpDkDFZWxiMh0zzsaKXWcP9KrfVTphgIZuthR1fl86tXHFB
KKaoZP+klj5Y9fmNViLVAM0CRIOBBQ2YVUTG+/e5CatXNtqisNT+wQk1Nwpf9l4P
14vTIW++RX2Kf7rn69LXvVkayubRTmJN8Z0LCtzcT0D7x+HiZK/6/NDQPP5QjBsK
Q9oLFKSPgwCsEjmbHWLaQyXwQw2d9REUH97FXY/toUWAn3xxmAQBS3H/F8Oq3B+A
DzWSm26XAHWe4kKn8L2s4CKczF+2gf817bYVtDYuB2p1PxjnWABVpT9iEC5Tqiqr
mkkBRVT1MjOFAEYaOH/q9QSG7Z7JR0m7737E3PFyNK7CBhxr6RZ81RDMVwXA8q34
Q0ydiOgg6730/kQhNMaXj+W6HtRuKuEbGmGV/wJw3iByZ0VFOVQVM0+jExGO3d8U
7fl1VvXOcunN9gdKIqSe0t9mY4tf4VN2DBBraeKTkwjtKAzViIR+TOgLTYxcn/Gn
5YcsRSlrEzwg0hg6pfaP2cXPNTycOYZlNvtl8ErWF9QncBY2O3zITMiyyLBax+Pk
x0aRGzGjEet/jN6fpR+lGTguEjHzDdB/lNsFM2jqXJBE+I0tn8gyhY/IzVrcDJnP
nKCvO4P/mBY2M7Wmv/icpAemW3OOBAyzmWGvfc6xvpgeyyHmC8CNVBT0/MbBBA3G
ODG9G+z8i08thga4i+jNZtIegQi9LRcrbakw2T92/EiOwh1NXQYjvU7wBaMzxXdI
Nf4uvbyJe0pWe3Bnbp67g0AvSjPaIxqfmdxy7BrB+itDSw6nwMQBjzr7YMAYjXLq
A4Wgzp5qM8s1SR2O+28Oe8ebXbjKtCqnYqYQ64LtyRnm0rmQhT0QXgFHHer0hhhQ
w0GgzxRU8AtbJ63DKb3OIptHJxonFPmzAKuDvrbxabzjm7gTeJ0fWw3figPXDwlZ
ZJFUDbk/5BZJaIfabvoL6PdXi8GdGunFI1eWRj0tPUCilNfFmbzD4upCA1jwwEHf
phr+hdhvifTS2/L1N6yVSlClDRE5qQjTA9ggYAftUHb9eUoQXR330IbI8J/KjOfG
/PR0GTJcdGJbXQpZM4vr8/dN6OWeagTTUZkhtrn1s+/Hbn9faySG+aOHjixyV5au
DcUMrjMPGDqBzD0EAcvdfCL5HqfXDoIBuGzO+gN7UbNh7z9onaK64LY5fXejqVWr
UdS2/X2Blkqe9DqXuvw5uML7Ys4OMPvfZ4LP1Y+/GwgwgAU9nb195kCZlbZYoGeu
kFARzmmd0mhFK/zhodeFkMytCTS8Ms7mZEt8ucevASkX2JRhI2Gn1giRaQi5IoHn
P//oTlNU1ikwNasIb3It6egVy98auSRvPo5wU2U4mlY6r2XPBInlbIx31gUanWxQ
KYP2namtJ0GnFw6xRs2YuKkhHCywBFI8V6v9ENOTdCIx+1Lv3lpuDKW2oscC9XV5
hb6yLJFEIV94RxYByoxu8A==
`protect END_PROTECTED
