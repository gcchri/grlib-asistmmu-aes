`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9jlSRNUnsMSvKm7tFK83isMiX/Sa/qDtIJSJn/7VBBA9LoDZOnnzqR/E/QwoCUh
5p0+fdzjFlOtxF0o3tn6lFlB/wvwOOaaG2r60HyMyOvhoOeLVHSfxRbNJJJXLnX5
PHGExuBG5wLqOPF+C0AvJVJPz5iLDPQjo5dGQnBr/7oba5oemsxlUNNEb7Lz2zxh
6x0dv0UcA56R5eASJ33G3BcjL1wEYMIKXL3fwK+2Xaaaa0itG4Wvagx+2SnbnX3i
hwSSex0rY6YMVEg/0bov6YNm9aMomoKwN0CjFanupxNxvQTamHkdWooV7K/B6Aak
m4DCP4R4JzZwZacS2CkGdw2gkO9y5lIlUEdQ2U+KjdfUAvdTjnuvCw2hc7ntq17n
Da+cYr4oK/Z+k8IZEhoTtnHAWZONPKMYjC6Ox5kUcVKPiv8GLg0CsuJQf/Ol+W+U
Od4bwQtGkinEJp9ZKWGcRMkqGLcjliq/5XwkgHEErm+2JhhP7CgoOfnJ80SO3QKi
UT12Trd+YAKHmkvd9a+PSN3FspAZFXorjkqss7pEu1YS+YBuX6MLnbT4ny7Ojfzs
M8GEpOglmARenQZvVqTTm7iGEci2spdQtYdAzBoWdRetKjmJPnHpT+suJzCAiKgQ
WVNPP7vPx3yVS8G6r8lbtyliKXODVIp2kj/jTRCsygDkWiNZUJ6xfxI+IMMSoiyM
69dbeeHmDFSo3sZzngP8gck/4mh9+aeO+S9UcdVtvQqCBLX+6E2RY+wogoe1EkjA
itQlT75OZPZFPArTis3yWyCjJzBIsxT/5zwEjoTMXJd0CS7A/BKKSAgRboDWvDi4
7qRaSYfHOMa7emxr1A5Iw0yjR62TnM2K23/VQqjOLU1pN2Vl7SYp1gtZVgNUVK+C
oN1Z/kr8LANBWx9ncDWju7IxVd78J2/JoQ1CHLkXBhi8tbcTO230g5qfRI0wPzp4
ZC5aaWW0aQZVIRaMTbPocax2N8W8YryF0stxgcEiKZPJKbSIc8PCQNi8ol4+PsOh
33xuYbcYHzxAtTHeA5RCMGRJtFuNrA6dKP8JvGufODCvX2JgNMwVknfc9aIlxa/d
93QyMmrWymUkbIuFbR1JpI3J+XN5gRVOZBWDMwUqaOZOqbGNuJjjuztqiV/Yzqpc
eUQRC30+GrARDrAlrXLZbVZ8Bh2y7+KHD7vVJyJSpV1oFpVaBPWl4vpUI8u2sfdD
qLS91wpfzIOIKWBbWTAKuqn64T2695d2GZwLh6hSx1JWHTMf2rycNdulk3mm5qpR
BKEArBjn54yA/V8xz9JOj27b/8ipDI67y2Z//Mc0NoaqKFH7MKS1w4YhKZTJ6Vvq
xnAZ1ZgLRjbZp1egHMovh86T90QvLEdHXquPrC4YJWOp1wFXGVfddiewio3Ir0YG
NErVFavGsNGBPlA+w0MkDNAfZ+ulzGsPIXigYedFFC3uVnCaLZquH3cnwjyO/Cys
nq8N1TpQ4rIhIstiBtmH6OVpZpRPWWB27Gma+tAROIhkTzDzGi/xdHfAOyuXZhJh
YUdy8UWK2hZO6iPfizAUP1Kebnf0V9UkrES7kItogtoqpqcVBq60buHWUQpmVJdp
lwSIExKwfeei6LjnnxFCemVVmNzpPD/0eGCUq+hmJquzjE7POPQc7d7ucjjF5WvO
RVm/pn/sQj6izg0a06C59B36ER7aU4OSM7tOfMQ5sFY=
`protect END_PROTECTED
