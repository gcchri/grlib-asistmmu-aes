`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1JXsk64bCDC/yrpccQGCKL/+BgjDsrEec3RPM5RPAQWYqZGLN169DQPvwfXEkUG1
+skpc1fdS0eihRHtuj1d7YB+Mod8rvct7t9fQDCwf4V3ZnU/USIVDDlnkrGesgYQ
vbSE37o0wt0tubI3sHsRLyo6YPR/BFd43PRns4jG0c3YlUi6d7dnTPJjg7Ut7PKM
rnFLzHtMOWj5ba4SlZLNdBy73LwWlC63DgWD+lTvmd3n0GChzAFm/wTU6j56Vo5X
jVLEFPjG+0+6cdNkomuwMpmEq90HH04aEoQ+wU+r5rzLUbcr7dT5b1pkCd0AT0HY
9MOwOZAUojALi3wxdklr31K/ImjaI9+VN8JBMKXNmh873vrTopiTmc3WHUA0W9PW
tyC/D9dPC5lHmZ4DJGPoHkurwj+CojAXcOh+RPFUDHMKDHP62/9pFsIMGzN6VwiB
IE9LhwjpbMNwZeS+QZ9TWHYY5wmLvZ5DqOC9sLeg2Uk=
`protect END_PROTECTED
