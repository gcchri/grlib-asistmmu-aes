`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GtBITHJsVePdQ1HTOPBzl7eKsgfTDQ2hTxBcMicZHyiex3jv9Bl2MmWmjsOywVTL
7LKXqNCp3WrxAPaNIn3gjTIROT1UIGG5Yh5tyEefj8JexFk0s6oXYX7uPyryEbwY
gw15EcDKHUigg5G9M5bSHWxZyXrAbah8aKDZUm8rCReQzIR8FGBZIjv5L3L+y29g
VtfqVc5kWMnlv6iYdEsaYLij1ZAZqvYSYFEDEn7MEuA1YJOHTSBHDxdBP2szlZHn
AsRkwlhpo6HXMQ5bUo5yQjLbc10nh+4ubBgkIH2B0TJUeEzz48IwofjMWNJOJBOL
lUzCICJa/ssHJbrcUNWsWFaVre2/nAF2z0K6o+CCzctOppMlZVVd6eBHl4ozbeZy
4nWXcJRrYYWpMq5Ml3uRFmmqy64YDRXMyBHkV83YMtUQ0IWaZiscY1Vi7Fd8O1sX
Vl22xCqn+Oe7F+rvhTzeZNq7q+rI94Xy9Pbl8YCx7sxNdsQMTKDyoaOYBQ2MMD8R
GvtGLYwDbOTEl/QU06mTWgHUKRlOphDmyTx/z8RzVdYI620D4Asq4LV0If1W8Hhv
VtYI34N6i19dTtuizEKxfw==
`protect END_PROTECTED
