`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fU0A/5Djk77Ai40bwJNEQWgNWFLE6T8C5OsxM3R8YC2Bgc59BP+OA7wtnLoqS6lf
CWxKc7NdYbt1VKvEAnyjOobmhwFR8z8NR1OGQK7N7Rj4FcDvXAN6NmY20X1NE4e3
kKNM13WbppAuJxIDyz7RnpAGLne/L8ctTQJxiUaph9NX/B46K3HoXQAUt5ZhOvCM
9bkS6veSG/uXEuYsvaEfp8q4//5xYYOWEmODz2OiD5n38kgm2+Rfl0LYIhaeoBCh
Srw1XJe9fP+l9l9IGa5l6eIdGkiVzn52g05TQfTjLtOMIw9E0uTx14/eBo/5DT7T
sk9dF5K1gE6Poo5pzqdSkio/nVgncrli2thJWIhO38wtf540dTIYGS0JVShxGghK
k7dc5m7fmVZCHighVnn3QK5GQ0oAGFgE/uPGN8Q5iTzMWTJ1sP6DXS0N18blYdsZ
6C/v/R7vF0gCyhStiKhJgi1wvqzElRqomPVjHKnJxVj/C2fl+yBqu5eiuxvS8rMo
FvCdJAFj5RLvTHxq7sHDrRyi4Va/ukZvgEP69k2eWdMniv6AOdL9L5vxf1xbqpnf
mBuwfXyJbYnmhpsSEQKItboq5ZhzgFjGRKtsBejBvf0Cp29yf2e8YLF9tkcJuz7Z
mIWsFtauuKKdfhkPKCMwhJ+RoUfzNzwp7WKZeKm6lm4NJzA5QndqgvdpeOhvLP7h
s3OEEO9eJQZJHHLaD9A57xZflDU5hTcOo/Xo1nBlvTOkPqwZK1K82TlXw3LgTYDD
LDwKT53HCIzbgkgQBxdI8NuojeCXK4OEF9+F0BI53/7NhwJzqgq6H1M5kv6v6r9D
fDwQzxQYMGGEJBeffb3PlxCbzDyJhd6fHK+87jk0AvYKNGJzKyR6V1VAIydLjB3I
JhCB/7okTV9Nd4aNUr/ujIyDQkKiDHqGVEA02CGHKXTeSp1b23/F6LG4L4Thbcis
JRvYS9ZkA7jVkK7kR0tHED97vyFpfnqGqbFMfb6AbNv+DjiNchjUaxoWEg+yBGQL
7s5nxzThE0ucgd9ChO03eWNNKfvYFbOJTRDQ6Ei6Kz77ricP3gP8lklXUzwNZvfc
DVnJDEjQ2H7zp8oOpgj/ClsM9lwqytrAuDDyv4VUTTHB+m9u/cAz4sNC+8cHwJdA
xGUWxXUaA0lzK6sCfoQe2/pSPFpDK6C8+83h9HK1ugXRisiw/vBK1UDpBixMi7+9
Dg6VpgyimYIdNeCp1sXr8MjoVl7uRxDqrVdUseK9lC4Jr3nnb0HxQpcxt/D57iwM
bogiQrjA234GsOAV6XXi/5ibqNq+Jxg9Dbt27HroWZ3DcyYCbzDFbt2btCQ2a8lB
xGQj6xgnwSg/2bUSgT1bkjAmdmJBjtGnjDj1bVhkJz1s5CGvNSs+eVXfiS/rE5aw
UmRIVHt8ijb910v8PCf6yZxWfewFv5YTZ6sGPLCnQXF28i8ZP3Vv02RNTELeeMcI
LNv21TvfrXHf0er+M0eLMWibGTgHqL9sFLnJyTklKfKW5LdKh/6cBO7PNSnQ+FyD
v1QHLitN6xMsmxcBnR0fhlY0Aj2iSrfAC1u7HS2WpjcyTA/yJtuOaEJ4mmfFIqtB
2OuYf+LhN58ORqeJlcKgYPxvBwjSHOEDV1KiujO9v+BS/SQARNSsHXdILMpjEQDZ
`protect END_PROTECTED
