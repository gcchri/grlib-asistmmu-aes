`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vYQWKke41wiac8WdoE1ocyL13cvyhi2l9/J3F6sT9VadP+XCjJdkXMsVpx81scOM
Cr0X9DuR4p6nViMOMljwIQXmMRUXsC5GdQ0LDPUjTKkfsMY896x2qKb8VearuAKz
VAsbiqKmKNSWHhLuaKy/AdhkSkN43o//kpU7Y34yb/GteYhl/xp7qq5i3xy/GmQ2
agbChfeW9/JvVO4IE3pGEO1mMpPZZNnN/n70jOicf3FOowRSBwyrSJaSnT1nL+3y
0UxSgyOlq2ASUNdOEzicA1L67w2bFZarqE8iCPnqQos4uNerXVGyQfDGQZRXHdNt
yvFYmx9vAM5U5fI31fMWxW3uq4JAfQPbLCVGhV4xWdkYGGr5R5CQK7kPbElT/UR2
lmxu1DRavYs4Hk5npv760PawyJS+NXBFT/lX/lhSkUENEetQU89p9MYkDATg0AUX
Bg+a8PfwDgilsqsad/hqbqLuTWrXGlC9zOguMXG7toapjqugff0ELrhfLr/DFCCC
+CKd/xijgNZGXSf4Oocok+SADnJi5WAI87GG8aE1fjFbSXKjjfw5nAmhOeQO3ixe
sVkmXDtotu1+B/vxURAa7w==
`protect END_PROTECTED
