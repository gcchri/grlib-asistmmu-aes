`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y4wXaoBeCDFuvHhj8OL1ym/6TY9fT/v2plW97nHegG0J1wOU0kbJXbuzhISBUUID
sJLz55oCA8f8fvVv7LxoXeXCKvOGIeY7zzCwYWBcaXmlJf5fdZR6lWh3uqhVE199
I5SLyg7bgxuIUehDXoWlUWFr6S0TJqESNi0NN3hnAatW1KooAp0ZFlgOPI+qePfR
oirJKkOX0Py8m1ckRbnZLTGImaj5qTabThhRG5W4SlvOflxONZFuCAXnVrA1SHZK
F9f2l7hwmzQ/3kk3CfZSmvNK1Fio/zESKs4U95thHFMbU+W1VPdkg69kuI6lr/jm
q0mjjfRqUqZQEy0pnBf4c5JuWjHkWq2DXmnDPWh2lwJ4AI/eOgkS9/Ob0y9BvunJ
c3Q2AAp82NkVBeMktC3WyQ==
`protect END_PROTECTED
