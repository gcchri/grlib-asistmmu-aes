`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SD0E6hoM9qXg024sNPx5oDslt3z6HQP1erCZaj35PpPoczFtSHErGPHwEz8eNDWO
Im9Xbd3IFUxyMZIifGHkjCBgtR77avuPTKmP11kDWhX1A4eVTmPlk2NVb/+9QBGo
os+5o+SzcnseQjblupbphAun8e9n8AwetCVW5q0PYjZd3PnauevvMCZ02Ird0ZxZ
SRqmK61fNtD8nMsqvBJm0/RNWI1EhUpXkjaOEN4M6f6+se0xhXfladFaWzHS+xD0
RxbEJ30mlIrmnCbacWOVOb6L1R0LsL10J4X4TkiVi5pveuqZPtVHuvPhVvgtNL4E
kwsKZKem1ZIz+5Z1jEgo29ggbnojHVgUmOhpbraaduZsuufkDdmaFExq8W3PTjXh
x16nWb4oXpUTmXU5NHEvYA05vPHpxLnBJGg/tE2Cn2+2XMsVXMmLNQkHKNHkarh4
7i3TbyeIM0wf7paCIRh66hoqQ5s3cBLyl9+G4B9mSv43pR+q6COoFvosiuIqfqO7
WmAuyR+fpWEHh3AgPpSrAKO8O/QLJnJjYutrF80Y/goDCS6w7RoRqODRPmk25dcY
L8vRQ+jzCosa5OmygHYg0VZ+K5aAeEDQIOozmOg+Vw1DzwBeSn3/p16q5coTbbvL
6vac/AjiHqDPhmxoc1VW2gYzKtlzyZOuoTi3Ly1wVDLYbyhWzsetMbaXfD/ehQeU
z8lWMxYbWG6NMHs0icjhjFzhxygZ4eQBUviUkrf0rO2mvkL+QV49LmN2L4CGDnp/
zZP2jQVRHYlwqThb3fLlwPJLs2NKMNAydlytfIXZioJrXAaQciDFQlO1yejkazOQ
lmNa5GrfWXLQ/o0Bo0HFQiyEikCV2+JQ0h6/1/O9xvq29zowpr87gqA29Ccu71Pr
4qnyX0iTK20R0rEzfAsHjmCNV/4s6Aj7RCjYvG2Hz2R8KZtuSqycp6p7zaJwmYkA
ZLLq5A3EW0Z6rc9RwmuzE1haVx7L8fy+3zYyLqPLYwWgdJp2YDFCSMrZzc8i1CxV
9v4tPSUmr4zQpVxFAliscLZUTDoie4NgXNwZW/v7WJMLRp4bTWqZ0t9oWiLn3yA/
Ad8PmpwDWiKqeKU1EsKVStuQeiF1rE7/LeC4LCXFkwl/+HtlYLOIGTAH/2TCk3mr
VTwmdijtHrDPfWFA9SdU3vnC0nqvLVKd7hG9hfQMmNfpbu1UnEBtPtRkq6hrFwX9
ZxnoNRb5wkWRIdg0w0vETqpu/D/r+aScwVi88v4gHjZMk821M+nhbt5xFtZ7CcZg
FFowDFe/rG3wj0EL2goc8qehvYcTEtZ3EA4KzJ9VE+dCTO5IIK2TKZyqU/4s4HtC
JhItiuc5/E62hWnacF0vWqNRJ50BlpdJcKDfWFf7EHIuIVNLTmRvnaN6GIyuVYkc
ex7bPfiUsw/qRVoZD6GTKg0XdYrlgCwo06MYOH/i3b1bXVaf6de9Slz46NiYYDtD
IHwxRm1p8iFcfeHFCQjyXLhuKFgTkMdouZpY6nF8b9tQPoamIS5apZltnHn9UTD6
XoTkS81qs1IBZMVDaqT3dRH8yc+rb1AVosQaegW4MMdMcRAZ/vop0Ae4TQK0/AIE
/mFwIQqSHvyVFF5SH9Z0Avb/VkO9rsxIl1t59dn0PpjDrEHVrsLIWABcPzrxyMHt
f383NYAUxyQ2kfq81Kw8lKkK3CRCvXMowHlnHa3EP321VHDpo0UOBMLq+aZeuK0l
ZzpBd8opSqpkqhqJJnE/R3njXuDuK11tuKoXEKaMM6s=
`protect END_PROTECTED
