`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
08nFEj4QovB/FjIT79zpSHlYRu3mUqmiiIrnyJhtShuZczN5fsF358iwp87yzLAc
+lRr6d0vvP90Hf3AeGS8lNybDqrR9H8Gi/RGNuFevKWR+aHjWYH/6D0J3Y3Iir1d
3p6JWzNkHWF89vA5Ks5k4CfsJBSeN4dweVo1wwgbS8kddPrQnbxT6zg5AWXUnCPB
ofj1y4mpfDMFY6h3ztmg1Sm2tzUdwuQATjF8/qilJob4i9rUaSJX51F5URVR0ZGz
zje6WsXbB0+BJh3Og+AQ02bQ0qKFE/9uaKW1ZRsgLQPBmTS9NYPXcnFVQKhl60hq
mSgfHMOyqUODJfGFurRXotfwZX5rZ4Mkw3ZZOXOUv3KpSOQzxApjUNxrye/0ASvB
CbTRJBZV/nGz1ZSCufMap2zHmV3RrLil0RcT+ZToFcSv3bDydMSb/uvP0IveTiUS
NXVqYpionrabHP9DB4FzBh5LhrSTdv/LBBvJXiW2t/fTshspW6TjZBvzjfMzVBM+
H7RLUxN8YEFpKxikHLD+8L/xV/SbMH/PrwI/3R5tsPgt6eUIjAbBggSybVJyOIzq
mvvQI7l8UJmxvE1BpR1limWV8vGzc+uwlfolRWIOV5m/yqcbb/1ssOrV1VwDSwA5
l/cYE20fioPYutyV2VDMZZvnv2+h71E5QbMLBN4WlRJ04b1B3bsJC1AsCHpv72Es
SXexJ0TXQoMmMmW4MVehBCAggvRl4cmBFZBPuJmGSnxBTOaXauH9tChObEN9FYo0
7l88ckOxvMUB26QNUutITpRA9zBeMXqwqON2yvDdJcDDhuFezAO0QoBw+Qfdyamz
hQ3ndbCfFqoeWFqZlegX8sXd/NawDrfbRhfZH1L2uR8ajd5ZupmpAEpn03I+ru9U
+ETaMMfcssD4R27FRr1raCOOVi4PCctuDckYXDhh5zj6NA2CBZrl28PdF+sQHpJV
4VKU0Py0sb9u5zA1utvzGq82c9TqqED6nObwmocNkqy1MlwYqIrpGRppQ77QQFWy
vUKc3K1+aKl1SG1MoNhtRMffD8vCLYtqLMPF62PLhRdTNgGbw7pNfb/fLpvaEwBs
arveuSMtwXV9kbMvOBeFpiE/qu8uL5IYfkiIC+vCTrsBzte5igld6VhGlAKkSp8f
1EOnTF4iomuxsRphoFLfD3NqrVFRija/OzKL1pOsQ7KYX7sddl3rZmlTfbjDB+X0
nqmXshhwmypgbGWM4VE4CQ==
`protect END_PROTECTED
