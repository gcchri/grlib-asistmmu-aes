`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ONBMyuTd8A/IGVRe6krF5iqu2a/fMSmls9vao6GGe5Z2cq8XQRpZCpc0wlHn3kru
yvM4Xu+lHPXOKKu/oewa1wzmhMxqkz21biqWe6xkh4b5DUaVgRl3/1w7GtozsSJx
HaPE+tOYYVCTpDkuoqlQDsIIHcpt7max1ZYYbKrMyIYzHPqJyVxHvvpPtNtO/Gxs
2iqgsm1NBTGv0GHdg6OFLpz4/kfqxuR1yBQbunrK9d7JIYMN0zwaqz0eAqqCh5K0
MlItspv8ToKd9clzLZZOTqSCY1vDMxHUKTOL4Er1W2DAktz2jcqLeSE5sXM4whll
dYyDTf2d35I0v8jo9N0sInnHFFfSwAR5KoyXDQItz+/owgksm8TPp5N0nFjHqIxs
uAssesjRJIqPgwJ4SgAh+q2mbDVZ2bJwx4e34jhap/xjn6zlzm7zvAMJQLL8mzY9
73KhUCvjh3kvu+MpifVELWC/cSgjLrct1Oo/lL6bp/mA3lCIzpNovgj0fuiO70g+
ob29HMEXxUTHcxb9dmak+rq2BHuwGmhiIC3PwmumRn8prupYGdIDMG6hIHU7CG3Z
gyuN/XfYYlMxohmh4Onk0OR0A+hNPYCnNcgouw3tmbcAIttXhvIPXUn8eeykprHb
Cjsy6ajjEnEn0Z5MV5wIsTt/v5hoJ7e27kO2g2mx34fEUR7GH9HD43ycglcKBgD9
626PPOR2NXXj0J/eEGqfSg==
`protect END_PROTECTED
