`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nibN44KuEgup6NJFkesqFXNCTr0u4lM/FIzwe4NPYMAofI+bnzbCK99SxEVxI4Bt
qtKHogh+c3nxGm3ltbeqOlmDj6ddio6N/yNcA9FPfJBwxsxDdvAlsxwNjjtCg6Q/
IsSfiP7hXyxwkdZQj1OQD55qH5rUnTk0CdK6rzJzTThByA5Pd0uzhmS1wjTOfl2t
1Uwtg5PsiMozo0k6DazJf45/qlUWMFqOxIg+yIbMkOyhB8Vd7ZQdRLKO5n8XpkuC
0/tDfW7nzAh7rRyiN5+lW9EjbwlPsHdXpKUcTU02nokDDZgv/SG8yKgjln4lVg41
TzUs4RsDTEgCYlv3+/QYXmwjuz8Hi2PaXcONKLPRcTChKP5Tzb+P3Ld1nd89VB0U
dO4jmveUlEeKAlnz2ToGt7SP1qpd3oXPfx0zQE+Z/D7mX2OCJbUXqkdaeaGmbe+T
V6/OeHi2QhC+VQO59uUVzhaantQFZgPo1MDbsWrHH9rDaojCDDwP9SxHgsB8edGl
EkjR0NflJdnbmz1CqwXGbST2+qSwN7FNsHjKgLCwoFGx6Tg7tH0OvxtGUurrCaki
VBgFyuSPuyg+JSN8aoDpfEM8PKaVxV9cYXywkg72y2YL4mCsbGTADx/fyq1If67U
clMiS75UiXT+KUsP+eiBv4pb5IdTm5ULMnlQTVb1zf+/hdyWsisiOx4XzfDRqR+3
Wjhz/IwL0C9WNSquGBhEDIGSSlmBmQN75bMCa6NteG5JfCTK6DDHYoGi1cHbd4p7
W+y1+SI2FaaqjtW3CJeJEaxWBipTZAxukB1/hLBDx8ltWEc2fVph6r8ANk/i36kx
W2NI1gq4xMF5WfZ5JN9KjQrjs6rZqkCxQ+UZYRd0eYy0VQjLV8jSFrY5aoLnoows
bhhLSMMx0JDae5Y1rjhx3QKhdP8tyDooCXjJNs/MiGT8ejmPD1Vgd2GN76b0lcOj
WC7YmmS45Pw4nCWEv9S4ElNK0lN/hO/VANtwK0aIWUInkNs/JMfS44/hVKwbKwrm
pX0QgLm2jFZfJ2jNj8SDmG6SmdDqjp7NRS5Wmcyzsv7ELhE/dx80xR8VMXG1PvPV
zPYldC5MrxLa3vWcRExkt4DmlGi08gb9fHH7M4F9lmDCfTnhSRq/0CbEl9kE3Qyu
e0BV6+nkCk1zj6VwgcfE/mt+cbZkWQra2BYdYuI99r3U0c6z48ubuqg73MdPOLTm
RcFqLfJK6B8S/Vt6eG9kaPZIRC47xnXd3uQqYdD4QY/WkOEpBl3xiTQvveDJQBR+
QJVa/fvSZOTB4RoP266lEcyerktu6WRrwmgBY10Sgx8LhuAVwieJfd16St+JtkOV
rPD5Jfi7O/pqvZHlmubAdGN3YODzMRzdUfZD/3MQwGdZoCmktUhh7HquusXSurOE
ixT8CdFpBWMptAz+EQk6NKQoAJZXlutdmI3sAl39Lm4AGTIGtIp9cGtkdx+aVCi8
mbrM6/eye3i1WX4aFqyOdv8rQtFPabLB7s9Aah+4e1eNziCcaBtbuQ/+omwukjkY
WC4vigwK1UefSJm/JOyjXopi3bJqi72dRWaSBsjYvUZThQJ9cI9pvZNUyxQlxAHW
1zVfKXHRszthtw7YYxn9Smqqx6enClYVPz52a9VC3G1IUL0yRVIb8rwnqAfMtEgN
tOm+GM0edWSE2mKBgjkXzVBLvmLiWaL9GfyKnQJlII2ge2sRUijHt4Gt6gCfS6of
wsNn1L7LfmC9iK8+axcb3/TOO6Ko/ICkT0kCLqybof/q0DAoZ/eFzaaF0W/TETUt
ZHBgQuGVxhRryWUwBHTkUqUvHmbEGGU0lqcYZPswNqIkMSTRGTQ909K0ZTlUOMK5
eIe9sZ6hc1Lg32GMskrrcz/zCD9Y0bNXCBW/SyxOLvHRD+xB2HcrT19o5LgqI6wa
g4TW2ubZHUs/LBKjDcr52MoGghjABxeEPI8DcBj4eTAjh9M3QMOSwvuLw0qu7nvS
GU0nZ+uPkjb718AJ3chxN5rJPzrPuWVEcoon5qIsXbuneBVBvydZFdt+hYhNNfk/
NM3O6vNhCeJ5hinJLd/9flg/1N0fKXfJA4hYBilufQSH8r+KXF6j5srDA9LTzihZ
f7v8sMLjDjiZ8YEW1YdmhCIzbr9Jvbtd8N13d4AYwccTxPJVUqNj21z4r3s5pHk/
0loXmpCTKTykIuU6jZ0eK7C5mD1lc2iHfHs58LikfCd+xkSNmZbfxvJWWcMvB6XI
KSeZ+sa9WQ1tmwyEXTbQZrjI9MHOdHedHv8ffyx4Qz+TWIQ92Lvf+lDrbN97Rxa2
CvMBdz0ZveoReLPRdyerXKew0ofrKQ6+R7oTl35Wwy29N8qMGtQr879PnzcpYZ3w
1xl6QMXIsLw5NyPXTi7PYSiMK6oDLnCE0gaUmSebsMvFIxQLAGvd2OuxpCVug5eE
3bBeH36wDd4oiaexwC0yfCiJnPldDbERwQJqjdFKjPQsSoHB7/bRam5Rc/G/yxGV
afQy6qHM1OngNbcRz3sBWmjxDmXgb/xCYYo7CaCbfa8nUqQHVwcoGTjc8Np+qxCX
y0jF7eQXwA9LiDi515JCL3szwjRoN7s9QhyQaXuROSvKM95MLWz8Qxbt05HCONRe
OjnLasDZrPOwMquyFYqSVYdBMPaRubscFIbs6rUKKXBp3nDYDL8dnTrQYrnpg9fQ
jCx6byyx1T0ctm+T0sNlWOyk8OTYOU1l6G9fZAcpGngxXJveHk/OZPrdDKaQvxjK
YIn1TMDkr+yk4mwV0pD5IewbDwP0dDHpY/4I1dKyaoGqX9tkgoU54kv0OUdR+iT0
NIJZ7MvBWDNaDKsQP/z50BJnp3Fq1l/KiMUtoouyDatK2Do/j/gR2bVRZIHPxDuk
9Vb/i50f2yGGaRBAwKYQqdPYwE27dVy4FRjOtk0oI3H1hVCnzTWk84ePd/QC0AnK
UnhBgit6jdMCIjTCm819N8A5HeI20O8Of+fngTZ5ldtCnioaPqIiYHIHBcs7fovl
px4QYZRUfiWeX3O4lnLYDgTu2z43sXIHOEFGk3UlKc56qGEJViIb3IEbCDVoLvs8
er4jciXbKfLIc/4r9Iwtq3mq/oHLyCldP4s6+OVt8NJM/FGfYJERh+88KOptXWX5
wCDclwbPyU+Jji5vLA63FOQ+JwrQQCyJ4h+aUQ09nDcd7I+TBeeI3UfhI6IccH9Z
f9qn5s4r1kiAcwJlS5eI0FnlXQGyc5wGU9QyB3tZTYxRlwb+kOEHXbB/ftK7n5Yv
rWq52TRkV/zPN5o8P5ioq/sd2XHWLev0I5q7IqB1bNYPQMt8BsAMpN5ep2Y5UlGV
dq+BJKVBNQoBF1qdB5eMQU8LJQPqBaE5fDmkT3JAgSe7kfVoDee+Bpo2vCvdUIdI
hMdN1/Ak+niiP0ggr7MN0Cwhumg3fY7oIdDMNWpAnrHrLHyLzS1iQBBH6U5w50yK
/tS+JCLxRpTcPDQaJZNuD/a1vDy02ay/Yk8w/GPKWtJmhjsaZkVSsSg4079TUsQu
U/5wNI5t1Z6C2+6BCFSHJ9SdX6LO4cPq8XH1FQ6k17hPy8KMjl5wqrnj4+m4hwkE
yLJPsRy6Pl/UfrFKkrb5D2F0FOmx/VrSvoG/h2o63TF1oYCoSVKvYb0ppYJ3gD6f
erZE2WE/cDS5jJ5zFVItWgJTAYKOmYGxNHQm7aW2f4FLxTLegL9aKcmuhtyYSPZB
HORmWuUv23IPXATPumrsDCFP36o9wbyc/Irh0abDMtJEs1YLARa9CBN3ylrzVMe3
Km5ebVr2mY1V092qw0yxOAt48v6rg4A8eWVOCVde2x5U/BeEvLbyMNnOpLRthmdS
6DCpRYVRNqdt5nP3N4jFVWNP/uJibRD0HuXSRr8CG3ORf+lb1cNkxmx0btSBLpOZ
HDiEFcvLTxmPbj3mmzPi76WGjjzc0WXhtdFgf6qHE5sqxXCgwZ9QtOeqan4dLkxr
9oDtGbGsWzYX/xoys48KGjyJTnrVmSPUXwb8EIkkg7OCOieZx75YvKdqF/ETSGV0
DanbGoeN3Dg3W3ZZVwTfOctpgpJH9hgQfxSLHad7/BGQg7LYFLYaxpPvA8DUJnpl
cICLHUR5dsUc5Ls1/q5Ti4isHFbUdDdkH7FG5WO7cf8/QCKt2STQN7m1iPtfzKpS
gatew2h6DMNazXK6eyIu6LGV9nFp4cCAC5DNix0fPlgzftvZFogiiPMsuwwZY9YN
7CLjrIcXiDcEHFTDpqNQeg5M/7JWadnWf408+VIimkbdaK5a5ZZNqUcGMEpW43en
rzGjm29ASFM9i/4ekeIxNTNcMJg7XfBhVv8BuSZTxyFCxAsM8nNf2rKBtgbnfVr7
7d33o0bXAyXlScovWMQfywtYF9OyhsAvtzi0NTWpkOi5cot9d1/YcAa72D/pqo4Q
bnMU3AI8VKPhG2IpsKEYD5++gqzVMjXR+TrpHsDYT+jfhVbH11TRaoykD1JKwrjj
+CH5forj+uW3aMb1v/gW3sLq1s7j1R5ywknKPKamfgZuzaohQ6eSUKUSlubZmxe8
CFwRIhMYE/E/YVhjKGv8HYsqhhV2lsF92FLhVc2sx39NZXeuZDUBZj7CM7hr3e4K
PdQfaHB1S/G7U9RNJioAUdsY4BdfDeTbAAsqMP9Sh2pquJaJqnAXAcxbQlw1BOFE
HvJD6eZ33HEPb6EKWm00wbU2yW8wz29YgwQGB5s9w1cYqIUoH5SqCO7aF57VH5N5
D3VY3n8RivF5rT9aOnmJTNjo3aVxk0gk8QkUS5RA2vdzpSFdDsBqw7TN6h7dp4zx
+6I7Cp+A1lb4n70tfnJf30tY99qZqByT89b1wBA9f27buK7KwsYq8xmKzMwyVgrR
9mE7b+em90K1bzNZj0uKXB0NlDC1IzLuMhy9XojXiG2CzmwjY/XSJZBCD5UOSvA0
2gznP9Qx0Ao8KipmHbWjmY5MUZNRNCouoBcBmBzXADZU29NcspsOC7up+mKA1OxW
IqoHGVrUWv2j0ZrsgQQ+78MyYa+zgi9xOvdZZw275DGDLoFq/4gJV9a1Ztzi1Dxz
5Hn8UXUEQIP6aILqR+uR/+l8sbUbHKaVR3EBeU/DwOk1JvWWkSR4eBrc0XXIeWQr
slZwUo9xN4diTZW3C2ODopl+PMP3J7Skr9dm2E68yqET8VZ8RN0FS0k3BkxcChhu
lVNbc+PMX1zZU6verkOyV6KK7ir1P85oXc3NUX1ZXgTvuHr/2SbbTiNphGykrsf6
sv3Rcc8O2p8o+ySRdYWAfmIQkDz9hVS7S+Of6cI/GJqN0QxnLA2jkBFRrkFteHBq
z/GOkKO3pWY/ZdcuPgomdsvBuNeGnP7U8yGwubliRqghdwZDHdvQgZa5q4uwSAQy
RTimIJcohv5NhotDQQn8YrCo+fgUR65bwbHFCkpqBxJ+KIXwnsb0GtDRDod7U3od
4oUNTVTIpfNZ6590KR9lrHK1gdXoQEXzwEjWZ+yeGSGHSVRV+fy1ea94kHiv57x/
ln2WqYKQy8K515mgFf2K1WQtsUVJS8cxf54UVBMHilsxn6JP5eCeM9xmM4HAYDrE
ruxQD9qh9JDq2m5IQusHY0ouK0xRpNjknGrUfXXFAxu4R0tkfAyXUTJzRgQxKcPb
b6htRs8kMf8M6qWWgcsAuAG11OnHpHtCy36sZyPF4d8zWaODcHzRtE9JtIg2NRta
i5a/9Hlh8U1FUEz5vPfBxHAnrL/bWMqEbc4VSswIHnr4gGRnD1CGbx67Lo1d3p08
iv1OERxFRLcbBINxceTC6vuU3fRPEGOwCXeX+8nXqF3CoAU+bf5KBnu3LGdzzxni
+d9aHSGPZwhobJsBUqwQZPUEr5JTjMVSVzQVX/1sJgShi5HsuUX/3qjFAvSINQUF
XG70WWafA4P+Fax+idJCc83WepXonBQmby/RD5jEdVpNg9+yDrnIefftkecIdJ3q
7on56oVjxkiISLyocRgQN3ohRuIejZkT162e9VDKyyh4PbN4/1S4xCRSA+F7iQRT
l0CcUCt2rGeDtVbNWi/m6ErSGZ/s9nPGziBnCH5hdDitpeqlSoSkI0+7OUbU7Nyo
yYaBPaWBthunTpzpk/o9HqjL2FWxgawDYxaDjVG/OtcWjVtGKXPS/lAIBzLgpiF1
3gRELrBdoat1l2qJD/idtFoH1MRt0pZ/0SqUIxTieeZH7pVPzgkAC+5gGe40324I
NaHE9TJqzlSHPJF1fTqKZGUTdAMV/xoaJym588FBlgmanBOlEyORCn4YVaA9NXGy
sHjm4FoypMVEaTpQtJlH6BsbuL/3EtCVJH8GwnWzx+cv2HXRp9ayk+0bQWimPcpJ
yAW4kDsqCQDnkpl14142xRQGuBiHD3R7x3tpVkDu4VrzNfrjlvAr1zu00wbIBHfJ
+0fFtq87H2gIBK+Fgv33Wb+LA+qT+bvbpu9pw9P0S/B4PiSKno/KmPVeh1gW+gg4
rDfTah79DEiFm3l7lDFF4hDNuDlwAGvvJKeVBxofL2b0kMIwUwj/YmmDysfw2xpi
NL3BdXOAEpuRIUGJlVubl1/8ybszbKRCmx6qh7vDYWNfrlPgdk/K0AqigvbcZgz8
cdtzWDMrxGfegE5MA93NOHebSEQddD0eJc143giGwraOSyVYzos7AC+k6ACoKcEq
kFAHI2LkBWxQ5VkTlvRolKa6olOV4qX4yOIVh7RJgANPxTVu/4DK9pRYCxEAbHqh
vg4t+Jm6JEKyxaF6P1U6yL+U5v1VNbtLD7CW5cW5dlPPM19TMWV9bMbfX3RJm/Q3
wXkiDQfG0gG4EE1tOLkzB+lwKwkoZOpLH0NLxnpDMM02A8oNiUzGLisZpXSi6jfK
dd1FWEX1OOHLgSoH6eXikUrkhSDip+gHhOJgD3hgOOgK/vo6t0+jwShNcbju55sk
CXwh1OB568VGsNR/D4K+K1sCsKV+C42mq4ipimSKeBAFfrvDPwovbN3vRelvsKpH
EwwUmTkJ+QdvUfm6zzthhNZv1aSVPpfcpP1MKYfFYk6C2W+Qewr8JTj/pEFYayev
LOBLjUDYagyzKOG6ptrQB1uf64KMKkkxaIlwj5RH0j+z+HLQuwrgY0iY8ROmNzTD
ODyTjEPCNYLo/b/gcfhIieySX6avI9qUaS0ORPwMplGLFLFPf7Rn1k8EBvQmtixM
791mgBc8FfgKh7GWlVQ7JO6nNCyefdTwrp8WMoaGE7vvLiDEjGOqujTZ3rJHHgfJ
+rsXaVFXKlZxT+xN1u8kWbWxo0WjY30tDXTZkTvkHfxmJSA8q9ak+Kdo/tPzA3Vz
4buhNnE1+yEq4272Au/v3Q6zZvSKJ9bqDSI4FqZnAEddyHPXOIVK0cVK+ppNJeOQ
3F/84iSSZx/jKIx46wAtY8Gp9sQb9Sgx1WHCn/8DswYuGEIv665eUKb8/zwxEXaE
5NCPilraj7uEAisco8AiPvXICi0l35rgGFT07Rik3cp0eVlzBT3sp2C8GcvBi0PH
nKZOX9eWWrq1Kfjfpw83Gyc0Um10YaWzrxBQLLRK97eHIlqUGNTSAtUmJnz3/ZOE
SF5NtK3mHGmJCtDlsdOR+Vl7ttJtYW8VCHqZ6jag7V/LsuEZCQUFz5yaIw1rYY28
gn3TcdLnhWKm6mUSYcM0q2Jnr5aESjHrPV7n1VbwrNHlFxMTS9vWlXAOMp9V6K+D
GzE4VDeoMAaVzxHwguNkwrzBh+AttvV39QpJuouwDvmfhS90Bfa72dbQI7xrIUd6
6kaViXbvRLLuVWCvQaBSS8XNPhwP4EBuAYhsizfsb6wbRW2HTu7HWWsAu4qsGkhx
dKBb9U/OkMDtyu90ARc/7pFeIeLLYXJe+JRYUtir/1MWlysTNxZcWEfmrnZXwDyp
sqpvnQu04VP8bBG9UX1eX5I4FC4A3m+dA4XF2ZpWpe17SCPVwUOzn5SHXjcWAyNX
AXRAH5EMXoanMejygCoqyfxQKYGFmy3djqs6cQCUT2EDnAND9Bb1EMkKl53hDACc
vL//onbYxvVLDMFOnZ0uLertpKmMadqOFhxrFS3dJxaicKxJLq7kRzOFgR06yCWn
n8Sz6+HRx67nBnhOsDQIxRjRDA/n8mUV+kEfNBzq30rdsKtJearZPZnwEUcR6sPc
bC5QnCw0/G8KeZjS1ylYmeGJBKqMp6zillAncb06RYKs4csG6oYInARKPwHXxUoH
xSsGHE30Ith1WIcqv/jwQW2HfronD0T8IBvLSMN904O0Zciae/GhEL7nsYN/mDq9
cKSYlGOkfjAm3aMGuqFJf7wRA2qwqz7YCxF576iLsZHdacrZQGavsdDTU8bVidlA
ZXY1SHFQQq8cSHKoycphyHkBpbNATV5E7r1cqYFUDbV5TKuScBUiyhw2cHzAugeD
Zwy4TIZwzh/ofyVOyOZeM+/4U1bBxFiw/K2/mf2lIbkB/62Vc7RFsPvaCikKh7zl
TdOVXx4d1mbPAJP2U2K1LdNkkS0VmDTWXQHsnqMaLViECUKwnAh0bLL48yX4bPE1
5dOB2ElTuSvezgI7L+0+2w4jBu6Vw343TGx4zDCXNpQRN9403JTaKOhfW1P71EeT
ec2IuC+QmQLIIchce7i6bpRtFb6sObvBb/apnKcSG+C1mfONUISgVdn7JcrQ6RiS
ro1DrUVxopmDrtEN8wW/lMs6QS2r/m9n04WZtXxYFmrh6hT+3AUrPQepkZJhvXUf
iEi9U2d4HXM+2jaE5ikARHYC1d9IxIuUWol/MeWN1rBh2QcE3bzgtBfJyMWk+Kk5
BzQDv3lVWKECSvAvw9gMLNCyMNNp8EUXgrUNKx839exeUhhEkztY/6hUVELyU5l/
cqLBEg0CphzQhX4m6HM1jpWGjdBrI/YsA2sWbJsNlaeInMgm8YWVVDMY0SGSk+1h
17dEoUz/ZwM4TsKOGuyE2IQnAOQsThdW0OgPm/b6uCya/Pye2lkR2mxq+IYHTPZs
zemyL1kqWdnD7ZcfZOf3UPBaWZ9rSLix5eoaU0PquQJRgvsdAGyDc7R2uxASH7kC
rSh1T6jwHUL7/sQI0uWWAp3ka3iz4Zzgjd+sttlSqawax5jZQvgAjUgNyVSZpXCe
j1GL179dyTOg5xUpmXoaONX6vb+0+mSGdxnL28lqgaq6EgVHTVxQhE4nW3H6MuX4
7ziQqtPwmm867COG2axeotnO8Hy0NBrv4qIasHqvgDZpba8B+9QqMmNGgY9KAsCO
+hwuw97PDr5bQi6n6giLWjr+BhJMA8rDEqxplX7zlNpDN/Z2Q59uESSBtPkUjdko
ys94GHC/IUUIXRqo22t1aYPaTzG+1HUDqUlozcZ+Z41s9yLSv2QZgZZKqiLCH5Vs
LNPPBVXLxoxXU2XrwwRq5pWr92IUonAXPnTeS/rKNLNYlQIWz9lgszCcHeUHfdin
4Wbb1HHxoiP5er3sFZwNPFcrOcjKmETeCcrLog+LYb/Dc8X3Wjkljk5cc85XdU8s
/eEJqTUsy6y7wbxrmi9n/FD4rSEamP0nDqaGaNYyDN/9ptZJnUURx214aPjO9A5/
g3EAamrOQd0aQMWsC/9lMy5s4OdnGRR3tt7BSUomCpB+9bdFP7eFkMdYj73t+lH7
d3OqW3DgcPV3/ed2n9uCokEbQ95H4k01v8VbJMHgD8T25qZ6Jx2EaDErymu//3gJ
NKYRTVCAydnJuI5f3MVDjdlx3/YTxQpEQSKXYAbf/zy5ZVCprRn4fY7iZKFTJqEw
Ux3hRQCqpIi1qq8s3fmNFxZlwkXd9I1cmYARF5Cg4tXVCyfA54e+tpIxdidFgrB7
oN2murZHDhqn5+LLPDVwOOQwZ+g11WOoXtBKhdZtIXIT1i5xY18QWbCMfuSN1wlm
RgZ/IJpUbF7I1sJtlGfF0n/kHTxrHfKyYx0rxAEG/Xfbk2oYXeEKdQpyjMIFSF+c
2mAlZIWPjw8rEraSVvo0CEN7wVHVDIsSb5WMr0sdpUQnfAnfiRxyHzKgOlRDnWoY
chU75fs2KdPZDyZUAUtcP25dR1Xl7ZXDE6dj5dDtRO24jUSHS6zaQaAxZLQszwrE
F+EC9DdsiqLWqGrcB40Pp+ccvZyKUN5VSrtpNE4id2zkj76VqdeGyHP1KsDBM/fe
qlodcoLTPRo0PcXnZXCkVAGUdmOEPgxUNZMptop8G0Sm6OXU8Ne25/eqsCJaeIys
pF1IZ2fKMc7BYNaDxAh7ouXXEWVmTPfsKpPlrUOoli8+7o7IwO+86eSEhOeYrTCi
HtYkIimqMILWEI39qLvBNlZlp1xvzlCTT54ha5jHynzpHYN+xC6IwplFRK1dhOE2
XIxEYP82KGiNijOQYoWNLOnNwf8ryET22BleXRa7s/175W0Qf+JUX0XmaopnHxP8
8awQsc7nE1kLeJOys31uV7OJHjUfCVOKl04ev0oWS4KnhghTk87WNKeLarXsd3do
orUPA421tD2Kpdsq3UBAjVoFpl1cbQuJSypvF38vAnsnoaIhMhEpgSgPOgVVqm22
EbTxh+Ys33zfDUjcDTt4eXFhpMcfCtdm39L3cZirDbYi18qjLYlb0lmlbP/vjzbo
NWi/jcaDLIs3vChZ9l+bfejLWBxSGKsssZyr/hxIw6mgQapQ+QUdaRh1xmx1ReRJ
6/yxdxY04qwTIM2qslnSWfshFS4a6nR603W0TEhhRf+gOaDR+MR1JOAbXbBC1SMM
gHZeBeH5lpyrZdv4DNGyVZlhzpUFI9T1kfc0KGSTKcxucGNYz0JSRsk0YH1KnA0F
TlcRaRUzwUN3J4LsgXCT6Z7eLZUc4moei9u4g8rtZ+kTLfSBjqX8kCKVJGKdHUZq
TuXH4s55XCUFGPUCkdMmXuokuS8aTfbCQzt/1UVWMWvA794gPHqFm7H0BF3GyHwk
Ewpqkjec8LItgU5cua5SZrbp6DiMUEznURvp1EavGLy6v9hnSo1+08xDScQkOzwy
UxRe4hK8kpElKxkMTDE5S5PnSjpATj9ejiD9Q/QtZkrrSMFDXJmguRCG5x8bKX+i
PtcAFx5XEU9EwC0ptq5A2xg7REFt3dZeDnInjdYEyqi69s34GIW4zU2sUnKNJM2n
PineXsYRZmfLqqJTlV+5Q9+mhkRbE6WY582j4hm+UvNwm69ETSN9ml0+5jFwiuQa
jLJ09jbcB3vylnkJwdTgBBhApTR4Uyun0mcD+wZX7DBwApRKs/83PVPFlrFVu3ms
lKtbP1C7Dr3KQtJWnWLyRbL8BsR8Srx4x50GCW3NrqK3qsalwmakEAZMMHzAvBD0
EpFowL7pA5ErxY5x5ujqFYOuuWeG3skDw3807nYROLvzXKbOto1Of0DcIVmTyLwH
AfF+fkWWISsmyy1IQ90BfwICxtVSeK9JpcZyC6RX4E6Hx5YQw8hdjVCGfGGL46DQ
ef1yPU7bw4Z+CFkaaZKPOnCswClEDVXk/6sAeF4JNEODBCsc7O8oRTxdJLOfuUVp
UrUTEe097yU149FZAWq2p1oNnPpD3PydjO8KKzUzryb+GYacZAH4syR5yUJ4tlSv
FH7pQNOPzVeQlzjztt6gy5421VF99lFOzFlrsCGOQWlfbdCDpgBMJPbFiw/+5sOM
p2jUS3MGj5xdKs3fJa7MocXr8/557EgMq/unigrMzRK7THe7fureO5Mx38cYV8Im
teN8DI3DepHZ48mzc1aGAPrDGiSmeLm4zOLhZ+PS09ydsP+jBTRKFcMmN3iu7jVE
pnk+U9EJN9H03DMoGMG3s+xyfszV4Y18/OX/X5ZFF2pPCi22KRfkZLqUrvNsgxXG
oyQcbEz1CMWRGwl9qV7fN5SBI+jospP6DSfGuGkQiX5UdsUlXWR7XEp3mkXTkWyt
IS4FVlDhq5j9+9d83KFqoMa2be+Uqgm/spactWhuUUwFM6IHVGU1YlUVWt8ARwAZ
cNR2yqut8+5MdKpNMd7fJN/wRY0Edqvy3bEFn3w/8VPf2SwDaxPUq0jro843lgPd
FdE0PLTyrqQY4PnueV4WEsJa7Vo6yvPHrQVHySQ9H51PHpGhgYN5OQdR3Axnsn6k
fxrg9dbkeY1AyD/j7bCv86qq4bYexrSkuDTbxboKerpMgiURq5+qurF/T7ONb/aV
eiMiPWiRZGI3PudqHggQuL+JWHN26vT8LjS50lHWZkg=
`protect END_PROTECTED
