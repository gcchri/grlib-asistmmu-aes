`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ue1RMIaNkMvpPPsBWjYDNn1KmWyH5xoIz+2TOwxSEJ/w9OFS72rUwpzXmv7t71kv
n3opubP5YpDioZWY6OLFtgnDf3f7TkGTK0n78y7N2K5QuWe9iWegvesJz9DPTB4m
WRvcf50JJzdQWDVyPrYgX1IgTRU6kcxyyYPaR8mxUdeiXJ+4PEix7m1+dg6rDIuH
bhNM1cU0upUiT2vzwhTLv2hFu44kD5Si53O0VyWlMagxFE7xTf/tpLU0JPkKeuwg
DfzG0J6zRckbgI/cL37ymw==
`protect END_PROTECTED
