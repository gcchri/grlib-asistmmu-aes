`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DGIkeBfONPBpbgjys7ZiZ52dKG4AQmouZgvt+f778WFp6CEodwbgCOEaJiYsgiZY
OOO9K3gyvE4l5kNWiaFVjb8m3YJJa5KPN4alA0zfG8Vx/yVmDXlHk92gVHQtDbw9
1twT72MqWrCf3WF7ApQTSvwq//ol9+HZ0gBl82NU4OFxeYHvfDZ3Yq1JadKwyYks
MSiLQgURfG+Bi1dj19LqhHFoLeZaXTrBcb5vzFZqhRLMpDXBCWgNHYAt/I6H/uHu
IPMUY9FFjNl6FCUVRtC7d8RA7pktCN/h7RtcyN7GdAMp15UAOCH+inqNvtDQN/Il
wfopXFyiQHqTQY+On2oPQlc3QR/5uAASJd1Q8AREuWhh+ylKBFFJgZDHtDW0b3hf
eZpekhts5YHPgIkurbk8fQL+BZcYbkr69GQwdxTLgM0+3sseGo8oHJ00YKY/2Qnw
gyKnP4RELjVDlyfwmVuGIHdtW+HvOqPzqnW/hkMiO9nZrX3BbiyKGuwVZ6IJbOSs
`protect END_PROTECTED
