`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z/j1SWiUHV6IKYXpIbTsCqZqjv7B/1AsaQUzjMdCTwJd3ohwNKOTCQ5PATdGoiLw
3QaKiQFRC6RpjoJvzzGMgA5qs2k+KXLujatVv/hMz/OZU6Mx4xBf/uJyUBo2XmPv
2Q38P+02iUuOvUXlJInYRMz/rXLrpA4ahN9/KgUqUuSEYa/A2b1QjwUUEqJj5IJ0
j6vkIAlkYDn4bsZ3IBR7FE0ud8e/1GVutptdzKg3dkO46lraQphNPNOC0h6jEUqx
lqFokhvCqD+0WRVBAhPCmbVTXl4LEsVkjdMu8nrMWS/9eW8NQjN6Ay7ddf+gx1OR
6W88GB2El/CJm5f3jSmtLbN0uPb1jmct13SP0IUZEG1Jc4fOmp2VFF37Zqi6HntB
LvqBYAMfo7xGXxUDQ4EnJhjIRJwiqylm/kAOxc7RToMdBBuslpZqpWCqlT7eo06B
QAe28WxJXqRfTuDmHzzDZqtDnzgrZiTufuW2R/2Z8Ts669TBw7+Y6CCrNRaCubgY
qBRdlYEF08oUhKndVdLw7Ld6LAynCU61Lyd9fUo32PqVZE0uqX6nUOQmGcaFE7ii
znm4YmmI+OJVTLnzYjOaw/qAGO5FiAanIZGcBu0Do37JDkrkxdeaDd+6ivTISyZN
8cJRIWDdBQzZyTbiYjRMCCjcw9TfLPbtzYyLIEr10l5gtoKo+coIMnu1mjZupPM2
J0WnhJwNu6jUiJPbdCg3ig==
`protect END_PROTECTED
