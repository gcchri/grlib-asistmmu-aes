`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QckqyAUlqp1xX4cl1r/0E/wWzgrVNxMVRXgKH2xaTaPLi4EHLbDQww6ZfRYxhunp
KDk/RWIKksuh2AFqJI8dm1eYDFXsYi1ZkUBvcZuBjQtBHu/xVIhyY6KwlQg/DJ0W
QMjJ/eHR+XeypBAsqQB1hfzFwzlrJ+ugEVscJ1YZPLyY6Ta3VCdbLWAx2BafqX3F
shpmB1d80LqlFXdd4TjPUGd9Z9NP3xvkGvuSgvu9aDm9e6MYoPNtxVGKiYynQy+D
onhEpdKSvzl+OZ8+jIqMwXvCNEdudvzj1ROT65blE1KJ791wCMqkuYBGANHzx82/
9IkghxExOjKBFNZUlK50t5UHpAtUufCNaI7hTEUCp0KLMbWsjcMqphbjPToXzA/O
Ihba3l/ClaRcT/Poggytt/YzAzu+dpuXf0n/nb2bSb9UrBAEl+/v3RFLyhrp3LBE
CEvEur9HE5WtriChJhUIfaLGh00DEo+dyiYHW8q8ns9mCyV1T55MnFdEeO66UIOP
UMyFMaSCo82U5+tCLCEtc2X9A3v4uwWzUSKsUq/S3JLs+Vki7UpHRPWhxzOWZ0Y8
x1/u499p6GZGhLyGu+fvcA==
`protect END_PROTECTED
