`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N7cENkBs6cJWcby+WaZSjxS0YBBVVi8fMehKMdXW+KKwtp5QA37uQJEV+WSnzXaA
bNdRgFpsMV8DTaysQ5QvtJZBbME9U3z8C0UgsgrVbL0shg4mVOWeQRhd7Geovms9
8Ka7DOxOmui1uv1z+US7SNY2XrWfW+mIb2sG+Lw1rF6ENbAmDJYNaEKzp5i5k6YV
gTYpYftafUCRAfZ8Eb7kHvzpcig3xXkFL9xWgbw9qaARQUNHDXn+3oSnAd2FJErR
yvGJoBSPZPs+Yrha6iAHal+Qw4ktUiTO37QwuzfU2t4VUeyYSpyfUMcGrxtsgupC
dwqb/nG/lsJK5DeQB2PKeKr/uQD1eqycwPS1o3RN4JRqvFHC56gySgX82TwW631D
df2ZbDZ+ouvzSeE5VDRHPPFNnfCOkuxOrFgjAVcF9pyiEs2HQU3nfZ+d3StLIHmX
bow3B4fhklTITjtumZ0riBgOUFbxa5pYhK6fSg9dAS3oubc5FE1vblqM8zZqZwBa
mvlQafiPb+ar21m6GyHTZTeMe+lFuBvVOVMKkFGHZg9yQ2JHrtxe7u+i4EsrjiXP
gYlM15Loi2o6tfXTYrC04jRr8LF88nfFSzSCh9KsdKEpv5xsYldlW+jzyOYjZU3r
Q0hoH/9jOqKGAVAPMeno3zu/mgZCvFkYi6am9wtmQ/4=
`protect END_PROTECTED
