`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DrLOwXhZWr1pxGDDrU2kQSAcd3VrAO4zTxRJTIzXqtQPFN4MeauMlG8/DnlifNnM
mH7vSIcKOLGenpJyHHHggz2m4FdnHaqdDsPNInIRK75gL87Sds9EiQwvZ5QKbouV
5PAhMFe/EIFbs1mBiStl9u4UcQeAMJ9rxCZlM/Gi2/vqrAsTzvnLrf7HZVx5lqVk
rOME41N1Wm8BHEJGtnpG8Wada+Nhk1vzRpgaJC0k69EsCHYPgAGypvUCqshY2QXn
zgjIcpVJN+HgV5nBs/Rr+CnQxLBzK8UbKgAAuL0tg5NK0BbYntrHgkbTzqXApPSN
JwBxaYhoSd3sTaxSzsUnPxSLbE5rS1mRpveC6wsLo3me78v0JK+KOU6F2+krg8TU
lLn4npyv5No2yMoHaLtg9CWe2Yzf4aeB9e4b9ACdpHGvzD7BoYSziEsGcJOdoVqx
ysRSpyXJQZFnUxckZV9JmmiMk8lpSrMki2SgP032rDNpHnf233nG4aZRh3TXqJcr
c0XwwS1cH+mJ5VhZGBxVcdVy8eqsCjrrmDWkAOqcUZAsbeWkrbB6Fix8eW+MjMd/
7zXKy71j+1GzXYh5T1MfUVy4Wr5oymh6aeHETQIOSgTPB/QM6H/J9vJzHOJjJOLe
aXO0UuQqHBYRxwLeRS6rPhcfgd27k2qIdCDjt2ehfDTXnIS7wKNW2knifr4L9Z2Z
FFT4OPOZ1d8jKe+/TD9dCUJsnbCTvwOGJGzZ/czXMtoWG6Jpi5/VFIs+Hr5+ClU1
QEjD1SJLkwlZenjMPQs5vp/KsLDbjxtw4KKVWX41eUJkKi1AKCeKaI2EdHymkTGw
x/Ky5EYO+y3clHJAG0p8TjGxHOPsm/C5dX/hkCU1H/2hpvfYCBIoTQjRuhNv0EA+
ZS7jVuDd2GQheNme+zPNEzoXdyIM8FFwkSt14Ktwth+oHPftyEfirDRv9VUXIQ3Y
fo9cwy62YrREc5jgmXTX3+JxarJbRFPpD0Kt3GT7FtmIb6bsU3OJ/pYEVfcGDIvj
IxXrhLDUIQcgT0eJEvpCH7s/JZFL73iPXiCK+ePriaQ481IE1DBJUY8S17y4LkMB
X0SFPSPHTAbUkz38Hxtu8k1nRv44fmBq3rQmrsZOsVvUNDcrvVcM49JM7FM9IuxU
amzBsOlqJgHWQiAu+EMwQwo1JuVY03GdPzlSGIGek0FxuhGYuHiPkESlMvPWt2iy
5eW5oZb+bZ/dWZKWvJeEa5dzg0ckHwzNkClKo6rDS+upx8hp2h1l6/fhVibFzxAb
/8rJ/HeOyHwvEtr+obRm0BHCl4z8sJspd8XprfFTibxd53YHb6JvSGfM4zUMn/Pg
GLqCuuuc+1KpoQ7rWr6Ve/Hry/lyCjJ/XnlNXFkLdQhofhag8NvI5E9/2Jaa65hj
3zBKBNF0o0LqxdD/RNlA7MpfdvZtBQ+Rv7myJHGKSjfIzBumIa9omhWbHgYygDfS
4FPVeoUb8E7IQMtMpu8v3wr/9pAt89lZn4kj7iQUm7A+c9DwpbmIlGQ7w/gmFGkV
OYN4GAYWU8YgrXRrZ/TQVOvFzJpzZZq+ecPcDJAclZPPzM2hbIweeL8K8nElnm6g
vU5QavoMf0fJzuwoz0FHJUrPCHMe8ggKBPGPuBhHQrBqKZTD7yjBDkBgvdmO/epg
i7NiQ/VQex4Mu0/Bk4xUH5oVBKiqQjCgekQSR3jZ1S0yS5dDwx3a5wQOimTpIOzl
7t9aAlP2slSfbA4zJFxcVsLRxnk2tI0hg4CeWXtK6ORI0rZDFSeI4mgjOVtKoiU0
iV+fpWna5ouHX4rFineSAE19xQ49mJIuTFAEY+Slfvrrr+sCXOTmxrxqFz5QHsRG
1e7yqR2j57ylCY//RqVYyA==
`protect END_PROTECTED
