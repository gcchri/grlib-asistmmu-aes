`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
19s+2xFBNj72Q6t4e0O1xJ3W61qyAuwLQoYVPHal6Dw7mJD+nLhn9uf28G64NScx
YJpp/oB7rbslo+cqyP6nfY6nTz8AbfgITR9Rvq1UBdlQbYvtqem/w1ysQppp8mT1
3aoDB4UGtD5vrX4d/PbeOYXSgwE3tzVfZpobLgyUjdiODEeK0VmpiL+kpXDPRC/p
LahVvbFjnFEo0EFn5ake2HWRuHRWiTSum9w4vcMpxk+ThkZdko9G0jc6RKjNNjQV
yQb6btHIjlNdbm7PHf6A+afiHZ58cZjdmeG+um+qQL3qWwgXCsZXHwYoYwWw3Vat
qfd+qf9pZqj3GeMohhIs2C5H039nTZdxwRtpEyY1H+aLkRGyVzH4TEOn4+hU4+Mq
7Pus77eNnuU4Ax+ExWJ9kbS9JL8NZa7Fq4ZnKMZwxEVn4aJ8dkP2ACt3GrmjcaQd
NBayiIJ1jy4Dci7s3qtoYNL/snsJdxz0qjYGC0mLwErP5xlIjHPqR82egMSCcR45
4RLwjnf6bw1TZhEEmSnC/1oVov/DZXd2Zwoh+iCSG4Tzl7phsHCLYE6+1VItRkXU
+2LIQK9VAV/jrEehSvzHq9f+ylXL0hwPDe2DhiCItA6+/6YvXSraNt9sV/m9S8b/
ic9mBPUfKRrHYYAWxsP8X+ISinc2yFCYxH7J/LNemliUTZ/vzyMrLClBQBk6kUWk
mxDnEQto7tavkr7cF1v2wEp2JS7rTcvKIhXnv1gVxFVxxmWt0iLThaBzO18zH7rd
89z35GvBO7et1Zc34UfDRGuHYI/O84anGgfhAmK3tNEq3OYxtnHolkzI/8+vGg72
7W9MokGOyH3Rh6WRo6tC6BmHq0XDzUFHMgkzp9zKvhZMMgpVgPq278k94Kdb+q4i
Gf2hMbliUNucsxJBNBuf1oFZkG/FmMSLdfbGviDfIi65BEHMdAmkz2SbsBezBCm3
`protect END_PROTECTED
