`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kkotM6WyFnf/3ZdX4TToQlQ4yP4sBJDpZZa1GMKFpK2LdAlaWyIZl21g8Xc1U/Oz
4CDiMbis3pFVK7rFeUNygaF43H3sPmP+L3qUJkmRfCF5W7i7plkYYc3AvHQJihBB
3OqgBD7ccnVWrYVhkcyjwZdryl1kFGSlGiguHmIlcNsiyr04kzgAhOfW8wcuE3Ee
R1jugHqFINjXV8FULYrxN4qw13+DY53JwN7w3eEvdBBVXRE6lGnY0RZu6Lvd/JT7
aJibN+T7BEp8nOJXJxJX1S5aRbsdmgjhfvpVVLZI2CRyXP2m/2rSFX0p3CnfNcBg
FWSAkylhTbQyZpsZHuKwn23hBqSQLizbc3gjjVMUAQ91vfY6y6WucFWBePbwKDTb
vh6Y6sNQJd0CDMx7nN9e1xWwi83US+e6wpOmVrTUmIwwk8u7pAllGeBkBIovYKDi
1dR6eulQySuQdDLAiwTaV0EMiYVgb28/M1UYAN+WefIOKV4eO18vpsqOM0cOa+oy
JHasqh/TLtKuo97wfhbSP4L19wFsxbYybOpaOYV2eaJ0HEFWSxGGnv6X7G9ydmIF
+CapXV6vQmQz3KxkV0dNdOra2iaYbrzCwvUX+SAEZPSjnnwBJzNY4PEvwCM3vH8d
XHB3a3pxJvn80Lox+NPwxXCT47CNHLph6qs+1yuvyGij5ikVHGqWfrDfourPgBcH
fn6n9zqJvuvkbigGhzmMndN+vccr5tdnUFNbXwG59PtYs5TTGI4NkWYwiXVOYS2v
dCYfEobmHd8LDppB4359+A==
`protect END_PROTECTED
