`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5urjwjbndDVbZr99ECnzQV1mbDdqNachiBs8lOx0RkKbKqE5FDDcqTrT+1qxj/Q+
lsr/pfASOzzi30uzh4avZloEoNaV/al59vlfY/W32gqrw8+64ZlY1cjNLM1sGcjn
cHAc6b7Cakc8G9/VKgzoCnspj9tHkk2jllnaX5wuakfEJCLWeZApeTrvu2dM2Wt3
pE+RQMdYGKckUOK+JW1fTTvMI9M5zTtAgXZ6Kmmj1kDG8f4ePNHc23P3T4243HaX
YXOARkqxgDu2CKyFpOs3WVDqGi62FB8rApu/GoSA0HIbVBwSpTTIBedKCiMlFEjf
Tcj7L7XSSUrnM++szB322XGM9z59TY8l0Q00T83Ye7zRyVL/1DQ0G/OiweLeWAFG
LzulYDn9bWhXVyE0jveOtFNz8JVervoHvlS3QD513si6QGtd4xMwOZAzGwFIfEp7
`protect END_PROTECTED
