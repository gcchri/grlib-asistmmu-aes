`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PhtzlE0t9NNZqgcDmeTCcK+8UUIwNDKMyD3GaQOR8Xok+uRBRq3jbzf0lWsdAh8j
Cd+yf4Yg24vyDsOzh5RL0nJC+EEbySk6r70+WyOnKAGHmMczJ0D7WXhEJ+k3u4PO
j8sAUdzIodvOk3wYV8Q2CTYOr7qTkmYOvAYwQ67wiW6QtJ3samRt/pDdGnBTXt7O
YjXUs9XfH7sMx/ZlkKD7kUqnw6TmZGyM5OOBhDhc9cnmE4qveX0PMQ5WmGlWsKeP
0sGgEadlfJbxf9qfJXt1IQ==
`protect END_PROTECTED
