`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mF2zjSrZhzDVqQu3oe3pxgUsTXv0t7te+geBJQisNj+YZEwPrlBCWcID0w2aMdIe
Ajdeq8Ll0rkXq9HtSMh4XCE3uroiCweEVd6s7xsUtlvNkeYFSbKtFT3IFD58s/eg
BdbekMoYbYQQ2NsQC/ABXYnItenRc2DSw17FJFmi3XSo4o5A8lITaLDd8ec6caFu
yp1mHaN/eFPT7/gO21B5Lfj6ugSVe3BU//c430vPmj8ANGxUqbY905qNgqlttyeS
NU/mchwSvZdXb709c/ok3edF3jvhii8xQ8Q6tJzHMoALBkl9ZCt6+3z+aX39Eyus
g+cnZTSlby7VinIhYxawCmp3mgYsDoSzE0x7RTTM3DVLFyEnZsOZcQ1ImLrLwHJL
vcllJ/Qvxy2By1eo8c5ndQ==
`protect END_PROTECTED
