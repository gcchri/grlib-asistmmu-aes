`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IWu3Q5nI8cwpILMLiZHEsQh4oqxxL8XBshm5xOaiZNIP0TWl0zqcbDMTPfGV9I4i
yNCOCUMRVCW8mxJ/iKHY4OP2zZYUEA8arQ6fOT0yqQEroHD2E/5t3Pw9NzlyZDTE
vSRIaQ41yYRelLo2rxgGXu7CvXTQbDnbPbKbqgdlS+O5arRObG3N79QHgCGGgSYe
rGUJZ4EnzeYjL+AeRiqsycQl8krTz2UbxfCjEhFfrgBDdzAH03XJZUWbLW4Ae1fc
kKdqfcV9N6iiI54kLGKZAEQM2dxLxGrSUQVZuUt+3G1XhFcVeNACX+cX4OlJtKQ9
KmMFDrWKoRPvZQE3L+BHWGOqlwvmRAbe2cE3inQvFuMc94rX9yDbjh5PFLYZe0Ap
qbKtMJrpRk7fy72wnu9/wIm6CdptPBFFU/f2Iw7XEB42eglKhz1jibliQCjUjL0c
YFtWR2aSszAKWKyhMBLr+e+GL7F4YClCoVjU97U8Su4N7+1MfmZiyE46MIIRp/cQ
jnFi5Jber+EIiALUFh3nXTDQl3wznP60OLPNIs8clthmP99Fu+SsC6aemxFQsQGs
9za8DpxtCsfPvtPYzS4KD0ofNV763qwpmZNhvwN5OTTCY4epXzOrQpxgV7bLUEV8
SFhLkAyX6j9azsX9X3pM4NREODeYKUPJNgYAonelVR3W3/6tNgOAigpL1/gMqAOi
V9MNo3+ktTK8wFUj94U1e5pfTIZuKHFzWBrIQMbNNAlpHpfmoiPxJY1RRT09XbjW
Wje99WUm1K4YEzrYsnegZLNY/BxIJ2Vg+SL8doxvL5o+4Ul1PSh9NxXqFjFBwAVD
7YnOswnl0EB/l8iYvfokdGKgY1WW/AaugP8enQsXrxBuD4Ghwauok+okY1v4ssh7
FfkzKO3Ly9/XO5ESFYXZY2vFQFnd4BlUoCVfaZb9xLbt2fhc3EERtZV6kMPuqYzP
cg3rJXQNTCX6UsSKwFqQkzLwms0GF7aQZKBfMw7lUhGAE2VYgP8NanisW00ekhY2
8AR4bGxgGQ7ZB/g7NPF1CZrWMcJbcpNiNkASYBdPl7lnSiw48ERUjGbBQr6dUhlJ
wyuMTtAOhCJc5TB9I+O2Aw0CvjPFSqkEakFQOV7B7hNGFRSjoEqIfRoRbe7z2mtb
jyl8hZ537MBJFsgX8gCAl4axED4vgdMotAhUYM3PunJGpbOGlFENyBFaxzIihcSp
qv6rUVM7R7iLABACf189XC7eBNEKh6jfCtMd2DGZLsRFOAheiEHeaNZtvcSLwg9T
MTzxaQeM/Xl2/iq3qKHTiWug3OUcP2oUX0zIrj+ENT4oYt6a4P8nmQV+Odc/5uhj
eIb60FHNSlAMpV3YSvtF8Nn7TOFch783YhJ9amANQ7NfJpmrfBhcmrrhgJRs3OQ6
ZO8n++5vyGPrtNpKmUzwiotTEdVObmFt7YfJ57OPxGo2JQ4/ciyG32i4AGGgKgKT
yg3tZbS7lS46U842U0d/Nnw/vpjph4EPGdpxNBbFqj0qEzm0HrpsRrkLF/S2BMJd
yZTNf6AtpLaU4SqUVqkj+CTuvFhVz8VEnmRVO3tFlyILmYTtCkbmSbI9lNI+VJJ4
1DTErvN/mDKXIWxlWzErqPyOHqeZmNdJ5bQ2xUna5rEnXQwICqCD+HTp8yCHccqZ
QmM7suW4CFrqFCH3NPsMLphLCUBVK1EtLIw6EFVjBjp0gSO60FppvCTE6G4KVtta
NTbP2wG1g0YBFJuor20rCNoVqGw+FiKhgjZOkRBGjQA+M2J0qdnhNO3WjfU/W0s/
NTBumvDpi119r/b1R5oNB20nRlWEokCMQwGsCa0kJIHTb83DDVelRSkafn5LMgbd
8phY0VBmxEuvZwk9GCkVUH0wkz4fXTd0xoHlRnYX1b6AG/wEBU6+ppn0TK/n+PQI
r/z37wZi0465CclG58CFRoddzSpR+JfBb74XUzpGCz6jnXyba4Mg3YoprOi8quDA
kxeYndvJLHJP1PYsSDKVqj7N5Kmvf7VyEddLQZHXS30mtMoC66wVIVZ90D2NXkyO
`protect END_PROTECTED
