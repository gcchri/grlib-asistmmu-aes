`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CbHaRHEIlF1ollHdOvvTDzk2UdJ0LAgytTG0X+bXCgLlqKZo3/xPpNM3Q+lRWckV
nZQEYPrXkrXonn1jeXGmqRRYNbtIXk0HSXG3FlWt2Dh0zLvcbgCEXrXhsoswl1hG
PCCRpyeGpt69LYczG0M3Rp6aPuse7qmGLCN6FnnvXH9IO9HhfwugRRT++SUNBFZV
9nAK6d3XK14NRtetuA01o1y8OHM77Vqg0OTIzX9blN4/x21lEONo4yAaA2QsgoMi
jThkXHZwV46rpsiPDdpbpQ==
`protect END_PROTECTED
