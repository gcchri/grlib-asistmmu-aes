`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CMsoJMuGecNWR682vEit0RMhumiPDf+EeVFt6vkTvUKP57Iom9ZteDygnutIXHca
q82edhIpWT1DuArqusQfnUZprr16Bd6ygjVpjZXLpSaQCiq/sFFKNvvsIuj5lNip
ZcnUDjkjs41C6xaw9EmuFdtYsakrf2yNiC36VfRVM5nYwdNEuH401MSirBkaMQ70
D6J/nghgainhni1MunFCLXaDptRSlUYXpHVRdzye8yE9PtXZJ366iYgTAioVk/Rp
v64Ju0gv0EJin86hSulYx91XTa5m2SeW9kcKo4j754QH1il7+eSxUBef0lAhDuZX
q9b6jyuwADsz/OUero52O+4BdYBuvnONUXonoPp1ykm1iJfepaKFAQLkvXPhtg4m
Iq+4mVWIlZGzt4UOD836IK8YRy3TZmppddD0GfcQKNiaGZPmnu5+OWlg9RxMqd+8
pj5Vogvy7nqgi+T4/7Sku819iVpBbiSnxjKV48wtfwYZH8TagFhUUNU1BZmDnPQt
0vcads+WY2Ar3yxLNNaGBLS3tdulF12UsHDEOuKJGTqZZzzmBdQ0qIRFVKhFoHJy
ina37yvGDJ7PXF9I8oDAZ37JcVrB+BiZIWQuJbCvMfPg4CmpU27ORlBRPuwPYKHI
VyWyPiD5Aq3FY9nPXydHT3XhFjBRhsa60uQ7iJPFZWjMziCnd+3tyO5V8h9Z5vEK
6DhJfztO5rOR0uQj88eOAvGfXQ9ulUL/2etDpDuSRe0qTIEX5m0s+MbcxFcT8MY7
NHEvF3qqUP1/pOH+zKlCzVPkdc+/2oLReelE7/Sf2UX/S8Sefl5rzw/YICyfsFfR
+gcSVMctx0W/xkyPu5QwHjXN08vMjawmt1zt54JUSWeFKl2x2n0mEsBDa48TT0Xb
ITgSi6DSFXSy5nQu07iBFp0XKH5GDYENV62kU/yWzNIgnc1X/eit9MKAMtU2eOO1
IS5qTmK3C++qyskPddhBTwafmEAwXAA3JzSisAUG9TB84VXWQI/JvYq0EitW1DoB
EZ02j0+ATODWrnA0WViR9yJioIkblrN//TWvK40addi3coquyAOqX5sDNdsAQesf
`protect END_PROTECTED
