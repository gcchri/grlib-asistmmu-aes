`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6FzueRCy/aYK16B97mj8lEo5u3sJ6xbUrgaQIcNMbnWn+BkkbxfQ+LW45MKpg5/7
utBRkwJOyxELaf54x4qOKU465XQuKkBRuTjsMDrptoLviaAOibLAFFGv5nn0/+me
5b7gb3wuJ5gMsoq/y0hyhf3luT8lGXz1vQBe5gtzXmsNklUEXs+0IY2Kow63wu5r
shaUEk1dEIJZQdIx8bzHB/oOpQn9bBcaceuFmYmpPzqD9L2EEJw0mFuyYMmN1X9N
tu1ceP48r1Aqm7GjN/NkIQ==
`protect END_PROTECTED
