`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P2EMF1D70TKs1aG7LDGpeobsbuBBbN5ShLljxfoPln3RG1bp1dh/L4iinw6TW1lP
vBiEVC6g3nzuKE9Rz9Glc40WTNgc5IsQq+EIyRlCBbfpLNEW0Nd9li7THlXsT1VG
6Id0Zl01A64aye3hpaoFTpWMMVZdao7DTUCDFRQcDDT6zV4hdO8jrNed40DSZ+Du
i4Wsr/3cx1OBzE8vD2peqq9Gck3YgiSIqtkhfxPrj8QVDW4JZGwiNOSJP7NsUHwR
EIcO93jLf2wTEDyVSW2M7CkZPOu/sEza0m3dHc7XTq5jq01AYIkeVuAU1/SKCg9M
NRSz/BVX5ObjGStF/F8BR4aGP+5LdBTa8GR6vwxntsyNNYHXiz+6gGH3LPqgfQv9
NoexHMh3Cm3/D5ispakaootH9cjHEKYdksPDWL6qYuDy5ORS1MIkeZTy1ZlX4Vnq
WMAZUAFmVeq4170QEJ3PQapoa65u840UCNQyeqxZwNSOn3qsOtBV0u49VpN2Khx6
`protect END_PROTECTED
