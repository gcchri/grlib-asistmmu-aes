`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a3izkjl5d8YXmYgCJQGgy8Kmpq1bCyZ14+3/P1RmiqdS4OD7Kt2EA1xdA6rdrpUr
IfVuWTW7/iKFbV2z97i4x9jXSclfNgoK0XYPtrOIB6U+mciibbK3Fgt40cA4Gh1G
lNbWGigQ0+4EnaP0f+SxVENowY3Npxow5G0mbkUcu1yE9emdT/khQIdNlz52zlzj
oir8+kqHpEUAOPidpJOCcYXZmes+6VxKNlywBHykLTd74JgDT8GNSv7QLFs7rd5D
DqdOMnK2g6vU2LDmKPk4/DzoZB8lpJF+m9EEvZKYqS4F2JrP06dHE5C6TQeOy4Zo
ja+80HeBzP5/PlI3gXBTJ1DlP6DgWzMJiYflm9mfl+LXo7j+G38LGf2wL7q7IxXC
`protect END_PROTECTED
