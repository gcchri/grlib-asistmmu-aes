`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kjnd6B1FeLmPEzyVAzRAhFQfLmPkssKLuG8H2bSniejQSAlkiOmLVNJA1vk2EOjI
qBr1wHbvFhyKyPOQy8Cs58O+bqVPyhvC510GeQc+n2SQs9Nbl6YU6ybXFAPj7iKw
pucN7uSO6K/h/ueXQg3lLQlhdzOYngS+f0cv+rIqNSmI4EAScVIjP2a98Edxz1j/
H/k1X/9efhzqZuyQjRicv1pvFB06yjdXzbxS84HmkBtdYDmJQWJGxfUGSVCssLIl
Vz7ETcsbd24oaqnD697rNjeSfOuYTPXOwpgC8BG5n0E=
`protect END_PROTECTED
