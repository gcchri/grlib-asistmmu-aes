`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lIYmpM6/qx4Xu5zqlaByH6baNQFGzOFyo6e1SZ8U5DEN3lfZu9BS+z5byuARt+w9
1T9Q7Ne6fwuO9d9ulUo7CsRYJCNvny0SQfhm49mfDhOzdstpw9axq/E+JhhMxp/p
DBHmIQ1uQyqaP+JhrHkREmfoDE7aOhAySgTPjKh/wBztgK8odQoUQ2NNcYN7+qv7
d63GtW/TPCOIf6QVOjKtAhk3O6qwIXv/6uCG/SgpOWTVUfqWcA0LKgnHCDGimAi0
tqPNtrX/Dt7Nqd7ESzc7tQxdm/cEpVtQAWN3LFc5vFh+nuiIHHVKjPArbB5xylsw
r7O9q+OdSIWin0f1ObMQdi99nYtj+ef4Y58dwf2Xj+uVXg9Sc5dH96eo2s6ozJ6M
qDkzQrBOVx4K3YzpBQnQJw/tL7PIPbVL3wk97r4OUKsTkjBpvJDucNk/BEp7I7gc
CQR24vpIvM/SCaF5JyEjmxTEGf4vy1xRvf7y2ELx5nKf0hUu/Rap0U2gc+k/tnli
g11/NdbzccuYdjn2owesPbjea9VarGNNbhTCZe2+VlzOyRUWn8WY7M/dccXhw6QJ
`protect END_PROTECTED
