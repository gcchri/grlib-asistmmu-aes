`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IaK1VkSBDK98xNZ+XDCI1sUc0Low4F8LBPGpcBY1OFLXkLJoDXXbJnbEweJSeQ6z
zDqbX7nodiaYsmAhUryFOobH8J7otF3ZqI73UYqUhS39axpfp7lOEAxtj0IYrsnK
6uAx9FK7zxB6Yk5biq0h4bUZ2KaTNKLcG2s4a0h4CsNo/Cx8azMvQs9mmusMQOnz
cJiaipIbl5G1vkBTmKUCwmawR8WMBqD4vrrttVA/00YMzV4n+9m8iQ+WxP1G5IHc
PWkG5yVSKEx3yOcvzUIj6k7RZLGrMIt+1RYQsB5IgaMnplZ1b2+k47TX8T93zu9w
0Jr57k/W5UhFUIEbLGo/8kLuzDAwWQGGLDr0Wk+biaLoZtA4kWRA3g1y8aLA32ey
d7apEv4tXaXvjN42zcdYSJcgfxZ1UxDf9X8VJovBkUGUeRVloFY5S7S43qLt311+
NkyxW849xhdY9Q7qFnvOBVcKhKlucR79Nu0+49IqKypKJuR58nNZU9ehc0sNSkCA
5qX4KcdqsAAYrxWatfWS1WtP5vltkSPjdn4kzxPRFmX+JXLulxRx2m55As0/j5yc
6v2wD+f1yHJxDTTh9AL0NzZGH5mSuEAy+c3JJoeB2Nhq8MHaLebxzf1Epci/22Ct
RZKztQUge8ucaM0PlSmdlUiXfZvuKZs0jk50+MvuLw5TpGDMMxtP1B97ehQpVBwP
K+bjEO0+1qTXNO7mz040GRZKxIArCxNY5i9Ya+FlYYvjhCBkq0yHqjPbb+AD0wJt
l2iyMmlisrdyiacOvPN8tgH/UVZVGQ4w/1EiPL8vvdhQ7yVbFEuiLNdO7UIT86ru
MTrpbvHXpVOgiwSlhK6zD5ymeg9ayWuj5v2Kdv4uFWKUsqvEHNLaCD3mN3tj0NVM
M6oVwVf/m/cqHY/opQ2KGZVx0N+i7jMh7hBKqu4iUcadLPs7naibam4Ul0ZnuraZ
E6t06peRCTqadWNnbI9CFPPgW2FsYHBuHA5FkbbENsROg8NOKcPEb8zfUPxFW2NK
/s6/z22mN2Jkif2bP3iO3j5pqEVvdEj0HQfuokH61gXKfs4PrVWEEZGIoeS202lW
bsaAeDieTKbpn7JjmIQA9DSb/oqc5hUAZqCCTBdPV9A1WFe2TakEA1iJbkaxrA69
ctrL3uakQzqYHYbTpqnk4ClUUvzZGxbo6CmTYlBCkVGrgzl6DG9qkX/RbJBbfcHf
pvz8sjCgJPUdAnHL04WuabBP5ZB4ib1GCPy5oer2dyvOGgVBusyveLjBH1CkY8ik
Jad0BvcB1wPwKV9KagoZMtwKk4uKAn6k8PatOPVcYPHt4sriKzbnE4PM4Qqw0T26
t2fGkVVeFu4gRD7SFNSfAuLLyufjV1u9Qk4piQ/HojkTppuATH7xnzKt62g0fyFn
9C8BnqXiGmflDt41yOSxQ5X8iqMQIIy6EPUlGmLWIFGKyKNgMtWGVM4H+Z/I23z+
WhLovTU4H+HAB8IIMqaE7DI6B1NHgYE5i47qYHoyaFLJiQ9j9GayDJ8yHVfWva/H
024Zbk1xerJh2CBcMga/dlhfpatwbJ1SZLVuCdGBHrL+F65HFqlep2n3WbmaVa66
Eg3EdYPDiAUGS09KOHDUb8IjnKa92bKl2TWizs3LqREL/mPsYOi+RcZxS5rN09mU
AECda32KBDXscPS2W9Z34G4nPeJyai8glJQWYCjpTSBMIMz7Cf38w/KE3o7JI67a
X1drR0Lpv8HevXHqJr5Y28ELtZs3mbzli9t75WlBSWW2KziG0z/7S6HYECVTymM/
cfY76Q3ZX5YGPSr+cuAb6SVn1pNHTQcwlnj1hMXaApheGoHXlhkO+QZLuyh83uIG
gFVTxEeImf1qoXrcX+GIgGodkyoMa9M22JZqHeYuVO4SQWPHuMe4dzSXDfRwWWpg
rp1zAUSfbJmrKXNqD6hDwacdSAjWE4t8AyIPmLrfte93i22C4Pj1UQMCct7SM+l8
40hrqoGQagbqbKQdLyp3m3jPbkEUZ3Jl5jmEh6Rsad3+lBw1unOkKkRNI6CbJSjA
GLwXetUTSYhCqvzLPiJ85QcSHhWvNfpdhNGS1NFHy7c6dfMxD/uoecsaWlF8XemQ
bvM6hnuubpnfe5FuIgUwbA==
`protect END_PROTECTED
