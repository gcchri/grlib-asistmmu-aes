`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KmGNCmRPtDnilYE0vQyzMXp8cCo2jF9uqPHmP99AGT7jUn7oUi9QIf7zP4MHWws+
2MwLbY/NZ5wbp7F5YilXDnZPf3WRyNINMK7HqJ5fD2J0Spy7czo5oxfxJEe5QB2s
SLz4RfPwnt/22Sc7jhvg+TVa6VDLvR+onwWiwUnst6fNzlkUYZD1/YIGrH38NxZd
Oo6jfks0BhLIvc9kQiOSS9HDNhZWf1h8o1WVqBXdP2KoWczSterX8c7P9YjTPZJ2
YjOsafG94+EjweP42KopwBISevSB1VSyp2BQAGyietejtgVStGLk2/KaGwT1ZTdq
CzgA4GTsUq4N2r7iRfFXjTyoXhvqcTtneIQcyFh2FzIAj4nYoruEAdw2QD/cEKS5
6xf6ezhod0V90NGfCWe/aD+QfUdXCweOWpKEu+bBj/CBxIUbRuhGerfwWC1+Puh5
6/kn3jfGnXvmG+mQuxeotP1da1oI8/l1ESXDInxTHT4=
`protect END_PROTECTED
