`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hv3K1ePCJ2jCsqPfUhOHKFvy0SZ8tvEl8lU3w2pNhK4NzEq6jc+R3IFE9Prxv7dN
w3SQFrBPWjo7F/af3mva9HHxvzfk6o/ij/CjvJDB6LtByCX+7TK1dZ8rL7ucT2tv
1FLjHl/SJz4KnORDs/M+TQLjwl19jo5HIHF6NGEXwONtbUlkFm+WqDzrHFX8LIv0
/pQNcEVPoMPZuqnnA9D9HRYjh8iwCTMTpE07MXJMNbJWhBsrWdDD5tY9VhyVfeRR
1fV4Zf1H9basH9lev8wHQdBeqXH9kDCky/0AoobQP+OiFxjtKjtXZmXp+NHGkcji
UvVWRGdFRYNNcHTfnUjbzo6xeja9y8Hj3u0xRvKjPq6VKH1otC8cttXAIfiFBsKY
jF+exiCOt7qKcglWGRKPwiNa2OCq9IoSGuKlb/24TmtIgAMVm01a9MTWmTnFv01I
m3iZkv1k1a+qf/tJCGcW8A==
`protect END_PROTECTED
