`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Njy+u1r7b/PpL4wnsvN9PIHN7TXSza/2QH9XMh6YVKFaaiw88EZ3U9ERsCL/fOq4
IRnqJ6I4ppUQPimzj5DhDqg241MFb+KpOs0eCbIdQdevQe0dH7ekK5Tp/5aVNcTN
ZuXX05HxPCq+OdmOWwUXLb5dlSn9Zaw+3lybI326dduDnvrFyQcFQGM2dKuWhfPp
kmKfnRV+39Z64mdcpcIhN7I7N1G6+O690Q55f4adFOlxqI8YeLQYXBUWZ9ccBcy+
OkyIk0pN8iFaMU1XqJTF1LI+AV14UUNeWtY5Y/hUzcaMN+4iCtQyG8x6/Ya1qNFc
orhtI/btDQJNQjr2aaL3YNkNcROxLf3x1hUowHxIAWLKloHENXz0tb7gnxm5lgDX
kIjeKtL6t3L7z7oah2UwZ683xwwbfX3QZpaoWJ4J4ArYhBebrOBXKdXJEUtujxsW
9PlG1QQxvrW3LenY9tCbmjBjoEiMVCZ8SwZgwWrnSyo=
`protect END_PROTECTED
