`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ZNSF+8i66vDGZDglgWUo8TPbXKi15XA30M/JkpAE+YL8oVKLCathO0YnPSJ3yc7
ccc6xnyyhZS6hmW5qHl6gdEgsXAQzY8i+CapRlzTIeaUvZszjb25ZgWRCQGAUipS
HJYg22R1BkMIwxmAQLyJr25DpVtKDGEfpEkL11u90CufpxrCpYCLehR4EAAknIg3
WM3UrwBOA9HoGgANBjnbJy939Yk5Wso3LlBqlV2TV534B9XeQu4pRzJRq66W8U6v
4PQSYUXBX7ahks4w4XjRFIHYyc/QbMWbGd9Atzmwew7WWOmy8z+Er4YqPN8jB3l5
yNbYGMcG3/oPgn/pGWsW6L2FQDvJu4b0mJguOXfb5zlwHT+NuiL8fEm45NvW5C0G
24m2XB73ub1P7W/HyyPD/9vTDDYGxQmxUBKRiml4+YdbxTpeHHio18/BYd6CjPI2
/mfy7swnvGy5Vwz37p3/5HKcdsjJLEXpbQnAZKrm+8IZmOT7pXOpbcMXYfQ4NFX0
yQo8h4cy6qBq3I7uayotfAP39ckWPj+oLzyGDBeEy9z0TXYJVsHc3lu3Wat4qyqb
QRYBBA0rRf6jjmBvs7nDNvnXT/K5++n0XmASsU7/hD+OEWeDM/0mHNsEqEKGgnz5
lXdNmdJC0dM4jElRY2Gvz+hTN1Cd75I5hU/09TWpXCguslEngOiEMCV72kb0DSuS
hl3rSeKL7XuFYEddalKs/QuK97hizGEj7Jd7vzNgrAF+983MWOKXDMjdGHa5tgPW
1uAssoTunkWDzcpYYqS0fAPp/R2kdlxOHDSITDaS6+14aU1CPSzK3cWJWcrBDE4E
fpdtftK1YF0kJoj/x1fv6cxYG9ajWb90kFHTY/tq7tMWToXHMCf7eH6JSRQF8aMb
B8i/OWMPE1cuWFAL0Bu8V6losua8L/xbaw84BOGF4kYrMF58tVZRrqm0Q7bH+jn/
vaQ8pxFRs2cnBno3hycMySLCNVIjjl2elrJ6CWDx9csRORkSylJT6p4do1RcmYwt
`protect END_PROTECTED
