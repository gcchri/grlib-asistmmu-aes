`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vc2A8F+bfkSEr52RVplujPxR9YETf1vVzLlJq1OFVsbQqCjBbW1XDqzs94LXLJtH
tHhqVYrmYoAQnS/Xjj0mMXWrf/jHmz34Qu612qP2S3MWOMPUvGtCh6g5lJQKCxT7
PDIBDhig6BPwXwGrBdKdajicFf4AfrQ4kbUVz8ZkjiyJNdmC8aylnL05J5H1YkyR
m+1WrmBdRAyddvTmbLMTEGGbKoYcROAEs5/vtDGhLLW9TbXxR3bnYKwZhvW/SIBE
21j+poFsQvxaMH3LPW2sBXd5u6OTj4ApvpSSXpnHyin3iUOrDipWJhKVU8I0Z8jA
yFtTJm3F430pcG59BmS3bQCetUEITOl+9w+zPEupvnqG54rarT/SNo285m5O1UHd
64Y0yFS0gx+1gdNifPgkEZOyC6CEnujpuze3HMC0RinnQpwJVH7cjkmYsgzvBkCm
`protect END_PROTECTED
