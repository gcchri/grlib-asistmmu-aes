`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SblkM6RfeZuTc3PzkQdYNmwhpi/WwORSG6ttJPzG9cghLWYXncW66cXQefYM4hMn
qCs85bSIGfTmC68nFOEitIBmRMShWfrBce8PSKeDjQXOlEhegpuPK0lBkcKK+VSo
PsPt32nG50JFeMjTZv1pjOF2ulfB3Xayww9WEGXM/DNrQrbuGqQzy/HODc3hrFKK
Rt4INSvu3tuKFM2ZR7NU8LiVqqoiBLQBpaOMRIcW0TL90D2ZoLGjDCpsnEZVSW4z
/EMONwhKpV2p0/RhflQjXw==
`protect END_PROTECTED
