`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xkohr/DRlMghz30+fe9DM0K5GRNEhBv7BkwkjqD8yTIBvtgsIzSBXl0CRTss52Ap
DFZRqFYOqmZ+x8iDzHthrtIvGcqlGG8fbsNWuPuqye16MlNxXYxeeTr514xSgo1i
ArdoPinv2tZB9wVNR65CYgopfaCleerE1OmybN4uQujM1ZRqBY7lkKeOFKwFl5ZJ
oJXbK2HM7oTmyeM5NlO/N1nrWWAx1CmdoonuHhQAXlKuXCe1fuC9fPxmPsWR8qwR
RnHTMT6Un1iW9zTubO8cscRUYQcYkcndBG30PjSejwH58A1AHXmr+HB8J7LhXJ3h
2D/DsuHOtugZSPRbq59VBYpfFskpwQyZMbfKxkmwVLqRr24KXoXDKaRCXIbnHnez
l5i+yqghQ8O8qldxpU8qKTY5cy5SxWqAKEa4v4QePFqOsuBsIPFZF7cQaeF/iOHd
12zCWY2wgHJLAg+w+PpkihpxTFT8nwH0rPSD0LmjmZPv6SUMzeiFuO7v3jAYsWsu
q/25nP5hK8zLRTue8AI2+70W54fzzZ1oKhxlCB0wCD/RrkZ7LwoSq4xzG2BpiJRG
Z8ICQrVSbhiZ0LoZzaVLrHYfbcGtNoxON7UuE8HVP7HIXAcOU7hgBuQUwGXft3q9
z3O47Cl7V44yFsfipgqbdQ==
`protect END_PROTECTED
