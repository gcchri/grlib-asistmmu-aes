`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fKFAsIeyn5brZ/71ryK9+ASU6sCfIbE5EESk6h6CinfBp4tFvOqcwpRkkgD+CDKw
sBdBY5tT4xx7KwBzAP2cF2WpudMAMrDArWIojZ7gHNyWDqQcj243rPlnOtRrWiGC
whWacPCyx3PQ5ohLFCehHCixaidMFTDStnIRUG8uOg7zWYocYh7pGF6rQ7ZyMt+7
rTnEEL2SvrrZap8NdyzEWf2UwQMSNlbbS6uPVzTiyLtIwdJk0TrRLjpPworArWCI
ydVslSt5hEb76Lo/oiFHDsAv+PaDSKuJ7xPw4wAtuUu/Hff3YOGfnJNo7O86493V
OmQlvkUJIeboOOn8V88DHLC5zHs5ZzLJoYa8eblrGzkVFAsEpZ1hCxglx90OrLZG
lzMNmvFpeo68A1+9nCU3TPwFSe5F/c3w4kG0P9aNOjWr9KIFLWPqpyb669TipAZr
OkC/A1pTPgdNMYbWVJCJwCB11cIGAwjCP/j3bpVtcfcwVmftfZF6poJ6Iq8FWJZ2
ZcVRu/jW5K8beWCl02myUVhoOMSswIoz3cOSuccUNLnclJFXce5ghobbCG4F3l8p
rYmC6vp/YfUdg9NsigPx9k2Vr/lt0te6eQwyARskrAr4SNxoeq322uq2ZY09cEbP
IR35QZgd2aHTnsrEKUNfNfgY0mYqurzqJ4i7Wjvpet7kF4adch6rWIiYv1cTvad/
knp3qib4RaGN+OF5e3lmDunuc4q4ZzqQOu1HeqLhwC3RhD/0MyKU9On+Qu35Pbc7
nP+WnHMWMvypt6j+Ob3di14FLyFDI0tknT9bq6dYW2xHUSAkeJB3ThKu6QUykPnn
vAmU9CsfYzwtHILEZkiYQqBAIDwCwu/oxxJZCyV7CSfFmOIVHZBN0EPhgRg8Y105
bKo2E/G5b7AMbL5KhQHzvX5dlHvlbz+t7fh1lIXoQjrd38p0T06fdTISAQ4gC8Xk
uimo2TIoTkVrcOqrWLMOpCtIwu8UG6vmMOgSgO8izTYGaoSBvXOBkrMVdUXHTLiS
qiHMrQbxoI2VNoc8Gl5/DwJDuWa/Qg8KZ5TFe8sidM80JBmqdrWLxBOqcudqyDZH
ZpUytV5n1PtjNgn5e7lqQs5ivjJTEUv3f/HDNY4dR6sY2gOAILi/mNdEvt7xoK8g
`protect END_PROTECTED
