`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
12YAH3vnGDf1ZW7//53E3mzLE8NfDRkfCTEfU92Yoszz3G6AC8UvfNiGytO/9FCa
ex8bzaCYUFruw87JJmrR3/wyx5TbtcyfF4ZqbLeBxDct4AfyNdDNMPxS3QWUe9pL
UUsffFshkbFgdcmTp9fqpMqUspggsjoIO0+BRMrvw4qcAsEys4hyYNxx+H/aT6YL
+FjrDYWUWMgLdLfgb/F9dgv6MUOmnezdZcGwfw/BbN9fyhVkiWNuL7XX9yPmEHYn
RuVXJXbULrLnohzoYzrYF3+fJMIWWqM8rctmiqmMJLNXBpoTxXBMrKcpg8ySLQbb
KuJ0Yw2rlpTpet1xx8Crm9M+kM9TysQIJrv+JyjsFk/q5C8xjHUu9WAtU9QnznI2
1+5Vg/eUEuWTs9kEeeqPMtCS0hCudOKc27DSS5e2tXaIlpuT41V/by/daUtZVjbF
VNsk8vXEeakSBUhTySNJ4rHMxnp0nWs9ZHKMHtsI970mIgIV0zVpuNqtbnZJ7SJi
zZcyL6wEQjWMl4sIsstZ5g4TyhNbIPTadI+6G7ZVh9LLG4a68RsvqaEIt/Fds+iz
UMSM++tI4SwrOIUbhVhf4UlRD9VqejC7z/9uUgEqOiLuwW5c5VTtPZoUzdO/LxYf
HR6MbGNQ40wIvkQBBDUJMOtM+P86PkPZalJo29YkG/kR22j2xs/VO60RGroo7r9S
Syg+0gHv5vmn1y0XGKH9RzjEvsVGudQHGFHl/6LVR1onWGjlB72ChcZDM12lA5u9
3NfVFDY3cVpLjr1y+UIXOw9QO2qijVAVlzVLy/CYn/kWURRXbpFpzxxIL4eWpamW
JDYYaBFxc45FsT+7X+wqxA==
`protect END_PROTECTED
