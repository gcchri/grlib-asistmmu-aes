`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t4esA1mILml1nEMneugJStNOtaEzBInCL6jjBqbUHr/h8ddBhsacnifMlSC63aAQ
MtgQ3yYRz4+swjbRcx7QrYNnlTOtYcwsZYLcGk1EGRqa97BNBkh4b4IAZBxFpnEU
ySbuCZ3pIhgBXGICwrPpH1qt8Qr7f3s0h8HGi6tKQSF4Q1PfOt8W9QClI13RiOdZ
hBR3PDiPMbVlvGSReCL0crqTl5DxyF8I8fsTWAmzOe1HtX7RIRciVSPMydOu5wT2
mIXzuzg2A3aKgWNjU2uak9mZNyRrLDwLvuGPHvDkdcymPZCijVN171YqfYLKFjFS
VVGWT8OqeNGtWPK80H0O8gfGny/bq+KX8pCNLRPwZraJvv1IsGvXiX8NNez2AOo7
w1PTIp+QMOHOSUEEj3925NxntWNFV13lX0MlTeX7UvxZOfWvodvKURlw5EYzuOls
xjscdc7ogEq+67jJZZeobK353Gx58sMCMUOtYoxPwwL2quqfXTFzokPzhgV6Sz12
LYiM6bOJf8I0Io4NcteqesYwjzpETwnEmtXIhfdbfH+1x3vGuEKIZ5AS7a3Y2CP/
`protect END_PROTECTED
