`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z0Ob1JMrYe1BsKbagm3q9UHyjDwWN3pmtlWdcdOkIdePbLySg8N8VPGp4SkQoo9N
HWdoTZA/nZpab4Z66Fdn3zGmFbCAstqFxZUmtVc3+qlSilPb64TmaP2hZ8Nc575+
Tajh3BmRbRcAQ4qbHLuhTPsvlxb8fqiuKrQXcKtirpSpH99pLIpBooSmr8/lGBEl
rt6wqiNzZn6FP/H05B3MTQ7lMt3zuZqDrvtCeJWQhSDZuJrwTGlfESCEcQooJFp9
u1FQKfAR13gZtZ4AU9ocpK0Y0kI0DqMPob16AJclJtIzL95tdM/lvfnqUNfncT3K
nRbauhMtCI4d5kK84iaGS0LdNFGMsr07VSPOr5R+JKW2k07qfEVcgU4/zaNXhQS+
XCeTOCCM5zfkHSxtxhyiSFa4RpvOhGiujCpcJNkUhc7Scb3hHLNUCNyF3fCYl4mx
HCTiNKDheRfYBxuCZp0kOA5rVjnC6ClQmmCIVmjgIgpYyveZ9ZAaF0K5GtzCWLtV
p6UY8F/nPOujG/UcH4eKhuttbkh24EEAXa7zfIchzSFA2908O4JiR+DDLDkttDye
L28stEnMs0NPbSP9Jt5ATZ0ci01s5lzo3wnkE0IzDu0tXiiTrji/uY2RdTGvz7u5
cux5oIswmUQeceO1/vmllVrAsR8PjnSrIBqAz8tEIkmGkDBGtPh55TuhhTo8N55e
GzWmsTRD/uWkTcOekkJQhMjSzsPxx4v/Hy0CThw7wVuRU/kNdUuYZ08V+YMMiiPZ
kPx6ZbDQzluWx4G2a1spsAoxnqHihM9wB9nnP6UXwYUhjqPi7Ia0wNJt93Va76CI
oxG7le/sUCRcz/AXsfM+DjuqLKYUiEwYfJBVbLU7DLfnci9biE7R9SJGUTeuucGl
VPcrUVjG5MQmKeKYG9kUxyBftvMDC7mGV1nReBn1zoTZE+suZB9fT68CL1VWPeae
78iQvG8z0d6Gsl/cOwkIwKJtCuuGeHWpdPkCDcZiPf/wXrdIRRbc9biSKUfVvCXA
OTTXSNE+YqN6BU/E4Mi1806Po0Rn8SzE6l1HnJDsOxc8eVbNPp96WMLXNBSvYXnG
b9eVGUFAwc/V4Apz97aAyl5q6mWuCj3rvvWfsmmMGn1bcF+dRtECq0bcMHFZ/6Pj
YBt65csQrSCSPKe3eJjDlQ==
`protect END_PROTECTED
