`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tlpOgsobG5G1OIhxGjsLW2gjHloIpJkLokAh/+lAJGZy+wTLLSTEMpQnYacQP4ng
/G4gGqdtmJH4fJdOLq/1KZ1KIwwJpyHbpoGKmKLjbvqdHGg1tFU0TQUEIoord87/
2/e+F0RzD1NkSBiYDskskv3+iysvidnfrNc48H/W0oT+jfZY8GumdZS5aQPlBoA/
oj1JxvsUYdkcTAbqECxJeN1n10SHa5vNQ9YMQzDBhWiJHhZV3vhL8UuWXKSzEYdK
7NSe79Gpif2IRj9E6TmuAHkqn1tfg4pzsrOlV94Lu87Eizsw9zs0OpECn1FmCjM6
J5m0zyZahN6LH05YnyQQjRIgDxSQB5mpSenBSekZChP4uYARbqh3VkHGhLHgjpk/
3LJBx9AM77xzuIHBQk/bRNd7ihirL+pK1NaCgcbs0Wfu9UFG8oZh8m/bP7cdx+Xr
C7DEA+BerUVwbCZf5aAG1Gc1tWHze2QzKD9YmVQmNjW3jH20BUsJRte4xy3VPUtX
XVQV4uvIkV4CXCIfhqRufdaL7ojOigtyAbTx8MYSMe1BaE0o4yQbfQpOpKsHp4IX
MIN9LqbBhpcUFkgoSu5RDxm8fj4Hk3xMIpxiI4Hh9BecWwPiIPQdyOqdmGW5u01O
SaucEQkl6uUmIx0+tBqfGQ==
`protect END_PROTECTED
