`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N88dgbNA4tbQwdnN76eDpfqwuXtMN+cEDUNsLMbuomTvUXZOPqQeTi85K/4jM6Da
3dCDVdhCapea21W/cFK737ymbTg4Nm4eX5r7h/PaBNfIUrw4X6y4fmMhPqcsZeqg
xMxTHo3DMu+FYjm9G8PZFgW1ozEyqx3NLAdHyYUe//aYAEK2cwbC8M1aLaSiRx+l
CveshG+N6wOmjq0rpRn8XDPssb1lMrdlZIgb/9rXqxyZ1LMH+zwXaF0t/a0+iHsr
1y8ro88PvoQcFAxal5Ke2fAdgpGniqrYLseXSKnazb3AOmDm4WmNvv1e0tanOYX0
9nLm0ujEsR39lv9oqRGOzxVJaugcyK1o0AK1Kc60IFpMIUQpvbQr2p3zR1gNP8Mc
pihrp+eiCux/Ib+CzG4DO0F6By86/gHpqwZ7w61yXZztOEXECXBilE8JgODyE6ZT
OgpbJY9+8We2xUKVb6OVYAvTqsgWFSwqkTg2cf5+3N08kOWA9vrDqNF3yx9dgBOP
vm5eKpvbkBcoecGMu8MNf7TgTYAC88G7yagsGDCGC9D0PZSURduyLuFBS+neLORp
mVpreXxt/gcLqgUgMiX/eXW8mvt7/i26ZzKjSSaUEzL0HmwWen9QD19wGaGNtyL0
jJDoNzfLPTjYEyTMYI0cfVPZPNF/wKwxkZO+B8RYHIDcmtHbN1+dbkNu/TbZJDLS
+NS6+Xz1LCkghJSJ0cuwC8o1kNnevsywautmptrGA/8ODDnQ4A8S2kQnyCOiMZjz
wn7bUZIrz3D9CGT9Yg6LJ7CfjqjMUdnmqLo7juWVAeLIty8vaHgmhayiho4D1BMy
zApzKrKHX2jaB4xEYor7icOExkkQSsEc2WKN6ewYYEGi/XatrBzckMP+XCz+a1aA
dqFGboyFPTgI4Rw7OJanxEmdwIT7RxTyCnn/iXYGgNjni/z/CD/KOYfdBPiK/L0o
xN26CvJo2wTbolGOX8ynwCCArWcJDrAyfhxPTyIKtbTeIrg1kRgos6suNc3FoLFP
hlhY1wS2ebwcT8m+UdPDtxXoqT+rXj1YNEhoEloVsYZfxyTcS2O9b5MEK1KpP0PS
SUfVltFZ2dwFjSuk8D9YyfrkwF39Mhjfd11ZZs/onrJnwiVCQrKVHnIdMlmzUEfZ
VdU7uILVFc+f+nokvI9UmW25CtJLEhDbpalAFFkj0obwRO8S8uBWbO0u9fi6zbpx
cQyWE4xTcZfRXmv3vVlnydiuxlT1klV3gR1gvNi2bdApBLWKpc/jeM+qbaJg/luQ
X4vt5dPJcCzpTlvojwtKg5fUFKnbLbBGUdDgSxFbDv8HjqB9JaLdRAhOMeaQDx8V
jUUa5c7OU6ZAA5fXeEk+e+XhqYIRR9N+gXyR6kUn7BrG2Wr/j90Ygiscg/ffG7WU
`protect END_PROTECTED
