`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E5vd1NO4PCQUTfpaW0Q7ebAwkhwpf1fr0c1b0bcR6n/zub89v4gz2FhFncncHcEU
7fytSyhHV/b2/9NgjhP5vbqv4tw3w9QgWPCSFhBkZIIEgwBcjZNI4jyRE54q/uof
aRWG9bMNaFqCNx76cZLgrRcs0Ll+SgmvsNSm/4LIHbnbwoAjeouOFHGWLOLxMMr1
7GTI+dKRy2rOpGS2WAAQcWwh4RjMvFiCIzrweBCbq9sPseX2HPIQ1EdGa4ZpNTVf
5yrJR4W80Td3W+s9neWCJChRyvHCtRLS8EpaaD/+FCCDLDRs3b8ePkjRM8Ycat0S
RIjov6GLXy/hZ9ka+v/n3j2LiOlth9th3YOka5OndrU5jKD3wZp9okEJMevsvhVO
sjvhjY+wWDivHfgJbHSs1b2YTH9WYDIvdixPlJYp5HD8IgUP7LztdWen2yDQQmMN
HkttAVilOpzlNuo7slkcvs3toaxPn4ZgJr3lpVQpJII=
`protect END_PROTECTED
