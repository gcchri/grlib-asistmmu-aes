`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bMXgVSvtLhhwVMThDpDTRScL9WXZcYIP89Uu3+tZizrUUBSukStXo7kDk69qOgO5
NibiBgKg7V35aegci8o7LzdyX+2TDNThQ8Rcuin9kCJu14B4PUlSrr1HpmJMbrMB
yMPeS33QpG5TuBeh54Q3Ps4a8PZD7M94cnfXAy4XzJYGSfDdrWioNch6HF/7Pa/s
XuLhWKArjQTephMaWX2YSu4SV7zrRAhojnr26IuYZZvC/K29w5Q/74hbPBisJ7rm
6sqI2FcfgrkGNetxgxe75ftzncJ8TzpY/Yj9NFG/hU1PDOyPC73AHwEMXrDJxhYZ
ZEsRbyOSoC9UKf6gtNOcnzr6A4222TA98kbC4nTOjkLrX64zQ6ZqxEixYS12SXyn
8URJHPrjvLLFH382uRcHe9JTBxjDhd7FC5Dwfo/ReITdwe6jykgPEHRkr3LI8cRd
GdU14IK3XebaqsmzLOJ5YrKdBSLGDCrW/fqrOg9YhnxoUuvxA2JtSZGyIAVhQHWY
zofN+vHFmmzxmnvv7TeJzuIpB0nQtg7FAOorcYgolgtbTC5Uqjhh/BOy9hOgzFJn
B+/jnq7YO027eAfUOXnJ9zQWnH7XqTRMDtjpGuzo+hSiwO/2Al84aYhGk2fg/52o
g2b41X6z+xom3H0/AL9D2We9FdikOpd3Awvh5aoKNT8ghj9nD9giZb8gUVjRuXbe
Or6czuRFcLQp37MAX+poJjIV6gSpwtlJiwQHV3SDuHgHtufKYC0whjqYRmyt3fmT
Qx0iGu8VlXqFOrdmyelCeIDBgkBAAIF4vge4qv0higYpuAmxZPUqkOfj3WHXhxdJ
x7z8gK2Ypn9IDvANr+nATblL6bIEARPBOc/8esIEzLG0VyW+KChoeddYuN+xRpIe
6xreaMyF8X8o4XT9Rk1Gj2I6Ecw4ft7EiGX/fZKP6ycymx+e/nWr6uALtYpWVSDR
8PyLfHECwCZcjnJmqY9BFK1bGA2CwYryCp/w7cidY0oK0QB7SKYzEcqaFeGlvmBp
9KOyG9l9RPC6BlCAt3c2qiU3eO4u1pd6CVl50yUC0m3hg6oa6J2OXs7fcFrJKS+P
9rdlQgGr2UAu+1ldnMOY+X9QEkZXSn5bx4RF4jW6kYCwV35eAlP/N/b09HWzd0F9
KCGdaPpbuV4NP+T5/a1u0BzTqumKeK81mnxJ+y17A7MoDBqYo8iGVq+xA4DVCdxS
aqtrJYUrUYJsRWVmuRI9qeCuZgOh40m8QLtG5molOBcjGAjaMVzPX8WwVTihv3Rg
`protect END_PROTECTED
