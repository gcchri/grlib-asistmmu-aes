`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yUOH0ZwoeegG+qOPMz42zmXOyUvW5WkfOAKyxh9w9iPElkLnRNuIUfPYxjwT+1Bx
7cOEjTVZ/2ikRGnD4falV2QsJZYvTsBTe30wfWXNEMHiXlLGT3QX3GMRaURkWT2d
7nrkCshxFGUB9newy04+JclegC/Mz066UewXiyLhPLPmZtlN64LNC08QISiqr0z1
+Vqvdx8NAXFcDzcAlT5FfSUiBV6pxw5c8WPjFgYCSGY94QTFmxfihY7WZily9/wv
clnwr1nKSZKA1WGqzdkpb3hBvjj47L478lhRf2iKlhJ3rijxR1DoGWvtv7+zH6tc
VD5RbbNMp/HaXopLbeQxfSMZN7ORrQC77/dCzAx9mX/YTy2ffFfvewGAQfkd9O+3
ja3LxqUL+oKQvpl0Q1XwP1MRB4plsXPcnxkw+G09GIsQ1Hr92hiPQiyLuJQatM0H
kB94DoXmqqlXu6dAwJsk4IDz9VKtNCJ+Lgf0eOJzLKRXd8sBFm0gopYMi3C6hOi+
kdz47F4CMHAm0O+i5Z9eLnGUab86a1Y5SuKX1j65/WtIgDn0iJZhwbtgLTKVXCQ4
Gr7/lZO3XmvN9hrZdoQv+bCnpTlLdxK0G20fLsK8stSWr+3EAN6e3iBFKiQjmzS0
OF3Blmf+dYtW3+CPH8Snrjfm0E2KZbotfLFMPLZt6NnwrUfkV5sxgJvo4qfhkCJx
UmTMCfzuK/4hHV4/MFrHJ2j030KxGemmboayIoFPP1xDNREjNSqgO1G95YK6bU30
UX6vd/HEIlts3RO5PDlgyg==
`protect END_PROTECTED
