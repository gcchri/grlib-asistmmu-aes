`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6YSUktuVaF7orTCaYCm4ZQZZF5I/AN+MYn3DXC5vtpSTLpI7OrWaVUAzsw8jru/w
Dazrx3Sy0iZ3DiQBFTRgzcL857HCzjPhumO3WMy/g86GUpoSUvF6AGeERF6YW0cE
GbbyVrU0sibVjrl0dIeb3vcOgz0Ps4mLIwpU26wnIaWSlI8SloyK2hESpo+Ft2iY
LC9tffnlDCAQYQEbyBB0t18zaXKoi+yuIVm85RzHIEW8A/PZ52A15ChXkRK8LVXY
mTGCpy+GeiRQmvOHyYePtKT391UNIS8MM0uvVozPPBGIBqWAAoOADemK0/H6sldy
huza4pgwY7MKk8rUI4om6Q==
`protect END_PROTECTED
