`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BX+OXoBGQBCk1/99i+yWk38XmEp5XSnfVOrDCXknAtq33I/IBTOgmNYe0v5iAQK5
z+MJ2SYBhkDsfEST0j/8rbvDqNbSq/6gp8aUEl3bdeu9Hj7D0HfvTMSBwM/r4lHu
kUWrVOVZysanhBtF7n/TV05WnDGRIbyNhGTaWyI9icFyKLGPxfQOYO1nWvP5G7HD
yx7QApR+1htdtVjYx5oyubqi89IcWuEiUzO+JS25/QSDA0u0VqFDckODF/txBdfQ
4GLdEnjqieSAebxOoAXstgoItmUexsfOVyK4+dk6Q+4WohtOj2xERcoTEpO5I8Au
KUlvwqMS0dsw+AH2vBuWxNofyvQCTSbXXeUhBdcT8twVzjJNEdmUgtZGy2yYzpAI
OnmPDgqK3NwRBFjwSnfdlw==
`protect END_PROTECTED
