`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V37N/524UFDlSoc0VbDApDrvi9zZkS6VJIhwm6xqLFixLQm748y87vcjpcxwF/UX
z2d+0z0WzUaIOOrg6FuLSUF3bqv5VQ0nKi1PvYyc+NXY0I1FHsVisd4Ept+B2hgQ
BiqtbmoMWYRI+hDvF0pYb8ygjelcoRizAssoHHgox5GgUcmjpdUYD0S4jfsUUiQJ
Qr/iSQ3RB3gEdgAmVBWzvSrNoYULG1jwBmHutDJh2f5k9zeHCAUVtwZgSnQSsa+s
aBIKt5ptmxbZ8LV+LE6PYnUtpmatqSwORa42llTxcVb2PTh6PBaWafGosNJTtaJv
w2aXrHh2ELkq9B8bct81E8sMLpot2Vd09rcKOPL1BFeFbpQ/PxgDDSVrHpJnn40A
gIpZ3WCHenXhGdhK01+5MQ==
`protect END_PROTECTED
