`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fEu0lWhrRWASiRbBkLkSwG/aMbCTWpc5HXof1QzvxZikJ2zViGEsXCOm3Gs8kDf8
CnsUzeNzS6Zd/v5M1ND0uU7w7ChIOopm1IL7HAmg5t2N+BJnsN7yQDFqJcPrxY+M
sXFznP4DtRJ6iGQ84g0iApfEPaqMk4/3nkgstGIrlALoomBoj+VJaSRheGGr2RX2
A9qVXYFQhqUACmj9oh79JZ7qi8zePjRQ3r/gM5be1q7S6/keSRYD2r9ZVte/MoxN
lSyvDXxracu1OBZsDB/5DCVq3uA1jzQUDvtmphXMBSFgCeycKolVGScKOw+F/BgU
9bzKbozrf4NEYMEXOm/4ssYbJtYmv8JZDzrxhcyijjPZ49XRvWivvUTgRel9yE6z
ZmrS3DzQqQGQ2QoxwH4wf1+rVFrBhddw6fUrDYyQZ5zKYKdk5wjxYRsDGR2hY9Vp
DSP1+MjTOOM/ZF4LtnpRDcm/8+Wa9KOwRrmbbsHtIePv9Z5o14A7HK6durDHURF+
f5O6IOpChXuFH3grUms90tkaA7k+bh7AmeUqdfa+ouDADIFIpX81PD1xB9UcOIa5
kXzQWNX00FE5l+eePLyg0388vlJfeYh/zk1iu20kKOP2lmmWDmPWyp4ZKc5l9+GB
0GZZdg7PMJNqfp+RLyGLBtUTfs4czcwZk2/ICjMTpwTvLV5QG70Y0jyAQtwSGwnK
1x9DDo7VgLA5p2G2+z35qlkQcUgJnf16w76mU3+BZY9ItClR7YWwv3D7VDv1ZbP9
pM7sqIN/AuuNtEt17n7XOZs8iLyRmUlzjtz7emztO2Fv4jAYL48PDkxJInawveZg
xFnZqViU87cpFe7Mf2PLcz9fFoYFm5+gyF1aLMxYWMBTigpXgKEf9VGvNVOSsfGG
6QLgLo5wnuX62jBm4EEmooC5K2FsMtoYQy7GPzAxdZABNTbZaYvWH6xFN1xO8g5J
HwUPS16O9lbbwX2VKRPfPwZAiXSjBRGkoSLmTFw4NOmFlMbDXoahrlJExIMc9Usq
ulo77VvfW+RwRUPJshi4M7gbS8K69KacKzgsvyhoM/ZEIwxmtzMw7TRBTynWEyn6
vFOPvf3RZqbpZ4z1O0bl5ziJ9IgaclJpVMSL8HX6V1J3u0m+POyKvx1aWorq2zYI
/mPl2JtaZB16MCf4rSzQbx7OtVPzxAZRIjg4kwDICYurrCcCEnThEAbJC6EpIa06
WKuvQJQRb29NVvAJTq2aD1CtzSj14YGxOxmwTbP4fXx2xVXd0PjAxmOVyRj+Xmwb
VsL16phIc05xoUA8+qVCyNw0ebGaSAKdFsasUk+uXKSkm4X88vARskCmyLirQycl
JpNmFafR6sluYXsjKFOod6B7bIop5SdP1Ym97sG0OvN7Y912+mrk6WsA1zbVdSP7
sO0trhfsjcvnET8+2ywG/cZ5Xt+Zu0/kiexHf9jf5sXt4xoKAT9Xn9Jth1MfkKKT
cKL4wzfzck20XGVAjVVEdCr5GccR/OGFvkeEF03SD4qH0NGNaq3OhjTr667SV/Dc
Dx1cTlFqoYRmR+jBrlRKSG66xb6wVafcjWYk7uREmZcAIz+eBNumpnKC26yTvIFz
GfhC13p+qvpqn8AXAv+9zNkT/P5itTaTAiFKRowmD6rPc5Xq7uVXAw2rZprWkXoC
QjOv8vKOyH7OVkWFYfhL5lfolfk5ngp3+IYuo/qgq7AZWwWzW0Z5habm5ZQxIZD1
DplBdw9KptzH1YS1qryTDMKxM5dLHQgGYrcYwbmi7dmN2VpxL6/jCHth0frmY9QU
o2+6Igv8SLlefSZIamjFiHWzIv1zNsraSVYZFr2L2xaK4tcVDeaX8Br2wIoJzsuR
N0CKqijs6fHRO4KW0zq9zvzQq5uTKjvYLsvLkI4eUJid2+hoPdVLnHHjINNNS8oa
DCh0+eKZGgTdBb7EbOLeoBa+a/nrfjjvrgWUWKWjbv1xKo0RSz8uxOXtDp4m/f82
By+KSGjJKqHgFsukw6QjcoS+NT4FRgcaVthoFvELzi1ky3QdfduOaXp9Z/eI9fts
8G9/RhPfvUNY0xFASKh1kJ7VLXp9bD9sPAhj3thzS7W99GjWsJSpY8sWM/O2EZzH
5y+FkYIlA3/Hkg6qfnphRqRdTlmkXe5Pue6xkH5AsXE79TfYslwofl4iICsOZO7E
snsGHPRZVFKhhfoGEv5M1TLTqMmAU2b9zMs9PqNUfln3Hk7CprmcWTrJN4BPHALm
Ly9ykHdBk9hdnq+t98GiYQT5CCgTeVdb0ZiUddrhos+nA3dJKwtdWKg/FQC1BF1u
fi8NSNVcJGzHkaWQh+nqsv8TnH3R+WjNEaoTpE0hdXpBTlG0Bx0cDl1rHYR3FAT6
`protect END_PROTECTED
