`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QT4MGje6H2RuQ3senvivYDihtTD/lH7yBj187M4Mfap8bWNs0GJ7ovcBnIEu6z9X
pv7puJvVkYTjGc948GRaazRGsJ18ZPqK+9F83uC0o0f7tm7BODvPpUSoWWK9Q5LZ
mmHAhOwfhiOHnXP/qJfGGHVNex/8LSx49bchnxtS8pAcilF63el62GO6saPA4LFP
K9iWxg98imhsqLCQofpxDl3XmYqomx1+K+nIuNRKSNmSGUcw/Y3BX0Xgo5Ye+Ti0
kYEZNvyZlmOjopT2k1Kmpg==
`protect END_PROTECTED
