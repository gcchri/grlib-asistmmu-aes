`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e40eZzw9qDJ3Hub4BxTY+l0VhAVMpUSTCj6y/5uC7dyKFQnrokM88g1kxO5Gv8fW
xxVjhRIw2Ab89pAOZ3DENdtecg32iF05pNwLDmVFEjySX9PVm0ax5usO1yzyIPPv
3sQMCV42ZYNRllBAyld8UdPXUGEUWEFJRDJjL/IxQLcHh6ociAUYPDsKJjsmgk7A
uC2Xia15DFa/GN6hGbK9fv0nveLF4P0pz0GTtIbtHvjdT8KCoOjrinTm+pMfKA/S
iARrwBQ2DVR7p0B7bYy5Vj8v8n/uH/Ijvj1uPR88IRntVIXdheUSEWiiZ+BPIK1b
uK7tmkFlJEGEUWcW78Yyz56/Bp7O/uif5wiCWAlYw+g5TI70lzAhkk89LaKsHWHX
8OO2WvItZJCOFOmt7P3nyVU4tgTFJ80exX6pRUTLJsBlYJupKx4gQYrDUzEmcIS6
`protect END_PROTECTED
