`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fkqUGgRZsQlK54tHb+8QLRmW1e/3SlBJUIonrmdbjDzrKtepy6Kh9TPFuNkg1P0D
VlilzyDHfgBYzXfuKrR1COL0n7L09UCBZUn389fxiV6MQnd2BvIpVRHpvN2ydYJm
s/ci3su2iZcLDliMP2mIYjtIR3GPg/4WED1lah64WKgVt/ZK9qU93THYCPpANQJq
D5cJ+DOX6t3dB+IUtlQhMT1Xup1JMP4XE7OV1c33G1SUqoyttPcMDOgLypvJJE/1
4ofEMvXDpd7SkQsggpjHkRYqRQzYoc9S8RqohXR+A936QQOkDmPsjKRAkcUrCHNZ
AFzDyry2VuUX/tU11yVSAGPkLYUJ/AaJ6bErUB1RzJiCWxLxMhdD9JeZszioF6Ey
2KiabVjdK3mqEywjRpodGuBgLgXDv/uFlAVZ/Z1kx/kP3ZZ7de0s4SKd/iO/mUhq
cHwIoyD9RMKoFaruaDA1PfPGDIEnChK76lf+3spukg4/mtJk82vCWips4D4AAaVU
Zw8u74FG9Hxx4jm5NYAEhSiPLb5a/4eAcToBhs/DbcLw2ZEXGnoeB6RD2A8V4eZj
fEkj421k4AuTn+OijdkWF9rzftmeVlGsxWUU+7qOaodNdU1BdzDjjj6RMAT5Jo7+
fnZkKwYwHV1UT3uF1iO8RPPLf7FbpbmYxIceVFGOeku5FYWME1GaR2fItC8IXYgB
OXJbOojfC44iIOWGBzUyNpb1w3MWBHlH83wk7tWaFd8+x43WndtKmRfHrhg6Kdrh
VYo8e6MI9LRdMyBJI2vKe0U9fS29Gq7Y6jb8iUvelfEQ65hEjbjVY800WYYt1Lpe
MCtsOtEQMXlTOgaIMBSCPJ7NiI2jgcg0ixn/HPyn5xaYIgh5Q8/XJ8/e9/Bly5Fm
vnMUaDAjXICvkVUjYEiRLDO1GvWUeIQbyIhUz6BNzaYthm3rT7dPqyoH8MyBwd4e
I7wJ/Igg3L0VNyzZoajTR2Ltbcs/TA1Lfr/9/qlFq7WViwlTOJe0D+FiKI/ySYgS
epPNpnmi7rmq33xx96cqqRV3/bUrpl2YNz0owfhWbHjeHja3xdOamYrmXU2qSh/3
nYY+5M3qOBo5S7T1S9Lq2BmR6TkRBQjDLPSY0CIX/M4C8MDUxwz2af+exp7MKlN1
bjh87qfmANDT+HPEe1/J9Y7SWnxmaQ0rvDPTKqBeGebIqe0kUgWGCb+43lxlEBjA
t9vODsDj77Lr00fi2C9XxFqhXnIrcN/ZvSQ1Hq2uvFoc/QdVnguXqsibzcBz02j+
SDWhqmIFX9btt+CRtEF5fONn+RiXG+br1urJXRZ9MgC0VkfFJpHIEaGBRqED5+li
LzEML7eCJSkLRaqvXwdxnFcE3fCDGaQ9zfZI6YU+GZXDLKQcrY83zz3woaibmfSR
tw7WOCHm5BYLPtbMOZXAEU+s75iwhhtsa7p0b6wki9lgzTxN68DClsuflFuY4Fz8
ozw+DQ3jn7MvyBmr3fSFjRowRwcZkqOs1EwFwYmUKFsB+6CADlRhXOgxSOgwdfYo
nherZy/JJuyPs2rn+0xQXW/XYk1f5v31SRMDozEoHiwe4YJXfA/YiYCdqjpNowAA
yjRbpJXdZBMtHBhRjPvAFy51e5/ShDk+RmtBAfbWXZhelraWyxEhADwchaBCEInM
cfAimhR/VyQWK1rKBpiyRAS5dSnr3N1CvD43QTK3NeXhKrTp10YI4nx+8Etsmf92
5iVnETBIJ4XLOg754Pi/D7mlV3tBBsY1Xks1g7Pt3l9EGnzoy6Htin9aHET6eJiN
IdxxG613VNfrTIGrkVM8NLaC4v3xb8q8nE1tm1IbrsZk2S0pqKO0YiQngHw6A8nz
Wmnb9eIWp/RrtrFBqc3DEAS+mYsGX6RliwW+ZD9wwTe+rXLdYwWdjeEjmdc6w/7K
I2q3BZZGJ/TDaS9e/auuaRHftaGFIMlQEzp+WvWQx70UtzdjlLV1hAtcCesYORHn
rB2e+bHHmYSczclM1TW92iiBd9yxM1jJvLfGEbbRylZKLhoIWxgUd1YRkPLs1+sS
24LGtEgbBIhEXWAWmTP/39R8Wc7Z1EbHlqKHLkgFWm54Bs8DLO5Sf3RIznLUKUJl
ovs9QjFjytYV0cNY9mjb4Yt0Nxxs+u7t1O/fv/i6hWK8rs537p3TznuI1S2f2GLh
z2FOEpGDp5diHVaoxSUZgA==
`protect END_PROTECTED
