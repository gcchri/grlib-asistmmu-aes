`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yhyz5SVIkxZyvlmtaOUoXG7zlvj9t5sg/rfbtRhdqCu4IwUtHbUgJFsEzJ/ZjxMf
qBoLW/A1AdBJp2Y4Zxv+Qk/z4VlKIFz4j3qtXyPJNB3ZHBl5Gx00BYNpXWg7wvLS
ceE2V+EQYoRM7kiZF+VYDbScoCPo9g9RgH6MWX9NA9JGbNs5+UVqQk3mAG727f8K
G9mxRBAudhqTphOqShfcpRFmv36WnZKLd+XE8M7MSVSJyb0nIh4050GWZoSjbhJg
QNVf+93XIyf3HkHqdbjkLjabOl26NPqFcRR30MC62vCQ/VsABW5tYwSHZVbC6Y3H
IcRqnLUx4N/1xchBQF09rNcCqFb3ZaW+wVIKKNY4wVdr4Km9J+gxSwIX6J6vAd5a
U650473pBrh3pDWpO+Y1PqqKkoB8xgWjBpgal5q7ssrNjuX1Pkx+AWclWaMHVK4c
lkyZvVqMv/FvhRX2+Kmfx7Ndi7wZ7sKN9lKU+LowopAp8boVugU+n3AcCIqo/V1M
lww/b1ZcFdWRCX3TbhsMX4F/C6nGuXcTT4kY0J+XBR6oT644mkZSWuz1rrmmnIAd
U1mzO+R0RQ6AVaUfx0MGA1wRSYY7PSNi4tupZzgAowDw53xQmV48lROQ6FXPI8wT
IN9RsWj8cw9+iWCgHnNA5Z15H7NtG1q68sE6dreWpukuNDIqOL+7OKXJjyLlh/Xx
DAn6xUNf/PaX0wTN/7zAZIxRRlDnYBkR7UbylZ4vh/XlQHBEZdfB6mqV1BHEk3oc
+LAveiEO/F3GPIE6brSJeDij7IV31IAF0gy3fUQrE2uHMEBt8CyJl3Nz3BBl7WL9
YqWgSBaUpEGGeTn9PQd2F3O9PsyJv2Fy5GrnSDez8sw+N31vg5OYTtOfti/7LmUX
cstE7M+wq6uuZaBeBUlut2TiE9gIdnZK8kqrsUhqTEubfGEfumWldvvqe3DQaVKg
VWTgYYAB4grQMWw4+wd2KfYIyqFkp71c3yC16F2S4I9w9ZUhbO/Hgz22mp4h27Fw
VstrZIHDrII6XPs6+KuYbacU6RvmJPo0m72O9J23ub+mD4ih1ygixRthWSxYSJ2B
mle8dc9pXHtuAY4dSd6tMK1y7vVXZBUMdIJCHFJ60mzGf2Cj2s8z3hOEwusrHhWq
T3ETO62IHMATEGBDy2xOBOyHI8sSY21NkdfpF5pBCKc1CKdLM9ejNRHEJ53SZ99R
xgRUp5XO4XRaxcqGO9i1KKD3BR01nZuMTA4dQgnNm4Vc/ajgnd079CJPvKmNAvuv
2WorrLe4SclFhsl6kzNEK/e3apa7Vymd2M/Ugu4Cr1GwyrOCeNfvBHk3BtxqGIzT
X7+NTx3sM+OnhxXBYcXDkAbj8fDz43xMk4umLY7Ora2V1sZa9LFIbSea9fTCFef3
mImAUpDJBRpz9FTXQjh7GrRVA5IPhZWupa37H29HefXJKW+p/TlVQaTsHaR386DP
Qqi89hB64nFCrAeA1djHlUBVhNg2e0PNVHWEfwR4NkIGzO3DHevt0A/z6pMRdM2A
zN5iTM3IVZFLHc9MJJnTcT+z+nAxBA0IL9RX16tL0Pw7NSUoZrgfJvwREbxrNkgJ
A8YBbXEZpgculUUACCUyzQ==
`protect END_PROTECTED
