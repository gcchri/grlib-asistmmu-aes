`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D/7PjUtyhVx/EHGUndMNBW388Iwaz4RXu90i4z/TStokKhrNPa+inGr0LpP5ZsI5
BmL9W/Jweus1yc8Khva4aAwMbaGUMniDxRxkhCZn3t1kzf0TD50+UJhYtmFnf+eU
kK1Xx5UDymE8m0tc2XkaepVey8Xdf/iKiEfXlDyQwARHDT8TXIL0BBly/J4lgAJp
Bqw8LVjDzXcRQJVQsSPD3tUPFm77zYeLxpWo1UdwGYN4Rrj9kNr/IJ91+QD7a29M
t1QcJusYrF+jP0M5N4GwQllYNRDEw99xua3lC1sR4p1RL0lAbW08/JeWliMLoQPE
3ejhbzG9SCA8vyYHkXl5R2cyU85R240aZMCg7Exf4CqboFm99gI3S7Q9hxUirf67
Sjw3VRjSZWtkBD42CiuAdd5aHR70b68RaNusdJq3rZgOEooCDoOzggK7kNZmb0vi
WsH89Z83IF1+NiEKklg5auUaFTbCUxoEOqn4YCzKM4hbDKHK/z6MScjKyBDsNXxO
Kl9sM2A+7vfMH9DwYISv8cGVS7g1eNm0fNuB0vyLeb080TKcnRJyVIHpsa/ELlPx
X08j5/H2Cftu0n/q/Am+KO53m8LFHYSGcMH+quOvwSd6XlrS/g2ePh4IQ1fOEnPu
kpVNqvR+nkQlChe6YF6pnL7LANUJalVFhkgwi4Kq3PfPdKrUDSJmEgOUbjolJ6Xq
ar3IO4KiWzSt5LewYKEV+IQ5c9+I2q81RG67bBjGIFA=
`protect END_PROTECTED
