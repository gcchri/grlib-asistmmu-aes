`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YOl42cmmRbc2xM/YEp/3DvgKCD+lR073nyusY/ErNfsA818mn1VbYQuDc5TI/+jU
rmb0pRxMVXUXCLIxv4DY953u+NI96E/+DYBfwglYjdo+FAkvoscFtKZHl4awe69P
23tgFtz6BI4zPCX20WR3Vvqf2ZzzwPm0v63rmvyKzOXvJqzMVzjSfrjTNXP1uEm4
pNY0XoRWpppMdAO7vdZ3oYoetsyspIwDA0qKCuQ0Qthrr7iDjAM3w6Y+aHm05mF1
R42SbIZb5kxPa5XNHXcmHAWR4BhwqctLENbECbl0wlNbJZQPrWTrl5V9FcfFq+bR
uF00H+SrkPTjgUbbt+TFOj7RxEDlpYHc5mZqkyIjffnRNsNxAdSSWOo03kHyiafl
y1gSChu5Vetfhs9IwJp2yQ==
`protect END_PROTECTED
