`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j23yFGOTvBi7fppkwofMBqLYIddle53ly4QVUYMIF2rFjhiLldognGinmxR7qGUf
Vhi0GPQi+z20sZ3zwJoMahuweWohM2S5wkmntO5/p79IcReGTQBU7IW5g70YfAlU
292Hq0uDsx7xi9h3ObGiKyHz6e5yai0UIexeWvc7/UWN0SahPXRdwLbPxhGJfSGX
19i8suaiE+2m1X/Hnq3UxOfJrd6ZmoS2mzlCkDkzTNiy/W4UO1QMjU+rLQodB60j
xTUKBoUeDeNIVT0EOUGgl2+Dni5yo4ISpM5BVV0mEACiXKGPnF05wxGrM/DfZxsv
rfD4fYITZu7B2B6XMAExyhneyZAHcuxiS2DzadkU/Wt11M9fdonn5/KpyEX7iZCT
DQQHKL27sOD5ux8zXhWz0yykCZdTJaiHRY/SMKIvRlFIXCHULBfIAfSGHjxBKCHg
W1Nyr9tC9sC9MGoHM8tzxG7XscTa1MF/l2HyAQNmxaoXqGtiCB5JpGLt8WPVohZj
fnGvfZzzau4h2ISaWb1c9gOo62PJP3WK4LlHY5qqf/Dj+g1o5MmYKAjaP1+fuw8I
bumPAZVL3os/OZYaGcb5aHxYoyPK+42SjUp0j0oKMy94dFzJx1ejmhqtnBs/QBHT
FB8pn9jKLv3gQbyUIkWKMFFEh4DcHPBCR/M9uSMCnhzQjkVdqCOupdbtL1ojB9f5
WaS/NSlj2uSvep6uu1TpJqOdLLUSYR6eWY5Go5s/IGiaRN27yUT3j0h9wVtXLKaz
8rLJEzx5nSeNu8uMJ6ytpQ==
`protect END_PROTECTED
