`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9I8G4Vf7SMclk4wnQpoJoHiO14ATGnQyFmAN34M7XSk8btlhSKCMC3aMdDIM5kO3
JObTGTpD6NaIwSu+DOoGoZFAAAs9xFnCpZVu/fmX+8xGxR1TE1U7R+jGAjcCAJEP
UYE29/U5ab3G3ETdP1hRqBhq+rPbRIsHoAB4mB1YVYILDprPKr9U++s9aIx9YhCc
2gEoCog2c7Sn+X5Mt4juyqY9+FPs1q45Nwjf54uvcMXWoRBNc0iO4k8hB8wXjmJh
kjqeyDYWFORPws1UyR9biANq0LSJ4rz2QPXtEA89QevtHGYDQYys67CT0GJsSbOW
wYKQ2jY5gjwWS9p+3LLFZ9AsTcCT1/3kmgAXlFsMi+u/AgNb33EtIi8tnYfut5JW
NNOuDkAdOTpplwSu/Cndwh4fKRlt77dfXsGYIKs8iwrP4AP9BsUHMepURDqPNtFD
QrDioUuw+UOif5rBvNvNUQvi80e7Lm2TvmocnEktHW9PKx59R+kOg6MtMQKnSR4s
zsoz49/abhWefMZ84lKuKxKbWyz0g2IQMOgQkm/NAY5SoY9PUCBjPixkSMkm7ix4
Fa01YOaaVeCU47MKVcmiSEf7Pz11bZLxS8E7sEAC2qD4p1Sdow34QAKUE1a3AyG5
RQ4ukyKeDwaU0iT64B27RYlDDuU9kmjeHwquo0Efr7tuMHOo8rh5wXF6pOqsQfN2
qGD9uJUNMo/HTSnq4q1Nuisd/XXaBJKaLreEf0jWbKIpbar0W2F4pdSZbQHLfR10
JB/PxkDZOAuMl5/SdJFIsUEJH90aOIt2HeVZ0hlcryQlo5CtlDJx+Jahkl8MGsrZ
wxrost9lNGg3Ox0ol/RFsPW6a3EAEigvx+w6SwS1o4DqAJ0E4obsUX2n1PHMVk2h
pNBSYtspuOjMzxGYUKut+CPTh1PWKZIPPl+doRrp6icBi7H3PhrWREbpAA85Z+U5
T5vqigMNyBulHO8ePmg32Sa9h00IHWuxDfTzBKf5x7cCVYgsFf9Hwk+evdZZj5MS
`protect END_PROTECTED
