`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tAWr1p+oWo8nYtgZgbKFbBxMyfRW98Tz4KXaKQd3ZwFmWN/yxZ3q7DBS4onvwjPc
k9kYfkVicgrPXcDJSp7pjhtWjWF5C0gfLLmsYOW7XuEYNGPAETs299XYkDJrcPGn
tO5dmd6Ua+tuaMgNmbXDtckWzm/H6QrD2KvGgB9FxisvAjMzQMneDmoY2YafO1Am
5NHhBewUBxIbwBJn5sNcrlrPy1TcFNNP37XU7vdoCB2yOQYlWLV3DFHqrECUnzX7
eDM8af0bijV9xgPJNYdNhnDmfEQGA48Ve6nNOJkx4Mw8gfdU+0gH95Xa2dbiJSbx
2mmgG0hHmZlSixH0szllJA==
`protect END_PROTECTED
