`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lPcEfXyLYKz6BdmWcMBXKPREklIf8Fm04cZ3/uS4m07HCz+v3ijqRib1yucjltr0
RrgoxsWTckW0vL0vFWkYMNtN47fuEEOiW3A29K8BNiEhEBHM+OIoqJb6a2lWxAH0
OZDfAZBXrk/2fDN73jBm46oOk1NZsaGNZYdFk3S7XXk8yGbSuWUWH0Nlk0SgrIVX
eKZ36gLjQ4YqcvjAtFgJj+0hkXkitDqApELEjfnl5/n67iTcsl+7k0Hm+gbk0mVT
XxwVxNz2SRsEtwwchnZR5zRcwUYsQSpslX4Y3Fs7P69TErrUcjCUXpd/ALA5ttXm
k6gZo5Q4CFm3J4tgnj/rIGoQPqhV1pRtrdBeVBK5be+xp9lYEsQKbaDPGg9V4ESq
cRArBkvFdDwMNGXr2/ArvGhT/9UnaSPvScO3mug7FIyjqpYixhfWRBhE5fuW8Wcv
+bQs9XDh8ZRQ33B/zKp6nLu0hmqy5fUdCJjZtTRaPnxh1c5rS1S9IscVdHOhZihI
OjZ3ylzsagbe4sNxqk/mmnnlQfqG4XpNWrxMYWjL63HNIau5eDzMuEpXCmamjdtU
yDLAvH3JoJHcWIPDrSXprgwv0RMi/tArJosUCoLINUNjllgRcpiAfdBoGfb4clqC
7fVNVyHEJnRxhAdGylT9ZzbxVT6RJRsMcC/ytVC4ny+x0VYvtZqpSP42oG5cmWs/
I9+W0Ony0U32m6X0IvGXmh/Xn8KS8gIVWIm6VYTX+HuArNgSfe0HP4c+CLElaoFB
8xagb5trrfbXNVOYechb9nZcYvSsaDa3D9PqSDWypLJx1nwT/SlAsA27Osce1LmW
SfqRxGR6TNlA1rGAbHRFvw2FPvuvBDYxN1OoQgujmsEzoZuusGUtLuhahXQ0dFCj
9/Wb5WcC2vSIEWJevJO0N09UPOZqxm7UnHILgnG0YsCQzEg3imfHUqLXCEd928dj
`protect END_PROTECTED
