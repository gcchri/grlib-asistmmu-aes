`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FDhFEnGBFjUldqP70OYtJsD+Zvd/+4/UTRTFGsBPvSqxH7QDIV6/AEoASz0/sEr+
n96qbkGMcs/oNC2xdLnvYw7NV0eUkvTN/zZQXgatMBrA91fWnny2Yp7sGv8IQc6f
oDiRO7yjmuEgCjxBnNzcoiCliMgV1ZLhe44eK0T3aSzzIujPQ0NTuG/equxuL+JN
m7YWZQNl6LBC1phTEGCRZlMpwBR0+Isylwee7WofeyrSLTHkLtEtBJfyLUjPWpcx
unOn9KD3Rh4jSRbTYwqfK70qhwKB07wu+O1ARaRg1hYwaVzl8ALAIq4K5xEwWt2+
P9HtSWivc1pkK3W1SXNgUMs/+tEqn4ceCukQgyxAm0/MXsKBtO1TvfdfMNyFe0yu
DbglLUqqdYX9UlnPsdFuC7VIS1y+IS8aNs0iz3PQewEtd5aCZvHPWDloq9mbG0Z7
EeUvV55atsRQz14J7A7TK5q1e5es5Hoz+mUeyWOTTY07xHdLPm4r2ZxIIF+7IYDU
0T2KBtxfHzsL5mpiR+e6l7QpVQC4ERF+TRowlxe0stskTY0QJl4YXY8UAF8Gd9PC
sOCJsXjjKnmymnsEsNYqBtLbhanoqDOHM6XuqA3g++Kx3p35KuOE6Ut/Sd4hq3T5
HKnk338Y/LU0OTH9/PwwxGaINTrhQWhR8TJt5dVXd4U6Kfv40ZnWvEAaVBbdsKVa
LuZbWtIicLCCNt6WizpMTYicfL3fGwLX5+rEvdsiJqCMgdyLYeftkfIfasbh/Bvo
CLGJUjzkdcQIXPOGu2TKcT9LweZnk+SXhmV1ACJkeergn1ZnlpEkw1l73iBuZX76
fF0r57Ur4NF3dcM8yGeWisZEBMahfcc8XqsZSYDFRIZIhfiiwT1AN3cjFYoFWXj3
/X8u/tOP1gNTcdIaM9Si1bi4qPOupv4UYdLkKFCOIOLiXxcmry0TuH6Gdq1alk7m
n0YlWhiuZNCRZ1RweGueW0jhdrm5GGjdZYItRmaKacnatF0NLO4P84gzulOx4Qgn
xGjgPsHN/AfvXh/cQ+vNJXEiSeID4HPofYXALkhJ2w+FyJUACJPqc2/4HMgCmWw7
GoNPg7EaD21gQWRSBh7N6MwgLy7xv8jlR9xHDcOmzRckjkkRHr4nR+md2XPG78A5
u/C4DfudswjvxRIuiEijFmsv2E/7ppiDpMa5KGaNE/+A6xfSSm3D3by12pA1fH32
cbeHjskA7iGxRECovIbM0PuwQlmVDBOfMEPJJiB898RR/eOtRyVvTqpZbpSvf4NN
CbHG8GmUXHPYVApCrP+5szp4oI9hpkzSSEo5svGzmOpJPStb+gKIITYxFlLPqSzZ
/5Nz3bwz9GdxCCGfGVLVRVXGP3Y9fV8lAzR5qUowNPRsC6kYCLC+3NM++LVKEOwG
5NQDyJ9H228SDSPsGlecHP+StyN5/vAKIFBys/R6ix6V8pAqO4HC9fz8iuoY8Efl
FenaIZCwdws5igRLB5UdaLsHaDu0PO+UmDOcYPMggANcYGE42LkbM4eStXAa6fwn
oZ4tC8D/ts3Ief4+TGqMc8RrqMpzxIqhYRZt0zWRR4kMWgohWefZzp2mzYjSbcpp
Pf8JwpCE8XmHwXL4vyNfQ8LppnbQX6IFkrMbtdzXwDwYGZEDBw0de5E1jP4WK1F9
zidatpfFGmc2QMbDWKbULKCK7UfvlLR/nDStZCa73xXqdHuzKu/e2PqjS6O7CcVK
/CT0ZUUFSzqobWiw8ab/eeWBxcESgoyuGJgPqtZO9Q3d5s0SPxwY+YRXOvPxvkaL
CSue0P6HI+sB/6Hxg2KVXnKNCnos3aQrXJfVrRWlVKjkJBKfmQpOt2AzaRLycdhD
FpNfssgEcl5UjDuNL+R0p7ghsUsn6oUsk94eSPh3owmdVEMy15x8igNo8auRsG0r
OYxDWvKJ6Ymsi9wuG+Pq7Q1406U8wU0kF8rJiLlQOjzeh2D1lRFlbqEsZY4Ci+ni
BFXINnrw2pp7tOyhiXGgqv6Rg/rgsH6eLdQE99mkrYGmsfUSBPPqoM/XclfnA3ML
yRGH9YedZKJC9AD5fF6UdXJjtdf6CFjlfWlJStlq0Bl+1oRTpXJRaOfb+D/eInBX
lQ6QekVvx0l50KzSzTGT+XgH2TkWIBxIVKTEuNcny43A6WCHgnKGV6+G3odFgz2t
vglmWRVdX4oLxWEKRsLBFAqXryY0o0Qn8RKVSidtKrlg4cZEtesiklR1uQXAdWOz
TkNElS8D6J8u/kDfoX1j1BWGPwXBfnHLfd0bYhKPZnL/9R+nXYPFK0/Fau5ydSUr
KD+RD+k51zc1YHQKAt/XnaNsRlxm9dZrXxcQXod8dyeUf8b/4JKqZj9PJU9JCOIP
DRToseP/2oNLLb1+yDPJaCsj/Hs/PJwMljOnIPxoiTv49/7OmejKuHE4Lu5DARMm
`protect END_PROTECTED
