`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2pDzYWzX8dlt078p5bCkn7AcrUABmxCnTcfbxbbAORn7BIupdjXoIofU58aRZCro
AhIZcnsVCxFsj0bDTfMHHsDr5UNh7oE5vWmOrBeD9ZVq42nqKQ6MGdDoWpi7uEIM
GWBKRBntPU9EKBHWL9R7xqnA9q4GxsqSw+6D12hIJ4NfzmHP2LTRRN0GdPEd1gbL
58wiNg1lL7migkK5LMqctEItdrlyJqkPtm29A1/bgYqh8qBNyIzk6kLkHYaGXzRX
+5sxaAkRLM2DNfxiz2qTDz3Z5Sq6oe84M8+ml680cFNMtOzz+ZLwpSNpKQLcRTWB
Z1k0G+JQKrsE3wZPHxtswNKyQbZU9fdJztQ3YQIdqrBC6rVlNHkRFIc0GpQIyEXU
HAUNv8K7/YHkamnESpaUiuQrlL+fBZohZnlX0KjIXKqE09V7/QvsSX7xjwGCgZkg
L9NfRg4d+Ms0P8w7mX+c5OFe0mgKShoDERYITLVJcNDOHeb99ydYlzTBNRS0nCjv
Ux75dRhRapYHiXZcveRd6mh8dWtb5XZ/N2xe0k8huO70Jtrq4TJmNm3bRPmpoP7x
uWDbO53XHvBa8WOCiYUmggnl1bXdgbMyPyRoWkoEiwcJYFDaLvAtYuFJaI3fNNwl
hBpTP4xcigQeBgKT16rpqQ6E30OINuX6eI1xYucfOi3OikTCio6a7dcnE1KOThTv
ZJzsJ0XTufFnu/QHmitPoFoVMJcf1+uH54b0nNL40QqW5j2so2Crr2fhkZ6E49bA
IQ+h+nqyMsH+4mV+GAfK3lPhvvPHN38h/RLXQWMIL6hEYpJK7UxWvOU6cSmqF6sV
w0GGkboU/3Yo0Wt3q6pjBpiBiR2a2az4APsD4yfvfaineHtve6XKHx2hhxbJx6E9
E9NwIaeQvyPNH3AW2PwaV9Mp8ito/fih9MkVIFjzCJ9ewpZ/sdkA0M3mBpbmIP5z
2ZVIylaXwD7jUm9VZ8QJfSl2QdT5robfPxX4fOcyjyoU1UwTFqEkGHaaiN2UBnXD
wy0O4WxmyyQVkFIgc/JJa4TXj22PmDo6Nt1OeYnqLDe+MITNDMKQWud4YV1PeigW
wqk1XUofHOTtQl7z5kihjbSoHMs+m5ghxwAkfNmWm0Vw5OLsNlZSdgvaNgbAomhc
wdGhiC7Jc39rmAwqMZxbhqj1oytWDNEJFqIT9dwoNXKnss/RuYNRWzN3MRbIzqyP
nfD+ftRz0aWQeXddmm/CSx8L8IHZVMba12wMtgLhHlbWBvT0FJN61TRMK8DI7vMn
UjN/HCb3CA5flM7XXws/+pzPeYSAn8JH407JAvI1OmAJsNknqzCLs1hS2wW+XhvS
mXXUBFGpFulI7jtxLImRVX02NCCpZt78n8f1akIsVbNZbPBFJAihnhpw58CnIWrF
cY/guYHy+WfX1dxEX1HpmOzfj2XwcKrfbhMnKWZ5xxwYl994vVPisr82xyptS7Xa
5AXIWx7XiSRgGBFDGMp7mh70cSH7kXTGyTuIDlTit37Li3f3qLCAIgNejrm2ETEe
lFo7SdCjObJoSMwHrfTLe7xHksLWG/Lz/QfEBDDOo1YHXxK0bDjYvrJbe/fqar9n
cbXxhvj2GKAi3S/WxMF64vKMMblnJ41YMZBQ1yHcMaXA603XSPoRRYV+HxRtIosw
dqrc1hjFyuJJNQZQjbaXnsyhPlisHzF/w5haEcnq02gidcDu76XTzm6DGZuBYxwv
p9q1BpOOP5P2YqE1i9xDI6VX1rY7nL1S5YqtX/d0nJecIFItlfrlma4MqxnGDrkQ
vKl9WvbH1M3FF52NsLP+uO2+YcvtcB30NvXR9aJ1r1EJfB2R/3Amffqwta3FCxr0
LDVnZOfP026JlfH82pitAmM1tNAOubBJQ763XVt/HOrSvbnIhiW73wVO5Iq+ecLF
OhQR9UFXXpB4GwJpeMU2acOFpnJD7NdjdVfK7OJhJm9N+hxv6HsKaa5uNV6X6uWN
MaVghpqLVkbj2WSYW/AOc9dSRp+tLVa85/86Evj2Hx3GlcC5h1u8MRXebwi8A6A6
QfdD8qff2n1LSGCGFUezzWia5Z8xIFVhGlhz76/M2GwRgcZ8siOSzSh2a76m6aEQ
0iU80lcydPf1Rr7jqZUQlpCNHfE81wpUJJ8EXgvA/NpVO1FqYLZt8jIujQSpKrUN
H+wf8ZphK/kdt1nL0fQeX0OsScHLPF2BTprSfC/8BWLQKuPpqeFxwAierOXiIVC9
7mQ6x5dON+gw+AUQy5Pd0RCFeWbUl8LvoQMkrW0XIW2nn9kAudv8PC6qDrh0wzTj
FCx5oQyzWVOc46TR+AhRMTQpDAsuZcLtv2MbY/6BDU16Pcjmiml4q2qDxbF3MyAE
4WhaXh0FN8XBspde7QsuD4CiqihhhQSzfInDd3bpo04=
`protect END_PROTECTED
