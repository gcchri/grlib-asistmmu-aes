`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bm9noGssujqu8zxNbR97xbBCZLyCYZQHFhXCPgwq46AkrFvlJGebkhPvCbiuMs1v
EnTvujB1JVu5eGIRW4bv6r1ubAAmWF5Hth2JvuaCNcYkfJjAEMVIzWTVPGGNnGb1
0lAI2PS7cDjBJpFEfBNMItCVAIYrgcyClC8K6mEBgQxR/q/FnVvxmGcllnN8FBMp
bw1PJTVwm7vjvk47V4E1rgCcCkvcLqSTM8W6+1RPM9X1sU15MIfJDBgpCtLZliwM
A2dk7Z0RBmNH8jXLGKit5BVlGAxcLcjU1YQ984En5htcPBw4rro4rwNKKiEgjAD3
zuO2IOW428PpNR3VT5o0hSOjAjlNJlCwANNwoRHQ+bAVQ/sdoLuFqDXDZLUdCpHK
IhWgPEUaMpVhUE7OxUB5jQ4R/tp9F2qq7LmqHf8UZ7MIfe/MaAglmltunzKNMUeG
KeiH+lurURIfuqC3ZLJhUU+3ChF03X9YokhKZxDYtBHcNJKDCwVNAxqxmSq4vtIP
K02Y/z4ckO+TUnH/CgT1ljCeiq4WbtbldTTe3l4h4IyMK01BL+rej2Lef3O9ywg7
0+d3iKI7/No7Hue/AtKVIwfCsQNGNJCkHLuIx/eEU0L/TtGdJC2adEKnVkXvMLbT
TEoluB1zWbcNZM7PPfEO+EC3KTdgnH/wCglOg6p6nb4=
`protect END_PROTECTED
