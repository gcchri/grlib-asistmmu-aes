`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
suOA66/6Xef0BcbqUyQyW17yyS52kxVLc9HM1wKgHamBWncZ6a5frBdHAsWHkOhE
Vo36h7ciRGkn2tbfoDtwrekXoZokuiVTCIIJAQ/EFSY5MmZzR+Vaav80Vq31d4LJ
8dwoxPCrgkSP/M6sYG7+xMV2McFT2Ssf/c4P3VK0tw1hhBx2wWGP19Rt+8grm33u
j9b3v/Jap2Fkx9868DI7aiJLpTj8qhqjHAuCwYrkRPcarVwMQzcwX8rJLCUjsmIa
+CLbr9BkieIRn6uN8E0TsXrIVTWnlrdgVm1GnUqgVFhSUb0r6zPLc1PDWOjzMNrK
d7btQVlxMtnWyS0MYck3Njkwm+zwpc19zyR6IkeZUerWvDbc7UuNc8pdqVkUU8O5
eaiXnlAtFvqbqVVzoB3i9ebNr1Dzpp7XwTNqDv/ahuqa+avOytbYZFU5w/yT65Q0
q8PfUp08Aw8jAWDKuRnlRM4dk5t9DpBxgpcZSJMC7a80DnhZx8V+jN3v8/4pWlrs
34RaEmP2jiSMGp5LgLDQj9IMPr6kEpy8joB4iVjuaovVrwNXHxKulOmzbfYL7S4j
wLiQwLMETMEYTiU3Y5ElnrdXts3gOaLwfSlvM9L1rP2rTwCp4jdBEKwcgzD252ow
oScR6NetfbQujsdhUn42J1r4Rb6vkAt9qdS/xrPkcdAAJg2mhy77lgZhOEGSTXrx
ZbKsTlyEAIqRq6jxGbyZ6ma81+lg7SMR82ohgnCCjX0Kx2NdjtwlXSR9wevZU27F
I7M5lfNuWnjpytCcUB3aCWhF4Ig+tbv8lEUoYyuui/Ks4N0G3DT/OpsUywsP4ILw
amG/b2SIGWLUA4d8YGYr15FtZ7lIpMgmMeTd/25IrpPc4k8nigQITnHqdsfzwR5J
L3Soc02yxvL/xoXY9OIR/O1XHtDMLnsFk8WyMHok5ax24yGxthXqk/I0VV95GTCQ
q9ZK+zF50y/miJdm+OSm5BHH0n02uyxTswMe6nneSsg3XYe5EC2mrBw8h5IXE+2E
BNZB51JKO9AEgLHUiPiugU8oxFlAStJfnsid4QD43mOFQ18sb6S9eUjromCd4UCe
P9Bt4UmCmShkBI8ghU4PwlkO2bszwB+Mv98slZfRCYQ+OVmR17lGXPiS8xH++13l
cRaZuNcG2OLkvpwD9VoQmtv61rwQLKkxWfy6BqREAVQ9nh2OGCIa9YGJmmVf7frQ
6sHWk1e6IONa54dJRZUsq2uQkVwKgrFQKILcBmOpjBQBq29f/S8gZ6tcSNfYYt6k
UPppDDAto6UA0P5o5hkqpS9bQzIi6MgvvyYZtVqgGU8k4k19OcluC0EGHNyP03gH
3pgainXxWnigMMJ8Aun4IHccx/lwOPKuzqpZEjHoSKwbgCjEsE+IrYNa/LTChM7e
p4e0OjOhB8ZZU1OsOYr5dOalv+vU0jXf2oTgmzjqE/qKh2+K5hfYQ+8CTr3v+LR7
PT8pWae5tQ9dOuDNcOLlTNQ6ZJYMV4uhBQB4WSgwsQOj0gDpN/buz16OlpJ9U7RJ
mDi30BP59wtt0LFnPdr6okEr18DoxnkKmjiV9aPYi3RfxSURsFn/XN6EmsL1/E8y
1detkZcIhShx1BH7biq/aNfmTEUO2+Il36LhBOw/UM4oHzL0ndcGLnAGIoYGrx/h
CmiIi15iGJvlRv0KcedSe8qCnaa+U47se2/qRdVAATodbqIhyh9bxrk9MO1TGEJs
4WEotPE7s1c58qW1E53ZeA24vhGE9jZkwOpm/EVt3HR52pXFI5NeEVfO7MkCOWck
7/B3ucQaod4gcn4iQUlj5hu8BofuGrHK8pea7Hwd+Ai0wpDmYqM8qb4jggi2rK+l
FA4Ymb4wK/jmwRacQWwWru0gwV3OBD5WfzS6/8PQQaxB5Bwcm8aAjuE6KInOlorm
bh/ubf1WxvGN0HLEcv+Nis269BXiaavximvxbBFfC1j3QpaiVfb8QMjUtUTmvHnj
fJX1Z9wlxDfMpfvMyP4ZG+Ak+qlWJDLMiGTMhjGGG7Wd+g9i2gTmN89Snny0uhlH
lY8BQ/gj4x+jKB2rbGG3eJS/VzghqCJW9bTL1h33bOEHYscmQGHhMwunCTEko16c
dQ6XdbO4icolLQnTMAke0wU5qWE3edwRXAZdYZ3Ftge7NYldy1nEY9az6SHRgtIi
qD41CojPsKJF+bUOi50cQj/xWim+nRmpFjeRvpgmRhBlqtfDaiMnLAFDWG78cOBh
pGaC72GASG/Gvwq33O0hoxv19UXIJuO2Ytfb7O/UM1FKUpG1d8C2F/uqmpaW0NLY
BgWUzIi0uo1JiJ3FS6tNhovXsEJzTV+SCeE/GF5hmDqXXpOYYbVae1uC1mbMB9ED
ObsDv5/icO5oVjfhpDt4YZTtDZ+aZENzpAcMUtS+NaDcBshiVSMi57EpZTjPhjjP
8zdVC8SEWWSgHdNgoV0zv1qkmcHCJDDtfZ7XPLTjG0++gTnBUXVypdRces32lpeN
16rzasMeanOBVvhKNopBfuUHyL7U83F2IUWz6aMR6lnjwEGZgr6lj3QtZQeEFb6k
FQ+X9DHaC1350ixcgDbqFjtLEGOu9AnLUN4sP5UNuyxmIMx7lYwQJ8cFcg6+eSw2
g21ASSfnxOmdxNbUevwSP5e70OYKsRuslwtUMzSCwAucgnQEc2LWEenokZ61rkZx
YVwTm78lWjCN7bLBlqanUc8GVARX+WUm9ItO+UWKo6fv7O8uf5hHuirfDWO3ad9b
drEByIYjcs4JlEdufm8ZzNLpotsJPgOKPAJawQGncla6AzdhUFP2Yh7HU6mfTt5/
DsgpVkX/M12TiBu/2MAx0aAMErAxwN7KL7gD5GhLwtR87bhxBZNUFwCxRa8fk6wo
I4G3AcyoXrLs+LYnGtZbGojj3ED5Kh3S7Yyw7XloOcPDlMIJ7GaWDgxix748+vu9
2k60d0feTf6aYWcJuKivchtD5lM9glFoRQQFGhnfDGArge2gnhQ8DXnq9xvYjFID
72CUGHta/YU8aveY9ho158YAxiHzX8Y2Ukg9LIeZYcx/2hy33PVjtMkm3u1dHRIW
iIYSlxZhkrQ42/JTIh5ewv93RQFEjMjezOm7tnePSxj1rpgkkytVvkQqWyeSoFEL
SQCtFz4nW5SwEsqS2cX4OZRjQdUiuiv7A7WAk1r4qK9p8yqbRFOMj2ixuhJsLTth
0tl4zp4KcNe2rXr4OqwLdNZHnQ96oL8x0WC2MjgShBWJw2PL4OvQf333U6bcUL0x
TxRh3ACOvXCdRExQM6+9qQZVn6srBiZNySwH7MdH4R6pmzKbKgf+IUrwLVp4EJ/Y
aR7vLTSc0gAInbZAp0izEfw95OiihT4mg/bJPNfP6vg6s/+nr0dCVh3cD/CqOSlw
bm9sMGud7+BxgzCR14cFIqq1NZNqCDm4Lsdx7f0OyvP2mapr6uE8uzlrqRMt/9oC
rOktSCaM2DlT0Y2RxWH31hD9+4tofSez6r3AmWNTvGsGiM+ZiYLa5P925+lyIAvG
CwxtPGetfX7mp/7Pxgr8VC6QX6oi7ntcTCYQEf8ZzhFjRIiCUIhU8AqqWLLNi6ff
`protect END_PROTECTED
