`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fF3phaBhrIgbh+DyYJiqhui8NgFmuLnCjkT/nEQX1dwS4sBf2PvTFZ8R8WLJCIZ7
AMSoAkrf4bLFf+7sfWAUYLSXsXRlLp36LFJRtg9CceKapLetPiODcYp5rIYmA0xx
ob9mHbzZNy1QHHQAob9NM55ByE91oZIX10N0nJ6sUvOEqg+H+EDpf/lXARaD32l7
JiBU+UbkcVFxRH2KgLCitJys4deBcNjOG71AC8AHhQJ0oaXgX+kN3yPPK2Sxj4jL
2j0I9Dm4IJWZpLAetxtVMJvNEkqa0jZuuXrmhB8g9Ucp9dBL2ELM/SrvgNj9UN2F
j3eK2iT6hHv6efJLDab5lQcDKmejHWkZqVbKccCYWBmRpnMwSNoTZXhk21pN71Jr
c6GaJFfwm7ROKMA6MA8eiQxFJuflUu/NsUkkC6P+/ScqE+Q9QwRstYmY9UY/Igau
Cy1PfpWWOeeMKwkV3Fv9eOBPD9lW/WjlAP6Sl6vvMfCUoYlNGLGMKnMWMp38ZQN0
ER+Mjb0CkbbYC1O9cwKXJutmnhoX7ka1mEd1s1Ed3LCrcmFUoVTCOIfW8ba8HHbC
I/AjPOpI5LGa4zYpSurin4kszDB0naGbG2IyQdZ8RxCpiYKfMv6pplq0GR7XQqhW
ldrANtsbsWTHYBr+Wo9skNwgK/TQXS//8GWZ6oFBhxPb4Sq/SvLtdcG+a+m6CONm
D51lFohpXCDAExS2Qrjfbi6mNSUyK43z1QK7YRq6ZbkvzkLSjFZ4S/1hYN/5PGUY
ah/m+MQPVLE5EB6xMOOF9a2wv4X/zJpa5ircHyLxK7c6Gj0rL7B5dC31YM6HgCrw
OW0wt0bbMK5h9OOwI95xUJY3jkec34Ep6wfoiqNNpZm3qtmd2Totkk8j87kNC8jt
ry3XeZSnEMajpErK8DuLs5nZp5YhhXHp1NcIyibckbmVM2M+RwWLOqZNnO2V7Hwa
`protect END_PROTECTED
