`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yWoXK9MA25MlI6Gq+L5kjs1UwTgZ4Uo/my8GedqgRdg94RF6Ii4vJwpgFaixatJ4
xV5rsK/QwhQY39FsKBh8LxQrPhj9qS9P62Z/m7z7ywA/tZUtrzPPqc+QL5GyeqFH
90AkUSNn49hqniWGP3pBzfRPRCXrijGVo7Lert3SzFkq7lkgCMN53GbY23EX3Xpe
OWEp6q615a3PEFc4UX1WcJMUzJyqYme5v4TffCSa6U7xwZ5As/6vFRg1jloTXWom
aPM9+zxawl4UNWwy3X6g8W+EpJzNLvlNdtGZFOz85dCZiu5IwIFclCuuJe0N57Rp
qOeHCfNdQutjoS50BqeIMA==
`protect END_PROTECTED
