`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tFtHUSLI2za0YTxsnZ54GQNaiJTXHu7it3kv9bu15o9GqLXCiv8EUesuRX49/MHi
3lrL5nU5ONNovKiM9vMnfQan80VK4H7CYPysdYGuRzulkUNTRAMYoUCL1mTuCWNm
ulPU/GSyaG7u4h88nePotxq0xtgskpBzhTyz9Njp0K96y5xyz4bnyX1ulPPn8Mt7
bEB5h7B794gD3lltczFTC1a/RLZXlDlvp/CK71U1KqMWZvSoGBzgiBQhb7YTh2ZA
laTWpZjKvIRrkXy7LnjMw1EWKpN2p2M8cNzNhCXbuT0L2Uito+E84c3fr7O24Uu1
n6be1e2Aj5RVPT2UbywImj3fwK17yUee/7L6VTdjDFTOZk8O0RWYqb8KVr86D6zp
iWYcAUfdXV6o6FIqHd4Dl/IpYr6yKzWC9bYxqwbm3xFhM6SZF9eazW7mdQe7scfV
dBjR/TMaBJeWU+iNq0EfqqyC5bL4eiJKzY7zeAl5MI3of7x8a8ZXevR9Sa5qT6id
GSfH8gY1TNbJDFlASvcA7WyqcQYv4XL/HUWdsigVd4cLmv+JFCvucRQOHh1vtQ0R
SwQaL0XwxHyxnCI8jRZkH7pRU7YxWfByWNVZHMQIQxV+yAvA58yrA7Q7srlU7iq4
guX+xDPDQZgEDvGFhthDl7kqFHKlPmBM4noDFv5Z6UeUDXksJ6AkpNcn1XbuFYuI
J+sgwh9nlEembC2XxxxZC970n8SThZT9wtVP/WsDu+u5J3wVRmt03ZSsNSi5u6vG
sqtkkaN3wJOOps7GMR48Gnyt+Gta1hXhbNbnHAIp9LgB+HuqXWCvoiLCzPcujffb
hlDbUXMV9aJjijSeZ/K9+kw2yHMXDPuxhuyxD/9o5Ye5mStMBoJ4B4tY+Ql5mhly
lMfPietyUUWCBeQTQfKEpqZTkJZo3ZH4iZ12vruJmXjUteuKTS4Dp6dJwT+2juKR
Zkou7CavJV5+M47PylwFG4NL2+NNJG00UiNuNQ/yP6gqY5SNhULkh4EfuHKyE5ct
U3NKg2lHmjBdwWTH0U8e3B53rsdVXVLkmSahmw56D10rA6ipygO9SdtK6jnaMZKh
ynl22EAcrs9vG94TueWhPEz5iPbXBNUI4EmB31NO14riqysVkXj0wXjWUMiNR/Vr
7H5JCwijiJNnqxrHuv8qfXf29hJUm3be+CO1+QYbkKmlTPTYYk4EBqa2Q2Bzy5Hb
QOt/KKVvPnLRY5pqHaxbOJryUbE6t5vogJ4CBBBn//mZD2z5FvZIjANFHKWr3q1g
Bcctm6uhUXED7Rc3eI73Q9lOC0RY1vv1mPFBJd3kwj8ZqsVVhtAlncKV5ShPQSu8
1JjUrApy+snbxNR35tu7D4/lnVXf3K+G/KrQ2Lxbsh23LVtlqXgsjKOQFFSZeqN/
kipt/AtpaZVDM8hyoLxSKPIrh2Eb1fPqd1FigYqbiwN0enNdMPiLZoBzqZj9MCqF
kjeSpsLkzo83c4g11IrtiX83Yc49W7ur3/FGL0YoY7ns/tScE+FidTGMDA4xsBj5
vvck7cdxg6Hyuzu1X2cD7ZKHGB75e16nemuKv9DnfeNENJLY/JOWbyfpZo6wAK+B
A2ZwJWm1OHFqk/oXvesfHDgqnEFn5HBOdb5wnsGb7o0Xf+kOrL/8/Mz2tCTfliTT
GgJyaOE4sdxCe03kAoAILrff1gs8/Zvpucq0+UCkglvusa4Fulcsnt2WSqKOl/OF
NEPgFIJs8gCBIDf4vjjlZuK1HoG1KJzdudWuTpdsDk15W+TPa0fwDOLCh+5oUVp3
rxE+FViqxf3Xh1gcISb4Y8MWjQ+a+hc/QGhJP57kXcvOQPzYg0H3c/NyiyYCKrbW
sNBkQBQEgy9Uwkr67YsuD0Tep3sMxbl+x6BqdnUJx8cgdzs399YzYQ1UgDb+2B2i
YBbZtnazBYpbZJ+NaqGSzqiTnbVmrX58huTSqcufitiEMh6wjBl/jIzAlqDK9vaG
8SKEgvQys2YIctE6WfU9L2Zwimk7wGRztpCl1T9cIU1R1IaNsQd8nkqPahpr8rRg
uIRCN5O11cXhDxntpydL3DamLlatlSUExxCWHBQGo4a390AVkdWcOZiEKg9Cxq2K
MGy9IqhXkVqe12Hl8vmoZjBAwx/JHAxBn2zOQG1CKkDPHgZ9bOlW/pDkGL2eDvLh
Z94WXBtBt7N+mcJQ3Ib9E5LPL4RsC/XCmlH2CeI/LCxFfHVQ68A6m6rU2Xufus6t
ctZWid+h4yfbxTtA9AUlFpdrEFkYchdXlDMN4IvBdxlSZfvytHePDx+qGfGYOWct
wEINw0rTDjKpvvRXmTZegLLbk181Jo9mEbUOH4nSNblZl24pmofoSfAo0oz2dwhG
aw6txpykD/FGmI+mI3+Ztc6jV/+Uzs8WD7ryPSaZviWMVvm/EH1P3WG6RTvybjUd
sqDePBCOJoSK94AuUTpIRP2kKfyU7Zg3F6enuVBdRvigfXq2kk4ikHqi23mr95cW
pDJI3NvOf6zFRVoes5XZnzzOZTMrOP4ARDFDyAtmPqXjUI6c4nXVREIAX5uEI1ks
jFb7u0uZ7ufnrvT3+N5afcteu11m0UIcbCIcrtuDYYnwXyJ/s+C5sukDZU7nT/Zy
BE+Ljz/XfMk6UORUgPTJLDYE3bkxYbUpqhUA6uNj/vQUiPO5YjOLdwOzGN6iDcxW
B/klAXOs1qv0ytsQjBrKZUn9+ffFkWrowVQH0Ss229bpG5YuVDYGCdYeW+wPZISc
/U3O5AokzEkCuJJiN5nj36s+aB/lLTNGufLg7iXmlXXaU7LlZ+IgowsiZvLrhLt5
JVsEg8vQfoatnVCEVTm/MSdg39czozt0npRRwdJV5Pna4fnZ8Zeg5DgAN3PE3YQO
+a86eFxXSGKCyq107IrvqUKzJbz8pwo/rVfl1ISuqzLcgwcIhK8Hs8TmNAd2QGem
4N73P41OrQEjKOqGtQdDZfJdjn1BvmZpaze7TTjUoC21pqYtl9g4clDi5ezcinTI
iKJhnhKxVrXxCaz5116HyCnHe8xwAXgAf00JXD5EEFUm+MFz6S0e5T/6dzF/w85T
EAx9HW0E/TYjtnQPaj+XkCZAdLlcpJ1g2kUydEnDZBMMd7D2jDH4ka3fJw6Rkede
upcsOwj0LcSms/A7vf8Rr2pAVol5teqUoXii7qI6Z1t5P0z8OvaxfsJhrfdHejn3
07UorGaVBwJV9+UIGEnyKwXYt8RWXZzG6VGPtDzvMXz6LxbtL55yguB2/BhhfP7g
PCAwSZrGKrjHr6/ZWw/CpnSNttx553Ig8YCW2h7gwwmlLyZ+dz09i78eWd3LyPMj
tZETwPejKzaBsDGnTrZ2t54Y0x1bVHAYPqKPX+tylRclFwFTQXKuwyfvlErd2hfE
z+27sB3cxUW1KMqrBldzUVG3vfyUIBJKFnMJvwIGUziwhmne1t7iT9N8A9dordhq
w0JVvGJ5JP/L/Mqadtje/eSn9yc9wzSILFxTWDHKPglY8FaGBmHQtUCu/xScDB5H
2FEmqM33Ur0ng7eA9rVV/e063Fi429vEjOJjopYxDIQP0AZ6sh0Iaivv7nyqg4TO
zlF6b3awLrGbm2zc/Takq2ofeovll7yCSl24bh3U3C04PHWq4YVHdJjybWBHsm8G
v4bo6Y4gloQNXJ0mMcNf+hxr30ZcYbgqUTFg9muuEEM+Ran0lD6pvDbfRBwDNiwB
0KXpVTBCGjLJqbkjvU7vJBT4jsUVqE/bHDtCW1re1Tvdg2glDjn7EA0ivqv+Qb8K
c0tHeQ+T+8w1kxU72M6DzaHdQ8CIE1tw6NijU8s9qmV/9fZxyizs7Hu5F1F4UwME
oYrh1eYUy3LOi6Fg0q+VgLqEfU/AOwA9+GPJqFbxFzTaHbPs9B5u1r/SKpQbvYNi
Bib0fIBseBm7q1/qa3XcCo//DfT/dMQ09q6FLrlNgWmidEyKED4mD0S1mXAidZq4
4yYsWuw+nftjmE1A0SYT8RFm+itEKoKcK9hr3vSgyxXWCO+6JYttkpdsxq8uMFL6
22vvzKSgOm8WntNfduBsrJ28azeq0VtzuZpZcTf+XyvPxp03EFUXzAuJF/hKfJ5m
gXqbpVRSF2rpya9wCbu+39C64OVNOnN81ijZrhkuq9qk/QXv2H/2TNa7cBHI3Biy
MvV6Td3ZsJQpNLoZmJzSBsmZw4sh3LO+iKKc3HapWiW0quX88MkDfb+aSgjkMqG5
RC83pUxVGz8X+ymYC2eHBjCFOQQ3VcjYeTQ3iI9uKfaNpR1PmGbgRH7oA7zj8hSp
d/YCZJUErQ8b3S3i+0VyslZiYrJ/KcDMttG8mL5PLBDDU7EuhhmPi47sVIRZk4bK
uvK6Av2UgltPGrwXC7ltCo6vxdbmjqdTiGmrFj0mw4QIeYNKTCuJCzCLPcqR1NNH
chCl50ru8XsQPdI/tqdxcqatW5sPyQI83hPMPDM/2flHlDYRtS5BbI7O1Ccu/M9b
uKtT/tte8ubMXzP+wGlHwmHk0K04H1xRs2zNl/TpRR6lbILIyvi8IbvQs8PVWrx4
4RXOilNZCv6hGIZBDUYSdlpsAxTGVagi6GIKKvC/fhxKle4Ir3phDaIW+hVqyqgo
sbT3wjxPetOYxaceSpehpIKSGG3JplqdTQPhn+RS3hh8lhuE7RLjK7xVyNtZIbCk
sErysGednn7KNGW4VUhPFqjUoxjyCATnWzPpZWTt6vfKHGIEv4960t0CSB5o70Vl
SaOy9oqtd6Tq5q2XH9nwLPZkbISOVOvfIm9dbTKNDzzJhbFVl+1rEO8wY7kAsaUD
q5Zd99wf1kRx2JHNEiU6p8zrfU259QUm8wBCULhTX5lnv8kyWXALRbJbPnnY1u5J
O9vC+JBmRODjpIka7TJ4aET64Gq0wIJSJ9GFJFGAcgISpgAgmTKQgVjIEUfyer6B
n6SYY30Vhm6szcWYF8hE1ET/LKwBZSpjasgQB0m9LJYIOBrATfGgXzv0QpCyLaMD
3xyIWtG0hLoVgUK8x+hamieVjrE1i+DbU4N44AH11+FRs7AC/oDYOxx04WWmrily
3+WMoFpW7vyBBoGlBMDFy0kJ7+5CROEKuaSuvNAba/qfkFOuLdFBDP+UlmmJljI8
uzgjgg/ZizMEgp6xX0EUeb0oqIPdpwksBlM8Fkcv6gjjhIY8nTNKW5lpJNTrqj24
W7x9RamTmUFdWncqf64cwG/JIIxFpdjUyWG2Tej5T+KQZnAMn6zrWKJpEGJ3CfsK
EOnWChk4MaX/aml78b3R83xnYYc/YeEaKi+O+R2G4Y1lebzujnx4n8ENrCBL+wjl
TbedyxwmHSi5I7fTRtaaVpuu4Ntf05ytG467eGNkeujOuP/ZGipb/LcSB3lATS3r
Ethx/x69ZNKYe11KaPaErhTYlTsfitzlB4CYdvtE2g2mXpAMalOw89zWHAQsOuPg
xLuEYIZwus2KsYn7cJnpQyMBeGc/D5b2FkWGfeZ4kG75nOi25oaeTHIw4QmRZ7OE
aIGctx+WWvqU/ldbMTaznCPLscN5XkzabiJq/kxdi//+0CPUy5rQQ50xxOp7x4m2
LNqWMBM41psiSsS5Za8D8b2F+6+OXvKS4D3XdrtP39JVwwt5ZGza1ohuBC3Y1XjL
k12JLrsk0eftIafSFfDJMRAh9WJqAiCSgg6GaPA7X8Uqsm4qHgKAnh/A47HZliYY
yH9PinVh2yMjqqcEtHbHx/KrBIpHycFD6DJE5bSOIx+0ffUHb69Mmwex3n3gyenx
sRzDjtqur7vpPot4xvcRruHsB/cdlyLnsiy7c2mnUvaJLrsXMdhxwUIiODwa65s4
azsaRylqAJlkCSHzetXYZo/TlEKNCaz7a6D2wNFkgTD3nZd7qfTQz1Ao7kd5kTNC
TffsSKHTrIMMO0+HDPudzeQGWuXWlImOs2u+12rehOyjQn0x2aWCJ+T2cA3X9tu5
mjc6GY7a/t1+TyPrpdHcgxb9DubqSY+lihRn73tf+o45ZWbOTBmQ8w7ovBT1fGh3
3SjunfO5pE9BdyQspw47ks9yKoQjoegUXpQPFG9agig4aHOON7o8skK+qKMdhxS4
RruIM5abLepGtzZlkROiMmm4S8eKWQk89wrQE5s2/whN0OhHhA5ok94Xfuu9uXnD
VOwpnSpk1YjgNmFFG6u/VdH7nrTdSI2OEv78lCqX33rbkebIUOXcmKDxHL318cxC
PUj7ZgWBnebjtbNqKOzeYZrWoDjAZ6iIXYMqFxNWgO8bhCPaBbtgRcb8pwJFAkiz
jv1J8J8fBPaK2GYkEFKwA0PmoFiSfpk/tyV7xtMxA4w/PvhOII/PClhClh/t+/t0
o1U33ydbyVcyVio6nCFmurrxGdCJU5anpE6BE2TD9R251pnszYEymAxtUXedzFkM
KwwDVn3hp86VGI8RJ6d5ioRBKWdkv2E25wlpJIYdbcHaPC0/NScRYlT3aTQOdf6b
F4pLbLnEbkqD+hxw/7vLZDeqD9ZQdjd9VMu+w0btcyQgr8odapkyil3MTQM9dyXW
n3blgDi5Ojk69779ygNj5VjhxqIBHyXJ6NTBwsO1zTUdP35VxrWBKz1oogpCP765
6y++3ctlfaV8+VBO9qwVTghTiVdXkcuGD4bob5mv/vWrgSj39VB0ZeyXHgzIHzlK
48lQ+MlFGcuEpLaMXdEonCw/Apg9akzJ4f+0S62IQsokN8CtJPMrIXSC9DCkUuk7
T6ZYRC21lH/c1yjN/q+s3XS3GocLtH6hkSWvgKZqrTFVQ4OqH48Ypa+2ITTk4zOR
YUaQMYymByjaS84uMCMnVWD+HP/dX/gw37/haiHWMfZBvUxfXkk389f8EfNLt4JJ
FWPaA3G4fds1nf1OY7pU1w6Du8VfyahFJoK7+zCOCD+IWllAke8q9Qw0MVlpBqC0
6tgglOGbpuxGiqkZLH547A==
`protect END_PROTECTED
