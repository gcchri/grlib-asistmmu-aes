`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z6hqvMS8q2+yjlcx3KFb/rPAYBMilu2qw67cd9VIavXyEFUYpLi4OZlCvJWKYGFS
dqPPaKHyAoZFppwmEHevpV7mxghTipx2BdPs2Oa6O5s6VTOghQdGUyu4MdPfGEfo
1CbusdzdPfc887GGTmt8csccWgiIDQt6HHd7MXG3NI1cuQoD26UiyJJ4b/izbncp
bstTxS9kJjs5ZRy7TVU/RckVJZAGuEQMBRuXZx5HBXKZCpN80ioDR0JqRFJF8JJe
ncFZncIrJKCmckC0xy/DtLmY4X3YAsTSCjKik38cMGDBUnI2zhZJvACza2gkKl9G
iFoYzvU5KQw/7dnmT78b2/lbpoLqzcfmifLMEMQD2EEnaj8dYlXUtjM1UGISU/7B
bXRSNL8hsnUTMn4LHNOhE0ELWVHd4hEtvo1TZQ/XF7W/K1mrofkz5NgEtQP1r8Li
v48l7HxucQvRAWHpeeFNox/2v8EYOIJ2aks/7CXFxiNwPkCilCrCOZbvMRYMBgTr
RNv//cXj5eBVhYVQNTuMkuQCyzDaQ4Os8Yzr592ghG7WRuIpvrjkVLRRIHoMaYT+
`protect END_PROTECTED
