`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VmYJFCRgQiTk7G3qRvn9J+jCTzmTuOKjW98nQS/aypM/XPCwMeTVqiaY3UyShCcM
FfPo0oxsN6QRs8I/Kr64OAYFveloQbl7r8AGKzpear/tlhZUVHBWk46fm/yy6Sxr
3VnefdUvd0TdoN3CKupa7guxt0aZ7p90MHG2Dqt+/lCCGd4+li6Ew5KZdbOy4TFI
vwEQELWat7GpGVij6/oF6C8lpP5BipKTx8/rvfUXROnFEP2CPS6oZtQmE2w3NQ/F
vA72MslfDQFBL/w4lelK08UBgd7ya5lZZtdjCwheRvo88Lh8w/OiA1TAjflekOzE
SzJB4MFdYprC4iTB4EBn1wzUTgGqa9/J7cpzmib376Mg76H1b4p5f+JFn9AjKtTf
OErj3bKl0tasTQzNPqChw1IU1EtndAvAnMMXDe86C6iCERzo586jq0WtnTlnauMb
C/ciYH5RtLQaE2DKq/TDDE4tnTNMVmbq6Ry3bShTH+qCqF8iXY16WApAn4F0+tAE
XT7YV5wCV15AcPFCLWFB5984mvvrvdrHGiuVxPO67sdV9/bbFEVDxDN2HzIgnLlj
tFi0s7L/anN193Eegd13mBxcc+Q/C5gF1Gx6TSTa25KM7/LlrEzWUmuJpn8PTPza
w9Y9HVKX94ovpzO3uv8xLQv2PN/DpLk//jGrxo6RAGNwQmMzW4veVPNS739hYR5d
7a2tLi9GioeEJyMyFajL+1lANh9XGvurO9FB4fHVZ3+h6iE/I5skKl5+cO0cBMPE
awYdWoRQf6SiZ3JBAzlYu3QXSmur8gVxjClQ+Gii34/spd2x+vhj1vBzEJdGuqLN
x/h8/KJpkw/GsUWN1h4OpmZuImH8sQYh2nn9I1AjMjAGKejJgKaZYOtbTB54III2
Et4V7iHB34+sJO1M7t1wrL6vhV+/mOLmLxohtsA8SWL+xCxm5wc5nqh0nyQrrLLj
OT0KXQzqNgkUU4w+bbryI67hvYUCnxPwZlGUbe72Mtc+eF64E8PC3IPkMGMB2LE2
I1aUPneZlEzYErPX2DyHyH7fy+IB8wYcLM0YQudQPQwPvNjMongzhd+YZ8EuNfgu
QY8TpzwV+2dXpbDsheAnOjGqUlo4BkdK2sxiD+F3ZfCaUtmEr/wZ5jRU+MYt+s4X
3NCrGcn5b5feUpemKek9CW+XhPgTFHRWvJuYE6f806H5P4LX15xnzZ4UHu323Vx/
6Rc6b2kHH5w15lhXeuY0SyOSuSe3/Bkmby05xF5H2wqQ1VSIPofpzpEDPp5hTOv/
fDuY4wPX1A07dwOSaKDAPN0z6k4oRtAG5CIhWOa7NNR1Cmk49b11SFd09XE20SLZ
5+qqlMIafonzg5QR+1MWqc43IGDT4E6qwHz9QlK707PHRi3zeSFYgkBa08lE6K19
bMNzfZuEn0x8NxAQVB1C0uvchRM9W1XUnHimxAA2FuhtIxUjy9NZaEhSq8VM6llx
Mf5md3jyixvQ4j2RmGzH55eZCtPIU7nuFhLjiPKBdO4SY35HPsgXYnMiSRKEJ2sH
jef9jFoth+NDG7TNTYvubNyIzwonAUw9Pbpbhr9n/HOJRSpBGnsbDLInONnUkdGr
XmErmhnhEyNonWoNjCVeJ234HX/1FCM2qO/n66aew7H7oubYI6H3SXHMO6oBpGRT
FnaZ8CTvyUCO0Lrra4H9oLf0+11nAuqc8ysc87fLN0d9ExhNuk0ItPFZ2XLQjDXn
6eoi9q1wgKGLWGkm7hHZiEjgLJj0P1gJPAzHWRlrBR955vFOiM85xNj7kOh2oHJW
Y6qdFzCGxyB8zIIuN52kyeL22PmLvnjxbZjzflOVBbtvQ9vFLarOJwCsOULs3np9
aYMJXofLfBAgJy2m5IUe9wO92zkGAW+K/cxAWTEwSs9U7OYhibNdLXvsFtR8QKcR
//HjRnXxcNQZjGpEV1+mM8VNSgPxajuRjPndUm8x+vvdqX8WTQAAP1+3PJ0Lmo3M
LXbpBR0PV+QUUm041thlNXY+d/1thDS3DhNJ/ZjqmxXa9N9y7DRTmn7BhY+Xxn7w
zXx0xpVTiZWdRk4nFVc3GuLDksm8zccAWuDlQc8tVDvGiwa8etezshnGV0n5L0oK
Tct5CoYP7pcyB/1bFsbdG7e0LBMjPup2FFms9mIrtTzNXzB4BRXyCzsbPHZ/WhsV
P79WmgYE1m5qhDLBgS45tO3tugNuCgHDTyXvz3ZlOO7etyOmZF1fPNVhWrecWyRo
fjoE75GCMNQS2yWUTIgGaTMLyebB24gPSMeE8bZFv08DBccpmYlQkTUTp6dNkNls
2au1+SggJfHntm7XNY8dGcEHrLhfe512hdtAKk/s+uDCVBPZI7Y5lhM/o+9cHoYI
KG60bPFHJVpFb9idWIDpJWG90attMdeCoBywZf3/kNdYBQ4zsM4pqPWLo7zM6ooO
tYxSsdP6fez51VimCprkMP4XSjNg8Q08UpPJR8n8sbg5m7GEUumAij88sF14K6Z/
8Cd96lCx0y3y7W//MWkYt9PNSNGvzSGwz+AhMQLDL7QyXTB7LIFRp1+vJbPOe2+b
6OGRf+NCcnSjm/u9K/TEl0ukHehYEQgMBB6B115PZUwED1WpIUMCIlvrU7+5+vOL
IwThwVD0y74GZibmjFfCow==
`protect END_PROTECTED
