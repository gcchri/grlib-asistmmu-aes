`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZdvRTZ86eeLOh/dB0m19toN8GDqYC4e3rwso2zNwx3I4RbVk9JiiJ637lwntKMkB
axLJB/JhT2cuLV8iV33s/A/kkmeRzgCZHNXarp4eJOceCwj7+9iVg9M/QiMFWIHu
Jz+XxQyo+VeLPXwxKhzoOQ6Ohjer3Ieh3S3rR5QLk/JOTlpreI9J4U4oo2VYrgk7
O8053HcCsKaU/1ioLjyUKJLYoQZ+66OubwV1d7FGFurAsq5iqDnAE5/qDYzDLjJi
Jc02x2IhgBG5Fp1psAXWgqeNCmFn1Ag+zqR8GZgf/xnpdEvcqTPZ7+1rAYc8kTz0
vwWeYzOutajAkZ8deV3s2l4XSqbDSuj0LT9E2RSh8j5Ms+CrcTTZCaNhuRLN4/ZB
FVCdl10amyy3YfTM1VquohEcETV3acIcwEWonYGnjDg=
`protect END_PROTECTED
