`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uqQ2t/7nvx3U6nuoBlTiftn5a9tG6lp6UpnlQO3Wd6HgyBy52RxnSLEhPbmqu0hY
tE1gAgCfnpzbEjfcn8IUdiCbFZ+zieNGIIs4epLGFXZQuEMZyQIjAGG4pjSZNYR3
qrnhdgSfNleg+WFctbb2/SjCA7h2MDH06fkBbYmqlUjNpX5qvoBgIj0PAghYv1zb
T46EWUBFHfcRiD1qyqZfKoTY3IrzZeujQ5dumoPvQHVINynm/waejQxHpVyD7Z0A
io/Gqte6dC9jYzpwB08nUEiSTzD07mvZV5LCbGW+SOA7oZN9MM3UtwGtTvtBd5Xb
c/mSkMmiab5jP0hO7HRhQpY9WKKkmtGKuEGTnJsoLVTd5RNqk2IbyyHmJmuJ/s/E
aTZIwRoayEdDVdzx99HOVjjUJgEqhROup1WADc8Bw3CH9/P0GrRjt0uHdchJ5Wnj
FgM+1LN/pK8HgKqZhNH8x2q+BR8okkagg2exSxO0/qoluVloOl1hcYMYVncUpB1C
aDqN7EO/2R06nzFJetXvPslvyokZvRL/5OSffIH9FbqXGl2af1G1gY71w1ZtXeGg
h93tX6ff338xiUuxonYFe/c7NpIORjNGDmUTIGO6wKgqjCepMxVj/7Vy/K5vDq/9
`protect END_PROTECTED
