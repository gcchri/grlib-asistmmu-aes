`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y0tuLyEmvpeXwidbuWmkxVUqs53/txxa0h+J1FfWRwPW0aeHEpbFT2artvD4fwC0
SmTgqgQ1q9E9nqHmGfFZQcby3w0xYvgW5sCe5NgX1qxLrvfA6A1surxVdzqW//jm
GQwMRXeqGbPskXT6hcpC8S5Z29IAPzxZCWasUtkcs2e84rs9wFhKhosgq7oNtprc
tXLRE3GvlX95RJ4SL5R618miZ17VRVeX42m79TqbmMGY3Dw1Ecu325C0I6hx79xw
uM9h9OReNZOmlbz/yknaYHLGlltC0jzTAgYXBP7MpXbU47V40RjAv1PBIY6drYEu
+QXpfES19NA0Pho+ZGeKyOiNaBO7Sk4YinWGO1bs5B8+syxgfIH9kxSmKO7QR4Gr
4Zu10QqspKbYu4rtl/Q4P6FFip4NErKiVbn1+lMg+BO/RPkWHF2MWmsw6kDy7Rxz
wwpvWzQ+5KShZDqD/zYSORuG3CSXgVD0V4yl+Klio8QbJwVQ6hwN7s6HMvl1QBbK
V0HdZ0/OZ6ZzAPpTjwL/MXm3ywrWl5bMxgWzbO87ZykmNlXY4I0opa6rRwcpxO1K
QIXq24+64h3toNh7i48pRS6WnXWfzRChCdjbknDgwrjo9EusRdJAcM8KpLgZSTBA
VXdPEEhx+B9dTilBM39sTshhX+XigogcgkR6v/ITBsU7EoP2wWEqSIbrGBk0OMzX
whzDWc5ck3SyhPbS8xkNHeDx9Teb1B3Wn2Jhlef5dwr3+4Iw1H34OkB2mcxP/ZTG
l58V2+f3NJlFDDi5deIOz6Z6S6m/3Ov3hE2wS4yrZm9Z5bOXwEPpim4U3/F0SQw+
BJycfLQf73DWaJSIvmdI0fdzVAdt0yoQneAdfOyqqfpd92dy3GvM+rV+g0f+6aLv
xOvN8/2gG+vZkP3CRwSI3tgjjZzSYb/sQx6uhjJyS+7JanZUNipul0NQKB3XW2Q7
jamNSPW3FMAfAT8FiGqqmHGn5Va9Zf78ay0suqSZXP6XTEoLM7FWVolezITujWko
4JIzerM+1/jDgCAO2LwKtnR84YXoap4MDfx65IKeIz4sqfE4+vhBdmhhThP7XRvF
F9YugkvK5IKHCx1UgewoMlBTntMlNYE0O7PyuDz3fyp616i9uPjHUCIJ6Z5Zu9sK
fnVh7sZ3LcQHsGUuy+2fvx2LAT1m0ndq68lOeo0+s1fmV2Lhc/NlVTgd/gfe2ygm
JFVRr4QW+dgdQ/X1I/H2EQekIyXrCzCeXwxS5OlKisQI8K9wg1nVKvJuKkmQIVdh
uXnAUaZD3BzqQbXzvi7u7gCcvJbk5rPO+zn7YC4PgRORbTvbAvTbf8M1V9upgEC0
Ljjvme9Coq6BeCKWnA1WAglm97dR1lov8CJltZLADAW8O7CSN745kRWX+P025hIn
IooGyN+tN1e8t4kLQryjSUBpmt6oWWoJ1oasqQRkV0tUklET3gFBdGENKZ8PmrHi
h1y1o7zfxcKLsCctWVZqwCe1WGJaAootPDki7OH+KcziPQNbYLicEoFLVEOlVH18
XBQjRitg2k/YvwCfG6WmkunJGtwI+SvL81Ma7bX2A5jepqQpjaB4Teh9y27jtInM
m/rDGp1WjaMLmGAT0Bhj6RtmMXnfsmn2uzvu0SYjCH5y/slu8fqncIcO4YiOY86e
zCBZIkjdaJUpR5ubWTQn8JZCBedsu+B9ced+mghBIyHM1VwD/x4+h/smLDULHMwe
3wxwhKneSkhIICvhtS5+EbpuG20965F4ltAz/IxyKp52rOGrQA/eUzBjcRQrbxOz
9YXNDeltMZM7cSfecjWtGdK7PE5GjsR1/FZQyrXF/RM3idKon1wJlidG3AFnCGPF
r+nUsnbrxyAAUpFjDEGdwKlC+UHeKS4GUyKOJPzYt9M=
`protect END_PROTECTED
