`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
03sDGdluK4r/8oTEdLjDknPn3FXe8DaK/tw1uP8uOPxDnClZBQCLDdWtl8dnl1Oo
80dcNcAj1wfEDzn/jU3K4qf4m2PmCbck6XUIAKUYh1g1jzhBaBg0ki3mbx9yZIqy
pTpSIu1C+stU2xPuCsWbW5wZAA2MPAt2qzSC8WQDBwyLESn9EHL1ZZBp+1KAmt3B
GQWterhi7YL6Y7CYwa0ndBQx6dO6BLgABTQ6h3VDDvydI/aTE48Mh4Tp2wQYQ75E
2RWAjFC9mYF0dqQ3d/iRKHh75mM/f1jhQcAgkiUaKQiySokO9AHX55ZTmdY0ca5J
TAJnQ0Sj++kWV4X+ScIHfIylZWhK8gnYyiPO4UveHdjwT6uv/7DaWVPUVPwP3sKD
+DmfBrJ6VDcE5zHBkDQti1QNg6ANuBGkcUqfIRwQ7VU=
`protect END_PROTECTED
