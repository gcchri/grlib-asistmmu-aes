`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GkIADu/vRGU0zbIm3d2BmGjWqnQ4t9q+cWJ+svg3x+C2Kp8FO+xec9kGTdtlr53j
8nBvnpSOrrkUyk5/GzKCYcJfCjT5D2+wB3hhXFOxozfSmiKxqA6FzSsdOV4s8mfs
WMaJd0jmU44kZTHxFf7o8S1SAvpeewM8Z27H2k28qWsNS0BbACHkpKFmeQ+iHFEl
iWsk74+w+yGeSY8xcKl2gZlKVbDqk+sYAz4EfEld3cjgtVLQkp7unvQmes652sBF
V8yoC/mmr/7z0wSXD9M6K1zXvC+29MDQCE7TXVeJYoFebeK2cAgPeYA3Fa0kyHfP
CMVVQ0TWDx3Eh7XTZJjSrWBNhsij2zJgs/qyaapD/bFCSaNsam7WbLYUIHjUPM1Z
NWo5WS0hUWVZnjx91wrBxljOzMoubzWd8xWSuEMlgUy/Y7WolABNn+XAhM89Bf/G
un7ExPLTceSzk45fNMaS4aedV0XYIBbHVQ8gNEmJDRuOANC/Tar/3iDYXpPcAoUW
+bc/QA9j2YZdj6haNSC4dfwUSe3h1sgK64OBG119kXRhqmIxB84E8SxWzwBJlnQx
MMXFQVs/GRL9A3lChBflr9NbsQdYUmgaV0hiqIeda5uw48g4MZfn4yjxat8Qmk6O
Y3XP1XBIPUD7ApmcWpUGzFCqqzisWBrF0BWIasBhGHrLRIy+U/l6bxLYVsslHbSk
mNGzdidw9gZ2ViHquJLtkg==
`protect END_PROTECTED
