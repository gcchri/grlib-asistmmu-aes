`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8zimrJEY7JyMgmtYVzzs1yifrzkvMZDKbCBwaODzMAmjqj2NokOivAGzDQTNET/8
4R5XA68V1Fi+8G6Vga41WtSo1WZ6rW3rxDzbE1zOmtqxTBz9TCCm7vUoblvxPFFA
GCrK19GgDcMKIoZNq8pZGHhv2brkltP/ymCYtJ0tInKOQoB+zp85w+XKTwGj8HwM
DZVQ6nGj7L+mTHZD73OUxkq5L0V0x/I4PxhYBGS06UE07WxvNl/L/OTB3IboFGwX
6DF7aGIwcTPAkGjCOZoV4fADfDcvNnryO0qFW90ZdOo=
`protect END_PROTECTED
