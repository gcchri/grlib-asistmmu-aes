`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3LHEtzjBmxzOfgRcGsoNwA7GkQ/V2lr15+ucDH5KJ+o8UUcUH70vLFr71+okybav
cqCiAmtTYxK1MbIshu6vC24zusBH1EyDYPiuF884NECPM6vPJ2STDV6hTEy7R+pg
JwgIWRqnoA0NlzoDyRti/skk8InB2JTuq0ZI3zmIfz5knm1fhsDGs30jyY6AiCxy
6UrMOc59tjO0rK3kes7mURSSGYLKK2j4x9U/p6PudXZzLM49rYuqswEX7bVLM4av
N3nyZ6o6ESb7Qz4jZipVY8F1FocLsoxOL5PZSweP1Qz/25TsjFIJHVeaANOAQum9
YHcsgn/jjQ7SDv4EHXYfPkbQ7eO8Acck3JOSvBUq8HoStEb3xFRPnk/oBtxfeMjj
aCyJPPyydGtOVUCC38MEGiYIXcQt8KwsPrWOjyuq+PHUvysbhb7cmbmsnVfzdUKa
XrGd2r1o+SRle4TgzsCthbIQ9iH7D78di04hQjahPn1G5XiCDdz+yOMAFKpoAgZi
Nb/Ydc5REM9HzOFABnBkZFfTEQhncRSuQ0WpQ7k20B+I0RkYM5Yc3odBtsBeNvtn
ePeDxnlWFrukYHORcZrUpnYUqaqyNpmNlZQUiHOa/7Voav3UvhTegOY+cwAxd0Ah
XZ7XU77RbBUAiKJ0ac/uiw==
`protect END_PROTECTED
