`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b945uqbdYy9SovS3tcBXr/plYtovNdwtSXzk+EK6s1AGUUcMS0MQSMq/CpaXiyCz
LoS3f9TyuuCGIaCxBX75XUbjIb/qJslNKc+W92jTCBd03oQwpNWxr2chn9y7IAaj
j6hKxuf5MNSu/hps2HJVa5OE/lMW77Yw5nfQmYqNRZJJZ4mrKS+AX17dddVYp2jB
Vdf8IR/tPKLKCYw63ZhblUiew/lTUEsEj16O0xxApEh/+GixQ8fYMTcXIoAI/V0F
+kGj0JZU+I7MTLiwfHvjtYyOQnsZc2fh9bHofBBgQwArZ3+dh65KDrkqhbAvFWzS
5R3mkSQ4Wk6foupDKX6vofBLdJL6bTeo8M6bg3LoNw2i9Lo4AKytYKEKcUFbNdAu
f/PlFRwoXH67OttFgk6GGmnNaFtQvEOv3GAu8gugqjA=
`protect END_PROTECTED
