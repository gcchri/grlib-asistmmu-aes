`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JuE+uI8gpiZSyq+zFaYIHnUwNgdPCbwfl7gCA4HemMrWdBd4e8Dz+oQVLQnPFPd0
r+oPC6bxywMMl20Xy1l5oZLp3+HxkXmBTYIPIlFEHD5y+S4ipDp/MopOILt7CD1S
Y64zuXSlo6kIi/LDMfO8RBZmh29ee5C+aLMHUjiMSPc8+afT0vQI+AD/K9yScIg5
OUhM1Jm1aDrmijICNrXPHeL0eAXxwjn2ZNW7dFuJ3sGPNryZHTpz0zLssOrGGCE0
q/+aI9yKXQ6Mdfj7L01DwIWlrnLXz72L0WBBBw+pw0+DVBBo0VbZF4hZui1wHtZH
xBPfYDrLGGpJqv5ASlvZYm+foo7JqD+pDGSoCBqT/5zScn2QEEJNi/fnjqIqhPvn
dXfGRvMjZRqB2FUfv8i9kerMLvlGAuFlG2ZFJChd2yeoppFGXioPRYUAqT82e7iy
gggmoRMA/gF3QgPWwhJiNciGuRLCGkrveLPm7EYbwQWprm5WbookxxxoqwpACrPU
y8l882VjxFQNvKD+CF7m4yPWSt31z3nKcDMIQF8+XcyUqXFaVEuyxX3a93kn4Lyl
6Zb+n6CdDSOFANA7JRtJUldxFeluZanJd5HR2rO3T/2ca3d92DsC5T3fBmK5oFLo
cnESPeCqMpW/8o2VwnzpBVH4QAapiCWebBc5kZFJoaycgQWHXUDBSzmiagMvtA+T
OJhEK7n/HS+WIFJ4s4slSWoUlpj5p5h1xgZ/mFUtdAVthwq/wVx3Td6PnfXgXLur
F3tFGtgtQkcKQ3PdRkoYES242xp/Q8XOf6y2DldH8KnDWOj37QQCR0ZF5zR0lAr2
Oj1M0AFpTL9wQBPaaepaDkuLTSYKD436r1UfG4qcCZVUKNkjHwg/4Sa+YH2zR7sW
6uKhi/a3EBwWjwyZIVza0Ar8jRrAe+v//APsamjXimW4NkIOvb4yjCYtTG0TuMx1
qrE83MZn2PgeJA9/yNdJR4+cgXeA/I8pdxrr98mbvUbzAg3PabQ35Eo8HswukNCw
8tRkTOV7uSXNFkWJP8YZYQ==
`protect END_PROTECTED
