`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y4K/86qGUQo5PWIxBP278YD1JuiYqMQiGk2EedjgOoCdkBsZ1c6Vo+mkRv3Rykjm
Pz4bMyEbD5wobGo2oUB2IIqsP6zzO7F1enYvpq6OE/NolUn5A8N6r24pO8Ulp4WF
h+5rFH21JdfDT5fZvXw3RiU4YdUoG7DVN+OkE/37Mc4mDv5HOPlUh2bONHE2xUfT
6kXFl29ftG0bWTmXLSvX6i9rzVXP3k8p8v1eXLGmNbbvfEPh8RanrXLskbLhhYxs
6FZ/9p8gosD+YurTaNeDzu88Nhe4qqDljOALWltxWFrItrDAc7s3a32IZ6cndwWe
MFPt5jz3w3ak5HQxOv9DpaTPvegfC/O09HjGeTnU9BJ91CoH4mQ+yvR6xz71qQmF
HLw7vhOMszwSrg0SXqs1yW/TPh98OGAZKMD2oLYWhqVPC9OvF0TNjmGJpnJNKBmH
mfZ+Cuj9K6xvSCGjoiu5MITXpZXjtJ5Ml89em91q3DTx3k43PWGrgJo+XwfnnYvj
0Vgr9RrMrKCGWMADtmV9eKjpOCx7xjcxD4bPDeizBt4qFozUMccJ+1oysrLRkksM
nHTE78lIaD2RXvcOsAvhK0h376tGFKIqTxmsIY7+xYevaD4woAjer4MXaqn/2nyH
57dBz4Xoi+3bJo5iNjDJMDIaW0SROt1PKLX/qlp0A5aZFx/qrRasWk6Cf3/PkEtz
OA2lsfT4R2l9G0SLw1YPj3JkS/epIIzBxYd01cOX2oernEm2dALQcmr7vyVW9dPz
hU1vXBJrO5x/i4OY/ynIdw==
`protect END_PROTECTED
