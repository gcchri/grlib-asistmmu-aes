`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
47g007xPlodwMmfohyqsAAr43rMcHyaC7s18sRsz2E3aS9SrQdsFHd6MZb6m1Z89
mFvzebQ1XBHi2rF3qTy+QYqvlKV2lG9urWndxmciDQCaNW1ZhcYMyMyOZ28L/E4a
RwJlQSr52DXsWfxAb8CHKcAY1fl52+G0MjJ9LWyCCFzksmHJ/UHW4i1IbthLymen
h94LGlrMePG6j0OS0dVYAlGKTj75bFI/HSRMgmy+WqHbyNMz0KPHEnZIqGP3iZDc
Ec8COqL/z84cvx/bXIlwLA==
`protect END_PROTECTED
