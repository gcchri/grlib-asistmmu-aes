`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EaqWCtEOIW0dL6OKzux8fQ0nA3coSA9s6ti05IeEsH9IVWBLAXofLl7JPpzu65tT
X+Qg7z6roAhsw/1ruPCu+cpjrFbFpzRVdF8271ULybTj98G1SXKk8SvnZgYGdgr8
Z+WzBDztmp9K4f50sd7jYKqsISAkMRbQGXTEqlwEN2wlzGtBlWeVzVE4WlroCxSB
qtezQQN8+PunAQwW2F3WGfABW6GtbhsU5oeA4+v/kyTpM7mBMdYv5wDPpZm38QSv
ks+p189sBk0J9OY5BBhB6UYxjn+2PAI02esKKzT3KE+EZXKkxMYtQAK56tj8l4VB
gBOLbU1gvrmEPa7+efTYa+DZIrW1PxIlVgmy2NGgDnQmrOoSy/sK9EVo5z6iRgVM
rF0Ox1BZj4uPSeFEH3S86qKtNHIzza+Xhh4J/0g2TKhsxkP7v0m+60MNyyTmVkc7
Or9dRcVCD/xQmmx0Rp8NbB3ZU6NoCxn6l4NG4LqF7rsObXSncfWrhb7ocMT4dTWA
f4Gk/lfqNr9iKG73+WYx0vlkkzIwNvlYn+geDEDoJVah8PhdY2GA8VvFtm2m74Eu
e3xrQzeAtToaMG9KTrqPy+PS3gJupcZnsU13ZF1rTEdHEIcx3aREU9efByxDngNj
2fQewkhX2l/06z5aSdi6KnpLctxzx6oo/5m7BAo57EprdvzuO7ZHHrJWUcITlNLu
BATGgNATOKtLUpegliAojvPNBRm0VEPbO6NLJXWFbPRXBTWjJOYHDzpiTaePrUhB
TBzRiVyZVPXM8yZTtCQF8mR5qoHRyn/zWwezTgn1YjgVYCISamBX4j5rTFSYGuus
+MtzNiahPJwMfsbejQz3YVZf0F1Qm94v/MZ5SyAKsGQIuEN+/X9dVAEUD8HESSYU
AQEGi0X3S9xmjekcKuHHT4a5qlxNAZwLCd3nfO2r1NSMwi9kD31zC4DF7ar4BKG4
fPYPPFTs0WhT6oWbimKuCt6WYuGvVAZQ6BB4oje4vuXtTpSLKmj+A7CVUH85tf3+
UHj4gn5gwKMoBTGb6zKDucj24ujraLeNklLjTIT8syv4ZncKUCeSfNu0uHmwZ5QA
JVtpArL9bKtjgFK4nLNdaXHfOR5B4e+T7RnG9oZ6UyaKQRfZIp8enGY09KOhoqWJ
urI/2ViftFdR6qDrgLNIpDEoMpSG6qAUc1rqYpqosbvKJkc2sudrIxrH0RccKjCq
sVzbtWeXei0O2r6X8AfV7mel57gYCTMWwgK9B/rMhNvH5nvy9wmfha9vj12pVneY
lDv926zhhuDRncE5GzKTsg+FaaYDjs+PMtTHXWQfqh6DkPe2eh0srAIrtoU2ip63
yQSn62OM+diXJFPIMPte+La3l2F+MJSZHEOHr7aNt0MZ8yV+RmdXSMtRtk3l8hy5
a2OjWT2Oe7ZExUF0XEcghuCFIjQ9YUxsA9fqYK8/QtRotf4bozAAuZLlOXZJwnG/
cgm2rLg72LJyEuR8UeBbrQtTIms3ltPmeP9bp/r28ndPDO9xhfbML7RI5a4VcWRE
KbL8FSQQTOUSMRXvaP1rxrn0CL7i4ruXJL86qQHXKXAbEP8cabLJwvvj7GJGFnRI
K0EieIV6yYcJv1l8otk9FUplcn/rpJJY6iXzx3Crp1DZoNYxzhj+G2fTvtt1XRmB
Vd3j8yMkvxFOQs330+NUbQJ4mfa/rAW/Yc5z4kmGyz3Bxq0X7VEFtsYFzZ32ldmH
`protect END_PROTECTED
