`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xYEh4xXJaqZFOPxuHsRVTpdGL1jSTphH+Oz58aRxWcH+NJmYZdgZ+1CxYIV1P1jA
mc/VkqAlt0fYlTEfmO9kqjgwqxTenzax29swMj5ZMgVIWP2e9b0RQAaawACYpdkH
SCM5kE7H6wmAdQD9icU4eTv5EdPZfQ4CrWj7KXDHXoy/tPiEAnTgYdyzhnr/zvyx
qarWpdtcv9IsSAuNWekFFvuYsoZtanQ5Vs4JDtAalWFx63T2h05PAk8bb8hwI891
WTroCIBpTny0a8TU3GZL6pmVrweFvEGnfAyELcxffizUovsDzc6eg2WEs+MNaERN
vdb+qYZ8ARpkPMn+t+dJjv5f88j41jSUjPiRFPsF38HawHHssvOdpVevEIeZX+9g
TEZ2ZxuHpW4fg5Llg2hj3hm3Li/uhe/ruaHj/A/37H52i/WI5XP6Kh/ROBGw+DRe
yQh4/5zTwNwuoy+VfCqz0bd67dpvz1yvcjAYvj2MSj9RfwLXZ8QS/U9YYtXebLNK
iSDGWJhTqFTNiYCgCZyMDf29sN/A5tHbbpAmEXqKvS7SVvWaMGRJWvrViDc8gAh4
zf50lWH7CiiPre21Mn8lMksl4tuuLuegWoA1LsGdwFGCik0IINOVBUd1zSIw3l49
D4JCW2VqEkxj+4nC05WxJxVzOWUaM5CQgIBCErLbgA1kJp68bh6YHZD9coYkF/TG
FAToT/2g54wi3MsUgkykHZBt8lkZU+PhSDtrNerQvQTwJoFsUJufz/AdIJorvqLx
BCqvoZxG5aMeW9GtqYAmcNes5pf0M23QAGdGhUA2yZuAnb3qk7cAPQL3Jsf9ESVl
fpBVDQ5iP5IlhNrqdGmfAL0qViU+edcyDdDPvHKK9TWa2O+rO8NDqha5IXV3yhAR
PbxjtSVUy+PaDXOjui2lCEGy/U8vdRCgSwo5WIlCHBVAqyE7Ir3mt50xr0kx4+h4
uh0rPskuge1oP4Sp2KXnZtMFtdynmKpwq2cQRYUAnT5tiO1ifDz+tgxg6JOei0tY
`protect END_PROTECTED
