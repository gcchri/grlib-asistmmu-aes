`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d976Vc+LEKTTH7oADW3loIRFYpMdGGFPD1CNHumIQKk1oJt9INO6B9ofFGQaH+9/
gS9rMq5yidq59q0RbteQpNjNrVxzlcgB7LRlt3iFHQZVof8wgtHKDcBgsXhVjozh
Iu+QlngMI2K+bkXUsi0PIiqcRrQw9v1+z48ApDWJ3b96XA4JHNx7d53Iu8svxvD4
yQ8UsHjAYsqHbv1Q/oicFcOSdcvH0q46g6E1aW3SgvNwvhdTY09FINlF33u+qreK
Z9JfapUDsu4TWM+zE0qz4UtqzejGRp//HkIMihUZodbK7EJwQHeXBeQAul1JjOwd
KtTAHClaCZ0apTjVCO6tXwm8r690u0m8LoGntKiZSxs=
`protect END_PROTECTED
