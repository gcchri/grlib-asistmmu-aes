`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4bztfMhchRpOX8am35X8oRwyHxDAy+EriEVCMPpou540SS0UPzKh7upCPG7SYhXH
7Ydi5YTccXvvrgT40buG3oZDVi/C6xfzYkIG8ezKWwg9IE8wy8fsc4xB16PeneAc
u+hXjHhwq1SEeB0VsE3BupRXQIrEhQpDTIbFsMyftPEgahRumZG/DDG83Ul5hBBD
Vm5mmel7POnVXL8uG4I9zIwk/1GJGVro2U1XiHt6PDFOu09BgQPzpCks/GZo3Gbk
isCva/hrYx3eh33jwV2N2f5HdhZ+R97I5NlFaD4031xlEEgw4iLCm3MN5vhtU7B0
BgZMk7B1GpHtm6V5EResaVAruT4wDpiPqR90Jy4K+/uftIAheY7CUzqzdT/qHGJO
J8v/2Y/GFrZ/O+mkVy+FqTt6ZCQRCQzE6V6RZUafiPDL2PVQ44t61lwv4yodZ48Q
xs/99/2HnYQfiLqtig8F6hrrMFxQum8h1yCtUnMDmF91GWiMyjY0hkmMTW7OdW3a
PQkfuhLKsvfql89fE3zKOLboQ5A1tIormCOelJ9TkLSk8jZzwipAcRSccWkFl8tu
E7SP+6UuJZSX7XkiE3c09fhzFiYwxBNGw/Z1eDiE+rc+XTaIalG6Ess4beBYmRLG
wI0oWKzao+0Vq3NQhOo1Cbgn8COLxyd9fb/wJE+zaiWlUkjLBCrEQIh0KA5HJjmE
walaRxA+65BbNy0YZiLsbxnKKvSMgRH0PU3hB+HIK2VS+edDlk/umtunCnhJOZ1u
We+vWE7YpVrx3MLS/BOvYgFC4gmxngKMyiM2N2C4HIO5Jj9Pn9eJzNf+cFpcg/f8
/glqpEYUj+s4fw51G8OGReSpLul50DZHgPXzT2AwSrJa+VFCBdMu7jXV5VCYjMRp
1mK+qntAyCzsN6fifqsmNjaTQAtRwh74zLnBW4Apyru484HM8ThlKd2sVgykmjqK
SuV3B1Njb+9lri6kkyT7IKAbcOm6GNXKLyXTHloqOT+8BR3TvnfbMc8w7+7Ek8mj
K7056T41PcYkpNrkL7Iwzjjw+urZPDVmSZIt759ld0lkeMYEbuVwQbeJSqB8sSyl
ww0PA5OSC4f6ZgTaYagBHw==
`protect END_PROTECTED
