`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n1Zp4zbPSI79ClJqopD1zX1huhhV7ODneVKWMkDvfpin8qwAgsKVZusgpRpREc0P
wxxfRz1M26tX1OOLG/BkSsMmElBY9Lc0OUVM16N+EOX8ewE21WFpnes/AYrCY8CK
Lj8i/ZH83z43bEEDj3NrfHxaQ5KoYjRO21OHUQyJB/fhw2J7gbkcuU3iyfVkrn6j
1ZjEuOO8149pb7g8aDPNl5AAY0iqNpEF63Q+6Jxnx011VC145loOB10qazRW4zgL
HmnzBufNBm8rp9p3pRtal9UJKiVBU+Tn6q4X47QqApQ/Yu2/8iIrMx3H6SsEOlV8
Pazk09tNpFk3AsKe5FKPa/jUMm/xwCjKyfQFk64j2Vo6Ud8dAoyXGLt8IsePrgJa
qlBimkZxybHY3LP4QAQymU2RFbwicUHTYBTN/nyewnvTPbVa7IDQKAEPmYJMNzcp
1MDVmgqgg/R4KzBRDLuudTXQtSdPSuzJ293SKfcV0ZHR4X/xxokbQCiA/CLLwwEb
TCvEG0xUoBTQoTt5OivqaHrzM0D8hnDtHPXj5zljpaV8Yk3JwqhMSx/jQfhzxB5j
j4yRMH68HJQVTTPkk0qUf16lHLFdaheWwiqZvZ34Q7nTMPkoehnStCFModFnFrRE
dZQVDhu2CJQ3TrAsWp8u0gbTeKodpOPpTH0L3dcxA43lrt7OEXb/79BlczEMJUvF
0aH6OAF/fK+o7sizBQaAPfibZJonPD0Qz6PrRn5NS4VJojHiKLnvlCTWoBPGUQFl
SJpYf/2j7sIVV8e92Ujz7VERbdVQRpmx9XNO6UFKNAwfhF0HvZ3zX709axwBk3WX
wmyKEH3e20IIGF5lAZnFPHh25E/33jaRHhYydhWmPmy19yNyoIUOfx+xldsf6SmD
HgtjRdiX4t7gQmha2L1TY7xD4F3VUOGtwFJMZ+5tBpIkPcHTfepy9eee1reNjFJp
`protect END_PROTECTED
