`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ih+yqvqL2qTRS4X3mXWGIYuR8g5WcslsPnN9gkVuh2Wnt6QsJzcs9cCkDGOXCMZu
DdoNusEMF8KlUIMXjnr5AHH3zeg9K2KtoE6RR3TzUnAezdqo88+5HWmNWoVC1cNU
wBHZjlyO3FL90hVEjHghY7HqmNhGiwUaYGkk0JRgXbmATS0+Tm9vYZWmio8mll9q
0RVMRM5fS6heiaTv4SuzcF90gOoH2mLbZJs8+kDBmYaRJr1HdY7xriNjOiowb1ol
PadrQO2fUYvPZ/v9Isl3jUDQ8nn37b1/A61xeuBpEVR/BYWPVN6YsGt3CVatqSij
`protect END_PROTECTED
