`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9ppV02Qex5tjkSxkasZ4eZm+pv+LiKZH87TNCMzVVSGd1T78YCDnnzamY3F6srpO
ydSO3WDWBFh+bufVKOAYN5Cy+dkqhMxXOa0d77F19l+zuKQiENNh1k8Z/BKSmWDl
xMB6Rb+rVAEVuII0QayhAFuq8LVO6QawASXU3wObg0eLRSAGHNSBDC8BxVmvgmZt
cOh6zlLdDo+qzLohNVkOIrm7H5YiPleFUBQJ5+2/3M9OojcZbdt2WNpFrwi6PnVx
qXeM5sdOdP1WHsUoKL8QJUKLQAZ7y460PLn9vuatDdQGotvvokailJ2lsOvm7YH8
mvMrL3eAI9wGLP1ajUhCyYQwsHbMaPkGIsHnEk2ldvt07LaeKSZdH6ZWIHIDwfcw
qLkU20G/jzx06OBMSZzLaPLwZx0FlLyhvQ1ZxtbAOVtYZyCtBn4CJZi1Y47kxVmV
fQia3wi+9b56f56W5DKL8YOxwZd7jHGbci9o3bBmE9CkdlOxJ2DGYq44abL3xF/D
qhNXJY1RIpxhXSSWAanLhlpIw6WejjB/M/QEiv7QLYtEjK4zB+vBr5a5nTV8WilU
lGp4ZYK4htSWAptQTxPk5W2Q162X9IWqEdCe31/PpNEKcvsnynrI81Aq5uHwQAKB
BhB22Fc/tQq5BD0E+oY7FTYHaqxHoaVn2Y5Zc8OxPdofc1FWXcM3buTwGwi0ew1S
4XFNZ/lBkb6Q7Q5QILtNiV6P0XE4NV10RLob346M3+t4yw+GiyO2gFYg08jIM4cu
RGtT/A85sAxlwL7XlDimvBFsgsAk0f6oxnvH2dnZOu6GohB2T+L1abpxpRXB2tuW
0lbj4lIUgythwK55l/gsd0YGD4mM1N+0x3uCguUx1AhwFN5dqQ5aFtPRHI+XiCJa
h3qoXQok13719g1IhwsXug6f4Lg529IP1ZQjwsCU4zVbAgrIkBdDJs8oQZ4owX6n
62bi0tVl3uVixMFOhdbZJJH0JMLC7lmqMwyIgCWLYoasoMvka7pfz6GBKXzGIyY7
GVZzSdpiorv+LsNz6kiRCMdazFkCjTvb6TF/H4APoWa8jltDeE8Kh9bXT6jSCvnq
XzS8DkEETSdx9zM6g2TUEAn1fjVweCsPitZSny01J0i/EAoetRoYsRBUDQHcKZl3
WolH4rVoyddTk6xkh1lu+yfCn/uFWaexhN87//T6xRsGxfRZOQzG+eghXvCoSKTq
QSQTh4a8veFq2N8ZUY9EmoK1MwdtIxKdMSgCt6ezG+mk7LKAZwBJ8ly9c41TmHeK
N4qDEM3wEzD6Lt9jSLVcFi5Ekwtf2LOaxmNrWPqaTUauVwKbZxTlQPk/WktBzzYg
VL/ZrNAksQWfLx2B30KLbwi5UIRnmPssJwjSCL1lb7b9jAd5EdiC1hvd3W3Tf7t+
IFz+RNRXbaehXVJraQv1zm+zLP2FLhUHkrSkO/e/MaZKWSTUpphCj5m6DgZuryOL
wjmIjf4NgiFaXy1IUT5KtZmY83tQNtqcOPLQpr1IXKteDqY7cLa/4PCYNMjPWKcN
+tjASl/cM4mFYZ9nQ9rENtWT4X8Zg9xjlLQb1ClxZ7KRp/unWcsM5uVq5GjDo2Bn
qICZ/w8lsGpBvbRyR95/ylkvpf3tyT2eWf7qq7427pyWgMgIu2a8jabh7pQ7IeYy
U6isiO+VjsqBiJ32nLEI2BNrHXIbdCpZ4NhuY/QAORlD8653fFI31FMoA/waMb6i
VAei9Eo51LetziO0HOB9OEAcvAEIirHg8RzwdSMA7jDhgnUpXF15iTPYqCJTmt1b
AhRfQTiV43wvGVm00ezaREtDhYancNw9LJub7J395DXE36gw31CtCdQIZSujArfF
ge5eyplMBlmQXNmHzTFLA/WfScLUWEKKDemkFsOZwsWr+GMUzXPwT3Dhu0G+W68L
6NzOVkNXCTXh9vq9HWdGunoU63t3pMw6Elca26ty45yVleoPtEtLPzrQEs1glDGh
RW0KGuC3AUlvPSIyDMsRMCNURHrudb6eLd7UZN0YUQcfrcOjo3fI5lLBnA34jul7
PMCrLzt/fgfSOruIYOi7jvfym7iWFFHx0/8HPtx0FeYmG2VdJLbkIZrUOv7RWd0L
r4KMhmXwQ8hGbJqM+4esjk1hNeuwkT/6yV6JHI9F9aYiRMfJAWr90Q+KNID01lFs
QquUBH6jVi9ikruyjBpHB0Wjv3UMqgXdpgRhJD6Kbb0L1hDvj+aFoRKpxTRPjg6K
GzLpkNlwWQ6neZw9Hdj19BPLW6bE1awYDOrvrBAtlX7D67gXMJgIp/8sOESrIVY4
i8B2Q3M9yXbztKKytlnmI9JENtFQZlNneGTgOE//IXgHiBlIVzRgECWKIi91bEjG
PjFpBI4ndh1at+V6QVGMUA5HyTQ3qGlwTHXqjHGr5AemrSfth0cjn8lCbuxaz4JF
fBkCbXueT6HmpE5sFajT6OOJ0Cy5eu8Sjh9HmwAMBRuYIkiEbqTvb5PgDGllLao2
8tchioyqeF83A/OIHjCGVYx3MxaP0rdy/jZ3WAQ9QZz/ECQ40K2ZE/pymdyTBx6f
JI8BGhby0+/vllAayEHXFdgMfqm8gRIaeROEtnB7N105i88p4z3v9gC8f6iGTAxW
2BPUdFP2XFVouZ+G5Z6lcciyytTsdhcGI2hsbOFUcFUWDPHTSh0HZ2hUiNCUalRr
UkgzrVIn/B9ed9KTFIJ4C0pKQ6hSv1CJkCgME0nIL+Y4+5b1osUt9KT+QJAEvf+/
KKXwjk4kLtpy7XcJU9XboO/2v649GdMMvrGjzR+Bker3VP2cl3iRLPhjmGDy/w3u
TIVjyjxBDZ1XCH8xHhz4ct92NoyhiqFWNA8HJiz6hn89jbCyLESQCJn72uopsmlz
VeBdGLnJ/yrD8cqY1CG/G6iJv5GckDQsoyLsAPfeF37qm+VkEpOXkQdx+VyTc+vU
o0/ipnTuKmPW3tzykUeoButc0/pk0KCcVj098ISYahyALNzj4tu4LcaQXW/didMY
A/92SfnQkedE5mXkdJ1cOyRa9oUffi6xxj9c8U6Jpy0K1GM/BhtO7eMTXMthSp/L
M0Wt8UvbrScyFW/osMaDWPrSh28K/mp0ZF06t1Ac24EnLASzB6izzyS608vKcGmc
v9kXC7Nil2EJSAS5ph16UJ3oltzBZuOH/cwd9SFxn4/XFl3XUb/A2YZ7hCFENF+E
bp+Z943c2X0GB7GywvCZHtoGlQ2N+LvmBrGGn01Drq6Aj1V3hHi4duwB+nb3/J/M
fzSkdAeAoDYQjGBYGrV90mkUFdItT78OPKCCuur03A4j1OofrS7OfrlEpGv4irzs
ZbMwg5TbyNi7p8J775O9QWbsWFYSQcSwKoH9iGiRn6XsJ+ev46qcNe1TxliBjjab
9Z/iu3p8/m5taZPwFYpvVhctAr5ovQfu0xURbJZz3HEA402UB8BoTn+xSOc7l8ok
gjWlKWaVBtrT7tiUDEpLHjmRCd5uHLI3MPV1BNk/w4l/DSihLz3DgYnnaTyL0+WC
r87rXPyXtUQ1PIEO3arusZK0Ilz5Cc+GkWfqD+2wLpxrTcFMAoA1xBSwxngqvQej
6HtTlsYrgvIO+ycz8nuuno5JhAaRyatV3z0EpgOkpZIhOKoKsVA270QKMVv1Mn+g
65t651/R5i9w/xhUQrUG1gx2j8ednMuj4PNwuuy1e9aoNo6SMHjvzTe3WAbUKxxr
GqWCiZXJH606fEOC3TiFtYMMkVTuL9BAINxlN50nRH0WgdypGRKD0BYe7GrOywWC
IjVxYBjKO9VuucrX00WkqFWkdsJg2Ql7Eun0MzG1ondAJKA4h1YOw6FQi7yK28vE
LNwQl+n677GEvi9gY5/WoWyXH+MYkJP7xrH6IwXFyt+YOaqiqcTD0iyhgI0YIstg
O5Phz55+91eFw+U75qel+Phgwt28AotdlF5Zp6aB6ZkhMN9IvQTlNrUv97pjVuAm
HRrfMwWjruqEIjyNkKlaUf0qmE2GibqQqLoiwxax8cbimMW6vtgdVw2mmoGBV5+V
2vuWZtXSzK92/yPM55bBGP0spGSLpOWloO/JD3Bn9sOaEDMghLClsdhJUSjlszKR
5XWUovYJFmwueJLf86wZdjDFzXNS5w9QkWaUSXSS3Ql4ADWfpYxTrFQVAs5+E+sJ
EK6wmmXGCRyp2m5i7ZnoZYj64/QLnHsfcza2H1rcKQdhAO2RXZx4W5KsIS/DMvKM
`protect END_PROTECTED
