`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F/sqnZh9CpsyThO926rUoVqqyZ588VrLYNL45fRnxdamLWPulvtZ9SJEqGhmHPBc
XhpHJdcf9ug+wDime0k4IZHqmWL6fGDGav3PRPMdXuA21keGY2jisGhKfOD5ql9X
u2F3Ys4x8HiX3kqrBGZuIbGsIYtiaKc0JXpZlTB7mpglAKEaFvlANzMNbshtCqer
Fu+NWZ82/F31fHtpFQyVqm8elV13In8zHOT+oT50TDLBVyrrtAYZtVl6TvWaN5ct
yKUHj1SmK4d02SExvnNWFu7Db9IRJ7/dwr3M9lvP+8mYX4dbMtmH9lWwEL01Oos5
faMe5RpQymVyqKJ1TajBJ72EpZyOPw19aswmLAljBX/hiZNBRoAMPKCKeMKTXnXT
ySunKpUMNCrOcn3AK88Q0Kl32EBrLdxFtgwSalwDEiGOM6j23kbQSLEOX9dt5Aly
Sd9Kw/MqElA5+6KDaclJYbwPNj5P+pG9QOCFCZ6TiJnGgnky7Wu23rR85vJo6dsy
YS2iJw8t0avmrLbN6oasfTGO5U0nUAQMjdbdd/092hSgbCjO0cpOXm0Z2x1u5pC0
NNQmRGiGeX83Gs3/ryIMGM8Iqtzg4zfWSt1iDLK6srZwrq5az11aQ/hPWHIXFBsY
5P9UAOzP7Ily7MoZIRlQEhFZu++IKVYU0AaQFZtdyS9L0wNsIRR0HkcDcniPNvlM
YDaEjqgWAyQ/aksJoJtvRH9uEUjl0LnmLvmpwzUEcV4CGqrj7wktIEw0GxRrvFH8
chIr4vF9u6PGvSYFgkAeOFxKXAYwqxppjzxGHvkw5xKtLRyqAUHOWlxr2NbEgck1
ee7J7qQeCB8xl7xZK9jTuJjeBPADh5U2FX2np0NZvPe8JhKHOkNETcHaFypSdVSe
mYerCbfTVHeg8ImSaBD9Yg==
`protect END_PROTECTED
