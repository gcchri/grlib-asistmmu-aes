`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ILohCuTwUrxQhVmAtb22zkSEK9l00FttgstxOu0UfRkXBy7RnGyMu754gmUlvkJa
zpdnTHjkUbQ0aLLr3tFnfeSQexKlTAqgW9C3/eekz1R/zpSGxMNR+tLs0TNwfhxg
N/gmGo2VZAD+uIgn9Sv8YqOYG2XnXhXyauhbu7v1LK9HtJdNNa1cyfvd8njwucb7
Ra8VS1NZlxr8HJIq8JKRhmlpCHg7P9gFIDoaaIHkKSjsNsLkfhdxV5fKXxBaewL3
YacowXU37Hys4D2J1YzaRPUpTXylhlnMcqk3wpivkZ5/GR0LMjC/ek8xEucV45qA
B5Zot/OufH3Q4Ie7U1ixAc/DPkRwd4T8GslRgALDuWDxfaNOyQAeCZut8Toora/I
G63t/KmAToa/CQ+fSPiloxqY641KtfMIYLpYlkuW3n5gSGq8HaeqEE/SJT+A04CY
auRc1ho82k7siubMGCdjY7MN69z+mbyhK6YYxUpeAg1kqGL8TqA7d+g3DzaPXaFz
xik5KGoMpDShaTRukYfkBXYhKKrUiuN2rUf4efCDUFvu8Imz49eIblQLsPTNr1P1
gIMnabW5UXl+xBIxRCHrKTVNedkYjcN4Lcq6ifiLNBMTXiNsl6hEBedUnR8gOqbD
ci/g79yG+PnLreknHDDsWCxg2jjgMYpZfDSyVuoV/N1OiUx47nBSsJYW9ixpeJIO
b9/TARJ9aaDnNXwHPxlChhDowc1G02pCCRlUOgrOA3omFF2dxj4MZPM0wavPmexw
HzONQP3xgBPjXIr35dANi7xZ7uRdckyorSwiaZS1jc7ZrWW7TD8Vhaacd9Pk+WgY
Q7spp3kzkSw8RcPbUo7ac/X83E+fxGRhvhxIEkMI1afepGD5CaOgV1onD/hKzqjS
pufoJZ+LBY9ry29abEV94w==
`protect END_PROTECTED
