`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mRrJmcFMOWyzH+NXWnBQbKv6EEEXf18Q+8Ig+VBe2mWoBW9rq898hoKzTToFlPmF
QYcNDjpMDqxHBoknWOljXQBWbxqh0bm/jz2ulnuuDNiJLpYCIGcHsrUuYhxQfLTC
7pbBCxzgZU9MzLCPDRzLq69EymIXarokML0L6sbZzRMTpvHQRJt7b10xsENapjzg
or4ekeH+7dYFiQSTohJiIs7qJaMBRJuqTNQ6RnxmA51XjDOBPz8h/JRuriAHXp06
GyZy+s02Aufl4341AlxRadc+d0nAR00Jr+lyZzXqFil64zwrVyukzJG1VbXClGj5
iSmy5xWt3p7p7ZWWWgt7XQOwjFYXMBgIJQhoFgde9Eh9iS29tGlAbMYAZqAE13Fl
Hx7aBSPEKCEKnkul6Q5L/hB81L/7KPPdTlBDh2lOtaZXug5adhMFONo7aRESJ3Ig
/sATwRtP8bM4f4tdmQQy0nX4jb/oaDAOQNfqBpV2J6aQh2gqQu6x40dglQexHMH1
`protect END_PROTECTED
