`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EuDR1jiO0+7LzwiAbMpyfbpXYvo6z8ARj1Co9FJp9ukPmcXht0w9HD7fyjuvYZZp
CDVv3SK39HpfL60xYkeh4MM+apZ9o7E1Xr+2YoB684aXnmATxev/u4B2/DwP9V86
kOPILUMlK8lqVtWb3yugo1z0RF9XM06rrIt0JAFpENH/qjzDCbdghdfas4VpiIbO
qgn470G4Lw6kaRzGbChGt8nEsrHLd5rgWtCfi7SCAQhhcP2OJ633dxHZaQ+Fa+gc
MPu9JBBa5wA3OBeyg31s3LJ794eV4N0vqooQoLkH+bPfulg1NTZpgDiNTbO1dBuE
7bWmxkl688wTJrdwzAEqN1gfhyUk8nl4LaTR8QDrqTm3X7ItdQhvqEf019qQr2Yl
3STbjFugC+zgAsPuHB8cjIsugfx4VaGHm9GPwZIIvuQ=
`protect END_PROTECTED
