`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cl71bk4S5KOPD9aGGaNrpjBMj3zQvN9ySnYrBR3cAaR55d/bSFR7FFwgtAJ0XXl7
6CLwtxjmncRFTyNEzwNXvAFsnuqLV92M6KynXV1P+SZKGdiohDrgJ6yVGY6j010R
ydmoJGnl5kE9cEkCQcBPNbmDacw6RYgX4r7advla2Lv6Qns3JTouMRW9GZh8QXF7
N3N6KU2C4x67USDlEDk8KxHEwiyGUVPc5BtQRTfwo0QoR0G+nwsMI7XT+nuGirQk
uPL83MNATDnaldWEMeroBvyrzokFo1lbeAAVEguXBrjsgwC5ivJQCcHnlgeEHhe7
diXvQA+yVzIPXstNNmPWR8p6BCCrSRYe+EREZ/UvRhkTTrAWPunmMNPaJsr6KBOI
Pm5cjrXNIbEJimHGwUenJsIUoNUM2o2yvFhwoHrXVFROewLtjk8cxd1sJ2T8lDwL
xubrLySBbYbHKJdw4lXejC2pL2Sc5k+odAeD/5lCxd9MlTRKHrnKz79q57tLxY3z
VOs2lU/sLVWIwJ9GcEgHAQGsuL2k1Vkew2tuk2zrPtAC+QoLTjAfDKgEV7D3oI5f
33awSOguJzMXbctTUXWOGSfo/SUsD7vUhZWPrtHglQQc63VqBbltk8YIOT7azyuG
CRfP7tgiORxyFGLPTDh+bBAXEYQ+YjRojJJcv3Gw5gRYdRbR8Zd/wuA1QZafS9jI
aqqqQ2MmOeGOpql5LeHe8D8A/kKrdNdI4LPsJFZepfAmmteDRD9gWqwWzuBX+RVx
aKqKzncRrJC4ZMIYgEpmg0f+c+uPkmBn2PiwjbQ8dEKpsGcaiUNM0EwuxEiMpb/0
MZ0dYsbzbRclbRzdV7PVM3KKL0+gKYl3pxFXic7++qbXfjDSunX47G0MJwcigKIt
W6EHDSQLnvlqMtx5zjc2HaMqhosZ9XTjNO+Kw63+aJwBuAkcxtVE889oZickdtuq
YoNEaW9qro3ltWZLnfzxn3AXy6o89QQ6xyPowsaxuJ90ejhevJMjsiCUTqq+Uj2j
TUiB6OYNgyOIc37hMor7ImiB2ZFrubf82plXX6090fSbiKIl1WknBvNj3fr5Z4UT
h7YkoasFcplnCxNXKI3LIedH2Wk1KJFSesJhCYoTQHNuIItrpXJBhU30ZxPM5CmR
JhoyFqjKbxNpDyNTDlaErg0EWC6wGUkOBCfEONPDBMad79Zsl6FKxIjQzqTqShSD
8h5r0Xhoohf1PLJNIgT3zHcGBamWjphErx07C7Gtgiu/2OpVgviZKYAHeyq5Aw16
aDoJCjnianOngk12QOQwWgxAmvogJvBJ1hZZMHzDId4/45lHv0EHFSe+2KbLA7KG
UMA5kWYZW1L3zq5lV6ZmP0869jPMSHprHf7JWlAI3S6U+SJICOdNNnzoQStCKDOE
RsuEIglGvNtsmafwTmtsX5iEOAVcJMjSYIObkgv7J3RwlXZMZefafb6sD0BZLP0b
pF/5cbn2Ox8gyGeB2rTuCCZjQpqui7Cp0JsHABa0hQ6/OZFTy3l2wiJGecTHiVvB
LTc2l8AHP+I5doSA+1V9nbo+EKkPzauox64t0avC+zGob2DyLn2QAYxg6/+wTmJt
6HdXZcQznlOfzOaEuJLn3pJQijpPNR96riVBjyaX2Ajaz3OVjv1uyCak0XXvhtN8
lSFfmA37A/RGZiLRJT0mYgLhqonUWRq9oaGrB0Il4fxZC+RhWTK+X7SsFXMwL8ni
Ps0bSjUaQGovCzZSG342+aJ12n2i2r9OxwDgG3rkY0DIoxNI7xgRf/rNw/F+n4C4
9wVpElaS8nkK2VEht7rPBfd/JYfM4fAJEfh4u1ZVCv/VZKogO2YAQgmeZ/3/g949
8Wv/e2vKy89H6uHR4OIf6h1U35xT6PbXq5CobZbX2EWAjfYK9uczCt+U0N0Jao91
H3JcLoyShKpIunfFxD4mCjt7Rir5zQ06eeImcLRj27Np1ZigM0BDYrAVqG7L5Zl4
uyoq3W733Jotrfls7WYUvYEpEye1FZLcLSL/2lC2DVnF0bHRLu4GdF8XIGyuxs5L
hPRcIFcDgrsf8O61S3nr8NSmy/qqXM/tC1rcZ4MXBnhDUxF1N36NnfllS9hcxlnV
PPGHWSs01TzLRUxOvedMjDD0oymAkZSSBe+0t5abiLObzk43ApBY1N22XcechbaN
mfe/scYc8gZR7Vs3zcrV9K70f/Tb/MUbqCLinldFIjiAC1WKdzStJ/t7/PIg/Z6b
czxazLThKqRcgm9vKHLpN2Jx3H5gPULZ9wjz0Ae9eqtu7KsWREYArjmMOIGMnrNn
QpUZiE6TR5z7zQsgOCLWWfDvLZ1ECAqSybXZL2yfvNBDsV0lpHy3SHUQEjXTrGs4
/mXPT/P/+okOxDfS+0gbmGjY89g6FyETJn3PmOnXHYLhyqPcBcHh0a1tafDs9UK9
KP42txHzBMBUv67RGBbT1s5hBkrCOr+atNUO+MNR9YXZD2bB9AcjtjwpVDYSp9zV
9VjlCKkh2uILDspzxaMVWFuQUwI3nzyGeSwyCGtceo4Q/RSg8Gkzh+Nw180JMTwD
sR6VQVwQ7LiCUlTYsj3kKAxaNtDDYEbOsmAYP+6dSJFvgrEvDeZRJzvFd4L1LNeo
+QoKK1xVlSWO8szTIcoHa2X7dQ2+9PqGBIMR72uKkB11KMFZEClDhX4VD6f+oStw
yo0HssqtfgBCMD2VpO33v7jfGdTZxETKwt0zWrze13Zt0SOJn0/3fDLQdLVe0++Z
OG7bfglX9ERFG4KCFPJTglxw0YOLgVdgvftKPtV5j4qpWNKQWShYn5H297KTbZTj
fP03g/1US8hBSnBtNyu69vLX/gCuA/uA+WCM2lyGnE81Qse+18OiThDoIhQoB9R0
v99Aif5IILShECRq7J3DyniJYGJ7Baguc4RkL+tcemC+jB3jLA0qbQqkxMF4noVH
a6EtDyJRAnJjYDYXTDyVi+cgVG+wE4elpqoVc8XxGxieKgphJZILBUkdCqmOXhoD
7i5J2yek/BgixN7eTbn250WT3Q4+94uCelbazIxSNZbKnyz7Slhf/C7IvMCi9Umd
`protect END_PROTECTED
