`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HrYdyrSgqVJJ76YDOX4aDheDFlnPhJJGPvwx4JN1xK6sSTQmsdFCxVIriOBVaxlc
Mi3BCB6Y/gM8CXATRMtkA94udKO8sDkWVwK03RzAdWGUWs+6tjgKRVJRkfaNIjVk
MJnFeKn4drK46dXrXmK4jxk+6n8v9+ZMyKbSnppnuUGUYPaOEk/55GPr1msEMIfH
kiF6yFDkr6u63suWLdenqOqGE8TC80czAN4z+le7GawpO+NYVfxYaVU/LXJOzNWm
oL3FPLTjZQlElBSRczj7yuU9nUy1PMxtY7hlqXMjsQExokWjsn884cMmEzcNG2vC
idTvXWjMtVjvtDTGUAHVgYX+8FEiAuy0IPcQYd+ebGYJU8EW+LzcqNnD/VDs0Qjp
ugZgMxBJXM7h1kjF6bOPZdKDQUQJlGDhyPh/7TICo9Li5o9cYauHy58QbH6AOPo7
/WDeS9WlmyiK14J0Jxph66Uzyt1HiVYHASbVn5rIhvrS3m/kjlOv9GnTd8+KGbW9
iYWBG52F9cHKc6qbdtFoXoSfhVvuiadN66NR2DHZ58RzA51nDRSxbALspwDq3g43
mBTcj8xN6gStk40CdyTSNlZ51FUR837JK3FjI0VvzFXtkfXX5EgEy4Gvmp/wAbE+
3Tbi0/tS2Kp3IdMkMaDT7pJnugW3SuUILMf8hU76D/2CjfS4Zj3WWmUOwHs+9C3J
kpKqSO3loLBRY5pIKhNI1Fn83fVm4irWj5Rp03NVuOc=
`protect END_PROTECTED
