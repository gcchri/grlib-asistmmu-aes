`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NmctRMRAdILXLG9bEqs/8beMe75T80SazNTM59+1JoGyPOaHp0oH8Xa7wpCarUbK
/9XZ1gRv4fZQGEfn8ZuiIu1UQUeeDr7g/G46bvR/lFbpKKr/WzJ87OaqTdJKBj0E
a/e6pm8f01Ppu3lYRGPoharDEdJPgA+Pmr87PWHyzlWtflHQXN3atUXBJF6tdu4T
RPis3T07j56deiuo755aGcakHJGUUMrTimp/5UN0j7AB/4Ok5NcXzQbgx6lRzYX+
UIqdBTFbbObqemkfI6+x0zk0BwvEoLzNljyzUKOCtbNjESR/6Dxmm7rxkBAZYoSJ
Glk6TbkEarkB4Zh+mvGiPwowHkxPCKMGBzfECX3YWwiXTOpEZRv135fjdAygacr/
wFPE3AZdJXflePqgObRoImfpc4jwWKTdk/03Vlsnd2zZr0HEBTPLBjFj3GV1qS70
H/WR5rb8W/zJFBvr51pac7ivYg5cFMnvW4d4NscYYmJebOC1ceq1r3XZp00kXW9R
09ZMw/WPbAnca7Q8PfkOibQqnOJoSpLKRJuLBOxAqRYjXXoyvRi9SBn73+1wb011
XKFyzl1SNaDGYXQSGOneRdvxoM7BiXmZ7uPAKC7hsrnxWT8VwLyCsgxXBgBMUrMj
bJB5YKoI9MvDR0F5zzg2JQO+igEDTPqCQxwG2C+iEksO+vhVXQGXtUoePW8g0sGs
kyida5XJQgGh9NNlH5vQbSujKG+YQZk5oamGrEq7e+SQcWUEt0G09OchAXcEKLNt
1/sxZqcaszDMgOKxNGlB/ZygHztvdxn81spjPJI09PfN+k9xhAgfDK5T29iqb+Z8
jXoBYHTCjPiwAhdi3nNWVGR8kpOGce7lR0rPbjjwyAZLhKQ2XDOHUIwZBq0zNpvf
kcJoXtADPcoJmqXAmNUrkFgV6odQJPG2OibFsKwSpmVIa8xxBJmGhdn89gVjmSBC
rUf49qj+4kg9eu9/5L0dtTRKavNBpjWrb83lN4Tg4PmJrBSxH7dFiyOI0MR13lgS
MoIOnEUU2n5H3ue0l16liDGkG+UuRPeM8Lp1KSULxfQ3cD1MQCLSHSYdZr35X/BH
iASi2uTjCxuIBt2UaIuXW8Uvv9aGtfnx6wtdOybFF/Vo2VFgmerdXasUqvuTx57s
+POEbFYuxzSXSk4afc5k58t8jIqDfHTlsljRETSpgfjok9kYqdieM744WU8f5C3d
5T9uCr7inQCufMwTZPaGSvTUnwDlOf9qMaicrfT1p0uyX9Q4omOlGNt3NzPX5qwy
0uY8zEO8qJ2LM2RzjNKjMOO0GfFDoWNh7lhONYY0rSfjtamdcHVIzGuewCtYxBC7
ZMuqwMF8KSsV/VIaOjPkccutRZMf6pHwuXPaxjUD5/LJVFxP095qFCg3rUStKou0
uuUTWIrkQtUJooYJ1JDkRpFTdxNjfAmGe0+Pwb1KUfpKfPaJhmtIRSy3gjWtpgUY
VQfBIJQC65LYn7aDcIYTn7gBfu+UlZILTbcQf6b6MPTSUBpc2pga/1AxczqXjX6M
gZeCRtZF6gDPcrWm9NInEMA7cDpFr61R2zaTKXsRmCCHztgDMeCKGaVQ0PNkO4im
coyYkWWa99iftKh0tu+YBZ25iv+L0jRdTrEKbhPgHaTbHM2LgkCHmk56itqutelY
qOwAUXgoB6sRsPkP1OHxFWgJ4dwh621y41qbrL8M5ADXuheEMNdSDjEQ2fKAxJXM
liiKb4jPnJ1FwWEYfmtGF35RNeT2XMm4Wj5JAaebZcOgfvF6iWLrKgjnSlHR5/YW
t1TilsdXrQUZDmA4I3IcgOBonTu1ySNWOfDdBU5NdiBH5xjXvtkYb2oWpJ5k7wMD
fDUyRLeI+shN3yp1c4yEnjIv/y+PEEnWhHkv8ffgd5CcSGdx9ncw4QVXB4yIco/f
To4dCIYYXIFvAA2hJLZPfjD/rFErxl/t796hzodECCNa18w2QHbpFU9BGSaDSFA7
88rSPZCZTjimR/Re0ERkFMMCga5J7vz9ku+ER6uP5U333gElTBeLFIPBg/azyI8g
RzCUGVoFLwE7a5nzk/m1MNlEILRfTZuwVaLqBJUnAaIsqS/U2f74gXYYV06vVpXD
xhsc9zQjl/EryiaHxcI9A41/m6IGM/7YFjh8xgQD/ELmg6AFL9rIME1eBqQmWv2I
PQeFuf3TxtBJWWKtwKXbLoGKYkvHWEpmb03F75FF23/EKux51V/s5MnSrlLI7Krg
HZvxBGo0iJhgrFuWycG+HRFLuRlF7GLja7wOmWjExE7BaGCsKVbJ+jeu9Sq0LiMF
4uwk/l354gRsH8TSwIn4rnxhImHJeMQS6gnPXVWH6IwMrEG2z+iiXSH7jzhJ2H8o
k+e7lB3o2pBtcpBHpE3buiQFgRMz5qfBcHDXPpqmHkyClB1mrHej5lwrwarMdjHF
BBwK1r/h64t6g20V8Zzo3kt3r2OQj+c3Wj4bYkgGpy2KhPVKfkdoYCPaspKNT5hv
q+zvwz8xZYwMOnrmb0Q7SqTYGqR+ZULLvpEOhGFV6XLOzmDL6wutTPFgSjO6i3rP
pmxscqB6KpvJfMGel0H9e9UB+jKOsXvTEi0DA9spPFZ6mHIt8PkkStkqVtTUZpGm
MkFEeUMDqr062gQiCsYQe6/jI+qW0QSkFoRF+/JomIQPw/bo/fhgPEqYt7r8r+so
3+9Eu5Ieh/n9fNRAyQ9ezO59KEuZq4W8H1/ix/mJgvtA/GPZ4/JMTIP7CeFweOqB
XMeI7mIz8HPbrr69POE7Bmqj59dkPBvIz53RJQ4hKplAeuaUXrJHVG23VMuaLRZd
rTZ4+QAqfYiN2Nx6Xetk4JaNnwLkO2AKFa3ZUekErGDA50RASnx6Ly8kixsTgLLD
ueOeB86Fb6/9b7HPvJ/SwOLt2XeXlQ6LXKx/CeBFZR1X4oty+gpywoC2RuAs/9IC
urPWD4rc0wPaCPSS98LqZKwv7TMbKnGvbhUaf9z+EZdFhw/n5qA5Awj2Ji12ZQaY
vhYRu7BviPlSvj4kAr1HFyz8v3kFkPjUjCk9EIETbAAtHf3cQO3trRy2FidiOmvq
m9Zb3eiZJcpBz2/ZnlYPdXGvc+WMPGthxDes87X5fqZCDtvqrgltP8BUCfwkvxTu
3pjRfpKorab+shoCTccLbCakSjq/uORvw8k+FgDiaVn099m5r3j3L/0E6FF1YFNM
YdUBrQNHUbArHxy+1lh9OQUXVWIpqM8n27PjmBcCX0n3xaTCw9phFcXiEdOetOBy
+m4sro0ohOTdfYbBYp3NlTCWUZWmcSGP/1sUHx2EPjZuNBhTuW0ORKxm7s2rYxv9
`protect END_PROTECTED
