`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
78BYnMcrxFVDBLsQGAXgO4TK2lJ7Z0MvgSOY9EdM5BoN235qmLScCK82A1++VqQv
xoqXq2hE41ZpEsZ/f/SBZd8ycsAeavJPDBFZT32Uc+OWH89cj8SQiZiyGec6pH5V
I4TVm3ZcQNkBNDofiB3ZSb0xknMJpM1sCqQ/mMmmKvQjgT7JsPQ7dXIET3XsEJMY
BQhVTgd6Dv/zbii0qEUt63i9Q7Qkql9kJSgzPWnMzgD95IPJ276fX+AOAD/IAVyk
TnPcNoSwuXAlzaGXw3SiaQ==
`protect END_PROTECTED
