`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
onAsf2nj7+++XvgsBVNo/FjUuyfBPu7SaD7VWijVJ/WQLF2sB+hrhofNpsK/0bpW
XQDsLpRMF1bdLNlcMbaW6J2E4k7IDAV+A/oLyw+McATEI34iUw1hXQb92moh617P
+jC7m0HWk7/HtxfhhlS81zf+S7OjEfDm2yk/CdsLNziDrWloRdb2narR5/HcssIG
/8QCu3fUWtU3lJ94vQcJhLaewY+4EMo/Kc8rEXO5xS2uB3bxp3cWBf5BlL9cNoUB
MZ2mvKWlh/9Kq+vhC78gSImdkIWv7k9SY+3SEf7rIU/Z4voS0aoLACc9vQHfqBTg
fyi9v1vAMlX6sZZlo/I6TARd6IWJkca+Tkb7JDluUN+gWwiCHyzZ6Kt9CX69HvEG
9cOupcO/zAwjlRyNSO0aTooSLe+H9TR+1t48nbML04QKpff9HhC1eGcA54lqU/rt
FfM2FuovNlM67BVPUGBSjfWquYSJZjaJSlfaoW5G3kwYZ/VsPZEhh872ZwvNuBp2
qsT9i9VBDj5jJhvp3kzSQcpf+s64zu3wZJUY8KT+8JlmJ1TGtTf97vOWgETb3bzG
`protect END_PROTECTED
