`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AxUt6dyRoGJzD13MM/46tDYhH0o+tH6mv0Ub2BH1inOJPBPuqK7avcqek2BhHKjb
2b3wWjc7LJjxerd0h18eMyulnoETJIYNIfbk4uaaQuK4d/n3NEWNClJxV3QdMh8N
FQ6f6wPucMF6znLCeI2VAKEInVMpqHe5H9hze7KLq65fcPMN0JRJRrUaciequ8pX
G1gup3iTZYwTbKHVTk6QdV1D8sCsbeaezIWTcyTPM9/L/yjQRVjDswN70/tixvi/
vlR6YrPVgRrB9kCcBsiawO5V3ebTqdLupsm/AKJrwWUq1wFsDdl7JvjI7pGMFl97
`protect END_PROTECTED
