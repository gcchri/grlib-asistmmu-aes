`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oG+/FUIMY3DEGRTq9LiPV///4XHIVNK8ntWMn4Xz202x40GLy1GHnfeS+sY1B7W5
JsJ2MvSniJ3QwkNiptFGRueBoKPLFKUlTSh63d6MMYV30HNkPqkMT/cqE9DMGIYE
jViSffo+oKHeGfpVtx1yGiPVex5XiZg4erCd9MSIWceBoquVusCMf19eQZLfu9Dy
pUlz3fEnkKTFj3Al5TuCiW9O/WfIycy5F2zkKXdYhIma7xLSCDkSdBJlt1oD985Q
5t/bKdRYluOjB+K7foQUl7ITZe+sRqu0dXkoC7i/DV+KSM7ezx7J8C3vq5kZ2OM1
I8ejicFDPz3Y13j8iDHQ6gXzxTGbCHw1w8kpCxeiJUVICR9uBoDnqxLaGcyJVT5v
4Rkfa1lzRUk7KxAlwpQuCmeDNbKg+LCogVsV3hiidelCCF7em/U80mdZ7MOlqzKa
eDzaiqwCjqLuiiUPCjyyYgWGJJ1stMRbiaKTD1ZsSPRf6OoKVAwHaTrYpt7j3dot
FEkQlAjjYimEZftE7BoJOpMuq2/c9IIcezQYfA54ASXPxTYg9Nf+ZTITacGNXXaX
1EMrzA+vazTp7yjMRpuklpK6sJptzEIGU+dzzza7T5f/QpJCBGsd06XLLXpfI0UN
6EZdVeGxRiL/+NHvOIquwHC6+wrV0TdlMk+xKvJ91V/92cuThrEZ3GuBdgvjf7YJ
q73IODf1ZdLKqu7PB2/SiLNzQJYC0zb+H8urDZz+cVAHDv+xAeuV3a1sSB4VGuiU
T9qaFuHwEflD/uk8/dJ61Xk2Wvj5KK6lPnxEyP6In6GBkydRHaTCOIbV4VdtEtJ4
t0XgUu/UuJyCLg2Wu6Xkb/1Ti4uv4wqorf0paJ1vT7rlcqcTVHx1p+b98Qk4IHXK
/reJigPK5sgD2ji2RCN9XUrdTisAuCmthz46vqlRXm91TqILduF4yGLMKS8OkQz5
2NQnzSRHhqJbCmp6Ncvx3iYM4HFG4v4/lYbUeBYYY80VkibErPfvNP0vQaz04Tnz
eUf0x+vEnq+OJtveBTYq/w==
`protect END_PROTECTED
