`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0I8jXj1zcBHU/sV/XrE/W9rIOGQMPu2IcKGbBMVoK4v+7wkjK8UioSGVcyHRhLMx
cqjTBayPyARTp9AXn8BGzb+F2jN4EsW5wpfRQpGMpTvRM3UGMkfr7FHVpLHFL5if
O65ZUsz4a74hauoA19RlbXhhKDtklDtG6f2RTjtzeYAu556D/aH/ot0Udo8JNsDj
Rg4SQtbkTgMn24YJpxmLyVOjiuvokP5NjMYRJkOokQO1ImmYPX8eYALhBK8uqGH9
Dt4w7RnsrU/fPGC8Eqb3C5yj9VetXa6qh8a6BAVU+pq6dKbXLoVSsveIrraUi8BX
OChtSAnrPom1YzTGL2/Jy04BP9NDZk1OhosqWn12CoG34AIv/1Np+KE3C5lG6+Gq
YXtqohTOspD3uGumiW9zQxoyNKTlv0F4LAkiYadVhBXIIANbOvW66b+E5d3GKGLo
lvZUE8vta7EvmfBBy16MM24Ej7KPCrz8rodcI3rpvo/J2SMGipvFT8PahrtLtxi8
0wuTUAiQKvZ1amoBRP2hSDjST1rZuE7Sat2mjkVOoXveR9XjMu5yi7jLbXPMynjD
`protect END_PROTECTED
