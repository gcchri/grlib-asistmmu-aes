`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oe862/HmSLxI+dJXh5Dvnh59+d+/oYL0Mri7zOYVbwZskAeKgIJBBjdCG2NYICuf
Nblzztxdb3oLwHB/+BuNxw104ZLXGKrdPY7SuDslzc0/jeQ7xAOsCjziMtVrx4zC
YK0eROcX+/ebLLkWCtzj+g==
`protect END_PROTECTED
