`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ji0INyGBBetRs7/j1ndz5EHhSvmd3dNPpQFZkg60Cxkly/aZSBAK7IT9HQhbKqA3
fEOawF9Ay5pnezNDEg5X91FhUfifQ7A7cfTrqZ7eq1DhrSJ83c7GDYPGmuhWWrto
PwYKyA0765Rb3K9YfgYK0E7x1XTGe5D3NT1HdSlEY0UoW2Qv4G8A8KV18zjKC5j7
ayc/223NKNFuJ6dS2/UntEevpt6DKvtWE3CTwIS997V1XSHNa0PimocxcW80/eG8
0DSduk8H8PJ/Ht2itjq09aNlgW4uFkEU6L/Bu4IPYeSR3AfhO4bMlRenI4TT0lvc
tZJ0FBcatmX+wsVvYWGC4foebhPbTBKqFfPbMAFrHG0h27qpD1MmHrMT+PlNQASa
qdT1bxVH/+NN4qSa8AsGbdDeB/IkkLLJTudjcYEAss2DK1+Y0aN8r19DPcXwpTI8
2D3IAPy7QxzFNnxS+jSsAmDDH/Bcjmud5MRLZA1jXauamHp+wxwjOLe3Yh8Cv9yT
2rCMtz6a2nWrQMY37tB1YRP4sIv2j2s18iY3srO6NMpDX0UWJpyFss34+SnOdRxv
EmX7WbuajXz1GUVPFJKXaS5WkMYb8SNc5W2ZlKY41me/xLNCMAEgQ69lmWp5+77F
czx1m7qdNLlI+96V25AWKCIPvJr9Q6Gr6tCF24MIJZE=
`protect END_PROTECTED
