`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rMN4yBFe5ewzhdCR5hmzdOQL5gV/To23lO74YeYXKNdAo+U05rlDXANWErdutcKh
2spADHb8XN6bA3Lu68x+P9JnVgRbRFoMCRrUgaknwE/P9PYgOX9hfR8WP6yZFGiY
S9zR6JFguG3YTDZQi+Jjv+XzrDjQDc3eDk5NnIx9zVJjFRqxFmdauer3vRM7d6s2
148DqPSUROC2ABujZfmDORi4jBBdI3wSOO6SK+C33uy2OncBwciONnGN5fNsEeV7
Qj3xBrgh5P4yBWadx+biwPO00PSGloXEZAcoBLtyZC0CraHg4//DQKycRZSU9dZu
6LrZBdLXhCPxcy0ndiOKDTv+5mZRHeXvVpsIM+AqGHtLDDWT1igoGrDj3EpZlc3J
`protect END_PROTECTED
