`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VbnCJ+MdbbcakhdLTK3IIK7bmy7lbV7pgPTrzEoTCE5nC7SSyyvY0zd2eJJZVNQt
cTihMRuvjT27gjn9DwLBlkVB1Xf0jrZthyltorW1oL3AOvWYHKVB+3tEOa2f5xRt
HCJ46wUA1TN5t5cmuDEAOYWFL0qPjmsqpoAt0m4C/vhVMz8qE52odSfDZkjHf3ag
+I+u1MEYwc3Osr0UixPdcoNrgjay9J61bfNBGbuXuBqn6K/a2MgTUJCDbHLHmFOw
zZdrCWGlG7dFYteWbDcF52eiRFKgjZofxeTzNLMTu1hgOIprwtfnosJtoROZmdu5
L7Ki8wKPqCNZxoFECN+nBXopuGFZ+xTCgZBYrEc+5ruZ4M1FeEFvMjRHlQJz2kUb
8QQqD4NudL2P0g5yrqRf/M4boLsQUZPX7pkuHUAlloslfkte1xUOXycleuFEWnWQ
qu1/PSQmROI7A/PHbCmXsP3MdtUXyH/Q5+ntMXSxv1xSaBboY8ENcXEcFQEDEC7b
ZTxuKbVmbwKhSRKVBmAeO2poo/Mot7gy1i+SIdm8j6iFsg4zoxj0WKIqFjOFrd6h
pBXlVYFoLQSijudTPuN3HWVRwPhdLR/69/fAv//95kKMqXLIo5ne+gw5j0kUcPMr
s5E+dYypah1Sw2fGCr2jYyuPPlboBvaFYCte+q4byCPaoQnYkC6R/i+//4ATXBP8
`protect END_PROTECTED
