`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VICDizqjuU0XYWV9RAV2hOE7UbArZ7rdQs5VByrV+w0EDfmvDrZY0V+M/K0Yzl2+
aBIcfF/lg3Im0XwuvGKUGD0E6Ms20sUG+Vt2dG8dzpctCxoHRWQLk5C6Bkhf8FqE
yjkxcMU7rXfjFwqIpqvmOcDKQjG34LmcWDgLM8HUvzHwkBSHmafzucLRNhLh3g33
bJINiA/cjw3NwDkp4SmmqWCQzJ7XRkgCEA9/qXo+5SQ3ukaq44j1w3XFrabiEsG5
xqvIL9wvjpkEOxdaO6852snupbUAjN50Skqqyo8oIZm0Li2EhWazQF/0uPp4s9Ea
dJ4cNCRCcdgnMMiDiYAizDnYh6KqxlnfRNKYRPnKRmju1rrUrg4UMBII1kVeDlEV
bJpRgudEtAR5z3TPp6OCJ50ZP+gxfW9vaYWzt2VUqjqYGhrODAtiWuu4ojnrYUZM
kJ5H+Vi4EGIk4Ud7SnsG4sjOaE7ofv+mMNUEaRbPrObe5EDJjMxN3Advzu6WF+PG
gHMaRlwqgLDmFMs85AdozZCNA+dbE1tMGVDqqzj06+dpBXWK3mFbaSQLtgJrYFdE
T7n3+BTfQtXqfEBKi+hf+93kXq8dd3NoExN3sG16ENKlQQrru6kb8et7lqcPc5rq
aXSFamHoBLDVXJPl2SRSakolaF2RHCnTRPY0dhNsTBC44i6TUFGZ2BhZhze/qYNL
uf9KI3pnsHksAxRzG5LALjalE69l8ExmD8TMpCQdSYgtMEh+GapCC9ukWaOllRUk
0dmilHU9cueTYjDyzxKI9/+Vrne3CIFRkDAWsYBHQdC7EATuKtb+BLZ2486b8DwJ
Rh/gQPozrTA8PW1v1Sy6bRIAYcsRAC7g5v7FDDv8dBFNUilPYj63aGx8t13vCLxz
znwNGMazrlUPCcQKWolOSjCU3WJYdOAOyz2tIsjfjuLtRT2aYinUoiwLe/cJKMcz
8Q2hjhU4FjeMw4vDcVeO9YrHLXuRZdd4fLGPrZpTSDRDuPov3INMDpqZ7Yu7MSYS
OLor8yxLBOMMwcXcHEXBbhjWtkXf14U4+woB0K/uenc11hxoRLDtsxJaTraBuMjd
N5PlLudmdtOq+6CWyMwfEWxTXwP7f2m4FKvkDlhtBuCHsffDQ+bJ1iWMVEgAQuzO
fN6X59lxf5F3BRDCmqXkPwQDfQcuDlJahp/c8OOoAYa8jDe24jFSkxapvMYeOTUQ
W0lVVKtWvUDh2+CX9OSbY0CDpO6SPPMt1d65QnU/IoV7cw90N43vqYpU9C+N+7xU
lb7q276oqiIfNn9A/iVOMjJB6iiuLve94vGKQmeyPV7WZjSGOfGOzRuCwz+rdHz8
7zXk8wWBlvIoW/fdl/JsNc0knyL//h05agLQQB9wPu4kHr5NGFj7KGQwxAv8LE1r
wmVUfPNnqmb1rwhhAfPNR+oEPQvykKe4kLroG+h6fHkWxh8appRDFjYvC1OIJtBR
aNvrmICv/AytGRyRtV0n6HZTu1zbYgT9tchhDPRsZIOtXKbCZ+lye+p8hlgplvhm
Y+h7SYv+Z944paQjm36yVGr47ugrg8ABtGuqGmrddRqMwf8N0XVxN51oBdBBQl/I
bNvAtmFeRup2vqSD2pNpe+t3qiDY9a6lQgBYxvav7JRXohI3y9CjG10Q5xQyoMEe
2KrnHXiQHfO6HEQ4iQNFbzgdwEF0mHHpXgjR4+23XCO1VfXg9bI3EqN0TiGMyiSQ
PEmJe2QvExC9oyfjQJZTsoJIB37JyiN+0l5IVIwrE4/hdVusmlNKDiQ6d3KPO6GC
tXCd58gyrutTWzQzdOvVDzQzk9vykH1ekvWTCSR789hzR0q1/+njS2hIlyN+RjdP
1jh9Iez68LVgTWLymiF718gTrwhRlYBqw4x6+uIetp08azPmaoj7lMnLY4MNIaeu
ZdzrTI9PU7oufPke8RwiCnR+6+2j5x3ADDOzbmD2rwL5duO0G08WkcXCKRf/LPQe
0bNI9sDPJdi6tlSAPZ0SoiWDNaZhBz7AQ9uGAh9zkhI4JYd/YctymaOPwrBmknnW
7w8n8eAUfpKXk48SENTBOMAwvp55BXXrrLNAC9tse+LuDGsrgi7789sE4Pk3tQW0
yR+BZJxEnGGD1cAdhHMLV3DYCNrv/DhvkEDtUJI3mL1A8bf6//vqmpfJuW2mRF9I
0SFcGpFsklLqe/FS9YB7DWnxtxfRUDzuQNy+QZrCWR+6IrBFYUm3cPoHbL5ji1MU
PZfcVqglGQkz3xrB6ENaEa7rH14/6KovMWKiOrxjMpkBF+Hb5VijI7oApwcpz0KD
0VYJk/1UOi0d1lBclg9xwGDGvsN+ULeN/Lx4IJVPklBuEByPWMuxnnLlwLGTxY1u
5ke+77CcAPunCTD49CvVI55tluXNmnlAseqn4kMB69+egeo4B/L65BDpugLMxVQL
w+4Rg6CKv5xZ21I7IB9w66X1smuhRYFl3Yxi88iVH379ATJviqPsmPQlWQtG3gwR
/lm4f2A8+u+Q1hEQVVw55gkqilivE7LEkwbGSqWKcUPEwjVQE9DOwhelgN071vl6
B004x4TI29AbAVtgU0tfQS92/eZoSwooD4yK5EMt3A8rLRTeTjtMH7KBhhOn8uKV
S5cCgPwECpVFXsE1BGDYfeIDkLzdUi9wrTuHct7jDS27HarWTKWtu6Klmx2J9yGq
Qt7ljj8XfzaRU1fX/YB2tv2KdGK/8j7J91U3Dbr/s0jEeI0OscCAPPKaJp3biLe/
gccuHnc6molklPYW2Zn+w+TnOxcZyvx97mCw7HgqLFBlF/xOFrTEnERVNZ/XoE1W
Rv2PgvGrqQ1uMA41Szvr4up0D9+yyRbKc0wl+eG1GsjzX/eNlwWxx4OFQwojl2+4
mtAEQA78TPINDJQBVGRrbzfb2N9Oif/M15R7AXqPIKeG1dUTHxdbwMbo2StO4ttC
iiwESlbKOGWxfooCvOLckr8TXh/vh1zBjlj7n96QhSDrHjuzXpJMRVbrpoRKQ9vW
0C+OdZJY66NcDZxML2HETkN3CH2SB3sqMEJK8tlRCF5PxyqneD56iNyU2vMp/CUl
adVqVS9MNSucI/chIPtZL5BQ7vHRZskLGXUfJpLgHqRZUGgX77m7IROVjMIj8dio
KYrqrjwGoOgQJT3ZIdpa1WJ50OeUNCzfVwhxqNvZhlh4Ek7blTRW+6TlXB2bPszG
vTC8BV6uijd7RY8k1I4YIJ9tIc9gxeaID0DfZqk2ERZIhpamOBAyuwExPLn0simO
d+UgjeqchNcsEvkOy24VS+Vg27tF9Jpl2VJ+F0/5UlcS0rjZNhhXJqyGlPyE49Ue
UOrg1QGqkhdnFx7sSkDiI+NuxCxrZOB1VpQN2YkEFH7oTXxM8VvR3/wsvndLSv57
P/KWkFyICkk3A8wrYL68Y3mWrMMaemgmpYj8BpntaTiv0i6qafytw98BWEgUjtwf
kzruI70/x3eWxh+xHH67l3/lLqFg/hENtICnl8GGjMuUdy4W7Wez3rmSEbjpSlao
0Gw4caYTKZdUOGybn7ouAg22PlemdLpogklIqNzxQiVQOCKxLF5Y+okc0wClatnD
Ypt17dkvuq3mAGMH9Gh+I0suJhz+ZHDr59TICMuYe6wrtQDOpED+X/HWMWRQKhCZ
wwi2+Fd/xccvOCS3xbD4Dn+OvHM3jIpr5sYPi65YAOWTm6/DF4IgNy1L2WICyjt9
Nm1PeW06muNRsdFJcJD2inmRRMb03mPoLeLk/hXB/aSaSXQ5L4o1x8odiffOFXnE
9ThSbqK3lB43+Y4xIRJzlw7MLlyouQBO9D/h02lK8HDzhbAeMWascLr+CkE7QXOZ
vG5z9n3/yPEAJbPMtBf+OYUY5unQkSKTU31t53GaD/1MfMzPstMGNvo8vy5XQoQq
teNaUCw+v0JMlLgowvhpeFjMpATggbTZ5KG3cRMoQLbF9riEScLkQ882QvO/Y4lT
gDQTSJcD8an9o9WRHSjQ60JPKpPz6aVJ61ybOrnKjzS2hlY76DOoQHOkpy+wwvei
25Cmwy+yJnNKJU2Ruu/IMU5+RlZHkP9Cy6sGPIb15sY7hgY4o2U0EHw5UsRpz3gt
zITkjDUuv4t8J8/hs3XyiOBTCEk4NVIIWSqCRjAPXX36DVbW4s7SObkwQAogBJi6
J0rpkeuZPc7rK5XSE6GYF0KGw2nW0iLvEUpbsIZ1cnOn+qhFJhMPRQuOGZ5+Q49H
0hE6WCPcuILMikXXS2AJXQ7l9WwkNY/bIKhcn3taXY8trD7HtXc0hLb3Y/xhQwXy
R9NKmaxEzbRMQ1j8JzXdB5dy9uA6VTQ5Q65ufKV2tE4G+BUuSen4oUx2P8Tw5VnQ
dDdYnJa8dZUZa6ZL/VJvcmLyVr7gDxWnN1HIG1CVq69LLzj4gDUteuHrjZbXz1/L
42/ZPpd4y9DFPVHFJ62jK1GyDfx9hzoUE1Ec0kEt4826sIGFtsatVTwTZD2WwqXe
M8LbDQAgmxDezE1AfPkmDluKn5ptTak5/lnOo72q4SUVqPJl7G5o9YXkOMKlfh6M
L4xfFXAxhKO3LhO2UdRUadCvn8nItRQbpEwsM/+Kco0nfa9VUMFec2khdCMzj7+W
EzFFpxuvIag796WnxQcf57Uf69B/8KekNLeZnHP455O1S//NLq++sQdjEHccH265
8zKUtRmJJXh7QD3mWjKQuJZ2tr/V+P4pYsEuU96TNYg8wXlYn8HODBxr3zzV0mwK
NNdB6QhXSX5QXQOf/fr0lLEAWgsaRbvIhblb+nvOs+DMgF9MJhCcj5M/6BfR5ICm
1GlASDXL9vWh7YEDDNWwkILSvLXLEc5qFkes6DCkRa4J5+rMqKpOQm9HzOtQ3GMj
4Gq7zqI7LWQfZO9H3J4P09uHjx3q2mWTfzTHWArc6pCbFtvrY9wijTrtrioxunHQ
+J1SdEwn7UnzSCBnfQdLGTwl0rxvTvlye4dlfTGjCL8IAokKt/FmBjAk82+qJ8zQ
HoKzE2AK1zurpZJ06CKEBkeSTvwx/LYAqnj7pV12Idm82trBG1h+FAsBhwzWr3eZ
oUvoajq+e+ME2iTFhlqFF+N2T9v3i9ZIJv5zHpT2+eaqcGTEmGDQJ57ijDlV/JnC
Mdzgo8YVEuCAIYDQV53PxDrv3yh5v8Tu4b8OfXgxYbIo883CNA/T4OyvGfunXGNP
q/19ze9sjpXldADd2dj7MIIJSONN30O68a3gfzFIhYkAraIwk58e7/ucoHgustYa
16V0Lq/CD7j8RDn7G+CPVDVfEDEmzEHh0sQMgJWrywLL1dUoTkAegUkNeQqNo4dJ
F0BMAx2PrBspx6jHNza3ufldi9wXdnHySadBrMiEA+g=
`protect END_PROTECTED
