`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ct2vKSUifDY9/wbePQrW8C3GWxaJ+hxDSiBkokWji4809m36d/PeCdBg5nuhU7DT
TUK9mlmZVFw5JKRrnvuWvycARLh+sTE/tH8g+TIaqhGJou17yGc3ZKerhs4V1QU/
9vnqqKuWtpdRDqQx+APR3FaSvCbE7JxEKaQWQ4izU904baOmgVBgXTte+b5se3Gz
vAlRDONVugqeZR9tm/MR4czQn8gJVodtjwtWpzDcf1D7gmXBhp6NtT+T7p3nbtSb
YDalS+tx0xFVcYr083qBewBdlYd34SJuC8Byf0FPaxadxE86/SUuhFqPT7wGaFqH
0MvURFeexHQf8oHz3LG23BCJ2JUrKRV8Axt7MtliDTL2IUSJbBhasN2dSx6tN8eG
yjdD5RtwQfD52wrIECecHxn8JooLyiiRhVS3lxiI3tebfWUUAWtRay4tuNn5UAka
RmNNb/arlbMPZ0rBqN46FKSgPmxEiXgis0xd42d8ejexfQ8UL51jJYSAYjEfr8bc
NV58idiq1wQsYfnjI+UjU0Ig5gBm6YoxjcDQKa1VmmFZ/g54xKfdqwLsZvLi3D1Z
lEyMRrhlDffGhTmCSvI4qKVOncD2DjjPW2HJdCr+fQloDHxkDWn4sVMuCWufXG6z
oMWBk6nx7kn0hp/BJRb6oJeEaIR7Gb61kgaTbtER+AvIZ2Q6xycQnrlkzrt1sx+0
3Y/HB8fFYTA1wntK3sSt4GSro8yaD7JvRRtAGWCxm1k=
`protect END_PROTECTED
