`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zxMI2+2BiUE70493Rka60s9daG5pdb1iYPcYQA+9wXUCjlEAj6PPwXc+WQCI4mub
E4WvcX2LaO/G+M+w/2spzhBr7njxQ2yCHmEX8CCEuoECHjwQRu4Z4YxgAZfcVISe
Kz9xUF/XKFMRF6GZlCwUzGX8UP/oK6oKCIT3/ZsoEuiXyXelypmgeQ4b57jZ4GJb
CO95EYc0mjqX8BRh+QA5Oz4mo3pzZltVlRAisRdsTLSyignTXV/mjHqiCi37uqyR
5ULqLXRb4ASCwPcKP49dItie4iWhm0YdfRfS+i0bX6ItGPBmrAxgz7guBRDC84BI
w5Q/HcHtQRLEAZ3sIhx7Pr3XD0owUc/iPmwePW+gUMRgXA8ahKLIh987+dZn+YrY
Fd2+Z8/aHVXW984XUJvTKLN2JiFkmeVDVATrzKSydJPmyKR0Tl/6uj+aFdt906bO
`protect END_PROTECTED
