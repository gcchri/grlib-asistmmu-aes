`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p2GGypw2DqYrKlnFGYQ1NOSYyykR9jDmUTjFoZZfp9x/oae+Bvrgqy40BUUFazur
hZHaoxOfj11kKdJZT21t0Wckd4iPpLczx2tG2gYjpyuIA5k+mwkoCXXd1eZ9jCY0
RqOHaTcksyZldyYB+XJ/+4sltAXV23FWSLxdI4+sslmZ+LxqdC3zLKooqqIQkSza
U+/Z6heKQbjYO7pSoGtQs6IDvARkiyhdl/XsGqMat6WBJg3QYZwRGYfylXw5oWue
yFZCTZV/2FwSZxMil2CrmDMDWau0Qr7yXanmRv/oH3OKf9MbhS5wsBr2/qrN3d06
tXzoldWqzvzaQrdkznor5NBqiZJxjQnpLffgvc7F3IxOu0K7UsXZid+Tq+NHRJNo
LAh2qdPjnagl2ckotkqVjy75V1pzz721hPWUiDo33w/dDUtwsmM3D/Tl9pj/K3Va
`protect END_PROTECTED
