`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UoeNTtAAlWBo3xscylBeS3P5+gwKHTYE9X0wHWm9OqdJPRmtFKuTK7FG1yQuZ/1t
Fi3KHP27r1RD1EbBRl1YmSaaNDGqQ2vHMBBqRtZWFJbPuYriG/2VMXQEM9ZL099Z
m/s0SwIJXwD/RTZMIF924vaa8eAQXgH6bJUrfSJsXAbded2QRqJjhBjiJpbnYPZb
ug3M8Tdn6sPhsYyOPQENF/gOgJoLZY7C1GiitZTiE0sNC33ljEKSH8DAEu3n1nSJ
wTXxR6sIsirMPiTTnNLPhbrxUURiUROuzhfWVelvzSsaNwfi65/t0YLjHvhHzuWo
ZNcPJSmG1ifU2xUG5RsmC2nl8GI0UcGdReoGzDenz7bJ4dqN+dNMBcYevCkfHgDn
MKPMAHV7pfUV/pR4/9zo9/zyt7tPVoVzKCTibl3Dh6k=
`protect END_PROTECTED
