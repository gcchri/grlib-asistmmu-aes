`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vuaeNe4qzC6R9xwaDKGQr2u0YXlBpHUFPxjyhqi+cpBUV612gl/Bb5W3rmwqkLen
Gctd0XhW8YpwWsupb5UtBdaZZdj1bwm4FhvrceDxYlVfBPbwOKJbrTkcskOWS7Xj
x7VKYp17vyYPiedWrDcso40o9iZvsLBrkJHoewxJ+jm4VdT0acax+usA/iwOEYVv
e9OfIrlXBSk5areVVvX/NAdQy35tLDF72KYarNDFgVan8eKHRQoFTUbZh0OR1yp/
lpq4u9qFuZvD6Y5FJ7JOlTpV1uo+SJklBYbXjvSB/ag1CYDpVnTgwNfjkhmlzqbF
BkHbWNgszJG9y0c7J5+MEwTS+4zsDe6Nd8eMBeIzlGfaGHOjBWMZRCQIYsoZR992
QFDZsIhKpnFb8W/5uOMF23zBQz0q2wIruvzVKehwvssn9uTOAyE5XIN0AuT1lT8s
wMwq3ev3BcJWua9+4aPSiSeXnt7CEZajR+4EkpxUnFDYDFc17zHxtdV0KKU8a0dI
80f62OQtLnv4FqRMFWPWsQqlKeqhd9KXNrGggwKPr8tOZ2XECucBGspXqZd4oNcX
nmj9YwdAK5Y8ZELHhMJ/tkeVEvd05anYeB78DZVw9cHjvuFfaktC9D4d7/Ldu26K
OtK2zfbmEOkIR2kWPY29B3EjlF+xN9qG5Fmg+2FQVdpHGSGeDUiowEJ5xZXK7I/L
GeXBECuOSFSfh03uzSCBPG1ivficyw114RToE5zB8WYEgf9I+2TiIwi5Cm2gPQHp
SDYnanQ8n87cr7CzDxNk74qTi9k1Nh863OWm1SxwoUg32KpvzTwPlgTGQUclpe9W
ghmejs63EMijU1a5LFREc87+6xS0bgCnE9Vx3Aw9cn2YW5Bn9I7aFT4i3QIoQgCx
x5QF1G1VN2RyqiH++CRec4oFTENMa6SdSajvG2W7cWVCA3ehGggIWlF+ieZxhrSz
FprBJ9ucDZ+Akw40rPrm1pW+g+QBoFs2231NHeBzVrl+1XRNUdKGMj6HAYo/yp0i
uMnMyNELGnTl4aPKOrWm1550DM6m+fUq4tvls7uqWuIDSQPRL/lOW45q6v/6DR/6
IzP9Jr6PCrLi95aiumRJ3Xt0KIWNv9rzzvopfJXfw4eaetfLftR0HnsYWhEBVT5y
pSEP2oW+Kf+Wbphztgm63xQYgpWi70m7aujetgL4k9ZF4o4BcrOeuB5xlgEd0Avy
DL+eAELCN5uWlXfOKXrsvkziUXol3EalwpDPxkH+Z3JFVef1yLrBuR6r26OfnoBZ
qxFMhYDXUmZsM5q5oTrqVj4a37jj3uQJzPAz/hGJ3h2Em6JDKJ3RbJAVlf+Puxk6
w7KA51sF/Q12xt689cCnnuLZgx5Tbx1gc+3xDirGAFYA43SrYIu2EmfT8fve/X4Q
pixXS8mu5xA4oIZC0pnl6uGjplXfoEhrAlm2Zq/t5ZcXQlS7V7Bx3Qhvh4jhS6Hr
Ay8LuGm9L1lp1Os1hY1qEwhp1vxG5KTEwOCHLmxOWniJVm/C+WKp76oVHfG/no27
cUDCJqiSPFa/78KjMe/2kyEvv3qNL/Q5bpzwtOXIH5imHZF3IrUUULirnGI61oYr
itpQtFGkdU08ChHC+tq+BrDXzeKye9URP/b1D+yhQEiVbjbCqRI9G239oAIDKcI4
qtCHmYuncY9UzhZxliMU2tDIYOxUwnywU3QZaiEkq4iRjMnVx9yBK927TGjSDi6a
XzGryxGoXrffDvFaeqz5XajLwxN3nmj/Sw84bGrRe3LKGE/v6qFHOvXRiHBxBHAl
CMZLrPqXi66jq/LcdMSAr36Cnj2a/nxa1zgxhikLz0TWlJ3YSH4OhEdMp1DYhTbf
SUxlU8EoA2Vwk4OAtLyyC57g8dFUV80CC1LpkT95GBg=
`protect END_PROTECTED
