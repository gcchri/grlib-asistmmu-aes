`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/xaz+4T1mwmanojCVv5snjI1R3N3BpXmqLiY3roW8sVE45GTCuP5ahjjmWY2Jv62
EgZIjPc7ppErKT3buAp06eDF6NDnF8gUmiZlfkmxFHoxmZp3u8zOu/NZFNkI82xa
C35ee8DxV7ytUOIa6S9kmOpci+fMm0J7xo0EZj0pooIh6yJ+y6576zqwU2jVM02w
wTcteiOYsb3nJ0ux0Rniqkslef8uTYvZDkjm2Xbnuv0ZOrRVS9X2fyvU47v6Qpzq
y99OoXyAX9B7vWp6Mzxwax3CZzI3nEYXPpn0+dDoQhMqzwMAIbuCJh5/VOw9Nm7i
zJ2Ui5K93QcFJ0wnRjp+hjYIqZ0LI8wBQSEydfPK/sF5+5ATWm//WqeTrc+OLjGg
R4p5/bpXOIuzyu3mBbtzqV+9nkblMeP8RU+14lK32FSwg/Earh0nTTm2uEZdOYMR
5s+giFDwCycoz3XmNguW30RCYBZY6t4KU/2au8DMc1Lm0s1EU0axfYcYtwuwVro0
PuoShJxRYdW6gyx/RgjdwoqYsLks/f1bI/kDdfPYmUjJIo0zq9dL6zR4SCdetw1i
Ut+bQe5tGuI0ibdS67fV5KjJS/bQGWWHBs/CxOyb5Zemt1WXryTQbY8H36+ZIWcw
zeSqXq9lJurN8xvrKTFzbNPG6cBhiYHWHzqHy0zLjCWK5gLrNRVdDWnSpOD2knWH
IG+2aCnQdqhSibPPsSayEA==
`protect END_PROTECTED
