`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MLIES6jt0SSPFrgWoAtqwroDEHV+/l1n9bEY6M4vOyxdbihCireXsVO6u959xoYk
+HdSTNC8QtYvBWybPq2aW7GAUF//E2jDNeRDIrLe9NAr6zQssu6qnCj/AEF84E5r
muKJRV7rwnPEUMbntB36tFD+kw+KNHVG8SrvZDv8t14l1h9XGzRyHewEJ2ByHdeT
0mEEX+I0+XhadcbBthUOlGgZq0D5A2ZRER03IDn+0rQcpU+RGuE+Ye00p+tzRRQm
HjAVndBA1JSvR6Y9tYRfcu4n/J3dcDkE6+qA4w6T6OMXQmfk/8DtMCmoPE6iy6LD
0e3+MnrGjbq7QIexM8e4I29PEDWwpaj8HVbmt2KNm/8MdaH82Gp2IPOMX3Oz4ExP
a+lm2XA0FjV2f3HGWL53cQ==
`protect END_PROTECTED
