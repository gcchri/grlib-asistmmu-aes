`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
meEA2jmVYm2neGAnxXHMf7J2bPJjabkKfmFLrPuz70S9+lqZEEmSyzj3/hyCGSsT
N+rNGjjbhTqmPmxKvv9Sjgu9TerwVWTtoLQ6UNqXkiphT66KI82VcS544R3b6Az0
3oFe6pNoKEJmMzqDJyQ4Bq12uCXOybrhigynpBX6ZsnpejqeiJG0Yn1PmQSBJ0qM
KC5ICFNhkSq0Pe68Vy55haBPYygXFZ2gTUSsXf+Vr6f7SuBXSlJI/CQCNmsHPkUK
b54en6MDxcsJaccLEdvHZeo1SUKBpxuwMhvqEHEluv1WZkeu7fjczAFA1e1i8v2s
oemfK7bZeuhF+s7WWdLm38tdB8MpR6VzKv+iBvVSIUr9g7afNGtjBmdHcszAgfjH
0It9YUxxXpC/HNpehfQSdu6RiHdv987wvd+ulDq0SJcuIIVmCgsdG0+ALB6hdCje
T1oi1bniTYRf9iDRkO5pepQa/FQPDXqrQTwdEKsuQGWKHDQaUhTXFH5L6JagTotT
dMqdcLqUE1G+4OS3JBePJJMSlxeWQsnCdcUsUVN0h5A=
`protect END_PROTECTED
