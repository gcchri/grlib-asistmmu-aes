`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0dZ+lbn7H3X1AWz3AHELD2dCG+uyLpLuqsyUBB+CTYVFleoWaWfPKWBOUwqgvOrz
yPhi+IO+dQSojL11kxHFl4LcEjNe/cxG5zb+v/X9yVZhW/aYLrnoIyVVe9OMwnRd
4k5l2wQ2FJL6Vi4cF0vCtKIQkaHCtFEA/F43IXTgJnGXCl81c+ZHxAxjzYuXhwPl
MN4mIYEHx5t9ShnmTmWM6npW5FMrOYVKwVIIhHEOMnWJvACV29o7D41R2bkyPDtz
asJSzNsMQ9AE16JF4kudTw==
`protect END_PROTECTED
