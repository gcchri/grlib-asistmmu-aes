`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pBwhf1bfyBgdyKKq4qQaL7oPpvWIlsYwP2b96aM0YkCqdHGo+dPEzUsZCgEopyZZ
KbBNVnJE4xZyfLwkKltkHRcLQHVFfV5BYpbObf6zP1jx8qufGbK4zUwtU2AEFEOX
QtfZFbiMkpOnMeifIVlEUfeKKJbnVBJ7OieWPjF0ZJZ7y8DwwuxTGoJMgK9Vor1x
RlIdHI47YR58rfKvLE8UxYesUdugyosE4egt7TIe96t4ZO3BpnbWRqawfyXhdrxB
rkTwY998+FjUIhOY8Wm5HugcH4C+TwnrSfuUschAeAfjRqFQbrTo4r2OntQ9RanL
y4gEunCYavDHmT+e8SjSGlMXDPa1QjVcLFWKyqb08zjwvrfaHiPmLj+gsFcvflr+
5lgt92eJp1/ABFSOkrErYVMFymeralT9BxJgp5ZoNDDn/6uO8TcfHwMdWg91cbeL
Mbk/wmFdUwVZfrHHJxSK/aBWC1tDgvYP65U/h6MpnMDSKr5nj1CCT+KBnpUii3MM
yW/EdoOnn8b/ifpjJdLQRUJgvitFXfcrzhVdg4Q+gzpW0XYWmo/RFF0gEqQ2dQLK
fvlEwP5/50XpQNTEPu1LtXGtPpFC+0Uf2qjbBy5eokSLLjibICF3/degbfsD5hLA
xegJcb/BJM0U3OzfjxUBZRqsEJDXyve8lSxxjpejPD3o9znIsINu2jqftWSPz0cM
/Askv5yYR8jorMJURm6IrysP40DzT5UBXNXqYGDKDQqZN26qmID55CYE7UNyd5qz
KInkm+9dUt3oPj1ie5YAyIupZabk5/tyfKKHVyDWpRx8RUICapsiZJnAUhgwS62P
ugh2a6sKFpzPm5OWYeLHU9by6MfzsPulO7GdZ4hftH7Qc/UO8Vahp6VPOt7zudYt
cqV3TDRr3JT+BM/FBrvqisEXem/TrzQ9w2Zt2yUk3J69rcO/QNkZF5XS5qgxlZoK
ygPETWQsxBOIfKFcdnnxLCfr+f61whWFVk1AiS3rTItQuPYKgOWikNQ3SyfQQInd
DDEyM00ijmBv3gazFwpT17EUJkeXeX+lX6nIuShENy5Qbhp/yPtavyBuVRhxWr8d
UTvp8VavvSj1qLN0NyPeR3X/KDlbKS9+YOu197hBdj3iYvqD1KFtlCUJ/Tcr/eJA
YPoMuAClfQBAFPkeUPDNGpoHo96kJ6C1JgnNvHE4QMy88A0mAusfoFDiv0cEp+mS
nVckswZp6LOlV0w4FaMC8ZYFe6vgzadz+AbOI9QqFtRU8qen8H41JjBuObbZwf1F
9ktlGUdjnEh7rLW9b5vT8k9MkCEzkUkuOPqd8YJGOAkkn/9KlAM1/7adQdMB31Yc
Gxb436NC/pvJ76qH2uQMQtHtc5EYQhhoiOGs58xgIDU3pzQzsRMUSVzvzaII81RZ
P3M+NHHfFgR/IiqNnrCWKLA33U8Hr9nS8hXyaRQ0sBTcJzTnoN3Pm4eWEXam8aTZ
ENo3jSrrOmr4zMb9aJxmviwnm4xocM0cX08U+IkIZz6kkOGxgwjoocy6uN4JdnPg
UbSkQhwow0sJwHMIpAQKEdbyVhyN/kZai9g3MeOxD45SJ9C8vMq27wo4dulwYZpG
rvVVRXJLrCCUVLsonJxwY4PE4SQY+Bt4w/vQs8bhX4Pp3Si8iSy0HpdSpPriOfPS
a3tONJjPm39Uydpjtd2+Bd1EVwqEPaNOuei33lYc7Sh4dDBlUE5GUwQG1iky3A4n
7PrmIMH5+dsCb3MA9pp0PHPph80Q9EUE82qJ9JrKh0kloJ4ar5aohazlZRiCGpFH
g68KmI0Yo/XRyVJJkttQzxFb8sit8G/GmOQC2pDBzsrws+5xdyclcHFA2zAds8AX
7gHZnpRqD/3/eBhTs0M9YS5d1hcVF4DQiOV2ETJoI9ueTDbrQnwQ8m8LFLOHESP+
i/ucFFfkuNG8p420rHWI3PCFL0E2WUTHoxpR8CF9CN6yM/QL+jaDi0Q3pwi8Pb4D
KzpC8YDScEkXGzffj4PH3c2kNYDFFtPKHbRMHur+gGl90NVKVmVEldkhpaKRfHa2
wqJ7SIxWP/s5Mrr/2+DsriZaTOZO1rXdKYU0tnuO0nOJBhH5Fc8qjOPFomkZzc4v
AL+yu9sI8bYdWSs31viQormmXJDl7+NDqpL5LyUz2vsLSQ97Vyl1Vrd9Hdclv8cW
v8ldtrWm9AIAC4UIkDKwD6XMCqsnq3jN7Q/mkTWoHmyqYvGfyvYCo/3S27R956BB
gVe3xnAXNBHG2l4x38U5JkfUBD7b+Wvw1HmSvaZjUVZlCEvIWI82Kbo6hedPgDBK
gZo8HmIcxrhKa0XJTWiH37Bg8JaBYqRNEYw/491SZl32eJ0ZcMJ+rK9G6QC4TlXg
421411ify46enqcHxRNsPdGMKBOtFRg71IrrHSgyLO2KXYw+0IqqHBPenVg/vF6Z
0xjKaFcTElrSlfkaolSlSb4sBwXtmGt0YmNfzZfm/VeB0iidzO7XFoAO7awxl9AI
qWUDxVYN0PxuWBzOzJ7Y0HXPgwNq9zW6xj5M8KBM//kuN2Sd2ByUwujx7jrVt/QA
cCqxiHCQ17l/WVLy1ZlBUZnXccBg02j8SpJbHsj70RbjBeUsKXHKIL0keoQuYq+C
3GIcIOrlz2HoGlm+qjZiem/pg+wyFHP16vepOtGVSjd7jL43iSo1/jW05urxMpSq
ngmIM7GSTZRiBkG3nuMV5HIyQ/ZO/lSulbfqBgxEb07fE8oIil6Sy4CkEVJjku4u
Hiev01A0OD5otFLB9ghaFcdK5P6r9J5N8AkFWi49iLHuEzqH1yUqU5tpSijHDiHU
yzbTuEzMLc0Pzr7XrCnrBKBYPP2hdZNAOdkv6ZcFZq0Ax6j+zG6XlL0Mv/deoJQN
YCbYyiNEYQMRUejQKaas1BN/m51RlKzGoZst7FbiOyJQsHxy0ZNqrEjLOUt/Eyau
BxeCEtLAq4cHxSBPUWWAKxTiQ8o75FyTKHIa0RfMpqbbYHKb3+BMwoPhzp7tay00
fA0Qid10tnpPEvrKnYrKjbOnjUmWSjeEn3JhEFR+VLFqQgKB4meug8TsO2VFdQSc
8t0LrdXIR2XcF3goZANfd9izUKgpXHuvPfsHEEMEbf/TCstLk0k/5s/DpsGgYQeA
s9zlhq+P7ONoO+fbNAy0eKsBZ+ljWt+4GRSgOX4uVgP7HzPSVesuac4ZTOz6ENM+
Q592FbQtN1KfN+txvGj28b78PYbknrB/Sc5KC7nt7lixbNzTJ+Z5QEJZ94eWmyfu
28a83jHfZJ+N1nXXAFtXHIAhqe3bSEzBRPd9p1+MfujqqPcHvC1Yo+pfwweygTIS
KBgF+1JixQYPCIt9tzrR0Ed+2Tnh+du1BsJ2za5c7UBVYbyHftUX4KD2FrJfeKm3
1A8KHlBB5EDad3Fv6t2IH1IjwZRkx30af6xWw9ZZ6bHVKYFoxXCNeXanWqU/yStz
cVDk82qmSsrs3MKEzr/2oBXJnVpGYnKLJdkPgR8tLA7k4veXDh22oIDoqNxcRD27
cjDJzWGJ1UScg7VvMVgU06FXSlUfOQi0AwcGgMXPnvp9D06tSa0XjcIQ7DV8/BYF
ljxI5YmHZqjBE2pyXnl1iob+ctLe7blf1dCvanb4Z/czLOWCXmAhwtb0gDbLtxOW
U4ff9oZfKG5aYbX+Z5m/j3lE+SmY70AnacT7BVAgqTNv3vnGPkHMqEnCNM5ME7g2
eSzCnJ2z7xbZ1pnLTVhFjnz87T/P0sG75bkk1prP+ttPdYCL9Ckc+4oz32wTibub
3d5tJiXDeUsUfa8cCopkSxo1v3VmyzAlsAFWdR9oSYaqKzVKp2zYq+otQ36Dd16z
TlsRe/fQLdYm6LKMAGw04lgpdxRXf4kCPjPmAPi2Ic95ot9caQQNEZNsskrDhF0C
R0ipn3wrkmnW20uYVUCMkiWE5yOAv3qX3jSYcfo1q2Vg1UoWx3Qx90AT23aSri7M
QGIS6lPqAOEkyLq9uxkYWEDA6NO91LY3udVnBDYRmgeT3wLYucY29luMtvi+iAiJ
`protect END_PROTECTED
