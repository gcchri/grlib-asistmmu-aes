`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8vdv+xy4PE7fxLAdBRB+CBvuYLE0ZC0M7ZOCccPzQq9G3hczGvutXTiSrqB4lsW+
SBrklTk9NlZcv8ZdsPq4YuRtFDPXqYoS8EOhTKpxjZAT/NVBdYTFHhxomcjkzaGY
uHWqk+RcvuAvpAxqLPU3D8jF5bLYQSuFw9uVUDIjZy8ir+X6UWO5lMj74u6xOLZU
CjA7l/3h+AliFbBnt5+yeYVpu+6OvrzbvIcVbqo31jjLSoDQHKxItgKWnvoBxelN
5Hcf0vLmurwgS/ajiN4t9YSGplREPkGUkE7ako4wFNoM5AJVbVL8r7eJxXFKM7DH
+lA+kHyB2tP2XFKMLBL0phzRaJVHH8AR0u9x0VYRf4v2R1l7Rvkm5L9IlHyeXewG
9Z3r1c6pSr11LLM7S5ic5I9EHuY6y9UBU4HVSd8/hyWjG6p+JT/Qna4jKouvHhS7
WkwYe179K6JhOnnq6gsMV+5L/3V/Bcx/+NrWDvYPKzXYiHw+xf9H1tz4eK9+g8Og
z4p74enrfFp6o1yJGYKCCiLzSM8uh19h+cK316/mMG8=
`protect END_PROTECTED
