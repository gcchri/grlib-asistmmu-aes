`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NKOoM1X5WWm4I5MrUFi471FtxtpNJ3bdcA+4bu2Zd9HSrzc3A6qz2/W+Bkyb7YfD
k4feY+TSRtX5V5kv2KNTTtZZzB21jrI89uCqqyVC6kenpgB/iw0w6QlOa694S6zb
AgAYNdhAH6V+4EBUahTxEzBBRCKLZdbY3SLNsG7yk0x+WwHpUwEl2s0OhdzZ4qtU
zYeS1v8wbtYp4m7QuqePbg7qDbiIuG41wuS5Faaa9tLV3da0HxJ/SgUpmVy8R4OJ
qbZGfRyW4Az9HHGtcB++6zztmKCGC8BsS28W9kErnTJxzrXzt4ncQY938GpJwqnS
hKL7YdA/eEEzf5SVJ/ObsEOcXWFe5wPvl6AdOhzhJvT8G+zkfKAArJwHBnRNQoWX
PPnHp+nukIbzVzV+ds5AFyNtQ+9A4wMhHHrZQolWK4eHSkL/PPHW+IHLtErftpEQ
pBgAoXoVCMG5WjS82v7+2SVC5neSukJhNC6FcpLtcgquTdtDHEz283zDAIyMnMyD
+JsgAD4EDso4v8YytImnPMPlWythizE7HOs2fOm1/Oo5DB3KX8kcRJdmuRqWt7MU
KAIKQAKwHCXqbSNT9oEclsokL0MmH1s/BsOgQm2LBzz42whSsPyTCsaLPS7Kq2vc
2mPd19M9IC9TdPn6yZIqBeue1tI/TNmpWtRzPKNQHqU=
`protect END_PROTECTED
