`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tJ6zegWkI/UfAsm+6IgSKxIWcI0GbgtcPzbp6ZEiYWQreqBt/LB8O6ob0K2jysCi
crDVY6u5IVleRUF4TamA8ry0Hic1cmzLlGjIiw7+eH9kPZC3PHsnIBFewnvWD105
AzubcvDe2iaRU2+SDe3pAulZRMG1PR+sLN+NEaFRH8bh2BExdl1L6kuAundvBsQZ
ULrXs4BdZ1TieZ/v4JK+Dc1pjq8+HH6RqtrFQceXigogOsbWm0WdPvI6UJOhr9cW
MZsbza+YoigM/Kj8Q8qrhDeSWS/rs3OQJ5Q6GqVFIH3P3QdP9TcRiigu7OdNlgyu
A2Qcf+wP4GqrZsw/tX32Ms4P0VR2RoNLK11i5IMfui/BC0fvVo65G0o4A40QhNA2
iwOtpj75ifhkx8rkMXBCJYE9rRQLqjHKzi7yq+Yql7Gd8h8Ch+4kWE5lkYc2a71Z
tzJgljkCYyKFGHqIJqndKnrAwZvDrykvLet+oFdyIyi5RAox8udNu5X/gYav3lxi
Jwhfzg0tNuzqKQZA6ssTzg==
`protect END_PROTECTED
