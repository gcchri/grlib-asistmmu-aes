`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WB8PbHAHF6j+1O76WEnM+AqSLxY3QacvN8CflZ+1sWQ4S24iwIxgN8QqeoO9Omxr
LTdtt22ReY7scEsAMrlnHEILe2VzQumiH2HzUZtqzL3gmChxGnVuCp/cz+jK3tQB
HHl2DO5+WuIhaiCo5m6B6k8NVSIrI31DuBTM7Z4N6C9a5w9ftMFNG+YzvSSIabcH
adZhsqL/9XikidbGvx7TncpkrvCbKSNcTt0jVQNT2zXNU5wBa5j3sKQLTJtxRSr4
3Cra2hFM4MR1FAfpI7TVFhqmJAIglYHtlmJY6W7ruDpSe2YeMCJKLC3C/ujuw7BM
k9tNbYrpFLwk35O/WtOHna8b9cr8CDNjpXlWelPeglrZNIKF1rNvk+84DfXjoI6A
nPe+kQKah0Q8KWQkybbCloM4MDa53MVFKFt/fXQSoykPu2EV80mWFwlOjCK/wQcq
/0C8ycuoS39H8Tz/ST9lwLbCyvXblOQzunBLIxu+35sXVyOl4/Kgt8EDL3DJdt9x
CrBPuFpsErcsjp05BrXu73e8tQaHzLStDlAjaEv5ho++pZowC52jnMtjTZd2nSFy
5YLlWXXCv2p2RPjw6cXS6V9m45yaiesxDaMD3+riDkOAt7s/8ZmTX2XFUORhqWxJ
PFmNhXYtDi0K1XNkZV8EPzDoEPZGnmBrNlQXYk4EXGetXe8L7OvWbL4wmqpE02YV
UCSKQqiwKj8AmcU5flvWQBhlHC0wNAMHffOO4/CRpSAUC0v7PjB7LGoRIqwTD+M9
QYsOBTCt6hfcIG/CsdOqcPlPD/+WvnB3ex31xEkQht+z0t4dNhGLJqwgfXNRCdtQ
c7J+lu/lpfEq67lDu6t8x4ynOPvyazqw4nR2b8zVPTwaNMfXxkzfCyHWxUkg0xAx
tzK55ZwUcsgmdJ0ePo952Pq2mQ57bAtUO7nD1ewijgvTbPtRTwAIyAU0s5bPNLWD
m0mgD0jJ/k04RbCs0FH9h9Ua6WHPy3gS5r6tiAwFM3fFc9+mKdWm+KiURZxDV8zF
KM/jDWI80ICieXAa7WfcEj0+br1ZFNxLgbA77n544CY7a8kjMfLybIFS90BLL7mE
PIkuqxUcRxwyfVdInGA5bv4SQ+LEz9K8fRa77cgUk1vuNxa22PoZcEFXCBbi1XMk
aiuo3tSh3bcAJ2UzJEDSEb4OaA4VP0O7Yhd1rBvqKg/0FX9N+y8r640LceTuIKk1
p1eLvIdx+luQjI2eFFL0jPyHQJ28kN5qnm5v/TigVF0wIFF71NH2BWf4M4fYl51b
qekjKLEpSwErAEFTmB91ng0MgJJaBYhEUvycTTXVXfKdKEnDBJTvXg7BAmLzZjEM
lLKkPx2OzCHXmZ7I/OYPi3sPjXhnYyRF3DNjxVyf31dWElumAzEs8m6YAIi6vct/
ivPx+pfAXZOB/9WFX8xeDS0M2eo8h1jZ4WGK9NprruESowJwhK/sCpdRakqKMCDT
Ql9nbb7EryQs5+PEsQ3HR1Y7NaAq6jybtLaaQVYTn1k8rCTchNT2C+LaAgIHiX/Q
V9ROJy/eXg+ZB0auhQ1189A16BTq16cuHdyKxi7qziLtLeTUsi+/j80FeLNOxWdk
kXYr7ixxTiM4gQJNQRiDsm4pQ5yjMawfCNxeu+MTcMs1zBwaoDEEGbY2KC9S17Lv
QbjDetJBLLFXwWvRGLv8/MmrCQS+BBtLg2x3mVXsH9kbcg44TCZfUc+T6a518Uld
IWWfNPP1//H1I9TgXKYyiYBUwUCdOMjJ17LDJg+O0rTHjPCpecf6XcuPOye5Xmz1
dQmXmkvCiI4QQ1RM2oh/CPn1BjoGOhD+G5XU1vnihD0ACD97jfOsnOS6q5qzY+Vq
v03t54Uziqswe957zHNEKf4RrwCmT48dy10PN2XJZ3JbxozODkh/3RsHuj1xZ5LW
3R5YM4fDHdXsntmRMjhQf5eaViMsbRLrtSAAK3lXON/ODot5MVSnAHWlszA/Xm7Y
DIAwvQ6nHJCGDYpxwFEnM14kCPiOYySez3lYNF+s+STmLtPRBVsAaKQx/K8j9Gov
rvc567cO7miYd2B+Y+eCXfwDUlk/rTi1GdpuCZj+0A+oHMCym973jVFw5HhOPoa6
2G0mrk6OR9kt+g347bIZM2YTY4BamTkYkSUNVuS4pKKJ+kos10+oxJn3GmMRcsGn
twOkJJWNc90QsMc4JYYgLViBpj2bZN5LoQyJROdRAN0kw5v+J1YlN7SkWpqeeLLf
HaPejwkgZJeBmQBRrTpBpmokMEFA7wbLbxVM6nTQ+PfFXAcFuVjCG+7Sm5ckjPDJ
l6Q74tNft9zpk1PkUGg3VPPRn4Qt1j0YZO5jwVtUmvsD0GW/RuWcw+ePgX7CRSWk
jf8AnH1gjBC55BBU2LI+LjZnwwjsJZaUXhrTplbJEAo83vaEK1VnACh9qi74lEq0
EIb4caql1LXQgPfN6bT1PTykKf78fC7CCZtkcKQXElsDNWO3Ai6bhYjlkaJXrbw+
8tOe8dOs7aZSDROQgz7IpnOmvx5NofYaIgB93HwxgFToNSIRZOsmkzU+emFJhBDS
M0N0rucOGawfYDsZe5kRk+A2hD08zhcaYhTkCJHYfP5LQxcteUuPcpg3FtQ2xpba
d7uPjrbIGJCg2dP0mtvOfjGIenWKL4ww1QfE6/6NVmLzP5TOVZB3UIwhL6NWRrwY
YGMicmMcPKfAyu+DX0+7embTKhAOlIcsKtYNukoNwl3n4eK/UuO98KMLKjJu1U+1
1i+uXPZsxqAEttQ6kV9Uka7HyedoYD28djrfugHIkBZF5pK3b1S0gZEuN8sQC1VD
4HK0vMXZH95zIPH3qGnBzJlBMgDVZr8sIDqcunhD1XAI+DoAB+IbZsHHUOeks5Gx
cjlZ+ajndg0bQbOSqoEhL+XKqUDjG4yqXOfEnm26/0pGvQN3kyt7WQ9RJQSB1Bdo
Zgv6D02patj1MCvVrej+ckETMJjYtA1Uiv5/cSI3hnjMwCMdsTq33P94jGNUqKrS
NwHemnTv78J5hsFzIbfTA7vHzYNW9EK1TEWfMGmdogQPqNqRNdGTYn93jSYvaDmy
tUL1VC2Ndo22N7UlLaZ3g/dpW2zrf/U6kSSTnkeX1L9KvQrR5iwiLQVjRjYWMuS5
QYZOKEdsZypPDXD0r/90gFM7gyl3zh2wyWyiwoZ+JI3C9Qad4EVfB9q0yIVo6/eE
0r6U0UGf5BCh31d/k+QEIcH83RZWAgQlXbUN072ah/9g1ruSrbennJrIoXz6mbZC
N1LKQANSo6WHVjnhWTKCUyStnfU2V4TwNuDGiKVkmtGdq7KVTbyLhUWzctq3IM44
PW5WGDOIeZLx1Uv2PPk1/ATKmh0/8i97eGOokW2sER4koIvPCtnB87nfyRb9onJp
7dikS2hIH4BcbTxCfdl8XW5EVIb5xqDF1EzKsXGDKidmHrdN738E/hZNXfYGiWQv
RcnSLqrSOI3zIJ0oyDiz/f45Mw2vRfAB9fcmvVYDx3ABI1Ptfh+0IEVTnm0T/Z/g
l78WrlOd0ti9bOasBsT1TfnpRCZBVGNQgM7TDDzwUeZauG2zgwkJ40GM58HIASAj
nZgEgZbcfHCVAtEKC+LkeFQOaw9K4eIAXmCklq07YVybtHG/CQ7dCJp91aHgwYH8
CEr3VeVw5zNmC71hJtdyTQjt4bvleS4d3ZT2g3RpPyVM7r+tHL74wMnCpNmH+JqL
/acIWkGyJDQ/WQCYdAg+Vtv9nozJ0dfHsrAB3uWLyfKqD5X1WtZxqrhJH14iTMSc
LBqkjme7d7fmm/90jtDygxNJ21b06gPqZIKMnhu5mNw1Qp6EbBTDmMStJXeYK7Ah
xTNAtJnubdTA3GVatZ39oUeZf8FG105oygHyI8EVU7jI9OLvLIpJl9dOyVaIR47r
+pj5ij+aXNfRfd7YhfhhwEZ276sq6T3TiTVGwrMyG+8lLPNOysy/kY2YJw8BEVmP
W6+m1+DIlqrlibzo8Ocmf3bzC6MOsjHhmwDpYhzLE3nvz+31IKTUMxAa2RDiATdA
iBab8/POE3974RhVF2dx9iKd1hEyyy55GuBt3VH2HZ0C1sOV+wnaiwvuBClXV1CI
RbSDuf9RV0JHbAVlcrFsUdU0bjyZWj3x/29MzTqOh4jhevDmza3vHx80ilCZW91r
K/MfCQENDrnLuVDT4D1OD8y4A2z0KM/Hl5lQrpQ8OqMBpl1V1HV/8xAVCW9e15ln
pms6gS8lIi8E/qsPJ8JnPCZKUgL0A0ni73cGIsUOuqd7P50Zg0y1vtV5rYfUgXdz
quA7X1rvgUfvupHCwDaOxZ0suNiFqdRISMKDTiSBKcTiEvInxB9fM/Y38TIRNOQU
EtiWGjQLUP7P6l1enRAlsvuYz0dnJGPhsa8ReIViZkjdFZ7jLjZu4RPI8yP6RL/y
jFI/BH+4Le+RbgMsoe8IDkeCUu0WB4H47jeH8PfcyCalKioahWfQGkf5CJj5COpp
X7ru/lTVuFCvdiOfZz0AcPEpwWKVvTJJUm1GvP+XpcS0y51RCIyJiRE6o1phLVoL
gVl+EiHARkdgX+Y7j0vxbfcjSSBG+kikuCm0dnbCMpBh60oMkFOqpmslFYmtSBd0
+3+iWi3fCSEOcD2jk6WC0VT4DUQ+d09pr5I4fkZBu3GbxYyCvMuBicxjmE2ozJ0i
AOIehDvy7jIFrDEMAl7ASU7fTUtoHpAltj5pCHvchj6cPBAyPbrt1b1wSfKz4XV2
OrmQOwkygsJetLAg62am2sAL2Gv99Zta1YbMXIYCyRP665EAqwVJ/3iX67Zwn1nU
+BIQRQ168Yb4ylyTT86Xc4x8GcppnG53bX43hqBKHQAJfyoctJaN4h1fDiBDeHML
DND5jTQzsVYe+72TpTMdcw5GTaxsKH9ESwJcUYWya1SNhkpd+QLMbjndEmRuJel3
1uSbAE35ymJvB236lyRNrsJGrVtCCoi/k92XIHXMH/ieTX9Y87rfDx+JGn3LHGWV
TDw9zKM1IiXB0ybvJntScsUyo9+iZ9XmKWSG9bFrfrTC97lzjx5sJuyRBJCuKWr/
S6yY2FZfnn91Z6VlvYhH1QpguK8zY5Z2m5fpBSpZF4e1AZCRuFINGgRNQ2DMu9su
RXdRMiaOjUQJHQMQFe6b+mtwKZTRUMXXlGl2mb/SVJAfFBRuTSAmoqYAhWmg24hC
2jpq8CyMl3o6E4os+dMqhv3SPV1FcIfJDZt3i44HbC0tk6X8td486Q5UIE4ZEOy3
N0G1U5T6LRAqc5PNRf1ybitUewl7Gt+bVVeMk+QHfn9FXnHcCXVX4uG76QVcltv9
N+ESX2xQhm8eynn4cq5K8VXYv92NR2tij+Co5Hx+JtxeBf0jLCZbrEG40DDswIlR
eppHzz80PJj5KhfDxYtSzKNdNlFbAV9CXdDbNBO9VMG2Cj5ofDY/IoHXiZ/FEZA0
DdTZ9EnCy0TbaG4sVJTSXh3S/sqXXWKX8loHx9Mw7ow2+yVadlKzxqBcjsOF2ldC
SxAxVEmuHQINzzLcTxWsDGHmp/okK6I/vFjLuz4s8jVrCm0TbwEEQFnyy9QqVKiD
edGRkAY2qqQXgiW3QK0+ykHW14Ruq4XLtYBW6yZBjZ+1F5DmHQLbQexhamvnwePK
b8bl84ou9MKkRFrXwRGV3ZmoRcq788jpkBA/OOEO2fYgLJbsp43z099dgvsFsEZH
DJCI36Bf9UL5cwSmQtrpEPVPTQxcV5whKyRnBGQzI9MlrHwIJ2inthY1FwuYIOcP
tl69OapbV5M86W/PnIizon+/c00ezgSNAND92OoGbCD2mnUW7D3gXxKq1R8rlbXv
kk47eAiDGGuL9nKBlDwU+Y3cGuMiiH5pspTHG2fi3JkERxwLeDjb8So4pZC7CQgm
5/SJ8VvC5oiLELrDurPLWMqSq5wWZQNISS0KS/TYzJlRB+OFfRF1vB09UoXXXY84
CXkyTWI/YbmVBcldOUA8estbcKeMFjDJasptcvdAs+jJpur/u5hm/+s1HdDcw77o
skn9mgzcOpK4YtpWwdSw1tO9lHDROfvfV/p37FL6COvIhXsa1Rg1EUdcPc7+Az6b
5E45AtrGoP0ajipSmc+vBLJkuqQ+d5cm/5Gtn2OuPj9RnCjFJBkO9JS8zGk5mSi5
BSzTvpfGqd7wQh5UYlFpjTtcn09V/3ESxXVTE6eEzWNNFplVMQ5Y8Bwh5R0S/3eo
aUCqHMbdNRSK8HYP1ZTOvtPMt9lMKa/dpbj8SKqmSylw+vOGxQKVtvzrlpFQI/tB
7V3k8epsPpmm6Fa3gQkfVrPWJmw9RxULbyZBmZHtvbOCYFxxFqavhKuxzKNaPB0H
Ez1woVTiDGJY/fObxsLaSImQU9B3H+yOBtvTc/mFD2UyV3GipE20AwGVw1B8dVej
EpxHIUyO8i0gr80x2DENJc1kmhBBfvIiGsvZ2hqaryTC/OYtbJPguaipXLoUPNla
H1PKll7Zmme6x7HaPJ4SSC0f1GnFVimeBfv9iPotY2pAG0kDytDB7nCqgbzSClUL
FHBUZD2szxt6BWqXhNGXFd1oUSL0jfFBRsT5Ldeewqr2P4BM2Au9wcYZ6bDNlvLX
A1qV/igjkDC2T1AXr2ive1T0YePzYpW+2Ys69li9h0bjWy/YqWZF8xLB4tWH8iV/
Q/skoVIXMfBYwieLKHyeSVSpopeTc9mF7yIvi2Z2gl5G08c2rL+ofxqZcPm94U44
nb1vabPnYaHNEZh4HouxuBPXXdiupROC3zfOyBovYyswDozfI7Kw9gE7nKwapTBF
xhA11CwS/b1FG7z5wkEJPUAD20wRhIpQEYBvKntRyDqgLlYodrptWVvsgLxunos1
2X3nGLO9zl56U+pPgGzTMJ706wHyNjn8NIiq/BYcclfd1WKoAAiglHQIeL9iXtKZ
EZx5OuKiQJM+AD216CgaoejH2eUnLsIJVITXGqSh3m1yGzG2mTd4HismOUmWz+g9
xQZIX1J8YKnZ95wpFkmW9eMUKTLybXKWntps4iniRAhySVRKBBAgBV6SDF8dxMKK
MT8smfBst39gBRunCnJcKA6L8saVH6GK9IeHsqKd/OPODdca+cJd3wi3jdbhTT80
n1pi2xMhyTjHLpOB9ax4tqoTFhYngrWlf1UA6Cq0q8qfFmBF32QEwq3sgZQMLWcb
k+vwg4PZRrzIkLYMJO7Nov0qyd5QhAFlM1OgQfntwxsw7Vidrw6suuX2Ad5gOP3w
RLmgzUvJ3eBw4/mV2vKkoivplO33MmR997SGeooR4cBGTEhmAxdCrwx7N+EAc4ZP
KNXBmKsMqkm+HhEHhT3C+2AM48Opc5VItA/Pprmn22mFfggdrgDzN9mqE9o9Pbs0
ry7hng6y3ZRFdlIObAMu99jJ+95NAY3NmIKRdUxbmxP6DFZ7MTaIvuGTaOEtA2TV
Nbe7AgCmj9P1IusqvsGFcPnOmgVFv0YHMoNLTfwng+Wizoav02V/uYrSBPjsQHJo
2iMm4ivAp1fKqq6F9eH3tGgJpGn+39PAxLfWDtlwRIV4MK8qfvHS8kN0lTsb7W8k
YjuwzLbB+ZmHthvmdL1IOOw/oa3CR6ZG5Zw/pHsvXjGf3BaYNUIFI5Ib12QJ2DQB
ltz/2oJujzgr9WB0BZxwgpOz4+AdaMksxgNYPNiPprL80D8AoEil19ixTwe3WnNk
VaMGkIgvyp43iAgyEIMnFYJJiSHa7liGwUmffvdzKLNWZSqZVeFzhlmer1wZ6xuT
dk9X61r/BRbuyG74yTmSAWBaGNbXOADvzLuV1SDdH6rPkKqad/5z4GkqxWugCz4F
JSgdZCVGeY3cZ+WQHD/pQz86NT8Yop4mSJGQIIcROr14Zxceg4H2bfU0K6AsuX0q
uY2dXFSe6ne8YMMHkYtAFgS2gjLu+Yc7wJqY8X/mnQf53TRBPiq05YJpUj7hZ/io
bJXbKV/61s2IEcFw1LYEoRD2F8rluqrmDK6ho4VLeMubDVkVPvf1/6nWoBfhyX3Q
LuFY8lpe+ZOVqLx9TWevdp9VgQpYZCft6Dw3xMWSJomVr/iyIQ82Ao6E3N0VyN+5
DB0Ph2GKHF78mP/3C9EaWNADSJOZjbHxKN0vjsh0hFJdoriiiRU0Io7utRsEqAkG
oT2lqu1/rY+6hEWrfooVklHWCSly6PGzR/ThxDd2DWPNKLFtqoSKRVyUcmdNmlDo
Fo57iuqIxYd0+3F7H3racDEzmVql3TFYLhuvkU4p+X46vUDH1knEGBwex0Y3vAJC
V1D+uLDn7InRF9Xb8gVLopDET3f+I0NfnSTK1VoH7VpTa+AUHg8TBfRJDXMC6CQX
aC/bxWDO64sR7PhZMfIqC6ZtYO2mzxxVNtDO1U1DtRjIG4dSJhK7tqNovqPPMunN
iNPC27aJ+48YARmm4c0hXgTtSaG7K5rKaNl1rCz2zDbjtRIavO/JcmBP1areyhro
0+E+rVvKsCGmm+S2PF+baChap+Viu+pWyh23LR5cH9BhilgKdaApIvzEqZ/UW41q
asKqm7Fv+wimm/WFZFan2eTHX4xqxLApGoljKN463yGG9qt2y9sBeQxohn25iPg8
HT2LUcjV23rmHYdThxRnLD07gYC8r3I2PG+J7E5JfND474H3NTuOT7Yu74uyk9lh
e3rgpn/dufEv0YwiYhSMEy4BwyGx+F4O5LKexqSqyCXBTqoY1KqyjviG1h9zgqPW
cfGKlpSuHAD7vQvR/6asK9ICMqvwiJyTxJWSGFfZpNN0u2IyO9xYReYVMUMiFE6z
y1uuaTaO7T6LdOgzoYfuCAHWYoQBhizX1RiWdrxA/3kIA4y05ElAp6Mwvrq0Q6jQ
9UhcWmOL/6w2ujvfD4N30pdAXer8/nyfN7LmQhi6BrSzIt4IxqWclXh25Lpy4oja
nkWCZeApe+5B0/4wJosmbJkcsRwMwtpUMC4OTcg5V4toR0zZyUuYnITfiK4FQ80/
s7bnkIEiP9yWnzjops9GK0r4YYQMb1Wh1cdJ4juw4xR++fcYA9JegZGCJfAbLxVB
NSJrk9z5g9Flo0/bLbZyWnRAkrQI7opMPh/YTmP8ijiPXNbtNxfLm1DhCDwYW06M
CrEa0w8+5ZtGu+Tn64RZbHxr1o+GMTQRO2F5hyiIc1vvoRFPnOju2KC2DsBR6ePk
GQq49FWGnShD/Zw/V83IJV2xE3Tv6htFrTgZ8lo+6gXFFntRE6jzfVQ/qPjbVwdh
65mlneklA56BKHIPcxXaK7P0ozAeBVZuBK85PDQ7vHCA4mOi3cEbSvgEB5SynGWL
vlMIBqdHI6D27hFR5AhCLVZJgKeUal4oBDFjgRwA7R2WRwLIxn76ZEWJ4F6V0wl6
l7SYVm0LvztY8fjrWOKTdnFwaKdZevjx53UPT6rRqM1guM3dTpOFgrpWbzy3UaBF
q86b/oCrO+OHcIIRnOuAV/3F8Dw56WlyfAPNfFTTg4dTSn/g5dOGEfTNYQx1fRNW
KHzIGQNZsKTJonCezh8MdVKE6uxWQKGfOd9FrPTr0UIwYpvuTWZhu/m7FNaxvD0t
nMxmWKQnLOPxD0zmShxS8bkzjFJOBPZuCpiPc0fWozTOzGE3xSsD2I9Qha3mBKau
CKnBSZaY/217eJwa+78xmwnIWN1bMTQyHl95cuXVUvckBY4eNmYl/3S/yxap5iOg
XfccIa/1V1e6xcoHNlhwfXxBEHEcUgKtcLhTOXB1KCiTEgDPruXQQkcf6dAN9knj
h2SaEzuxucvG2FTkjxgVOrHMSLp28MFRA3bGbxO0AEfK7KXYv3CscOHH/NEbYHYl
dYy6xSUjFvy6PUSQ1qHPgYJOuvhOC7ptpPaVUkT9Uy/JEfwln+ZAfgSZAIj+FyZ6
Wsi0JxGPbltYxFp4guTM35/VtDDXSaOU+sYAxtF7PwID14u+FjBqOpIbJrqj5OTs
Y/a31a4qdqCqCXKX4rAYUmaXwWCL+ef0ypc2ZdvTzMskJdAtNBy9CyXDVgh+G5Mg
WNosJeVPOJ+DvckcCQGURkt0055JsvjwsSKpmj2w4NyLBMPlC/KZet6025NYWK5t
nc5Kp8Xyur1QqeR1YpUdAMOXLOyXWhU3DywecYACiJyBwLPIfHoKDQeFcdFdafDO
kH21Ek+Hyvwvvo1oUkotzoXZmNHINtAYpykWgXutBpGgJO5BfUtXcLQ4y49pDfEY
warpOQATJLD7uvHkCsEuMXfyh2Njj/np88VwkyyaU1TJ3cmB1Vzj6EUND/uAxajw
kSQdBVFDTq36dW76nRMj89CNCUjGiPtlRJihfVBwpNIEmQD7JCh36B2XI+mmQSDW
9u/KmJBjGAjD2t19cRfaCuBo6gAl+1yRob1e+KqPjcIWUehUQ+jDSguuAKD5IHZJ
Er8rX8DPgLOu9sGo9vK+rS/pnqI0ciPtwOA5Ko5CKTZyDKB5U9VxhKXYYAWBFlJ+
ed/WcsxSR7skejsIyg8DlZ0mVScXexz00avqnO0CuqfTGz+XG+HgAXTql+OBHf9D
1hZO7tJ1qOuesEbeelBB9sMr3IFU5G8QDb2d9kiQGZgRWB6VSQadIvsomhhELCS0
c1Ai5GWhQ8NVVO4EGc6UNIZN11kaBxMva2VrVTMZBKrzGQJqMRnCeVsCe9901RX2
MqxNNkkUU8W4L+DrqOD62O3YmHXV4bjYvKeSGdA82aRgpjY7KfEvDmvUzpf8N48L
CiFfXchf9y07gZ5XucEcaki4wh6//3M8YxYbf+aWYhhLA84rsWy0PUCHuKXHy28s
aRB5dRouryOGI75+C4pEhSm+7p5rEB6fHghbYMCWW4k0Qpe4GjXcUi2kZ5SsyLUB
cXM3y6boNkPvEjxLCM3J7rN6FSb2JoCcIK3pGOFSUowgt5GQDm9UOiJkQnwGpQKw
y+mRgi1gqHDI27bqomXKfG2/fzvuK/e98n1KfBcaA/V/1+ZZ4rXH40qKfIySNLUM
iWZAU+uX88PClNwyTSFbgT1092IsUSY/n1mybRa54IDRC98BStxdh0QGzZkTYBAD
ICyqy5WWnlYQOUtK69TnHpzZljiogrAfU6NKDv088H7GH7dZanGB7kdEErlkg2ML
2RDjMckF4c3kh1uFD764EUTZHdmYUaigCH2l+tw5bV3VSmhkt03CZF+jvpJL/aw2
nApOOnsLB05mCv2ROpGFv+dvUpa8PHg8UAoGASf2GRh2w+7FrTqXUUHygSM45tfS
1lwRnoYW43iXbCy3QKtVj+LFBU7MC6aI69os+Mh2ROXSmLTlZp+Kw04+xI5WZc9S
7y6i4YPVi5yyqCzCYQ87CbUO4/Aqt6GJHmTn95pSrjPpnnhKvgvTvRPIG/0UHZK7
18xOMVpAwfaCaWTjK1ijMg9Cx4U2JUgPGi/mDors9MZhfHnnvZ9Iu0MuoP01e5Kj
Vw3GoOEXvNu9bvHfDiYUZ7cm+Uu0CwwkFEaRyYnXbkzgbFA8DPBw7XZQZLXfopQI
XsO29HcnmXuB7egCWl7ei8V664q4SZnvt4eYT+AzfojBTAIAy6Pj5voGBBYtt/eX
KHwc4yFVhlSTeN+dIRdrVpyN3hXm0nvjyH/km9ZSNHKq4bqsblZGrqNmTwgJswxz
BtG3GKDaN/u3TQzvb4xA7CMc7OeH80eA2V2TNwgf88ARkzHtDzdvlZFfPq5Q8Ucy
KzPMrAfI/Wu7ohQPZyCD2fq9l1niqudMfmRrPXuw61dW+8qZ2wRLx+ngVmnBpCH2
3IVaLodqcytQNEewvJs4Q28UjmCq+sPpORRnp/U2kFj5sV/4kmXbEDlcLjamXagz
1ddB7mJ2MKqVyNF4crJOHQBuwM/ILMW5PXxUxZH5t6NtR1FiGssS4i/xcpOyoYlb
5zhclgJ3pU5wAv4lrUe3f6gdlPEH6S4L6HDAzu1LZSIyF1H6viHoxFcauK9U04sm
rwEqPrqaH2L9EkJ23f1p8OAdBKwdr8e9muRJ1UrIw2eL9U8rrg8mrg5AP9LhkWX2
JkYtPjzpCHSp/CHfqBthr55nM40iuL9B59uugLJm75NLDLHLRqeik0jdwF67sGRz
TCc6KyvX1IQBldlJaWhQ/vwmBLAoc1dsnw0bx4aUJpWAl2jAYAhskiLZ2bL2AeMF
qpu7RffQawCsuH1CCQ+4BZWO3Dye4xa4SVb61vaXhteiWi7LK5CV7RbD1y7x4xJ7
4X5iOQ2w3iaTAO6aO+AEH57EsZfg2B9NXHSbVi7qt07Rf2tipYpoB7159E491Ty/
QHxLIEj/IpSYxJ6qo3WysXJEVv6f/UU+0kL6iASWSpyQetyqnnermA0wf/1Hvalq
Nn7WLHrtRnQ4tfV+KRWAUPio+Z3Dt8e8HjWA3Ggzjy+5fxyvYg/4jqBv9/w3YwYE
tfSLSpfDsL48j92FxaHbYiltQJvKS7veasQnPz0AKWGSf2CbQ46JMF73Hu7+bKzt
fpCe5G30CGY8LU58TuAEDFhACRgsfVUj5lRSGAMKOiShibyImJV4EL7rIq8GnU5p
JF1Mec6kDzIlf5cw5fjAq2VvgdFMOdJ/Vaq06V/DXGhF8UqtZHk4QtzAqwWejvbf
cG3kfh1t+sJ/N5Wd98i463Jqq61OSHcFgPh4Zyr5JKx3jBHF+tp4YA9IPWANM3SH
Bo7aEnBNTYthwGNq8nv6gXZ4ncKfOc9I7zEpdIr1POWSGY7lu6VtiF5ZEepTnXxk
bf4xCC/Ry2KcHVj2N4iZvEF8mVSm36GOSwCmApdlm2shHyfVcQv6xLDkjozCznuB
VlFmo0J5MmX+Nhdek5LhrMyVhwtysgWK+6tMZt/ceP/ZcPkqbMCbNu5EY6q0EKs9
A3c6P034x/ek3bgN52OdY1EnkY2SjwyQ8l4prJ4ycgvlg6UExQdShbnNpSicJLcm
dZ8UhtZD74Ti6Sp6GVOupEaKuTK7UX4aqr7rmS893mZfH5Lzx8DdkNv6Ibo9Ckqt
bNFa+AGkStAXe/SGwSgqioNlDUoOC5CzPWbpzOGYod0O86UUBf1eWdWjPITiagqE
eR+XivDuv0SIsNfglOQy0+j7B7hphBAtya+BgbZ15aVpmFwl7x5uEF7axV13YAqA
E6KUGJSlucJ+An7zPSoyowbixbG8HAvhYUnGLZUfs0x3cYMwynVGYS+hxMW2fPnq
YkrzD7MrLEJeq2hMhFmTaq72ZybTNs9gZzcYVcA3VOYlh8IY9WQwpzBG5VzVQZtN
Qx2n8Jz384VkRzcfEwo+6PiREajrgQQvHxcvZu/6ex1zM667dbVd2obO3F7hMs67
zWr3Bc3cVfnsEXIH4hGPynRLorbwOMFSFfFIdH6c9uKoGgtq1vnE4hrUPGx52cp4
EAdNhsUmfuZee3Fj1Nqkwq17eHvkeDknllPjcoVvLJ8nQPiy1alc1Q/WaWNCy6tW
qrHvsaSeqPQ5+KpDyz8EVKu8mEfTpW3pRNCHJJ7ENE8B1HBX/bqVo/i0THxVgG6/
O0+HpFrnal8y9Yg0GS806x8uZxay6uoiqz9Q7tmEDtv9OohlMa5qn0LJBc93vLLL
dgNMVqsl267arPIDr2aiIhXlTKkr59zJXvLqTX3D2kvgrwZlerAfB/A1NwE8H/AL
iDGprWlJRjFqnAQumf6sKfrj9dBKkgY8dTkn0x/HqWmQzFm6fdMER3BBAjLUYgOw
HIf3t7yYEQgKYD7dcXDFY/8kvkGTz105rDHdtkL0WROINZ8mYxN/QmutP8SmdyDm
HYjKIjO2SnrUQzImD5k1aTX16D5iY3sxNzP4GVE5gFH60ogTq3JLrdm5Qgjwsz+n
KaYoe4y0KbjigLFgQLpl/pbPflj9OoPAj9t2Cc58AnqplKZ7vW0xD8Ve54ok/W7D
uug49XB8vq6opgSlLaiKaNUFwkaQJWkWVRRrswBecSltb2+4BBSYVn3h/FXQdLz+
YDrSyUifkQa7eOFKTxnD+JkpnBzncPlrgvId8X7ALco+IHZVRQ9c5GTv6QCTANWQ
5IE6V7k7jgO0QTCj5mVAnySzv/zseKYTWs/WQmIbzcElSBUfgi721cdwCQBjcPOA
SKXZkFSXIRcGWTMfFkM0TBU+uw26IQKmX4Ax6KB9dzrp7GljcmwXH4DZLFzOeUIN
JoBtU01j5OuWSDWuXXaWchjmFEfVkME8UhkX55d+QTKEoM2Pv23mfn5BuizdhlxO
0chKxQiZa/LpQAltqwrJFkhzh8Nn4C9V1aZ9gvJ4i1Yf8Tc8wWsgJGH7NJfFPEZv
xL+ikgijHNTtKBrdA7nEihGY+bTQ3oLjKIxNGdmyXGEziP/ZzIXd0/IcMPhMvXvy
6oH4xPiASvp41m6kvNFfCiJ+oR+45EcnBmvQMRjp1n6XFA4d2uqDMm0RTRGty5Dx
EgYNLk2TNVkgp9kR+xmNEBJM0ZtOe/lGMn79GnsT+oeoQt7u0LkeMA8q0R7C5qBf
ALbWTrqLDOVVtOq2ssi7TYkJYEwthvcOoG4wGQx0PS9v+0qJ+6xTCg+8KDTnawQf
kfF3iEJAzmzRErol1rP8EPrnWYrpANxqXLg+F1gaRBM+ibYcn8BlR2rC9imwxS9t
LBrpne/Zxjdr3siHkLnLVyl1jwr9EaegxYNsbzg/VTWCaahXcqauS1Zp/LAauSsB
3PIJdAhKF+mjPECdyxmaFCKDsNRUK2NOuUHtilopSomm+DARQZtdeqHydEsnVJJY
Kks+Jw/deO55EmQ4HJQCO2jyJQpRAWZPIFhKeOdh31CwK7KJ11OhCNTpyYTjVVnl
VVim8fhPs+rk37jiUwsfB2Y4X1bjJj7g5+NMC2EUdQSw+S+P+c/lomjwWzhleAUu
TSYPWLExn22YFMqj+6AQINsxbEDCuG/oOpGYUxNsny01EowXEw+ZxMYrJHEpjPVy
stM4CAdpHdSXWAjbKY3QOrLkR+QgWS+gyVsc8a+bgUX+d3+0F7yTFOGN1sbUKETR
QXFIRc9Jl4TkIDt6dJ98jebys1m+9uXDKX1Ywb7tEUdPNXN26J9JPKTrJ1S4s8uA
SP8xVSmkOUO3EX9aM1I9Wm9wfsIP8qAPmdLSkIWb98xtvKwqSYw9wisxWefXgokK
HJWfjdVbKdLMoioj/TpIfVYv/q6++2hTLtyggABpvKlo1KIXDiD+D2Y1MnLDyHao
UOO8Ruk3XZwrFrXJL6DKLD8R9a3uvH7sY7drqihp78z/HDMcpW4C/dMIS8ehnJx+
Sc8B/Q+BnP2LiRkMt54tau+VA6ulkdLHkPGt+AGj/oGsC5YsgFoSXZXms/7XSKDy
OebtDjECLJX4n0ZxKO0kqrxtoL5W1eLfDjf3mKhRFeQ38rFawsYbEQ8+Y9I5Cbhz
UoB/OIVa3aY/bL+5EijDs263s2F0O98PdDGdAtx0TAAHtt+tGZjC6JvO1xSsKjaj
mGgBgFP8zLqskGFi0h/zd6drbGqQrHoD7M7QRbxAQFnCUyU2f2yhkaCgiTUg8W//
qht+nreI5pI3bPrV82UNZxwUnTlYHcRlQNV7fM7onOgg+geyzSb7Xb8ABYO+kQnU
/zaJ5/nemXBZOYDDZqc7tT1JNno4hDLaNxW4zwCFAFGB3t+vLhVZ1hwHAGk8QM4R
d/YJ9mCq0FCNG2ICNPi/wBor8EVT3noKlNmmVqGOOs7Z5CHBzVm7O9p5/fFFSIpf
ciw8pBown0cBGEGsanA7K/ex48yrSHRtkpt9E9nPsJqt7lSB+Fh8HX2wogPx1WPm
+ZoMax1CFyaQzoPtbZuUbXqpWnQUV4RUMjYzNPXP++cAxo90ARRz73UJTlCcX/7H
8FanLej5GuLipBX/3HYv67Q4RUmTuSryZ23e5GdtPRe5LkJ6kQFOhRM5TiXXLML+
Fbcg93sKTP8pX9TJoxSn8dbEREPO/5GIUSIPf8vHQxNjIezVu+mpLi4W8fY8Jnok
lyEj4gHiw6zFFEd1WPVKLrJQRQjz4OnzIyWe4vSdKoeP3WHmd3sHP6b/iRBFZm9O
QjgWodyCWqgxxuklGP8ybHonLZiAGYtmQtxez3G9xSk4GOcojhUJCFjMJNcpKMAu
G/7Tn9r85VFU+BKQJ7LPKJ65BiTuTMXTsjycRaxZ7s5vfqJFDViWdNPy2fXJFpaP
GZAwYXQGRKtSwDONVdj7JayiHqhXpYSjI5tKfp/RoVaKIxGa8udJm6EuL1m0ji3H
klOQcrkFgCVJGuHdf1lU8ggpWf+PNLisiyxhbcLzNTj2fzvhIhKVOCh0FULqNt9P
WZi4A0xDCX3fp4SIcqA/NAPP/U+Y3sz1avUh3oYStelj3h7saWb2HbAWItOTP6Va
VFIdoLm+yrKSPtoq0hfPPp5duTwow+R3Q70gM3hiT8QdgX5D91qjW1QbBAqM6a3r
Yok4R3L32gFBbN6nAjhxQnvZeVY9lMjGDZ2v2vwI4+DWocyxEaRYoAvoo5Z/Y8RA
FjDpx3vyEoYJW8QWPt9FDq7Z30ybFsdR0Vq2ZG49sGapuePwYpmHjBwvG/fYHIzW
/pGwVUQKArYluJDb8xbe0P7ZxErbkuuV8O/tpKresCBzRd/wOTTZWMK1IYP1w7zY
296X7TNMasmxJHnMA+O/SCjNWm1XucxqA1swb0VDgSgIraXzyYqPLkF8WGm6TwN2
hdILX3r55t5H0fPnNJekUgO+B7scAKLO+iBUrr4FCl9gimKwfu9lALOs3hVUmCZv
u0O5zNDS1AE4iZvP9gwhCHV33CBJyilc6UP2vjsQuxpbBCW1GRr6L+HXa3a/wMro
m/mPmY220Qxr8A/xqZMDUoLNAe9LKCJLG37b3kIUIH5ilECAGwTh/YdWABSquerW
C3QuPYuTarE0FoZFUTpI9VMHa+d06kUtR0uajBvVt1lTsDEQpFSxeJZzrOOkV7l5
NDXsq31QVq4axJ210+9O21PjFPa6NnoTzXBQO0wuMJ6M4hDBv9VyQ0OnE850vmUB
aIZOBkM3aIWc04mWwATS/qRFmtTsOHRH04h9aR/mx85qgOh6njLJqsoiOKxpc/v1
pB692lXBEVhMMfhWyZ09hquzXChElH8PVaB4zv2pmH3haI8LNvvZP9yr47Yx5rCD
9MV0/yP4OWpT3UyTCVujeoOQ5ThkFqlym8p8Voo//23bBL6ABrMe9gjlC7Ht+VSf
fZm5cTL793gtdXg4Ku6Lq51z1AsolnuJSqDWUIF41pllLjYQbjvyRCoOqkufbEf9
/XYP1kbdSTumSZLlqTKrtXJhYa+EyUBC3tnF7/BuSixaQe/xNjMVsULTCcyBmU1r
OGK6RcLcjFwR0Ys3kREWw9BDKlyJqZhu/05RDrWEyMBzsiFdTN6yPgaEzo7AgtcU
1Y/NgjNZYI9R9D2TPv04vsIOIeAdi+2REkBgfPSiwVB1hJR0cMbKojCFKqCOtGtY
yj/sdEsSNT/r00mjDdqp5Qf8BZzg4cvYkhtLFYkSAnr4Z1ehzRNrWtrPXyyvKPe4
x/Pt3rrpauqerZWvLUMbynqYTJw4JRnVcqR7pNoK2ueegu3kW5ye7n3VNg/0ShaD
NT3YtFbiCk+WNdWseZMUBO/SuGkyRACLRrW3ncNxZqLC+joXRho7CKjcINuoCfAN
7LaTS+IBBjkufCgo7wCJQRIbzFsHpC+Q7S46FBXS3NFds3WuJcMl7ZfR/nMbj4HJ
PyX6S3RdSGXgueYgDxQrkGt1+1+2FBCzsyqiOLS5lAOK86Pd5MLn8EwdyJW6ueYe
RkDDuKdRbvHVMyroiENkJpO6c6VJpbCS+FuCxfyAlSr/XYXfhIhpnTg5jdIiSLHW
jkGbvZNjtqjBX2lfg3RmkyombwidvbQKt7DohVfwsFrjd/tr/7jWOMW/uHq+Tm6Z
QjwaZU57JsqiztwIQcm9Nji4/RTI1e79Rr84rQY3hWX69b94aveVCWAo0CGZ/DUY
NNBmrdx+TW7H7OuDXbAyQeMHyvZWd0foxwO4lzhWCthk+SKp1IGMK45xaF593Isr
NZkcT4u/fsZmhT3tYApBaoAJl3/cw+J7A1Q+hl4b+p3JgTXz6xy1kxnEFo8mUu3Q
ot6xeWKUg/hdHG0bjYWzd63afn5kk9a3T45HJHA+J1d8qidFsG9wo+JjMJTOCTSQ
QAoAaQY27tU1Ki/Kevb4DLihn5ziDFH0N6CSiHb+VJ8j7frFORAQA0l13lOUvTn0
6a8Z/dkRr5Fo8a8usBVEkceOZlYIUV35JK1VzPF4RNrSQq4c7HtMy4lffS0Z5QPI
l9lRUGwjMAo9NlaHpf3tdYr4lm9QWs30bkwr1CoPKHS7VDMydgEl42u6oGq6BQdX
s2s0sB20FRowJdUhXUuY/WEjUQB43c97PoKR9gUGOa0vbGWAiyn8BpPEOjpchc8g
2H8eSQ6dBPuBWcUkbwYbrVdxDAWOBm9iCcPmzKzbHsmkW+pF02nmSNqyTFnEBHrl
k8d1qEZfnGtkXXrIR3yBPVXxasaDZLBQ1KWrZ3xxfELTvfHaOAnXLQfcVXDJEf+s
w/RGww+E27roHZM5O/wrtOe61liY33Ywjxbsfi5laEchDEc8T6eFGImisTCwpy4I
I8pRyQ9PFqk2JyTw8Fvehvv+lXTzA6N8fCVswgQ2d9jcaFkWgU0EEfdLxzNJQTMi
KLkNRnDH2tWxW5sCIlAP7dOb6fN9TiN/TKIo+fooI8ctVA14X6jhP1F3zKwS9Uov
b8RhuhN4eWMftN4UHkpZ2/OjPQ5ufKB9yFmE+9astPWMR3YPKWPDx+xD2BypwrK/
16ECBhy0VevVSB8ctFkMxL9/Tncx2NONih9qfXEo/0R7MvaMR7LeWFViQ1nhencH
o4VzWHkq9u+/jxvc03nsIyNa16U6O+2rJWYiRMbhBxx+hq2ZMLnHbvBMmSEIYR4U
QGpjlq39zmMY8vlvgRdTdoU5PbadUfSH4i46Ir67MQNSx97NN4LS3+36OxoC/SIu
bDdZh5PByK9pPPKxIEQwTwuWmD4AWrLM8zYTn3dtuuTpuC5UV/i9csgx8UGWwmSA
Gx/8pGDj1edmDowJt/RSWI9fUu/SLV7k0SHnL+7pUoUAG4tDXgyi1WHDdwgN8PjK
NJUcJi8aCzTDd3C2eqbJGt0+RVtE9Jbfl8W55oYkGRKh50ABvTjr4FRHpfrjNEUM
/16KJEWS+Z6qFEb1yuqfInFUmo6zeyeRh3IMp3CLaT8A8cyV/8voANIfz9bhO3i9
VAhz6USqynQmbUSK7CFFvnt4YzR3GfHQFJO4TvyVlxhodiqJetMx2AsdkMeBYq2X
VZ68jblfHNPYSo9vdz6K9V88eV89MsC9o3NUTKDCfGAithKEB3W+Wtmch4DGUGnD
8FcCz3zMX10WwF0a1HXhynQvTA/Y+CclORPIpEYqjoJ/RcO+RQZszqEVULK0MnMZ
EeNCHWDp1eXRXDK4I8+19A7BuX9ihQpR974KEGfUQF1zBncnkji35Rn7pknRrec1
wNrDdYBHthBujuZWRLN/Bs+G2eKOBVt/gHmH7Z/qKz3gF01w4vBHQBR2TF9UCMUg
1NqxNxbxIYLpoLXvlKvo0/PBWu+Dlrs4ew/HZC3pDazkvGYF3OOdwF5zNoJLMI3H
WELgjj2FPlYnJJwEoWX4Nwln0UagXKvvfJ6zMYlhvd9Rq1gMg4cZrcuX4p1BE7Oy
3HuSQiXc6izcvBVUWB63pHw6RWXfogy4/quzdiMqBqstLJrANJfmi6VXxdtm12vS
cIsycp1EUyRE6BJznvDo71dYnNUezVI7VoZOxYpb2xK863+P9vqH/PuWeGHS+1fp
eLYgAPDH/7WO2orBn3DcfRiNGGBCEqufDPYkOCD3o0LMvnWkyLOPkwid+m0G0dv/
PlqewvNbssHK+zoLaRLG7lDchMtbrhM9CidiNUfSjFH9JXXn0ZuQswVgdq7NKgLV
BeTDy13gu03ZDLC/KBssj8mPmYdPARNghu4Zd+m7wzvbj1lEOxGX+nrMngol08sP
0UgrdibGDrapwspplSgkDHlznanJ0Xz4AnG0x1IFJBaKTMnqgoMOpOsiA79ptwt6
V2LB6qxpoZ6FqCEbzC+h43NDd4ZqgHZZdWLlFfX0x6reAuAyx0BEhLkLMFkLIpny
+cCl3xt09HSd1rWY3x+Gubh0hfUFKoP/4dRTKf+A72OTvrJJagEHJdno5R2YWJ1w
3Zvq/Kwe4tPBTuCk/wp86jiQZ5v8gV19NEzMZYd7xVC1u5cVJtBzyvbkzq8+yq2U
Sqo4mfvoPyqlW+T2IxSu9JOoieFKxzsKH47K9XrE931d6AcgKNX+HexDdU5ngRFO
nsJz6x+vTgBsX5SKmy1QsaYqXwUl3GrjPyMl09uRcVH0WO2ivWCwO5m2gsL6Rt+I
nJo5FgDkh3ZkPwgC8TXkty6y14EmBKJc6YJ+QDL1/aUkf9U4y7xj6bC/e0kZ+QHR
JrGuOHmnuceEsRPtsWA6L1wNSY/tuvA2uxTTHzAqQcQf562A2FDwfmJlMAUn3Rd8
/9iyj29kDdbzIVsdfwRCFeyC5fqYrA96bFu///GDXyKGEk40tIamjwMN5K4u5urh
hft6BlH/9b2exHv91Yyvuh7G3YmDr4gb5rRXoVchZKJjQ+w7haBW+FKUx4AM6yfE
v7Kl+4kYKWbdQzt2YhCeWlr6rlAtSDmRBY5RSsuPalSYvYlr1d45rSGyDOeUckDw
QecTyf7mn7yYGXwoCGrSXieWo3KgmpVPigayb3epO8oaOMWfrT+tDqAHpKt+LpOS
bCfBo7zQJh27U8a0oVPPmi+oZ9Sg09hj9QOziIKc8i+HH5P9PCpECYxSs2KABBxH
elUOH+o+r3L2zbN2jLENBzigjAskT14oco25GPKUunP+jCyGNMtWXUvLxSbAHYQW
LGV427IVCPy5oVKfyO7MxFh/0YjEgJK7BlLUBGcL/naDw8c9Kp7UizJBC+1lrCJ/
VCkT9gjG8AG587oK+bPC0aNgyy2q9oBi1XBwyhcXz9jZdolJFI2ByW122HpBz5Rc
aZVS4id76vAKrYIgMJwx5Q8jos+5nvczoJ2jMoRvTqufSVE4yp+glzVhyCHiMH9u
cBtysCI2JTmd0X1xtzpa43wmp3SoRsORpbAoPxaSigN6mRQqRr3TZVEex2oQK8cU
mS9vxpWeVjZ5eETjOd/kbo9F379cpGLrsmNrxLE6v8u5BN1UcttC7+k9pVjEKT2e
lRbocMMbuMmMk/j3rF1tpdoGc19lmWC72U3yLGVscApLaQjQhcvMeOdBAa6GiXKb
Ngj4Ino53C75Fsj31B7VnBhO9fdidqaSzKgyfl9/7jMrC8EmoVgkJJl//ZmpvXG2
hGtgkgW60G1aQLFfigv4vaqMyF75zybQX3PCjW3UAOwFfhGEAZVMz2fggsEauBzJ
LKr98+n/kJdVwC19e2ERQeEhM6elt8sqcwrB2ksVCburQ6NPa2qvJe02o0tqBr0Z
IL9fAa2KaLkzW4i+R2cL+m/Y21IkujeLzMt1psBSCuMB8+xWw5ZhgHhlArX0O1Iu
D2wDY9Gs6YpWHnXju4jGChNuGbYKUnRI0Q22BYRFOxbiveG4yFzaWYkgMy6QIO5L
Sjanxq5QOYyBZ8SzdnOl5F0PeKPuG7jSEbS9Mh57fGkuxoue183k62QY0IrmRZDy
8Fn2Hhm0uFD2EDic9kIfOTNhGzxJyBFenTOQy8KULTDv6VNRK4YMMnPC7PcgTQwA
KNUkSLHXURXTIqY1MDu5Ho0j3KcoYx/6oENYpcp/uoIxxgnlkCsvnKRlwKtMewIg
sPZuwnhvkmsd6s+e+vOYnX6Lu3V90J6/yWTE0g08clqrTTq6sS5SxStwadrPPwb1
hR/6Qc5zDe/mabtit4eeOXQr3MW86sKlf+UVunIoARNaTqNSyiqXAkAQFovcayuy
oZzy3ZlPADKOb5zWwlxx9r3BDRlWciUA6Sl4/LcA1VbPeo73iEa0s6ZVYfronfrT
gpTrPkrnx10JHpX73Od85ysBwHDR2ELDkDN8CPDKKwAoMd3/YFBQsqItZxFyzH+I
TQdP5lI+Llf81BnEmJshZy4bTeNKDQY3OI7O1XhDGZAyDC+hcnqGYC2Tw3/Kqimv
BSG0YxcWCYnz1P1o1B1HJqao0vmg9w72HAg0lJDPOrIEmZ2OUfc+7v7HphdzYYqv
Fhr8HLonqh1AxTznMNZ9gTTSpZAfyjVA8yeIEgpNfbHG0k6x4oP6T15EZyoHroz6
rh5Q50Pfq75MKpjEsHytVJqIDv5f+BPIyH/YimqWXXpMKIjAAQlLSpsONJTQaA6H
pwvcbuEQSOEPUHsZC46Dp4dzrzpq1dlu0MQJsrT5c3NgNrG8ca+MmQpJzKVfLSzB
MZEz+wiY+Hk5v6yw7uqHLE+LSMe4hZnmDPhgVMPltkz7oLg+GSsmx0EppPGW8jp1
SGFNM+fzYk7MCQhgqnyk1zMC2fDJ3rocWxiFWetNWF83BLaYqBgFMgeymHBE6Qvo
rLbdG+VU/BbkiD80JtxE/hELn4VEVW/800B9iYauAzspcw14z3pVw4bHrsJTZsP+
s+ZjzKApFrjkE+F2hqwyrg==
`protect END_PROTECTED
