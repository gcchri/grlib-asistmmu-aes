`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZnPg0TNCsA9haXC7OjO4PtPiq0VHX93UfHmCmYcyCRCIePhqmPNzB+wWHtIhnR1E
yxeBdr+vXWyyZF4ynBXVKSdE/Dp+ZS55pTdmS9jHJ0WWMe9sUoI7RujatOXrxYUp
9R0c3NMVq0XxzkJkFkNtvaIlSh1CQNbYUVMNGtFP6YGud/ERecyyzrtTjEAAmxC3
0pmKu4MoK8Zojs63QX72tfglJXZnpZemEeqcros6tuPycDq6neZ7wFJKvhKkb0sV
m+VvfDRGtxKTEl7P5SYrmIyityd53M8SwqLE49sBr61yA41X4phic61cV4tZPoiX
X6S2kcBAOtlZxkkrpPHCSA==
`protect END_PROTECTED
