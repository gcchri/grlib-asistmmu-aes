`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q3PStch2GmngxUh3YU8rINr8iL3y4wqxc6h/j+xvMdAaGpL/RRL4sFS81oTBB5/S
+Owp1NAW4n8bj7dZdYRAFfXIfTiZ5nl8g/3CvBjxQmBOOC4Ol5PslH7yKAMso7+w
1D9J+89dKk2tgZfczXpfoeBdSq43EJX+qCMDr3tlP4cpJMQMXjQlprTjO1G40J9f
y0V+/fxk5o5hZQmRF4jPol+uBtWGS+pOMynt7WNcro1V5e3Lvy54/hCmzfAUVnsI
cz0h4BLzu12EgNq3eM1le4m+woIPJHWdm2dIoPp5oB2T4yxEz1H1mD4rsmLn0z76
CGLc5kUejiv2kT+BJbeEthZpXSUftCnOu0O0bBWYuvHCS8gp92ac2tR2cvkTOVLM
pq+ygueJcUUNu9mE33AQrtuze1D6oD0WCdpjRj8uua8emJFCwXMaevoybPDZm1BH
`protect END_PROTECTED
