`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
StS0QSNKQlEeGWZ4vx2+kDHrYpKqM/PyXiV4qVP34Vqxxs7HDa+ibktN034ALzMM
JiMdAjxAfo1Fm/jsIZkZvXyzMiar1pD7f2Oit+6lS9MN0lua4HUyNYw8E3xoGu/W
Ekfi2ojVWtR07i7zc7rIfg0UjqPIG6M5wqtubQQn0RxGG3VbMsB+qFBi1LU3nDap
+JGbCxzVdgIxy7ZpvjTua3Doej8dlmlUNXcI5nWn8JYKyLCdyKhXcOrQIDLGNsO5
7My+ZSI5rh9yRd8A1herWN7PEr0KUb2ZZGgHkCKCVHlQgz4RYKfeowtL4atsnax2
Lbgumc8C/kdRIIpyCO2aDr3dUwcdsJ/1UOgafqJ9J26P4sRt8ysGg4jhnjsSr2Dn
T6QvcOco6Fv1sogMgLmQfZgtZGUKCv5w0jjMh3+hlEmPd3oY8fFTbiOPrn+IPDZt
9+cmFp9oP2B7+IMv26yXzHgS/3MrsXrUEAo+Rvv45RQUNA/tAAFLfjWkLXZcS4jr
GkZJGrR+0/Y1bsU0gAhfuUKo5B/WDeQDOLHqpFOp0A8tGS4WcaL+MFMIQvBtlls3
QVx+Vh0NByMxW9nLwPqTSoLR+Mqg9yLK22Khg5sLlwI=
`protect END_PROTECTED
