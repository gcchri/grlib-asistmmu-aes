`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
35f5QFM9LYefaMSfLxZGXs4o1bQBtk6GWAfDeniuY7d4lv+NPPzep09F1ePFuxSN
zCnaspgtkQDAlWsFC5Ow8vbF1fR2BabjVvVWSkiHFm3T6aHEwJexJDzWmgHXxXlO
1QUYV8uZfQ0VO2MtVAgbnNJsMakdR/JvsekxDgiXcGGg6VqAn2VW/MTq9Ilf44Uk
2BZ4iXaKHa7KS3hj5WcOPB2HmOIef2JjDJNfsnAmii/TpDsKJBGpS9EGmHTpSGbd
T7ZFRVWqqV0GjoUzTqmqofqXgoRjqpVUfdXFYd6WEdhRgedkEAmGafu1872n0kBE
jKCO/NVAq9n6zujbon+HNg==
`protect END_PROTECTED
