`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NC7f66IbKKxGORxvah1G7SAR0hu33XZ5ljXYnJZs300yWSLM0w3PhgO1f1FYIyuQ
5DdxGMMwCUXTMb1hvDeN5f+Cx38J1qOmeCL6AcsSmhUz4m6NQrz0oEzXGyRSJ6wZ
54ca+Q8JlXYz/lrw84vlrPmtv89LhuMEZsZ1KAT68JkJ6XIIktW5HPd8BqXkCcEk
YZseIsm5f8/EGkKcZ8jmBZfXW7B8c2OOAokShfVvtLa6nDLIIgTsM/W7BFZPBtvv
nDQmSzPpJXpTBERXz0fDhBrVePNukObM3drERxuRfzHkZVrBvac6z/+57zKR3JI6
VSMNRyzbyUCaRk3i+eqiPnGK3QMzd6EW+c72QNFVzy7y7hlPMSn92fTY1BFqEa1K
CuJmfBuaXslPQEpy5MqhiplFP7vTgEbes07FISIAoeDQPwWLdzYLa6Wa5sMxZD+k
2TsOEn1i/rdoRkeX2RW1ndOJvpSLgvqtaf5eBufCkWvpIbmHbSzZh4GQETiBwTX9
22pNBI5wlt3nr7zcvVdkxbPAGVgxxaLAU4U5hlspVedg91Q8qUnWCaCoZm7jyMLj
ESn8cYsMlp9ATs1rBEbMaTHo8scEvWgHOo+AoN8XTjXVC+r/7iSNvmDCjuz9hnmy
O7kpoCMliywkCjefED790nOsnvoqGusNHS7xaz3jeGs7mZ+qfhAHoqpEGi5Td/pZ
rlfSXwGFWGXTqwrID2wjfS79wjUnQ2bD77BAI7yltldpMqiuisGUy3Nvcp00A6E1
yabZityKx8rAVkBY740iltwnDK92o/tYs/6mT9RutYKH2t9LBaq5xmOzJWxZyDsJ
tSIkRPuLufcoPyAdFV0fCjCBZOnochdSBj+dPyPJX683jIw7PWWzrqQPU7d2ztcS
oU55IDRmHi6o9a2XFFM4kBEEWHdtUZVFT5m5nZSJmG3qKItEeYao9hpkr5NZmlPL
B5WsKReSTTKaHLajOwmhIGsUW6YDxAlyyyvHR8ndoS8ua3do7RvuyG/y6+AY3lUN
qROcxx6ROYldmx4TvJM5rDLxPDjGiAP3cQCLn34A2jolcOKIDErtCLJRT01CMNaF
5+1Yx0SXuQ5Q6MMoxs4IUFBiKz+sS9IYPntUnm0bqVthVSR/xfaURB1/wlwAwcNG
yQcKwgIZsHDjT5m6Ah6IUXoc7Lq6qBn2Dbbz4pJVycoL8lEJFF8a44epQ2GjwfYi
SVF7Jh64VM3FWYbx78uJ/3tbp4q2G+POajRYdq3C+P4GYTBwHufN3ofJJLiZAIHA
fa/PA0rviTkN+1IWs6zL2rbK7KNIQPnCCsWGwfeu45vc9ojhQNBNmq0kpWOp0E2L
c78FFH2tGRJhfy7Z43d++ewbcznWfqqZh8kF9yq+N5MIIrDVx6dr4o3xblk8mQqt
`protect END_PROTECTED
