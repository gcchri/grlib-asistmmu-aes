`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEOY8dqm8fQA+E8mgxtzt7FprNJz/icl47VoFg+heA9yqTYv3kvavGbhUt4JmkcO
y3LetIfVsa16tB1N8z9Z5Z2SVnwbXHLXs9kiYnTMWAU8Bbbg2gxHDcs+wMBa5C/h
mXu4alohIhUFb0yOirCNhNtR+E6GSlpH1k/2Xly3IrmdFrx/vdwTObKPCKvZ4sTy
zfDou4irjCBDklMZzaKfJF2WGoRrQVn+3BiY/wDSnBryP+oab519dyzLKR3W37S0
nvGwphpGdlWTlbmNNKCrHHW/UOeB8rNWmVIRkYrqruarWSUNgaFRienkA9IsH2T/
wbmehscCjBZL90PkpYOlZ6/i39X3upB4xDpU8Np1WcPw27Zdoh4kzQ8LGBlLl8yN
ErVWmnMf3tD9j2tW7TUd4KHrJwN/LLDZCV85xICaRatjTTD6bLGGhpD0T+q03z6P
TCIcJAKYmytfh6Zxg2B59KcD0ip8gGxcG7jbgxNEMj/0g/eGkSX1kjz2haNPXngF
ly3xaYQ3F03A/GjHz6Ir3vP6ZTSoGplgxnOxaNWYOI+ZjA/1g35akaKi1l9d0xsa
Y6WurSWoZBxxT5flacN0Uw==
`protect END_PROTECTED
