`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HAM34+sBleYCOyimHRfTGpErT/KxISfX+h4TZWwTSkNuJAAT936cNbLtF7csW+rJ
HQeHipmgmPHl5nDNRMBGQGy0snljahnYJZOscP7EG3xtFEx/0BakNqgV+9Fd8xOG
bIfFIaUfZ6nv3McYinfSheZMm6bWzyTJEfC+WpBQFlAvJAlyPBvoDFIV6lMviwwE
Z/BTfMPDi2WtemXUKvYw1OhSjvxcJvOCoQ4IGwGMicBxZeH4qiSXhMkPwf2C+fvX
d3zyqxgcDFtf9q1jIctxlDQeMgbAuOvHyKe08sOISfrKE6iRDZTKod661u/FR4vD
wKLRpyoHx6xNIfIyWQlamVkARnd1n+GTdaCyhns+yE7/HYuGSFx25W+EXmyZaHZV
cClLpMJOyOU2rd0W939lbpEzjFL3w6g7pR7ItQyWp1qhiKsuVWTo3KrY2htR+Z8o
IqETYIwjrUkGubFxpvzSUOt4RmwtzeP0w0f/GzbGO4zbZ7OctWnABPafbcJcOmU6
UtcrVK5ighZCnoQc4esG2qClIss38JlSdSR9WphDlrCNaV4omAEJk+R8HeemxZSI
gYdmIM8uWtXBbsLbqjfvNfjrov7jFPBSrf+EX2quJK7qtg9xrOZbvBXqNe09T+uc
Nt5vfrqG4fc9oPsFjKjhqZ1MBfxOsTAMeZGrpIcl6IuGRruSLU/ATXbbPV52GfOh
TqUz/iYi0W5GInXLwOsJtqWumdnRFSOWBpmDtdvRJBIul6AbsxXunJ5TXmhAbcPm
4JCqo6mN2KHoXE+pokzgBSyuJq/iepLzRcSdGx4SZTrAhrpdUBKzkvz72myo4hkK
OJ/XXAjJ1cYUJpFQkPawHkLnZil/oJlu4qNDkxojH10=
`protect END_PROTECTED
