`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T6/6f6UgFT1SglA3zaHFIA1dJTb9uZlAq0vgJ9A061N3RxVSQQUwrBuHLdGu8g02
sNI+wNWNt6DESx9gMPROJ1gMEDLEFroUIRAia2XloTqKaGENP1aV8KIn76IKMpUH
CFHCclZ6KYVmVb5Bub3ySHhrxhWX3DUXO9PvMwNenJ3MtWh5+NpPcS/IF0dWbxQA
m5xxdt/I3+7ZyMCoR2PD0LM9h2xPIQqhP/nx2uq7EJlVzJDt+WlJ+bW3r+rFys2B
Lb/9+/5LYViXe1F78smrB/yIN2hVpzt91L9VnMR3tl/bsXa43pME84tPXGpjw3Na
fmNifNLxOaXIU7QMx9HDtSvzbpt39TmGjfQTPwyGsRzrTrmqDXdSe2S/GqcMX6DA
myWjzg/rWkPvLxDdykDQ9p5Q5yWJLx/FnXE2HFqJH2xNIbTrjCOSGyEVlQTOrOfX
tl6Ip7qqPFW8Uqk/dGggeb8oQjJMytzkwD3JZV9vmjcVFIoQp+w9OMnxzEf+02D1
`protect END_PROTECTED
