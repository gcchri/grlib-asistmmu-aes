`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eayk2LtaM8gDXIMKW/UWsuvFlz203JcIAdVLiaVuxkTgdClaqtL68d4Xu8AL8npa
sey3m+pchIi/QAtlaA4HP+AH3A5IJWcwY7dUcs/UanJbzl+jpT2H4QOaktCMR+Av
NzKQKofjXtNNuDDiv3LpekDuzc8ngMfdK5vs6X5M7DcANoU4fl4s3GwHySg1OHhC
9rXEYt/iFfPJucdUN0yi6BCmxmQ+QTGd/asQYDfDyxiTngQGQIdDuW2R57toc2Qv
EtkYmrLZTLWNvzUUwElDKA==
`protect END_PROTECTED
