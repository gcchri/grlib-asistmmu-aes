`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FOrx3ls+AWRuuQ8dpdlMkjeXOC9Pc44cH+C2Od9NXPMJKi82PGAK6BcVrr+UCgkp
PP+YjXJu87ElgmiLlxm8a2ElsH5n4IQgwMDWO4PJF+voLZIa/qZCPlCjY1DqvU9L
Kg4qdA3XYy7DNonheHNs4bbXRW/M0o8u9fbN8GIwLwixcCmR+p8ibIC3I4KXqU4a
B2H+NGnY/3BXOtNB7XKhKhDTzMtX0RvY9n1407WtXFNB+7CMu0ys+8gR+yCpjV+f
AFLFnZMixuWAkDv0ExAp2+Etr9tuD56feQ1vRkUry0ly/eR/clOzNLE+msP37A9w
7ED6f8mQ8Wf7CTAmneZ0XYQ0DqntzR05iCCqi5n/eCDzMddZrJsOasbOMFW/KvcY
omIv+Jv+CaLqiiX5c9X+YcpGbhIzRr++NIbfybOM9n8cy/gqE90/XwTBZksCq/tc
NoYbEhA5QFggemA9fAvvOirgj1eMjeMYovwS4Uuaqa2C3UY+rbq8g6tmiZRAJVsM
i102FxQA3gC0XKRtrjvYLRNAAw6mbCaC5ifjN25TUl/NosSYodrTmaYZFoCQqmcL
qH3cXWWUylBfTAwQwYPBfuE8JisR9IwlpJvPqCW+jzAjTm9Q5Km9b/gBAT54Nbx2
u42WPpyqzWoXw91EkvEtVivxI3Sg1w4LqmfV2wpxI36YWZsxYsaekA4zWwGbkioW
8+S0Wp5qbap+pyoG0t0LNw==
`protect END_PROTECTED
