`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NoeBBL71tgcy5AFST94A08FR3vPbtm3W+wJ4D9XTxfgREyuvfw6WWjuyPDChFu4Z
pBupitlWJqvRyBAIUf2QHDnrdjh1ZusEXo6E/z0t6XXzZc0jnjskIrrZnVnyoPM7
h9hxj84LbB8Jwy33u5/Szy6ZfYwHA3muqDuJwlV+9Il0UBylNayKTSRvMevmRgpx
iHOmXSTHbg56Zo/V6F7Ikgr48RQBPd4mO8ARhA06X4TXN5dSbtkEs+iFEftwLAVx
IHfIP9E+K2VFJCamg8g/3n/Sb5csfob4vFR2B1hL0ReiZgosAKasfSr0elxnOov1
OIFVSFqFhS2QqK4pRyN0Z7BGYJBbEnCxD6HR4kR4MOdyvKh5FWZup5OdEnanDbuG
0lm6K4Fp0bmeN0i+4mYljOyC/v/xBe6dx8xsEc5DNDe0+QeeVZJXxm2e28iV+/oF
fRXfhD/8sgIo4AckEUMiIBxkS6YQJmfEGlNCXlhRKMSl+H9l2sj/9EEOGfhMl0ro
wb8qBVG4hhZJoSMhxf6b8T0m1maHG7Hnm8Tn2gkUmXyNrATClMEjsJOO8dWGdiwo
T6YqDaaAffCZhwjnDUNtjPpM3Uo4QWjTKVSOVkQ7X1CVjF8d5UF6LiWHF2upEa0A
tYe8tzcDX3Kf61K/0qBg38u/RCaxyHzVLqs+VqKO+bygbjzlpJpcaIYDwU9h0Ta1
gLQlltqNU5KIAd3QZU8OatpRQYyvU2vCbcktGcOmSVC7V+DuY6HyWCqPXnR9YehB
gSkW/SqMdj0lmiE5eQnUK8Z5I1YMftcP5vTyTpjpyx/DgJhfFp6QncOIziw3RVGP
QRhNeQUXmePRjawLcgEJJWDxQPVnQ0hcg4GF9Huj2Hg=
`protect END_PROTECTED
