`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iTE+poHpBQZaOexus9X4CPiBlaC+lEnzA0KDk0Kq62n8xqmwqyYFqAvruZHnAG6a
gMm4EwI2uNMXr9crRcFojdawnrvD49lhdu92zUZtrJ+S7BDthNuFGKX9p6bAtxrt
w3YncTJ4Rz5IG03WjYBhWxJ1Rrxtr0/wNfnhEb1wrOj2T9Y6copTcF6vuDz6AbTC
VYWt0eXsnlVTLrzpHez8EzF9xf6xhQ6G3W/kPEyFJkgw1hv2d4mUvk0w2Z3XeDm9
omOfPTCqjSDAO4ZbQaEO3srXE7MOlHCUPrRVOjWsXcvwzhvUJuiZQAjZwGXfm9DN
WXdsstB9EwVNlQOldrZ3GJoseh2PNvHQ5VJspQsJ9AQZ59zO40gEKzWETagUpU3P
xtXY5PEpB/AJXjgrRETdCn4vgGFr3M/vYx0K8qtfrPcQ2PHz3qprwqofdmqgvK2V
aNnR1o8KOimXlVxq3ozySPAfjO5KegmpBcRGfKVBVO5DskiXNJ8kh73pclz3iTcD
`protect END_PROTECTED
