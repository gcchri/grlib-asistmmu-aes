`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0FgcDVwIW4fVY5ccZ5G8Wi09vzqwDMechgvaqBZmobjCEsQp4R88GthZQ16A2lyP
L43+O3MoQWPbhEJLX1xpvpEMxA9WRybKtQP5/HlRM2F3SWhnjgVoVvcXbGim9ZpV
jQ8sCu0AM98w4fHEVhGmYr13Vk4G+obRh77TrvLwzHRJ3CbWF2UBk9dNhDHqYE0s
OVVlVHxB6PvoFfAEyIIu5lRaGWoBN6SRcxazJuVvjVlIhAaVXbNjvKNYuAznhCis
BF2Cl+eLq5y/u230pG3zINTpXqOQX+JCUzoUlxmcfDHIiXos5pTleLpqAhPyyM9E
f08Q6Shc7a0/kw3+7kdnDG8i7LTxtqMWHpyGx0Ctm+n7xxq7jSVZiL/nxCdesx+a
QC9iCEO5Jbav7eXHVckqDz02XyQBCR/etM/1xxO8/Ev6596dSWVDXbI9C++DTqAx
GSXgxmqMnniOsd6TREZZdFSRZQACykO0JZsavJBDPPU3DnkJ8a8yvt4uac5EVEDB
Zj2fybFPbiKlub3+OzComOHyfw1dJQDv3I4EsMS1s0wlSKJT9o9qdLz5rjyZDcxj
KjEBOT3iLgAV5s1Wlx48QQ==
`protect END_PROTECTED
