`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
21trC7tp63Vcxnv2X8lfUkh3D7DTG35VbsHRmzXPCLJtIw8KHkBjyLDx/BziJ21o
wjM2pH2Qq8KS9OlTAmNROEBr4lAqOKSgtetIy714GJU1gVCQ7iBVO/TP5vNqFWIq
LdvkxODaX5g2pLrHC2hwFe1Cv2JI5TP9z5TzVrjvLYTsDU0EfaWG+V8aybMvNjEv
uRG/WHsgygHirA2do3I2AjCzRlnUQN+yrbG/sBANHLQZvN1sdTVjKN2d0guPWOuV
emDYzxVq212wEY/4PSKzi01UE756Cls6nDAqEgMB71svgyShe0T9ITVD6IgVK/1y
JzEddk/42Nh2bn88rSOZTbfdKWJtAv2vI+7FJkea22XIY6BpvkITt/ZVE8QF1px9
Vwuc8xV3MEF7MDMo9xPF7Q==
`protect END_PROTECTED
