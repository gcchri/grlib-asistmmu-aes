`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jaOBfOjiIlWJ8DcxFX2R7IS1XK8dwr26nIZS0Cm8L3r0NcbQPsA5XJFFxkpg3aq2
jrDVofJEO6lht3vWC4/kHxkT01BX/uS7Pr0EAPu6BOpTipCvzc94DBtpu4uC6VR3
b1LUaOwh43afgXa2iDqdiXVFPoLYFojd8pHA7t5DCOw543vrF2mfs0OA8HN98R66
ar3q50ByxZt+PrQvRpj1VI9wJJvcOL6H4ZcwLw/WI9Qvh8DBwvz0UCVmFRCy2pZV
OpBWOkF2nU9fyyG2d9uqIOv1He+LqEayn6atC4VUdKEpiYKgzKCuPvw9tUeMtU2i
jRQ1NC4OXK3arm4UpX0muuZEXK3na2O6koeIkA1a6VKVcnBdbTqyHnRmhvf2bzI2
j1k5MDkEcqxCR9dpJMPzQIIiMefAbQg/clah9xFKwP1fKwlFTfIKG+Y+BaY/K34z
3dh2TOOU9jpxEEnUdlcCnz40hCpqJbV64uEhBsGIUxtSJDHyiEcfRin75Pg0Aw0N
gXz4yG4WKT9nyTY6LIpeN1oNjaHTqf6cZ/SyoFYVI+CIEaEMY+TnKocBi60SEDxK
iqRCISC1bKYkdepacPY3iophMo6SBeWcxYaKySQVhs8SnjvG7I66qo+58/p/RgU2
VO5+iXPmXwi6SZFBqEYBd4C1uVoxow0nWVf/P1FPwWP9X2DFV6MdDhcLJ5zoDQqu
Gpo8LNS2epwAsgOzAxEZPOByDxuKHNvt/1868wlD8l0=
`protect END_PROTECTED
