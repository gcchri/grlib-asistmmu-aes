`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5/YB19+Iyc7qewK3lvdgGh1HW+Lnz48LCbwWg68Jtv18I/EJIGANZCxabnR0ehRv
o13oKlBWwZGSrEWEciMu1HHYUT/MnQEenwSIzkp2TzPo2Nfi1ROna7UDQGwO7BRR
CD25Sy7wzSjpNdfc+NBOhA7ZjpLxPcDmcHAtzUJinCZFEz9UulB5/U4o2SuEtOZ5
Ez8LUjDq0xPYjNTs9mcSvW240dcYwWRi6XxiB5cSfRc7Tde36tPH7gzDPf7HA+vh
vXCXOxhONXygQsKr6ma9r4ReqYJh+JsvzKbi2eI6arlckUSEHDfIteIjqKuuSZ1u
UpCCHn67U7P7Hh1mNw8Vrg8B7eyiAbx5QRjiPjFhcf1zn6/gPXYhzSQVkDITZQhX
cYlNemTZ4kxvisMTm/gzETwzbeEDcnI0wDmd2jFM9vmXC5GmYePezNUcf23EZEIc
1RKdoXFof054JFgqz24/s3mDp+/b6CDhJdMFmTLbChKbXofySDbim9lJTwHWo0Pc
UJnJk9yybazvSUcreFjZiwruUPPtv4N7UDC/LaUDqoj5jpaBPO7++DEtCBwf3eA8
SHGKEYy2OIthqqAFf00H0n5T6W7ZatLbm9+09rRTYtffpGxNzosDuW2JctrOVMdX
AQzqaN0hYFiT065bV57uS2/nN3D/kjsjZ0zy6GmxJ/5j6MO/XwxC0xvLbPs8LD7K
XMyaFe/Ln+J8iD4lVm+urAhqAfjdAeDayXMFZxlgYwL2i9lnj28EansbaYLPlAuP
zOKeXe1//EBhxYyIhrhcwOipQTnOyAYKwG1etptlh2tXzdNKR3czm4zbmeUnznAt
dXPfqDqkO3w0xGhifNHqUOXLadwBPjk1RjTaTPnzBqaInXzz2PZKWoWNLC9zBjC3
64fZwz+t9wzldsVqA9be42zlGZAUH2LdgdrXwdj4VzA9VSvwHmI6staBEj1n6mDs
NKg+9U7utd/knra/toAbBZv9U0AK5iiHn9XUdowxVc3/r18j84dCBSpgA+A69AK+
Vh6Z0QmCITzk6qgnICqXtecs+eU6dk2Ia9X2WBdSTyllPvOS1HNLm6OnY89coLpi
eJ9q0a3+TD3n7NaCW0csFXaIFsVKSWfhei/K11Vjtks9rqHnxtik4ggIDnN2qfTa
rQrEvNiiI3AvQm2TxwTkp+6kuSEk3YVEofx1+bV1TP7hGHS7x+6g3Si6JcfvJjJF
VsxAzvSDCX8m0zDgFVHZmjpFSP+k5UQOAEVsp8Loqw4qkExItlrbWwAJ/HEfnZFl
/EC68GfwRsEFEy4QmAmz4CZ5SH58r/PBpFN4FQAO62O+SjegonPdvF7dMi1iA3rG
9LBHCLl3ihxvqCk+udCy8+bbHbXLIVDnu5DxJlJrtVHvH0bvF7Lzw/toJTW8FKyp
BOs7RRuEoKVl4+aLQ6Lcg8w8U0PG6UjYmqy0Iv4puxV2+XZjIIkpKlhBlm7G6Ejq
Mb0tc4GA9MMj+aN5jVAlYf+3EkWrMH7iyuh4I4xVrV6HFf8jOhBV4ZFt1fJD+csK
eTqpk3HzeMIclKHx/x1tb2blIyVzWRGNXmo03R64CsLqOpxeZ1MkH0CRYBJIrw/D
72Yc5xyWIYdH7W8WR8LM//7YlhVbKCHZoZsfJT8BLWIciq35kkEts92GCBBPIDqB
ekVt26hmgu84g848rABCmWMMqqFrZe5ctaMsbe1sWxOGzq1iVKI+g8QlhOqifRQQ
6XLxWqKRXvkxdzJyZzDHlQ49Tl5tPOKkUzsGkU+KVceSzw80K7cpkqyfS2TxzbKD
k8uMoRTyQ9dmPUb9mlF6JhBnrZQYiNfKiYX49wL+PB8ixrw6W8fphq8lipPOj6BN
onQv35sYpj+T2y98M1RdGY8AFUsG0zQsclfwfaTcktusL8r08i1eW6KxoxHv4dH0
+woE/qaSSIJ8BIu/lOcZd/+y+VmLyPhP73CjuRDDT2Yh8wYfB9312KD+g6t106Kj
nszR9mT8iRYf019h5m16bzHUbns2NjZtgTdMl3Rd45A0IkZs1XxBMMAxA21JEW0T
9Oy91PkEIwUKyKrNRAOOtXnlT6ds+ICPzgUoRRC9O1Cuk6CB5E2JqnQS+8dJf95l
tUFQexhAUq3EPvlnkaB+7gZx/+cQR6kFX+RBdOGd/oljkdk5lOUHuJdGffkXxMiS
ttWXK5epzKmLov8cqXly2w2ld9JnAhzYqX8zsEMzUcP3p+0YAubocrrDqZ+pkS8X
+G4XuaVMkWra4katlvUed9wjOdWk0krqpDTwSe3l3Xj2HlbqQUQ0V8GpaEJvNZdw
Utx7oiFm5U29WJnJCNncgP1wNKk3vu8mbRh10NgVGvFldeiOtRIMkfDzzJphbv2d
TaPY97BnIGnZc2gr4wTIBPPUWQ9HHgdWw4hSoMw/imvLGDdMTrxE3xReAEDUGy6N
+eCSXP2LL/XWcQractPyGCpmWCqiCdb2anMsQopt/qb4pAk1SDUh4KWZe86Oai0b
7H+7rJEqHMwnpLbVAbs1Azgdo6J+Nu+aw7fMbP1IcJ6TtMd2fwF6OA/zLeHm9aCu
zKvBX/A7YT4xXF4StEEn5JhT7rRshWiP2XJPGdMx2K2pLjSsK6c7hWR0yW1ExhZH
oLhMzLNsi0H7ZfKz6aHHsRA3d/w2bLui4S2Gf38I/dPtssftJzmSWFHWeZF98wHn
NwpArz77TyPbX35TWvOxyM9ShEo149kfSTYkn3inrt8q+7QftsDfSCGg9cKwIAXX
iRWEtifJyu90K2uCci3yewlYm217cYpSTITM0Flh7uMXDiz1LMAk/bQFoH1tMgo5
UoLdDABSgBA7XSWESB8vkiQrr48CHQlNmU7onh1RrmUeWVs7r32Zuxir6N+vAAnE
ZoOLYqqkw8uT1aM79k5dgYjLQmRoAHwkDQHR5iAy76BtNllGX1Y0xNB40HB6DG+p
pX3Oyf35eWhQI5HoWWPa/ppyI/fVo77iYy+3B2AwXAdcp+zVNriIJe81nDRpYnZY
7GW06VpuIcHBXJKBXkEncbcVljIERbEQ6oDlSRbuZbu3ZYR5Y8XiCbtL8A+3BknA
IFbg+dBI1JEc61sOenlH+iJKnSyQs3GOjdl/rV+WLTvhX1u5cstfzVBE7Rvm26t/
RiMrffzqijDZuA9qP3u+aPZNLlM4gxQqmqmL3DAzeGEHfu9vA5X7rMtRbl95PnMX
S2CUFb9tlJMfbHSepyT5ZAWCuC91GinQAtwFtetPpF81XE0+awZxVW28gaNQIji5
55nxwnbCdJA9/uZYmL9y74qnyHPNYBov3VRdCqXagPh/MftiL1gVmlabEGDkVcXG
HgpKE86+atjjwOBH9iHubBOq4YnEf7hp8boZW0y8AnEamBEvucursL6yTQdU7GtR
xHZd/9SlOlKUZQPoNt/QKsOEr3Rx3uYen7082X4wp+M/1nJWen9LMaE379rTgOL8
WS/lSz1U3T0dnvqwqJGDUBu/7YTLd2UmY5hH8OhIRdQqfX9gIxEw2uscBOg5bkHY
7kFSEczASWUerxwNr9+C2wDqbrUWiHkoKQsEiggCvmoIxXDC4kE5UDRXE7W71ExU
Oit8j3smhZWKCWNsy75Ciekx5ENhr2Q5diaBtORrh0mEKt/rAiOPsjTdUKjLoCf6
XAAlcPLU5Fdt5f7bYh5+SrXzah5jAAkSSN9MRHPe3MXU6WstocIMUnJ5L7imYDB3
fsW+WOp+MHwYw3Q7YDOBkx8A1fQZOkyeGyxtfgBfNQGI4anrwld+esIecLmhTKzd
JKeEuG6e7yfWlK66gv7VYHqXf18+A85uFCDfbPVaQRfmDa1L0P7CXeTPMsGaaM8r
whSteBcs/P7ya195/qB6Tq2fuV45xBg4iPsZUYh0J4kS4gr79w0eTqr9ikY7uSj+
a+cvwjQ1Z8BkEP1wqmkwfOet9MNxg24UhT/PYCLE+xWKtNMdjTIdZkgsqSyz+akK
vpPotIplu4AGXu54XIK2iLXIUHw89VLM1qUQeG4EtvyHgyeDG4BgwnqJvUKZib5+
kmRl8QThzq4uaBx9iZIxe2kb0USmVfsC2ZsfytlCBrFA1lAngCwivPLQwbAziKov
ikcIoHdfCu00LI/xaj1vWyTPm7Yj6wRSj10YdwkI3nnqmf0P11Cu43s3vNYTJyNQ
dKcdGWkerN5iA1AEEbqPFwijFZOaqVhkoXZqGwUGFKDKgL9iW3F3f3vCaengfR3v
871LwColJ0gkf6b274xk/INM4JcwUcywac2W2sV03tQP94TCIe/GOIRmBXSsCo/v
27GUMpnjX5XwKPwI1i9y5JBkXD2MLgJpCumF9HMUvrOfbfrLVJDxfDju+Woqsj5F
p6ljbuCxpT0Q+hhC5E1VaUFtMGibLSr9dB+kBM1Xp5x+kuJoMZO+u/XBsPsZXIU/
eLzjLaouCsiNlkmueISx0q3zzv0NBEqvmyy1TxETcpOud9k8oor00TPk6JIjtZUx
pvc3sDs6PkL6MwVz05sm8nCeIXgM59uuDliyB8EjGi822MwiPz8PhcnEg6jh9ND8
LMmDgQN7/ZPg8BoJ0oT6tR7IF5C3MKJLDT8oegt+ZN6I4a6LVyCH1VFh85AjSYR+
HYjTucbs4W11jRGYlfr3N7xTs8OOSHzdmn6F6j3VuxsW3uRh5cWV+O8sZwDDy7ix
0n6CoQVaENgos0T7ZuP9tnmrwJMFktQXnN3ek+zgd9rpCD4ud2r2sE0Eb8aVCx3k
xaFvNOpqCEaGpfMrYq6b61LsxN8nDU9AW5TX36ZKso5P2G/TG3Dw6HRnqsZrRtfN
/tf/qJjlWrQHWIRfnWMpLf7ZJVLIoSx82IXjlVIpUTD+F9L2Id2Qd3lg+PLszZ4p
opuZoyQfuEedpZk5GYbOHyE1krbAKaGbVchsQSqWNzVDjzP/X9VKLi/rPDQoDC4L
XohNQTevnu3sLKP0AfojQ/RDl8jdhOjp78qrBZwafoCJX8QDSr/ZoOJwzKGxy5Pb
1Y2xTfRfox8HW/5DrxL71rJbcdwwNglx7sRoefxGOaf6TLce+p0A3rn2OkH/bkja
F3stHpPD8o0eK++FYpdAVJ7RgOPvwLbeSykFL/w20QIrJ95sHkw+CYGCohzudgBw
n7yBjl+pJp4kmzG8Oi/tBV1lpriZd1ImsUDOzznxQhvL3b2G5zfwdfxUExMkJxwf
wlaCsw+12QkXRoOFQB/ofwrS9YWSwKNDFkgRkm8KPookIRBqnShzVoM9hqrX4tsi
og18etKupgWp4avxsmrUh4ADajqf31OmGaWvgDo8LhTpqf95GozgdhyKqVH5pboG
bXTTko7pKGbYQF45Tvq4/dduU5UUD2g9AesV+85npBqlk60sI0KYGNm+xALS88dy
braZI2TFuHpoi88Y9GLIXDEwCbDsS/fd2k9W1hhjz8TnFHpe+D6lHaLkBZzin8yd
boat4Dzf5GEkovBtwQaB+vW2b27uAiUiA1tUI0A5CKrof1H2PFg/wpcjrA6Oj4vI
jrUkEchlB5jiZcmnuE/B0eeUcFkiMrw7tpyJI7eSsUJ7+R0DOueaWX+AzkxLCmqE
pOZvs1RaDNERoR5YSKSb39V3lmjARF/ivQUJ++Su4jjOvvVUKGMzGX0zCsqC17Pg
7fGNoSZTfluUfWaiqO9hyQet4idHh/1JbLItWdX/5yOmjxQgvuQXd/ui/Z+I2uCJ
SXnU15E8RIbev8h61y0BxKZOTt4IXJr3pG2ee9ctGrRpUp/lIFtSgDSHsicFFbL4
Iab9EfLcsWaS7dh0stRFyn+By+3qE10eeNrIGmescDuKtvyVzoXSrr0m4vNZdycD
ePL6hUNtzWzDqw8JeN2DIRpuZqW0jBlMTsf9HgidkH4CurAyLcjaDA1I0b6LrDpB
RyjeKCC+CF/r0y4VFl3dy5XmR8ou18TvlJzRtg8LVeV2P/NK8qYAyq6WMoMJ7XKR
r68gLF3naNM2QCVG4Z/CX7RDe+x0vpROqEHi9L6UhR3QVsXb1SyisdFWw86uij8I
RBdVF2DSHh7kfBXM2uEcsz2uUtBIwKNgDnx7p/8m4jR/gw4WaxiXBM+A66MbG1r4
xYUkLTCR4mixi/OkAUOh40Tx3Apj9TsNuxpp3QlaDX3wfAE6vjPHrbMdBF2mOnGH
vp0CZ4Pj1stl9Bg9p+4i/LwrPIkky/+QUoIKiKHalET1ZG4uEwW1VsC/bJyvKYXw
u/NMV0RKt365nyxoEAue23pY0SaPL0JmklYIeLE9kuoF/y80PzMejYPh6eyNdFpi
sOI1fBqb049Mi8s51yT4bjXkfg4XrjGj12x56nWzQ8UpNSb3vKEJZyXGgsUYbt6E
ws9wjxhmAIGLUT0hNcXBq23H+wuVig+nPWIQOPd9sf69hVJw7MGSaoqEcar10Vn6
uvXNgIMYIFbFlQ9+0VBc9BrkPQFQhaSA2bnoFLeeBgcpBRs85ziyA2AROPe2IW6r
8ERGBcUdzoT+lWDKhcXTIUYfcccUPKfbDrc0NRG2Dfc65arlcskDd2D92tOZG+RZ
bPs/3jGozJgJVYBxM/E9F752+sq/0/p9LJWmv/S1E4+i1HRhmCtR6VaPIMtMjPDh
6MVg6UomxUWdOAu89q4QcEyz+yYmzqt2ZzD3SrYaF0vcjrqvr+mrkVV0dEGNRkiX
+TbVzz/I4sfXEiZwPeMZNsHaVHtNsQ5RT85qvnszwFgNDguQZWNsytKsw++y5qrb
G3d/p+4HKB6JCPoMvjlBDzRj2lGOoOVdCpTaUSTbswVKeQiZHnLadZkmTOEBXXWR
Yp+WOXE3fp+Y8NBRsmAsJEdXhPZ/S2pYjFJf/JBT24T/rVomgpnXjkwf7VxCfMWu
nOzq05kzE2i+A56JgriCMT67QvmPOSQWvutb98+TM9KZZjACo79f/mw1ByjEktA5
ndRqUJ450EuhM+FHMXMlApQClySBxTg35xgLb/mW0l0PhHSsIyfW9hrTFKCOYsKT
0RtaN+bZQTkOSUpLHrwUcoL19sRYxNhcr6QH5YQeUHwNtAuwAgC/EvGGc4FrQjJ8
s4C2gYrIBu1DRkfR7M/mTMr2cC6MLoChOrKqsrV0d1f8T8EbwNwiL4t/4J/J+DXz
O2ThAfkceBC0Tdm4KI0DD4O0XxDmDO1BX5QlO+bXVg401mYV0PlNO1Ler60W93Br
jZZzpnMUwD3/d+1WW5MsgYoogrjwiFrFcC1FMcmWX/09IBI9GGNMmMG+nwwz7BzL
ZB2ufYNom988ULS/siU3J2YqBCMBMT0KC3NuEb7/2S6feFLA3MU5HXiCzCPDJ78I
m6d8JSkQI+yKPdbMeoBl8FYyqq+KozwZQK2kc9NHrB54d+7F9CRuCWKKtw6W7BQq
vy5RRGbc7O4CUGUcWRPOtWMaF045sVQBsgNy2AOd5blQOGoAPIzYoxGW4omimg1e
ksp0H2huIowyVCjrxoGv0nr9OxgjnrLsEw5z7gtwUhnPyDzQexOwcEcxFIClO4OP
hmtxAHs2OFXXr/H+qmJVvbwGizhkcovMrobPVKx6fiGKiaFQmStR/11is014Vci3
unZKmxYkdUzp6j+NEY+nRntqsQpwY+JmA6cJ/IGyJT9O8Q0/0FurpWCvn75hOaOg
Xm9iNW9FRE80x6/uKtg51lhtZWa6RVzM0SZy+l0kSLrd3IVLCMXJCDX/HZkHIV2V
OR6fmGDN80oInSp1eOC8eii34c2onMGcBAqxUmUgDk9z++xRw0diwScCLMjzEkxC
SdAGcXVFxUT41R5zf1NhEFfniSkQT3Lba2jp8zQEpZSW1Ko6fSjQlFOcXGpR2No9
hiuDxkgt9paSY+RblXaqr/LtimPpVISwbWXcu04ZpA0HD8tf8D2LKLxQ5Udr/g8K
FcX/ecuw4XloBnKhOcXGoaqzYEyqvVKzaeOpAFkYqVwWUo3fbkVf7Cc8viPOfQOC
P97HM7/y6joxw+6VB3wXB6yaK4q04Lj9xiH628lugPl9UjDTzhVo/JGy19YzSwth
KyVKl/y98Y9h8FWSN9IUEiKiVo/wwI3T+uEbjMUWa6OulHgupFEZeoC8F2mYTXRK
0D3OZe9T6TZ9qc1vqpz4Wr6jYuLejokrjf4SfHR0LbH2GcsLtAXOJYe/Rz6EvASm
hjK5lkcrh6qx5opZ6XQsr3ibt5G0Xv6g/T6r6Yzo/MZoCiP3I2h+fVGxtOYPhVmq
LMSwu+Y1oxNkuDESPebOOE/qj3D6P9cX3HDngJRJdzVPpK4Pyp3gMfhYIWPOhg2c
JxeG1LV6yjJ16/dF92dzdgbCC289BMJF1DxIaI5u7JyQ1Rwu4ljLAAYp0KiZLRzf
dTuSrK1lborMx+aGHhH30KYsh2C1aH6jTnIzkJ/Rwq+2DoidsYPK27l/29MSAyPR
495EE5rqtlOLkbBCVSLKbTi6LaW8DVduHbKXKb9PWZhuqMZx9/Hn0S7q9pGCeXlk
fXkeKBgKoNr5J1nyTNxLUrlEdYPPPnwq2AC4tdRilex4sWWoT5hu/gkKtzXfwa4E
xGhTNafzA1WLa5dtn0B5usMPtgzRep2t6n4qavWg2EQwwllZxLxf3OLA4Sk2M3Ld
7++EXLrct1bLZ2VUz7AR5y20DAJpOwX3Pb+wR1buzF4sjq2mGC+n81/YcPCW97p2
92PJuL5u0XpfMRgruZKhrUf+W6j2BAa846sPr9hobg8rMMa1BW0fV3XOL/CEdlSW
dCUUBdcpzltsQANJvUc0ZiRrau3hB0Y5yTLIysv4hIca4+8aH8VMrknC2qvG8Roq
qHfNHzhm7u+/GQ0wxOEJAOhsuqPuHpZYj8LWYRvB/eYeaqggPCRpgGpeyJv0NxAM
Ekk5clXVcvmDp75QlbNZn1p2J2M3tSBUC9y/JOJ+2FmXuqu0MBod/rYPpvEP1WeJ
cpKxKD5SJuKrgtCBolt2I8IotdoORNPXaVScn67sOP69MTUuTUdS4udPMurYPxlG
gHvpDgNxQn8Pe43TAClG7grCE1mNotf0QH04ugF+cMjQ45ltf6A8PhekPqdJHOH9
2KMn5TehUZ1mD30i2MBVvTcgacUM9BwYrLI6PSZPZeN1TqFiBuyLkWRVzGn3As07
cUxHqyWWqyZIZDIjKvNBnKwmyvaOqibd5D12424caRdCdYNA5rsCh+JdoBTMN9Ec
zvXkp61eQRnUhcHyVb5i2Yf130mPA1I3Pyhkjo45lbg+zHnOdKfy1mCsiI0+Tij6
c+ng1Ci8yk9dqgNek4ZrzeSezLAmF6YA1JWP5acZ6HJO0AswOQS02/Ck2NVslb2Z
1+/UAnOJWT8/0NhLduESG8BV2Ut0sk1MRubg1+URr5pt+09hILCrEJIgVr2D5UKt
v0PBH696lDa5jY60Q7RGM2g/gGzcLUMYjh1Q7S39Z1JnEF3UPgRZy+LzE8+4sS3c
cKCGGRDMZVjdVAY8HEUzrRfhjlAAx/2tFvnt7s5gcvsSA7JSqS5hYtS0D6cJ6XYQ
MMzjoqutsFOBknzIQXnNpdD7BwO6o12gPpEmKXBI4XkpHnUjIQSIdXzsyIUXeawd
LNCqU7Ti6n2UMfTdqe4h0ksWeM1nE+mfZ5gcA045O9/DmHA3Ip93aTUAVDzU0Du2
MeLF7p/c2a02qmsoxspckiz1Tlg/Y2wK6+MDS5DCj0xBjGhCqwAZok0iH1HPjajc
XA0Y9V7PGEO4L7q2givMztAkCIeWruaiXXTDCYmZ8lgnL66LLOWsmBymGKhaqn35
I77jN4ybt6Nmtq6rdDf0jxFmDjV4QiRh0wPjs0paPN5epL9UvkwrTrAwnVEk7VAt
igxpEzooG5w6JTVfqitZU9FBNkD3IxL2CBuGKCTHNmTMCD5oqDv7rRaEX7tkZzAA
ZbOwvRBKY5H2KjUyzbFbWSLrq8PkkiES6TbHAUseRx9Tn7CTDZSLgNHAYLweALgo
ue1dOr8fe65RKYaPfINpSMGBl4pKsEmbRKG0CTyiwXNmLbQav/nAqTei53ahKH/I
dJpvOHw1feTvEAtJhykntKnoM7OLZHEAyavFut21SNVvb32SPJVU2TeA0U+cc73O
UyiX4Ggi0WKm5kMjKaBItcynwTLh9nlXOZm4ksB1joyz5bv+CrspiUyrU/L/6Drs
C6OpHaLnMn11D9wSskh109AYD1b9LjTRs0CSRgd2IDWrCqVyvePNaHGw0k1Zs0wy
UgnC0cP89B0FGLC+RgWHxxs+MeYlHGPi5lPZtOIFqqLAKfQ0jbJRe8JkfARunvaf
IbhTsQr+eV1UkIbNbWxbKMAcNw62iYF75jwCki/S8jUzQ5ZUD3PxYFK2pfNI1tK3
xvnwQgG9YXSMBkk3FNgJiY3MNe2B6zAuTn6HHNqBuUX8tezoiWp1fKZ+hKhzlLkG
+slcxVP9o6NXfhIoxsKsn1L9l9Xg/4oqUkMZXDbBeVmLdPpWcKGxL51XgZndHDle
xRD8l7W8Kjht4KlJtQCgdUQhLyaEiLx+ZCOm0ss82V9jUu0yy5jxO5t0e/yOc/q1
8P9Ynrl9nzUgXyOsFqC4MItOd/9LkFdhrTFLy6w4dmcfaAJYoCjgj/YbauDcoG3s
yXRxiIHKepn+zgzutMACL/gLFP93ikYWlWjNtlrmX8mlQbE6rsXUMRl1KpZgU+nU
5lu45ASF+9YgTzaAEx4CcMAg0m1YROQqMwn4qedkP2VkaT8nLmvF0TnXKce4SeLR
1Lhywg7aM7R3gk3HLwNSmT0p7h5d8jHp1Bz592VItN5sfa7V3MPpNZCMd93hAt3q
b77tIjq3UrZLIIOavXOgqbsDhRN122gDUgo5yh9GxtwoR1uAAjpcP3JtG3naDi4/
MFrrgTsE0qGZUIMJrRpk72Pt1uwmNvE/5nGUAIIS4l9xR4g2zaM6wXcdHCBIrC5S
4UjQ9XB3SfZdfz6zuZW1bXCtTPX8Eh574YVLtLsvfTxo7CEN+aeFy43j2aeaVf1i
5WtF4DXkCdhQHjTHYrX7Q3H4/tLebVVbx4ulS3mzBM6Kp1xxwDWUn0EVaJ5bw2Ns
IKaPQ5q1tLOIKQUJCKxDMK4JUlsDb0TTk9knyP8c8+sw23FhS7yeP5zWXkrKkSCD
uo1Oiv5pXgVI1iwRje8kSPbieyuz4PpOZfTVRpZM9oEXpFK8pBVQ9FZ5hT5b2e7f
ullCVqSokPCoiHAotsGthzjj6XgsJu1jZaISnGIOXgn6HCc/f+CVAr10K+GAYNCM
ZxuduXUwf/mWBy1LdpEl1PntxlZh9CpMGVvExL/k4iI6D27GF243r5kGGxxf6zpN
flTOXPRupCwugw+QCI9A2j4Dfrck+uEYJeugdGkbf/1Bpy0XrLR+OzCYDdR1T62M
ekJPhOY8WfyaZV65qwoXPQoHwvYlLMXanoxwaYKnDq71P2VOzGOe+Iq5QeMSyAWF
Ryl5ijFdnT1AdO3Fc0nbXSiHetu32UYBymgn2Nr5orRuJZekXbSXf/kfULJPlbLR
wFK6hObsau2pBt926f9UkFO0iyjuNQhWhzqG/RcfaSILFm2CHPE+eDvsRjNmAhR0
+nL1D90Vin+GBRWI/p79cWomoz9BLmnkUL16AnJOF9jXfe+gh4OJJpZc9E2QFtke
Ru9nh1edw53R21s7ZW090y1h1OvYsCwRZNXr245odRjhQjzJ9l/PTB++PBfl6ax+
8FNQzid5r8b8NJJLzpjZryA/xCp3GXkHoGO3eCjueZlq4xNpKvKxOKXxyWEUTBzi
3jth/nVlVzHJZPO6FoPJ+Qhxwf4h/diBNRFH/xdfazc9xxrCJpe8nqRVHJdlIjN4
l6xv609nMkrSFTA9ewKYb5iGSvdMwlI+n2Umb9OuKFA5MmUq9KyssonTh+83tmF+
g3weE9JETdSsSvLbXvOQjgsaNe3rH7gTEXG1F2gG7Og3Eqr+0LQ0zgdrEDlp5mql
vuyzgeUu1MFOBOgMoku0p0SPG+qHNLZb+vMi3y/X1m6WxiPl+jweyx/hwiM2Q/DM
pczL1e0LCkdgyYznKYpgCTEuYw24WAbzmdPyIfCeM/xaLkrBenEQPM4GnjpQtSy/
1GH2GZUD8xCXsjrX73o3KxvIJrsCScblaMhyBP0kQ+WRxjyNcZCXmkYl0VYwR0j0
clcT465eI58jgYrzvaGfCtaHljGi3blTk3wck/XL7dvzAap438UvOiJGT+ybfByA
EkRH12Dju1uXilMLiN2aFDOQjxAnSugLzzRCmAxYeGaQoEybQxOY9yLI3oYdyx/A
x2Di2dX/1JLBqcMlOHeL90toHCaDO/Wp4/2uc68e3yX0DdlkN/mQP3cjGhPJGUGg
uXBMmgbpOc6X67ODDYoJgg12PT2CVJOCcrwfwGXsW7wAI9RmFQusBudJ0GlObPWz
a/n4Xm9vtY9N64FyjEzUx5OX1/dvdTJCqWHyPxwGL9qwoDFpZbiF3sTuh0ODzBeQ
VR2EmGd5sUxydDc5VaL6zqisXEgQPItteFY81vgRyZNUErNvN8dD38owsTxEMNFN
M3coA1O3fJKj9Vw4RFQwIJQ+qBXHdSeAQc3JEyhZHFa2odwO1DSmtUCmhnfHqhnr
fox8/L1iX9uu1/MFOgOhytlghaDULClCTDTYZrH28u053IY5jy2VHyn2aGcmCwS3
HpoALJ4tmiJpoDkeqWgoVtzBUkSywLKXo3yIQhTmKiVvLXMv2z8S9HSenqf3muZd
3qz5/1sumLvOgRJSYliEt5fO+Uh1Kw3vBoP/3Wv3sTrLGiv26DhJGjG7OdSi7gK6
nQECkAH9MbLB+jn+8dxeCBG8QdDn+Qpw3vL1CEszhdgQsNr9UETcg/r1f4oLmWol
Uvzle3w1+JJn+cgIxIz2qxyp5uC/xjIerOHqdBTPpCrgHnu7IjetH7uu9So8yXxk
l/fZscI6Dej2QAezQvqZAzZfY3G1KAqQMQQru3PqhUMjKCwJPuMPCHXc04p5xjMe
iLKWy5ZYmTsAmZoGZzUm9t/Bv7w65eSsCnq1+h/CK9g6Pv5owsFqsaai99x7fKdS
ij7WHsYxTf0sdSVUS0/ZmcuswOSLfn7KVXxtWTIL3aj3RoVRzPXqCUJfSxcN9/Am
neIL+bWRSilIvxBBgh5i+R/OypVuhdI17GnlnBOTiq4AMe4DFLiEaogowV5EMGmE
tXgk3kA1/tJuQxN1H1122B60BvxS06EZDKIdv6LTDBNA4CiYmKMIs4Nchzsx8LXP
PBVMfOs+GFG1aySB6hrFGQoP5vqhkwQWe1dO1qxEPfqxVXikpgseSNmUzPRW+u5a
HETs7KVZiPWOoAPE/BcDPv9xYKroz5VoNKdnI7XJyZW4HX9sam7pwsESgm1ZlW0O
7bzfzBUm2UjqwDGl8meeANi7j20LioCITCCgV1PnVi2yr+fqRJxQ0ACbH7itfgkM
mBqu/DOR6TKkhdMzjucDkjPysrY+Piexir6VrRq4c/ldd+vAbzvkQ9S9/xTYO/9y
ONcEXWdI00ukdUfeG05qY0yZZJiH3Cc6omIsxm+qLtWib1asEpRCjf+0dNZTqoJP
V0wzSDUVSCBWFQGUgTYwIoPjm7CTfooEvrj30+G4039ZIpLEWm+9aQ55ZsjK7oRm
ZsP7kZHVLy2FaEZ01jyDp2kJt35Y18XE1mYs91nSAHfH+QlyDMAdVXt6g3nqsx5S
Xe72WSk56EtoGAQ97Qy53yH+m++AeC14h8XQvbGqfwlrYwG6K0VKFHalyvpzS+b2
zHWwylVwWEtpmwyWmMedaL1Bz32na7Ut2LNrbVFO03A1Mjz2s7NTy33h88RAq02+
1LAc1vpr0d+HPe/1WKEyY+whTRMiBYZjZEZb9v8dSosdXs+eXFAuXp3idCT6tIWJ
8fhHYcAeod5zwEBeIdzjmninxd9orFe0RXVZ6C6LTIAzVFOMaQ0m8Lj3XiBgF2IU
cDF00jHWxPyu/42Wa3yI6xYd6UXtdPEfFbJfUi9ybG5sd+pnAK6YP8tQIxsnknNP
SU6z0HOQtoTG1f/BsMbk1EyB+RX/6xpnfck452BJdXhG5ZZZRe5i1jv7zfFnE2YH
Slomx5aemem8i4BIDmnBZDfUzXMUyInOMYDVuzjsj3Q9+Li+LRabIeM+VccixPgT
agD56DB9PgwK4nQMAtgr+qlGw32QuBf5jmy2RusHS8DKZnek6ESI/ne74jDME4wG
3SYoWB1bAoq0Bj1ZnMQ8HI7Y+0mYcY20HLjEDDwcop2BVyPtdfizhzlRleb7wCJB
vPgHmrxNnlk3aRktl0ObBUBC7CAzgtEfsHjo+YYCAYSctMsFezBnrt3/6SX5QUzA
thEMc1+/sF+I0tnizXTJ7XP5syQWfUExkzitgxUbhKG+a3VJrcaVF11N7+TZspl3
a8ynmJwmq1D8bJAbLbxRY3D8W8BHfQsl/SnSuqNtbKi+LlMUWnhRVwD9qaqbi0jn
qp+YgPZtNx1rtespFh80o7yiPjRS+mFD840+QCx1vtDPx98jrFX9pu10cbTeH/D/
xyIeXpPnX5kkhS/I9qHgaGTVhuAnUPoqfQIGrdTHWSWub8b06BjBjt+Pi8wBvN+r
x9IGCNm3/90extyKGTclUhPigXty+pzEoYMrrD6GH18Xtu+xURSYjCPFDZBxvOiY
/kAgVU1j/ylLlslGHNU/HETsp4KwN1zTyCrO9ThPiSBQQ2Kaa/CQVLqw09/0vKyp
mDT/Xrx7SY5Tm07/TY/+T2kfK2/6WfeXKcM5AXmgjxKbz2x1OZlwU1ShmfsLF+60
GtryNmXMVm5Z1Z+OqyB3v4mFdtA5GGfH/k1KtvxyPhdI9Cl+RY6/ma9/YpDtO1PH
XOxXPnZ9KUwHEoD4uTDly/IBXtSl7PTV4Nza4XD84krgf8kH71B6sB3un/8L7FGd
CaGIffSIDUo29aGWEDL3hD/1hJONq9bmfa/fFlcguHWZRM2yLPUNyqCuECIZ3Ytq
KPHL+44ZmtjbSnmrUL+ytGQt5jY/iFRug9GgSZ6v1WWwNNpKXjEnndUjCpXrONp7
E+JZ89QMfQeptp914dSUP3vUHL3YnuxZ03Kk9q/u32ly2SNY50LSdzdiYlmVsYon
9yxqrEkEPKQ797HHqIKnbxaECj87OvvRfn1LuiYrjJi1Ry4q5kM/9d5Ax2VWeg3n
HaqX0OevodWFIPx70CfG9ucA5Vk/hM1YusNtes78kF3YRU4RsI7XEJZw06QoykT2
yZ6qR+UtC2LeDv7QPvF9oghAF7+oP7CpFX4KAzNfF7PYwstnN9WY8atMt+FwYcbS
A4yNXCOP7U6YFEE10hclhL8m0Akan8hK9zGX9b8D00OZI3DeAlBpanQpXnQNNzBB
EVIExcNey/aI5Bb3rBxlH7YYaBKvblkzM/MFqxrYT0KI0lDWhICk38X2y7iQMFHF
9D52j142O2Lp9m5mCFR6479//jYV1OhhfHApoBD5KADPhONdCcRtQ5b2foxjGNm4
6Gzx5zOVBbKPRnjVb7qqPMEKh4+Qks3uoUq1LOuQe+FhSV79ZpynS/wUrV5+E6Yr
Ds9hO2aTn73qGr2Si2OnjAMcLTukrPIHZ0whuClVRcbO740NzmERzIOfZtNo3Mr0
iyMp9YLmgRvcghmsmHD2b4lwA3zzruogsJeysvB1Ui/H9ZeHkWagM7Ep5Vh95PHx
9IsRxCO97P7DqRqYR6YJjhh/xAZa/Czs+vmD+PT3++825bjV62AVsyFxRcpnHU7Y
cVkxK/PQ5XKpVxkazAFV70hlZivf77qmkGC17qDbbddTOhZPcim3d63s6sv6AitK
vJumFDEa+ZzyJby16vCUTbByJdSUPsEgq+Jnebd9qhYgpUBesyvlkntp6GzigV8B
CDO/5DQJ2zvuRC00HKGq0xakiXRlzsAycJ7u/vgVTrJSs+sy67UeDY/g5stDOTW1
HB+Wj8YWj0iPk9AX3tPV4FCBfxpX6s0qsKHcXChj73Pqnz9udX3T782tv1hDEkFv
gAIx8xFQVov6vbfwB2optWezs/HKMILH51ZdCF52dbAuVDJAlUxnfQHw5rYWWu09
qLDdbZK52igFB8h04zI/GSN9Jv3bGqobfaaIXRGSB9dZ8BaxGEfJDDJSv2Pq2ayo
ntorWcyYSjZK90uoxyt3wVVGqYIIPbGxIkyQUZ1PGXd9V9B7zXH/myivewH8KvmA
soUyGaTxHBTFEhJTT8pmkaZt/nob/637N4yJ+XG4/irM2mEAcAC1gpwlbcSpD1LW
309W6mBOS7ELYrbyjlSS6SXVKhqnNrVRmx8KTjCZXQzEpme2Aa4ryjHvWaLkt2N2
QbXSM12Z4JiSSEhrXb3QPIoKjuRgQ4Z7/xiXQaELmQVCO8Kak4nYUaTO0f/RdJP2
ABvLxQJI48CbIMYwPeETO3fThiGulxB7nC3On1OXbqL800YwhvvTe5wle0AnL4Oh
D2B1xBo+u9becgaDnIYXnMgTEA2m9JoCvZ32TOIgbkKgrsMUiV9PyhI7IiBi/C3r
qwudXd9Q30gJlN/ORz6WnOU/Remr7C3UBWyZ3Rn1kYwUK0FUHXoqsSS+RtXU5Ur8
zSYyfxmw5yYZIewPNuGvaUNC3Hf4lvq/jF/aMs2ot4NKlHC1YPmumOdQV2TXoSwf
4adrV4rE29o07BfA52KY5iDQ3voII2z/kZLhDq3DlHUC/523Kuw0stYVkFUyoCJX
6LZpeHWKipdhcZ3QMSTp+nMn0rTACdzRa7Z2HZ+B3Hx7Z5Ld4SJY5IrMVz0MpV4u
1fDm/RWAA50BvwPL6ZS6Rp8aSeeU0kENyayGafxhF1j0c9yJZXon5/s1Slg+KG3i
1k82oIxFFDFNX8+GkiE59IURaOA2+CbVOsQNt/vchvEjH5Hx3B3GLg2ykXVKP3w5
pr4QUx7kNlCuaqmbe2YcdhLJSBE3rtHn6DTG1ItYwPqCC9FSIi2vQyWz4RSPo4jp
cNkfAK5cY1hs3PPTj3jcZYam6ULr7hHn5BmxQg8Clt002F5DsGBlfo6ejEFqTm1f
LoakB82SKo6/t4j/DSLVU0QDrnCbkdMQHEncBcY2vHXh7DC4+ylj6cSzIUysvIsQ
w9DkLCzWiTogCD4gvUFlt7ogsIcyUXBZQQ+qit5ftB9ufXIaH9I4XXUhJ0+8qImd
DAxx25YD4h9koOVGD1e04gu+ke4A8qR9UNxhNObB1NhLT56N69s4a+UiiKRR0Vp0
iKC5k5CgyaHhNCZztmqE+axlLeaH+d2vz3zo4FGK6JsbCOm4OTDD0A7V0EAUIO2P
gZ7Nu+GYqex6ay9k8yL9e3nbjSx//Bmu9TVnfzCoBnDOTYCrc9hF0E/ImUlStJ2a
rEaYa46Z63J562Egn0XvoK6dVULG/yszNnt5xtiEIGvQd+1QZzkNcpjkowJ6cCDE
VONEGBsjulyluGFUJDGFV7M0NY4DQ25a8+guBcoK3fr1okv+tHUJKaifNq8FzxF3
Uu6IG+IrL2xfvqdhGNonGzMjEFBGC92jQSaDdFVS55mzZM1k+Sw6JMsq24d9oLrM
QIUPdYcmP627DqSbd6BpCuwwSGwdrJzTd8A97v6TmPq9pQIyo5weulg3jSgP2UOk
iYHOkGHh75Mu9c3IuEuuhYqFNIkct+AxNToz3GUiCYJ11n6GDzS+ZqJ8odw63ywA
QfIQvOhx9Iu5jGZmea/lBIN1UuBA1JeLxWjtYSqkTWxkzOIZ+T9Ajrmd001TAuuZ
6LuK64ddBKBkxExKCZDSaFNZPHInav1XwPPGn5yfQsrD4sSXdbPLH8eIZxW9lih0
RLkMWhKRe+YDkmM2x4F3CshX+tNU9DpSJCvKj4CAm5QCD64KgcPFvCPTHrFBgApq
vwUjMXV3gw6IFjPJCIciBt2J2J1JmUL2p7yza7Qz0h7UipEQ97n7jOs42qjCR93c
15mg0jF86wwuCKewlJDTXwjQkMk1ILEBZQ2RPekpPQixYYC3xRHLDOwxENwIZFuv
z0RDbeg6TAtRj0dXkzTZBvT8u5sz9l2UpTWlPHb8J9SACiGDiZ1qn+FbRYfi7x2e
7qbtmr6c4wT4ds8yheOyWfjCEziIwB0Q6puQ7+hU2hRPWrRkvd5t967RHyTr6a77
zy5yn46vZmfM0o7PF4ff88QSyIvohmmWA0Vh+IMDrUegEupgqZNw9eZFNhdRFWpf
LsVoHRC+6HQuvLGUBLxLdv0IrD9YZoanuiPcY0q+RbSpP6FdGAlQipLAI/i5kK/G
lXvh//w7VYLlMGsLafjPSnuR+DvdzlCj7EaZ5YV/t86EAt/XNSssO+l1an1j8FDn
th4Ptmy99JwY3y/Y3sa3MPhXvDv9Mikqmf+bCNIbUJr4NgW5gnFwrS+fMxl9P2gN
K0X6q+UrvnWcTW6qjBRC187sHXddJt0iuEXZE+rv5TzfSE05qioy0xTuFmFHAXT3
2ZJh9tlMR4hQw+LnGvxBnO6vwlkS8bl09ZvIJtylg5MutUirGIHjAl5pnsTqNvS0
9161TBbuyl++ATZ0AmMDkTD39kskW8SYiXih0Wycp9CLBJwugiruusdgaAKULguR
Brq1Ju3DLPMr2Gcx1UeCA5VvmbALXp2cBXDzRa5xbs8daTEmRS8htpzN0XPUrskG
VuxT2YCmF0kPcvcRFFx48mIqm8pV2il97pL8oUBr3nKI1CSyKwrdhr5fgYIQ81Gw
HHnKxN7WKhvJqUlEQujkZ5yK9yOAI54IFmdnlUbBq62Fp22EP9+OstHCOfkHlsfA
oyHHvxvH3uXTUYKgE9zG6ckBZ8PKGDeL4RO5CizbEYkGM7kNHknLbS9iOQV4Exh2
adFnXkUZ6xdk5WshUXZozIJdpjTZtyZQc9TWS13PX9B9WSbo3rk+c41VKJr6/+wB
YEtiEttrxlzx7q+8y7obZFKpL3WLtNJzIP7DT9krhB7Za9jgiiRAAYM6JvT0p1QQ
+WFqaVD+oba9z3WecbSuB44veQS3fBdA5h/LkwFLb3By9CGnxNfkXQ1Wfn50FiIE
HsIFHPQKfQ/5hfbLHVBPLQOOk8JQO1QVGfLEvTAn1TmfVXNwH1kF8VryW5+MS9v3
0xP+y/OOYu2RcF6N8uCXRqWbnZ7vkKooTjpIQfAa0c+vKGN2BYHzqg9yxew6INwQ
mZ/e7J2DQ+V38XijxzowpAdwMsFrEJrafb20i0S1dpg++Xb9+BxFtzAla6hlQn1v
Lad2JGMi8ER79Xrra3E7qEKGR7TX4QjJmw753TL5NRFFan0ZkrZkm70QMcrrgRzm
xMIHig0y/UoCNXEb2kM/aHyKLzBfkQipv8VIQNPdmSDrvVXMj7mHT5WoigVV5elM
ReSPnYopkm9yiMNk1SXo354XPy4wJO0gVVwoK5iabrbZT+jI36QJLe+s6n+puQD8
V7ezhTvu/s/FD5skETETSMVtzQe18Q3tyvvxftVuCrkIviq1IrHBSYCkjkv7FKR5
D2OxhbX1ekbCOhTsKBA+U8HH8Dagahe8C6rIg2a9/1el6Y/3NRCSzFUwuO8j8MTI
5zaY/EpYGAX4Lgpf9SwLYBq886/XJzLsIynqQHY7poOXlzEI65DPcF+LRyrl9xEa
OdHWFfFDSyf4j4IuPQHaNZPC2r/Br/YVogocLIbldyGRw4xiJckSphUwUms7l0wH
7auvhbrPrrvjxIdMrJGVMWWv9A3IKcPoVqesFZQRr92XPdRTjyGbYE96/5jWiAvG
/ziMr2dT8gWlmsg/IWOc0qs7/hDfhkmZygZ6LvE3gdALqar1KeetlcBiWnMi/0nu
HZU/HxmHGHx8I+RE5KZK7ODhXaILeZLF5rgkHaauQqFCor1DRLq3xZKoSmLg2X3J
JAARgpi6dY2GfSZa3/0ek7vxzI/FDHS7VKlKEmV55L8ozlRqmPDwgiFIuSfl/h4h
dapxStkO1XCaAXeU0umF0y9qG0IZqeXxKeYxQUrQfegf6M43nQ1wKMdl1MPYsGD9
J8uLOPY++KfKji293fodHJIgwg7SZIdFELcQ6IpLXPxt1BMEJ2O4Zk6Lgkknlnoy
JSKrMWD2AXcLST8/6WSn05xKjCf9B4QE43L7vDyfhOdr3sgvM/8LiouyEA6+L9bj
c4NhHWAR6Zq+kq/6Qs9zwcMIs9wPhozPzEf/FtmLhh7pKMA6ZHPtSmHg9X1RV1m0
XyTu8qf0Hn3/8Q73/0ykc9ZPkUiUHUL0qmN7Eu87KQVBY1KFOpWIhnWVQDGxXBJN
sviC4SciDumCxzfxqriTjv2PSbm1juz9Wra+1+7DfQY7MU1KUvisUp0N6FNXdTQC
E4NaETsBcKz6OCX4JoHMbxXYJ4CYbTMSaCd7RWD1AtmKxUbhpWAp5f3I2EoB7ERA
IbfHQJHaC3zQ9NzyvjIJRzamqrlIoE5GzIoqIXjMi7GpsgcBegWx9w4xIliuvQH0
+UFxQXLZw7BTpYn5OQAFNtH7QpPN1Oxo7tVRzLuIJLpnHOuEgRtTo+NxFjTdld9S
QdeyFtIeU3pHF0MZOdGDTta8GtslR5U57/Zd1OxVeOuycWw8yf8pOma3tMcgskT4
VG3qZ61xG2Txshd2HeVh/yoh+d5dp5kwbfbZLh2+rvsZPGOUcJ1GankU0BeaxftI
VOlm+3wWOegsiQJj8mg5IWok5wh+ZBRwUClpHtGgZ+C1umZIYfcwrWjotq/Nf5ES
wE6n7cZTKZbxHFMZSH58/CUBEVXXKbPJy0oZB1xbf5RpvPVmAdCPGftpk6Uh0rcn
fbWenr872HP/wHIKHTsGlfJaj3lHfFeZwk9nRglIuLbdF6pXIthqDGzYkDWgQ+dX
NwuoflFVHwmzrxB/c7FzRkfo7++YeKSrPfi//8W98LtoKoTYnP2sWJ7KhcpZpWD+
K3rCqbSxQ6gASb6AX8LzNTuWHJ5IfPFVy4R7wHhwKC9+yTllR2v6xzzMwitXXCsQ
nvcX1qXmHAFB6pWtJHABpindHQQf3jAyzsvtynxUP9zwOjgbJPZh40g4elSN5tUq
NMAP9r/ZbtiqGN1DtJohAztNJYJJWZ+BmlgbgtgD3hhGNVgcBqOH7dkMh56hJBQj
uRudgjp2Q+mNroQ9mPS6dHcq2H1CLi9nBknCWzpu50D/dx1+wPrGZ5xENRnKOFkF
4sPXskJTFG2M9F/nNDC+DEFm9PVqBTImL+6BAWJDIV6PbMiJpAjTgi9W8zXWMIA+
huQk9Ij1IseVACgidOOqFq806qtvH5XKmfU6czVfrBIiLftfjwuGGfCOHWwWgavJ
V9tW5BGkDoBJ1M2KB1EG0FOgg1BH8WbNwjBH1vEYEuoj8Vi9KOcNlbZTT00YsWzG
pOTpw9lK/WKspA6X4PScNGxWAY56f9nI2sOMmRyIipRGT+EX4IZL5mKTfu58Mhdg
74O9T2cKKj5Cz/5rzP74tR36HchlWUn42DfxsXcEqKY0TnqFg9KBLyV2jC3K8tG2
MLJyle0gr4sLoe7a/bt2vFeqI8PzJAlzle8HLubaJmU3kAxaP2QBdDZWS8Msf42N
Lieca9c+HwI52NXIIcHJqouckpw4PSG2wiXJGhhm6hdysG+c2OjrR+Zz5DhX55u5
5I0aPgjv43uMo/ZhddKZHEi9cIMIcwUFBRyDe9BG5nF7EUTe8Ob9/4/xbGc7ad2h
EArmwQ/3TzHa+1Da/VzZROO/lg+8ic8OqA9MtP89AFXZaFxngacOYpm36HeAbebj
sMWL0Pf3OcePgT3upBwNROf5Xf9YUvlyADMTI9DFh1eNTV1akLapA3ZrFZnBoY7d
jTl8EYbyIjj4853D6Wj/QrejNNE3zg9mGzOijBmr2A5sop5Z0p3atVY/UwyHJhJx
sjvpbjMd01qb4OJrEmu00RBU0uvybXZwfkqzlHVHipRTjEAIQInXlT+t4yuS2qQX
bUEpiSEZr6E9NrYvGSOk7r32dAsI1k4RutkYbI3CvTetw2i/aEestFjCLohaz2TM
NPPQR/rOQ0ja3ejMXDtqex4CAMBRhFO9KzSHyTGnL6/nSZf8f2IvaXViDKfm86n8
4jsrSs/m10IRStEg1sHpsDhvKajqRyQFfvjs8obGPQWdXy6UdsekKolHtethQ0So
D042+H0Y7CyoLDYdV5OEd8TXFhaLkvCGnlK4ZkZVTt0ygtXWzXkCb1BXnfWIeUeB
gNUoWZhdoqGz/hunHLnvg3DglnuIeMce0yCkQtzS/STnSPNEPwmB5nN0o3jKOZEp
cuFzFjPUsiNNaavixlcpEMvkuPKjw/JFqvWegsShpvcaouCWAJexo/Zi5cmInA3n
ycRxcyew1Jz4p9ulXU4xT+qlBROrJASUpKYFZjBt4UEnpq76M/WwEIBI6RRieHN6
4sbGIELbwWTG2Vuf21GR+1uga/VIkFcDhJJO9OeSZ/JXT24URi6RhZPG8MD3p5jW
i6EUdL26A06h6Ui490hZduksKTs/mSO/2hVb58Wh+R65JVm6hWeYD0i2VpsG/DiV
uUixcMlR5DvK6XA+oIeUpa9DfOA7yVeYYcCncdqIym5UBFwNJ4tOy9x8ujOE0hes
61lalqSP8oijaWcIuMuA0p+y4tCJIl5QNJ41OJSIzgKHHkJcfGeVHHMdooBkHXK0
4dMBogEtglLbif11M4L8deRl96UnlYrfjbp1y82ibCiGkcX+A851yvT6haOwfkvT
MaVjUcnREdKay3dMa5ZS5hakw8TOHf0rRyyEegw5bZGHJsard79V8mmRwv3SgDWt
nGStegTFzlXmVInLbllq31FDbhI7Ki0yhjQXor8o9+SRzfh6rTFLpCGITkGjmg0e
BaOcbCKCCrughH/GDuDnvWddNf3+kYzjeF9dQLmbR8j0Pu+sE4ROXO7yaDUgfG9C
kzytLNPONu1JVq1StFRDLFEgAHC+sKDdvJjFv4Ayu2CKhouClaB/4A3X7+77auTM
6KojagxDxMfh30ZGLmOby4MQfHXaqwVBCcN9r7qxqGMgtXpZxDaUc8DGqRXocN+J
G/k+JtOHxxIkNimQeKoHyzwWsBq0y6bZI/8xWFDmG3FTmzkhS/LaQeSAAQMpIsa3
INJZl8gyNO3ErO6yuBE57M26YhAtozdkJw2C0W48uCcQfIytnsYkZutOnhCil/aQ
zhduyPS+4OviUzlNe1P9o6TMI+flQDGSJ7srE9jYuUfwpEUUO5ZQoJ+8tm/9Lkw0
h6YSjRy7dkUg/a5l5bYvCzMfDvjZ4BP6AotuU9e+d002Dg9sH1CUG0NKE5TsjK2i
vqF67j0KneWZUWKVnSuHh74/fzp6nariY4lFPAcjKMpIDyBS5wBgjBZgUE2I9R6y
+klFUcN8ZTvkm9MbwUdiWyGPsR0iuYeflaIIyesFfHoE10kjAi9+cQc7ciNeK/EQ
uIA/ZFOy1ugrvFOY0sBGHPMM4pTRKzpZ2VzuH4creJo3D3+xOQWEjqxwDHB84axZ
smxin3eCTMQt+7b5WNg+Hf9K7qxB07FlDfUQ8cs3IHCsgy/AVf6QWhTkesutoTj3
qUWzRizozw6PmOQ2xpLpKTgHl4sGfLiBlN8DIL3wnGcfjqkkMvCoGJ28Rga42fSt
ABNWmn4drRv0Srng7mm5OZlIpNCxPXXChoCWkmouT+hHQEFOmXrzgZQEFbkobzQk
buCOqS0JYIaVyIwlJMleKWa+lbg/MaozOPS8tO/C1cJtg+GtR3VEIt7npxjHRaLg
vjUs1YzUmCvynL3u6LZxHNfUbtwFCJouS29/fS+mTcjzHGzzNWNDR88b17UYBriP
SBZyKlPq0yJkbMi6RIRhcfax5xXqyfB/tgYwsH78k+1zhxszE2yksLKZx+hV3NpU
bOqlWaHug9VNfTwt3MbC3Z+oP9q0s1XK7s3AgeUitGaMr1tDFuZEE940naQCAcLI
GfNEusgZeIAithw+IuP9gH/clyO9QdjyZiI7yRIns2KnMwnBeyr9FaywAMF3/RuZ
k3GVfKINknZZO83QIE6jrbB+jU2ijMuP+MrfrL/8LjqKOXkZ69/1DudZebxl2R1Q
YXnAI9PQS8iAM1WGKZB/ECmyhUJpy/LLzNlqzuCXvMLVXtWArbK3VVUif7s2XBl/
Fj3TckeV2LRJspPzvPJipGnYM9eWH1ReE38moE061zWrUKHFMO+mb0KC2a/ks+ai
nGNiCNeAcipi275mzt5rdZjAWQ6wtu6wveh2aKKKzwxy1ClAZBJFlqXAohvO4RCK
/tUCY2p2nCgeFTu8QAXX+f59lzyVLC098yoEGsCDQh3fkmL9JsDQMKVFzo603kB5
PUe/TIHv3/srlP5Q8iAcNLae/cnqUnjQ8nPrTcaUHZU37dYM7XYT/U+1GLvwgO8f
CENWpU2T/zTA9rzFMuRK1f3FC5xTmD5imJLCcUfXMCcB11L0NppI5EYsDJyheyJo
1Oci+EuW6UnJXNDP/BH/P5S9uPx+E8hP5Dpg+Clj6S7Pkt5xdDUklkSRxJkr9iep
L6HtzvVNTBYbmggkE4YyWMdZAb7Nb+R+J+1eJzNxbiBNCmpTcuD5dmD5G38kkEVO
BUUnm1AiF2UM7yNC3uwHy2VKgGXZpX6W/94Jk/f0Cad2zt9yqrVnXZrltYK6zQ1J
+xCUHcFhYkMOt03QGHG0Hu4Fg4Za2Uit7bhc4ktTZWLxcHDgGQAr4i90ucCbueY4
q6lXvI99x5FHozQBl3eVuu8FKJZC98SbUyCXs+Mi6+Hk78I19uMYSV4NzIltUKXd
Yh93aHlfVQha0Um0mL9gFmQlq5jijkdJ7gieugVsYzFMLy3BCejU0bIUFIDYnAfa
JmGWteeeRvtK56a2uOl0huBbs/OmX7uFDzFab1xgi9LBx/MmCkStdsKKZGDqtait
WdjC5AQKUt9hR/YYRrxSVOMJ/MFphlRY8wh5LI7fg4bzMgc/GSEYyoBW19ul+jXQ
B++zCWcqzbGAX1DIHBPDAfBvZzY7Qq6JIhr2EjbMy0y6jw9k6VU9wuNfRyfavAx1
uNOTCyvFGjcZVILVsRE6XQGEaVu2kfQsMKbANcmCns6mIzKoWBxgl90cLqN0HOnL
Zi6j4rzGrFl9Gxt0LivEuDQ74tfUQrNGoNvr0iwEvH1KJ1fWD8XzbQ8OvQOz/jdh
TPywOHKRcl+h/1Br3G8FpUw7gO3vqeZ94Z/TKuNRWPccnGMXYdePBgHxmmOWikXm
MiEfPKJXkcHHDTqnUoCVIT9VlGeQ/jLtrZrlzadFr+EmhZkp8vRjFBH8Expik1bJ
JGqkDRwK6zsrMz+N0XXEV3nzEA6U+pdMSL67wAwZoqpVoflSxyPg+t+hA2sxiFYc
6VqUeQwEENlQttKDPMXlW8QMEffkubnqwp148pELUH9dxEEOQxFQX5ZMwPPS2XBB
20tEFtP7ZsUVTUe8TdXVw9JwNRFOqLTpUUHYf+Kwsjuet9kRWORDx+GChQiG2fTK
ZCUFym8jMqW2sNYd/75OogEBKlIFfPBBfaKBhNXtk76bxXp9qy0ZcIh6R98acCOP
dWEOMMMTMFSIch5CDqpxIj5C1BRuNk09rZnmQiXgeJW9iqGRerlTqGrT4TKVlQnB
S39PaXpoGCfPSeFmMRBZhKfg9XRgwhTTu/QZaAPrM+5QS595bKNw8z+b2lIwUiYK
ScWBZpip23tH751eioCxXxIOQKDJC8aCh/pz4oi78G5vRVgKy1uDIAAllxQwJ4Z/
hy4zVTTHcVyB61ZqwDZCKAZYCl42HzAsb5gIykrwaXrog0mOj/PSXXwTHH2+cG8E
7tniZwE+v4FhR10eOpfiKtHK+Pfdtwdn0LNpoZ5clEPuXa5LHfLHqnBnFuuX1PbE
cIuLye3zgs7E1aO15hIyGXugXap2IVehSWgdCLw1flAxxDGv1cvVkta7CDcxee9+
olW3vFLksEl0rL7mXUaXBr+1iwlg7JdjIAV8OsaoZEm51NTh8ruQvTQ326Rc5w/V
lkVsu3YoxWlKNbK93YJnNgEHFJ7P2sNZRI7A/j18/FnYPfEZQiiwXyw3TWQ81LCm
RceImrxgseGxtWVRmn/ZJwVBPqOPWEzc9EWW3bP5vVgX9h+pMmEJxn2Ez5totEWr
Rj10o0R626A7lWJzNqDGLw==
`protect END_PROTECTED
