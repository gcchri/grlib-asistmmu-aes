`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cnifVxxN5H3OQOfi/Xmtf0yuVDvCHRupptnO+R+zrSgBadFmelcWSiCV71J/bTTz
qtJpfIENv1SWxpPknta38UvAnsi2IoWk1xSk8j9I7VvDoDbjcAGocopt8EtAJoG9
nNlVBUm9kA892K76gJuxRX4J9Fx/bWBy6x/Fov3eWg/EaKC1PW1nCy8Dfv9NusX+
k1CajX2co1CDwQ8sEUNk0hOcNlln7II4cfxdXu3FQQ3+X3XPCs6iHS+42sEzAyKH
nG0XPxlMd/V4G8rSbV+4fQDnz2v6b2sSFVHGqoX0w0ney/NtIkNbyoXHD76zrilq
uBFcrA3Fe99C16p51e6yJpth42s65QOky+3wlXQCmQQEGgel7zAtsxIBf/ccQQbT
M12oLrFIn0TvmcAw3+8MXccSynbNDmNIYYu5jl6cPdgOK5gfuRX8dt7zMx+1zDGO
9Ax3lusK/bECuc5C5Vh+ChflVVHuG2SlaBj+GyaaUOBUmgX6yTRzSI2ffq/ranRh
0M72HefXylsSH1ls2bJvMN44Kjv7r0rSZBRpDnTfjZtrBHY8fwzhzSHkyynhSPEV
LQGGSIuq3sn6ryUMHcsZcmMegfkXnTWaE4EE79S9AF0AFRIsCVasWabCAHdmH0yt
7czqhO1+X40Iz3c/lT8uUQ==
`protect END_PROTECTED
