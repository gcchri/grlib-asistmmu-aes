`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
POQat3UJWf7nuID8uENKuRmzTwaYZffjzZVnfBsTv1CLNBB7nxr9HxtKHV3j3I9G
nstBi7LmrslX6DOQv7LcbdE5R/n/HH18roEne9v2O3+QTyOdPogdEG420lVOLR53
qq7KbLXOXd/AuDy2Prf+Z07JiOVcR5bq/jYY7GdaFBvIJe+9I2EV8495180reTwN
fa69KMzNrpJVoNLIshNHg1jRkWzWnk6O1r7B1ttgMm3dO9a7JZ9Qf00Q0tIlAvuD
6LAXlLRDvZEZ3RyyuKgZTpa9WrWcQyY9iquy3RGy6JeJrd2m6w3Whmp5FutBxKtY
U/tbq5VB6H/c1K3yh37sogBYyYmCCKva8FgXl8pF8JwxZZaUKsslOKYV6FtILGzQ
0ndMvasYhnPmUOqG0x8+hQdWgt7CYrKf++ldy8U/E0pR9WpndC55/gS0p43IwMbY
6vw2h8DIRen2Gcrz+Y7H9B17l9cMPVECtpRVr3mspigSCgISfD2gx9ZQRe/WRgfp
umus4q+hq45JMsUvWtDqYQ8h7/Zg8dtgiyt6hAYXsMKLZHgfqjOdnTMRGFTBjokA
Vbxo41124N+R2JcqKOL5zlOdsg411ByvHnwHzZ944s+GzVEiNL4dnu6F+amyYTGT
rGy7F6tsXl+1nkH6zpgnu+cRuZX++UvzzQTL8H7CDGgfNUntBClEyBYGF2EhnVkJ
mxm62iGPsc/1KvXuwp8xoL7+o4lhdBmIVJAR87vkRacoxrzS53F2uq4I0ObmBoy9
`protect END_PROTECTED
