`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IRjcGVFkOi9yT0x7Krl5vsK/vafqFYR/QjrD5qomNoZEIvCduh86B1agvrgZyBYA
/tx4IFAiRaRq5VeVVtjXEy03FpeGbdt9NXprg2pJtvTre8UuZ37fBRsk5qqIE/84
zG8jx6eygl5mtSCvjytv+3d5MlG3TBQhKuip87top+XZDag2APdeKQr224vFczAs
7Ke0MwoC2sGzkpX8D86J5x2Fwmg7aYlw2rUr9fmG2IVC0PKffhmhEFYNFRo9CLSh
9HzzAPEJ6PCm/Mt1VjOHiy8O1mOq2Gk5y533G01UPz7lcDZfkmOqV5XG1gfG5mmt
R1YXYQ+h9/8HsgYEazIP4A==
`protect END_PROTECTED
