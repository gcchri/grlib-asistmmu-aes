`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sSuR126s6bBJ0Z/zo0RIVrt0ojbHtOEnU5oA539YikSEQL9XIqynzJMpKwpsyUB5
iqtZxYltE4BrFl975s9sMvQ9r9brTs/D7O3q6uIv4tZ7IVQ0IvKx6oTP8VX1+TXM
iq7DP1EX+9MTvTok7KeAfSMJDsPSB4xrKwr3QPnUTtJM1Mh8V/NU3Gg5CdrVKndm
9q1FeXyUSpRoaK1PMk/omOnU8NsPyuy9/VwvtHEB/YHbF6LeoC9LBnWd0DXi8oWJ
pLVWWovMqNaoj3dxsZqInHr9IuhgPH4q+Wf+y6e+uR+PwAj/Z0FRymAY7vtvYyfv
t+gCBu7qQsGuMFmQDPOSINMaQXMi7sRqF6gcD6iQfGgEsBFQfqqL3dilJeCW1NRm
GEq1F4xjT43hdS8W74nIM0mRxk4IKrB5YdxHra3UWhSncK0oOmD7dumf983foMpe
WU7Jxz/TnlP3SnvPMK7WcAXk1JFtMI+5lOCMt+EgXbS3d59tFnOLVMOURZq3D9fa
VD9bx0ACWjAzcQ32/IkZu8TKMmE5plfFpBbQea/kdB/T2b/AXuuoGUUP6Bup+a/5
npQVA7cbOaQ1crwz7VvOC7YkXku7LjABaDVD+/CcvAqtx0Cx15wv+nKxiXN/yhmN
a6+HPdG5RFjY6UZCiBxz9EPAceWWO9F62mDu7TrfQ00eb7LqGTdwWE3rCTo7QFWg
kSEXJV15ceNnZt4hhfo5RlxShBbUCUz8RIrsrm0PvRcuvQuwI4ad1HTH9rJfHBQc
6awytn56rI/Lo0vprLoA5lU/38R5frBOWf+zAnORm0YCOLz18/v9WDTLuaPmQAHE
ZIYU/rCi4zSQLlRIL/hHqFosb2EFXXpDo/TA8JkNyzvbJRwfu5e4X8XIS1TUYswc
2g2v/4fFJUnMLSlKEctyM150RMx4NQK1ZBQnLX2pKJw0pqVlmK8wqqKkRvSoHmix
3zk5EysOHkEdkNaoIRjqKGovJQZLLis/vuDOTK8rwNqrtbIjPCSt6wlRqngCeTvq
3kT86I83kI6QZBl78O6cRC45CgKYBWQzVmUo7Hn6k9aHdc7H2Wx4jpHmick5izNP
AUTzdB3OkOYvyNcgZNuZg1A8MtZvpY6SPKq4EFXBBCXJy2xIwz0pmrkNU4QhxvDP
Yx6awYlKDmlrhRlpWwAoybwlZdz0oyEFEktYlQXUT+v6R9h4CtKKsSYmCOR5nWKe
XwGCj/VFsO3H+5fjeeyk6Ww+sfadYa+9XjpsVs+il5BSTmkbjHSa+YqXOi4/8pSQ
b5Vtot4zHoP9/UcecTC0y8mAVu9JgHDf06gNyllLXQ1ly1xWwSKFMOPahaRMRXlQ
AbQmYb4AUp/J83yYyIZb7xgGGRj+Pse7PbcbBMwU61Nbyusii6KO3uEP9DyPD2cp
`protect END_PROTECTED
