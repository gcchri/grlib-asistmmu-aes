`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MzcuEWHNLCadGKY2GmfZnKPNfp3FHc3q6R6VQi5S8uRBV3N3N3ijmPuAoK3HLNne
9LwpNWIUqNONNgpAHhemUgzzZk4buXrzNHrpMwMo4CrWLBxtwfQylz4jxmjFlmVL
wkEkH5nFxu/XtSVIakQcXgh7z8KaJiRSsmYWrep8mdhInFqBzC5wJIkulzDPSKbw
GPCf/L+vxvDeKWZ9yXNQHPQstQ996RGt9P/HlgU+0nckfWyrWgcZbo6477Tgp2Nl
BQwS4zUbC+eBZpgBh+0EsvVHZEBgYIlmgTmHSb9jzxE=
`protect END_PROTECTED
