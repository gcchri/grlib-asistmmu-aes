`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KIZgZX3shgmfWK0sEpasN7fwmmGcvfjwl+oiifPJZnuv6tpmtlTwwJB0zyn895E1
NhQTwM7S9ec26bLEfVoDEEn5GxJwN/4ejDf1QgLi9GuyXUsKF6A8VjRyXftMSfKB
lOhZ6TAhbOmiuXsVnB4YbiedGTLePE6/I2RDgy63gIFqOAexo8D9pUXOCkkYxI5q
kDYhIc/qSnYUFgr/1Vb06rVE/JwBN8RCnXG0HFKxg2xnrrkB0Rh6G4tfQmmUQZn3
X9vgMpnwAzldn69CNCB8l0wjj9p3MopPWPC4j6l1AWrGEMwPL1BNmcOd76whxJMv
cQICBftBdZ3kKGtwyXAytvFLE4ElAjR42EopZnsTSiaek7KiuH/kE5QIiVz+07t5
LRVUMhaaYQL7JgPCEqzg1euBXEOCalRWcna9+tzfDxwTbtloSUASWWbX+ajB+j19
KeOn8TwGKp1y8m29zlUr3tU2OXM5NPg41JpLWm8HbkL3EGB9pzwPTaSwUW1pEBB4
ukytRgdI068E5W5OV5l92zY5RcM72qqqwjS95JMNbUs4BqAtAtvxD5MjI3dbHDuC
L5YDUp6agaNZ31ruYN4toazsLZAyJZNVUfydvBAnKWlDbD1V816I/JEeS4rrCg+8
puKG0vGDVWiepOI4sL4kHbknyPWJmw4Mq44uxZgovaHfbQXTdnZOF0iy2m5D4MwM
vzWdVdZP/6AD0kkXq3eoUodFQ1RSBTz2n+HT9WjhQiOmM64TWxTdQphb06WJLlRJ
65VOsKffajPEhHbxXNiM5+v2zrASqpdOJNszCpxpvj5GRGtuNvkxS43jGuzJOW1f
tdZ3KQrBKZBdc9pUtl5YO4RE0OAw2sJGhrGYfBhRvBn7S2TOJyvO1sPf1TO+/S8f
D/l5myBJDXTXGgNpwIQke4/a4G+lFdaO8b1vodsEPzo=
`protect END_PROTECTED
