`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pL8DSyDIyDphunyjZ/bMgsPqCXGQ/rcwhEW8mpmSNhH8CeD3wIjmM4izESQWzSbr
NrXMhxpC/ytunhwJQt8mcO67mm0HqmFdxmKCJi4bkek2I0dmlgBewJ6quPWecuBc
eCsn52RlFy8cNMjezYwnxYPU0GI/vAvR9wnrrVUFZiYQQQlgBK6Wj2LVvbqMxnTq
Um8wEHYaaLvgDwJKmH81RY6fwGJGBajvGKmYjV/RS5S5uOUTJiAhextqBmeDAXtQ
+/HjcV78mdIgOYTV6KLP82ottZaX/TKkTcwLe1OzgMN+jGQXqnK9s8kGo1yIOSSR
4SvADGbu9oZ40jJCySiuG2AG15Wfzi2/u0y0N44OnGYyWD9+XL92MzKpU35y8Zxq
Pr66GTU4iApITx2oksL9yuarn57bqVcYGYj505tfFGi7Z7AiT8DQHnSpNZcWsmMw
xut7K5cJxAobsg4dseCUmmO/NdZ8rPAlnDMcccjaeAaw9/eSmvK+jb6Re2jDaJOm
KzOTfB1kzYoKKbBaX62PnFIy1jKLhWd7x9PIaRQexxutDm082WQoyG/Zpysrs+p/
frjN8R+zUwpV+4F3NHGVQL6KLm2qD6Z4158BmAo/CgrJbTjxkn4zzQ3I3W1iOc1z
rProfuSK2MxHipdI/BE5yhCrkdXj4PCsfLAi4RErr2o=
`protect END_PROTECTED
