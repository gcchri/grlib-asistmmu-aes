`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/qBhQcFTS3xTIz4nWB6xNW22ddNrHWaqgTVR/WQuZritR1dJ3/U8zreSHG5+rS63
9eETiERKUlMPFM+0NkWVVM/RprXlYazT8WZ/ZU2v/7x34WnWNsiQtC04Y20TJIdw
IqJ14h6NCYtUIziMpLvv9YChGcULR7fBTxRcTAKY764KqzBK1viRLhEjoOYvcvAT
9/ejv6fcm+OC1zYMj8DojQAL248NWg+A2S1Fr+tq3i/o0aPCkshUtPMIehgeWc4y
LJARQmtkyEZ354oCaWwa3Nob0/AQgfg0rFcpabV5C4VwvKgNZ8691lSd5v3mNxzc
3mOrTeMohMRzWUP7UOgu9J5wcZiONXoh5mgksuuP2eltPQRkWeQ8mw+HjNaXpI1C
Sn+glpow2M582rcJPKtpgIcenD2mVfIy12ZZ62/pzscpc1My7J+OZwgqfMhbpZbQ
oRD+JRmpw9EAHEdKaynBi0nLUpLSX3/r3/6wVP1AlG1NAuQCFHxr8mVqmmHdBcqD
4jZUoq2duXfxw78oDyUt0+e78xYFt4F/2X2OEGteQcEZ0Ee/q6cIV8AEoLWDeOQL
Y5Ty+3ufOeDf56pmBf6BQxn67ODXZR9GDIbVRvo2sp7DdAuSKsX9UNwP2zlLLOqe
XXTjQKgUbtUbwz0lm1FYqTacnf6s1HtOn0u0MOI9Qffubo8aUIx9EY9Ihs6yM8HL
cZzzNnOtdwQ2k4Be8Ub2C+w9YUnrpmQcSDs9fmIj25j79XG8mpxnqJNL73nPCOqj
6W4+mlq/PccmjRLm+4HV62YlXzrpMQcVu7o/XA5R58HUZnxXfwoN+5imPrWBogoh
AnKOxEOKQj9JQEdrVlhYevCXOSMnIaxigeb1EyvXk5QnUaLWiikOJLGGlPCQy4Un
nIGgJ/TmQTMWrH1DzMpTRTcoKXWZldpBuBUGzpd8Y6lfhtASt+8svg4feGd5UFEp
`protect END_PROTECTED
