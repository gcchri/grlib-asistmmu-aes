`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/FDwFInLwQYtqmYJ5rkgTIYhX23YVZrW2xW5Qe1lxyYFvi3CIKBmIaJGpG0627nF
rITkxC3w0gBmYQRobT5gZTB4FIQ5Nr/ktfNkEOimV8/SFSAQuOC9vKSqehQQS3tN
6k9AnayRckOL4IOWGPdQQE+RYtqzOt1ooQPJey7JyOeFKPxgoj6RCM/EgyocdDq0
e17IDKWbFNvegsVaNO9M5BNhyNBsovNzzcp4BVUwT9wf9oq8U9MzU0jy20HmHlEz
Tgert0jr1bzVxtoGrw0HQvajRuXOJSxPqTayVlLS8rTCRxpusyVuT2jAPSaRxRdH
RxyhUodWXEqeZph7dZs2Ng==
`protect END_PROTECTED
