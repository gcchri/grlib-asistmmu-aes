`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ltu2wvFK9lkmboO6UZr5By2FmJ0JAK+ubV9K4M+8zR2lpNQM7Pgj2OKSGDF4xRTM
CbDLhgopfGjN8T29KcrWuLiZjpprifkCAFLoAt+5n0zY5gq1h90RueBLjREuYcRR
CZTGxCClzgyG6zaJTUCw4MFAy7DLtJe6hneGi8mho+ZNHg7bg/aZ6LJ7/PNuip3W
xRTuOuJqft31Y0NMLmxwwDhQRmmbQmljCjHzuLfuiXJ319K50UY78T9ez3pzRFOz
Fxs7wpdRkdFndBQfvDfQCvze2HRKylFKhpISG+0TGR3zao5gvcTZFYTJlXm6pMrB
bfoPV7EDIjKwixT4h5qE8vDlUMuoHWIauvLAeT9THzu2Uvms+0dPX6IlmRpEdPqd
a/dWh0wud0HeMAs26YvT4aa9gws3EFEyp8+/OpbuCBGe9boS1tLA7XalF7nzR4N7
639TMe2sgcZtP4XXLSrs/20ZADT9guUfTtdcki6Tjo1TDxWgbHm5g1euN/dv+xee
6nfPFGlrs030UTKue5xHCqfQtfvTgvrUs0OTp5XwX7mZefhqRh1Ffwg56Gv094L/
`protect END_PROTECTED
