`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oEeNplPQTaV3ugwpA84zsZKCsHwvPUi2w29H9VuspRPEI2mn+d9ihYVf05YMQBEw
V/es2EX4pJa2Y4rm3LLbt4RchZAd4DmezH1LAFoS+jGad+U8VS3iz5mZ/DjcbHXJ
COGOLuTzHxG9TAkPIioL/LJlVORtW4JY9afPb5kEZ5hctbYEfn8oyKp9RlXgCFjJ
WrGzxazen4/Id0v7kLokxS2z8QL/dNtG39DYDAv3tmOj/rNwsRL/W2Fo63GE8XpN
hnznYkxq/TQyFtImv3+1JPexd2fyQ4oQY+85CKJUwNrfmTsg4Hu7qQ/m8w/azK16
U9UeqZR0Er9eJ5HOv1ceQU0VL0Sq6bld46p/YQxnYgWkcGVA9cp8OAoyKmTN8rtp
zlLqj6oglVNAo6Eq5mJ+nLaFQjuRJgZdMOG9H8ybw1RtQU59y4rqfJuw09om6pxr
2Dsa/NBBjawC435il4MCERE4CHEHYiCHJaFs9+QhaZFNFm+KtgyFHJdFnMW5rOf7
q9WBZKISq4r0gbwWx2MqV+92Uvj09v2/5yQX8BYT9/L9CdjJKZSuPw/uORCJtuyi
rR4idubwDoPofTsqGC5bpQCGzY/mkcKTd4PS2TtpGJ43VddtW0Dk9bxIbSF1R2Pd
CVAszDsfFBr2WVnQjyIjK3Pwv9lgPDtppSL79B6c/6+Oiy67jJ9UcUqgW+TIVm1U
J68ChCwyDyWC0GlhgutG5OTpHH4NehoxYZ4H/ToR5Zk=
`protect END_PROTECTED
