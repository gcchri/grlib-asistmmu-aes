`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gbORlCCOXEt0EJ3UrSM9HNjnpDKSuDTiXoqzVTrPZgCpMnu8+KDdWHtjqJnk7NC0
ImbgZd/Fu2oI6P2Sy1N9Pv9b/p3ATw3ZVppCFDNjrYQA/f/puTGSwUFK1uaQDnQw
Q3rKLqmZKrQ0EJUnHOz6+gv48j1kYxkvzbooXZ49jK9FVaIT/tP+XF82qC47U9my
WfxcYBC8BpHC0TBOL4XcWASt4BTi6SXf8QvAn3LsXd1UCQCOAJsO5CFMrWvXw+BZ
yO8pCx5J1POmNQoE/zH7g9Rfam4l+iuT3QV25HNjj7A+/ZQ8oBHLAB8UWwTBTrN3
qTCNHh1EL/ck4Kt93l708pdAktRIaJmM+419OMhgkpsLd3stGUiMxIvgMXUIcZp4
gjCiQFVrXB6zhYOsNE/n1Q==
`protect END_PROTECTED
