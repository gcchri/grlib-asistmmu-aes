`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tfM2bUzxTFEhscoJQuhrInUENYooiztEZpKLANexwG6ZM3/AOkpzjzqIOkcENZ1e
AT/l1dtGBOZ7A/ZCcHOu+T2WI7Iz5iHbl6JFbwJMnb4iBRfQn5eZdtpF3ZIDYCBa
CjHaS9WznJLK48J3vdzABzpRF+7HsH3i9cPGgZEVCopd8RtCSXNMzqhKqm8fEYbv
a/AV56SMYeixtoVJiGC46zVrceZatKHyfEqgTKvqaPmwsqGQUFyeM12VrAGys/V8
JjSyrO2Z2E8GGX2RTIyw7qgiR9CNU8EXbGlzIGkYGSkGkkQYbyAsbuYgMyFT+5qs
2QSk/edUAKplsA3mMgoRfkgcjniCnB8sd8Bc8y00sQIzYQcBEOX5Yt+XZ2P/XaAr
1ypV/2vc/6LzIpKAO+TP5oUnAoDURdtS51l4ZoIAddJgQXwsR/ZW7b+0hW/Xzz5q
qm884GcaAa09ug9J1dcAKDChqO+HwY5R2JykjrwvHs3Ll6csdNcMA/ElfjdVS00H
psXGpSnuKQvSsXubshiyj4g4Ac7Wo4JQj+xpWec+WCCN0qsXDLjiT3ICI2Guz9e0
cDR7LC9dZxiJXia4EuPkXguhgXOEfmrErI1oVBYOSAoKy2t+koltEbAQe2qWfypV
WpXoHKiCw5DKWVhwnB2CjC2xipO2oaNXp9oSbJSg5RPFnLesn01mGD9gqHjb5Lkk
gGAIYAIZdBXQ/NiaEywd/lpCw/sU92nzzyj3MDfi6C6f32RK/NqK2qzMqLKIoGkx
Q7OAGpt7g4/VyT2njObku2N7qrQ8Aw+nPlCOlwV2SjMrXHhiyEb2XRs9oTMTZ9ja
hrhlIP6bx9+Pa9nY1a230rtp/4mFrZsl/6T+6bCuOa9BpHcidOXibxctWTFwj9pa
mWyq6o1AcU7REq0zzR8hy0mf+P13g9ID7WcqtrvsijJ3fvIePUwRZ2ZNQMauSDOf
EQSrdHSDLNCVKgemP5ezqeyxjEaJcPK5w5uPQO3qQ86N6/mDwXqGJw3BP68nuG33
iq7+Ug7Yx/Hi+Gp91GE9hWtRo3W3FlX4hik/tADHHmh7RE2Fu7bRwdqBXiANIanl
odfqEH7csjQ5EpMxyKdQbRERpha03qa8+BozY++K6qAgQxVeySaGvAGW7tGXGlkP
`protect END_PROTECTED
