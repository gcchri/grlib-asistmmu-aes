`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Un3eX8OGynfH+dZd1eyZeuYjAQLkrLtI0v6PrWsv8V+jDqcP4yXFQiWUL3sJtOLO
s17o4Ro0Q/4RhOnImjplqXvVLS4fHMbAu+sbMqmGPqN/Yy7A29S+2U1qmzuX6rLM
P3NVHFhvMgJqS6oO7WvA5TJM8eLMdk7vLaxDLlvi3nVdahhXBeIB3P8gSP9pJ28C
Cl4nnNMtIKdMgHzAefcRKt3Bg1rsmrl+/lOc+HvQzqqF+5N4jKUQq7CjPKaj94JA
ikWx+JltqAeSywXw1DJWfO9be1M6LIsMUBvC/tAbgD+9muoGxIJgsiqT4bzzrqac
exSL135YuMH0dfL7oEOF3GedcaKnXfGjAUi+aNPPWwW4fJ9T75gH9y59ivqpRHhJ
`protect END_PROTECTED
