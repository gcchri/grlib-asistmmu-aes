`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BpMWl0uX/dgoxecUIoHsj1SOBAVvP+X1kup499OUv4iPPtrCrklRHdD+lsWMzClN
+TNz/JRZjN9dAaJipsBUHZ1epEeJfvG81zSoXZRqDSCc5rm45lUNsA4wgsUzL204
mGrhuTT3mHqXIs5YLqfCetHXEfhtYJ+E+H3HkU2+0qh/oM+b7mI2eAJhB/QI16wC
dclksgKsoELga55UgFUrEP5jtisL8FfxhDT4nnybzyiLarT4QAy4vrkmJFBbq7Y9
19kieciqmDh9KcOKswzu9OSeOds6bnw0DZyGg9mri+m1aH0kD1tcLCvanoOt2Uco
qlGAQx5OMbfC9L0c3aBLBdrSLvVM6JgCmSDBWfYs+xdgCJyFEC8grNksiMmf3CWg
UaZ37zXDSxeFdF5wxUOul+M8escMn59JyGIVUwm8hM0FLOzOw3I9hG6MleD2T5yG
Im08mTdVJmO5EUYkSU5Spso5tapUKGslV4uKghMFPhYp2t1fHvqToUIcnESRlJ9E
c32WeiD1wA+1EDSYTWuxc5IAykjMkFZhgNfPlqoVIRMvJKHqevHvI0ziBGB3CMZQ
JJEQgTop3X7U+z54obgB/+M8I1pXZN0SMXCJlBi4EF9mw2hvGa37xItpyU34zF9+
SgfaGYb7gZ4+6e/2K+GmdmN5zBa7r3MKJ/0E48uPms5LiOzyNZL02ogJoKktddGu
Sw4HQ0X1Xdc0FN21BgkxpLyRAuDRABDhzcr16nUFfrvWdaiQ4bVYol2j7bv9kZYf
ex9nwPrl3jm/6t01m+m4123Jm19GRd6NdpQK75yhGqDEyFKIqJDmojuv/m1Rgwh4
dE5sWY+PNyoA8WWzFiEV8CQ0p9WzFfGyYYxO+rRTN8LD5kExyyQ6ReIZPZMuMTO+
5RhWN0j3pMkGjkZwtt2FimFRbAmtfuKFAtWv4VB48a8lfVJz46t6X1llRJpQflRe
kmerI8BBsKIjp6UNlsL1MjM9p1f2q5yqnP8Nt+792oIi0MuyN4bTcKKIkZ0K27dZ
MUijVSDUZx/700RVgANpd6U/aHHJXvvfw6hHbmiuC2fd6fj/RHfjqhR+KNx0bIzB
dlO8LgFEUEm3uJd7oxPY9WCQGclGG6xqEFlzNaP8mIw227TJCGrD8KcQfr6ew4hC
GlBx13O8H6mnt0WqR0TEyRKV2WOcZJNPRGdG792Ecd86J0BhrHqtc0ZgbRs42fiD
RZ6eVHh5p8i/OC27oEiKfhWCC2VXufBCLQXdxs389/wh4+DYFvXDdghnS+6oxdTE
ynC5sz0iTxglasVhTNjn8UdEDQtcesk5vBnzKunFuc6dbC07jihYzG0HqhJ9+Qdi
/y4ZNuMN2vf+f760HThZf5pvAHq3UAMdjlWJVPTkJ3DNzB6t34LnOA85XgUn2hbN
ALdcINDCMuWJnPkX75VgIufzeMB8pBqlviEhFDZnbdQR2iIIgZWyAS31l6O/uF9Y
wnW06/rlLMBJhIZPvN6IDO7KerbHSUqZVwri/MAuNCrb/pivdQbDfnbwSlu5ktD8
N9T04kmq0F6KX2PbDbCP+jyJd4AZDkAemjrLBA5NBA7W8GaqyQSX4XpRhym5Nc6m
KZ91m/hpwjDu2QHoFCspxnQZ/AkjpoUgcPMxpcNEzg3DR6jGwakeJ7daOgtE6u67
l0Xj1CXek2yQnhiU+ZfOf6kvXVn0IAHAMdUtlSeUBrvCT7e6h9naikvpY16ijQ7+
OtgYZaYzLGVMWegD0vLyVw==
`protect END_PROTECTED
