`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W/y3Dok+8UTB3HNki24y4O5dPL8akyW1T2e5QA6CuZcOmiYEtz6fHpg0XNZn+hlA
3/iD6brt7HKYqSXWqb3FJrZWsL7epCizoNLnCDN5zA8tUIL9IPwq/dcrUkhL2g4z
3f9k/hwOmfou/YjQuq7m92k9SraejKnWCe+LcmwxyOVC7Dm8TkYLoMR7eDqanfuc
wIUdRP9IuTnak3cK2maZlTpyyqOSzA8JdlxHwWavf33I5Ls1J+GVzYr4EH1bgR78
JaLqSk5qJfrm0Rt4F0RImcHmAXZ528dESWMrkEHY3ElLSbuFI3mS6fFimLQOzGyF
cx3JHpOaejbx6z7chMylKdnwGEOEFmOBGYww/yl3HJiGZba4VRo+k5z9HxCyE8oN
cBjMKNkKMQaFN7Vl/F2VBUnXlx4LXycq/msPQjx90PeAfB6UhNDijcZA/J2W15YW
3ldINCvv9Ho9odA0klun6621T0b9zLjZ33xIIS+bkjRsC4pKA9AiwHGBmI6YAtpe
oMJYGXopaTd3p/Q5Ce4ChfUU/wDZ77tjf7E26raupGtblLtjrcwJEnCUqlT+HQxS
jIg8KuFQzftOoV2IvhLRCB8SV4FN8WkEJ4MYl5s1fBu2QIZryrYqL6UQTJgJ1tXB
6iw5IxsTZe7TAzuJeDlkd2ax9Me5Uxu3hADtCWdA0is6jMFkGt6DJWdMyzEVhZyi
IjP7XdmXb0XzrRtvLRu80vHus5tq8z9N4VnoweuU8xNuU32DCFE6wJ5Ju5Bvho/f
DHssJuTWDOMLWhU7VaIi3wxQLYvPc/v/5RkRAjdumYRCvNWAaOTwdMsGj3W5+Vq3
IqYeX1hcW/j8xNVskPQg9dFIsr1U9IqIRqM3lwGCLojV4Mycjfq3W8fS/ZLS/LX4
c14QyFHLCae80BPjbx6Nsh2+jjbgGXWikAj35I/aUh95da0mglMA3uQ2B2sudQl0
xKi1fXOmsoni7s4YhFm4lDw4f9QCnYrnfl2Hl8o8pYQcwc+iMOzxhULr4Ngw2pYX
9CIwUY3YfEiCQtKuQ5kAUfM8FhXU2prd4VzXYQjFOYgC0T/QcOqqpA43rwlVdWi8
tpAto4UilGIZnFbEvW0m2kBnOthL24d0asMCsp6YSJylZ+O/faGRl4qpEL3zkMyW
zpgWXE6cadADvFJma0a4a0m5yCLltvP7z1PeeMGmPdi54eP/nk0aL3iv6y+huIRB
ufQMpoqPs06rwbi5uJahfASDHtha8FDo+mu71MvUxziNf+rav6ChiXKwMVLBm4f2
S4id17IHaee23ur084GQWI6yKw2xd0u54eEc/YZRO0i5JSP7vEeevQmHRc1XElod
Int7wpdhUsAtKbAFje5GsO/L4g2YrXFuObg56q0P8G89Ak0OYSY3Y7AdgqyBUObG
FAFe8NREqtkS7tFXaCufPUbKEDNVphxoX846EfuLoBjThFAz0JDW+cy6SkeViJGF
xondyTlrgiOybQ0yZAl2my8RYncBItMO8SG5fgaljy/PplmPA0qWp87NgMp7umcr
+Uij2hOLfJUx1zVsIREuIVuhc5G1zZBiZpTh9jP5/geLLCTXHnwf0jrcCooDYcf3
ai9LniBvAkdE/cfa7qCNmgqamYLVzI3ajcZz21cypyr0Rzshsri8GAe4uz8C25e0
0I4nUBP1jg6qtZGx3WD9LesxH2TxqFSvj5NDVitwOvt5Bxns+8WxY75sFijN3B1h
VGPRrLXunoNqlrOHYE+dCFRUknZGZ/wwXeK2BprmW6kcU8SL7sLz88JxSuYQTjwE
MIG1p1UFp0pbKkv33jQz11ZLgVolHL1LDsBuhpwym45lHL6jOP0fzolKHb0NMj7z
UDpuc1ra+/pmw36wTMHq3bAwZoI5JF1vJnFVvuBwCL4hnxP7npJO0lJgw+YcHiu3
qaDclbEwRd3pHX94WgE5dPnAOQXwBFGm1B6bFZ2rdzjwJiZIFr6tT8KMwbJMfw5w
QGu3MtTG1qj/KL5MwQuzDKvGk1Rd2Mtg3cvc9ZJB4SjtR1AMaG+lf920XnGhpwib
8Xmzi8NvZtReRzAZ6e8cUfcg5mYdPO3wS4L7PGpsL/SgSJZpDr5bhv8+HUBpNKz/
tBubbsrff8RJNM2WhR84G96ss/6V5Q8YRh8eu8aQ+GXDpv0sX5w9XfbU18WWi8hM
E7WabmpENL/gV+AGbL2h3y22SEWtUluuQUOIM6TVHPWa87TYQ/o/vp9zEVGJ+t5z
5MlqYKcspeIKCYlvCuja0AzIw8KxKNxiusgTwu5XkmH4PVoO72Z29Ctc9OyHc8w0
IjYP+bQeY3wlxh8fPVpBPw==
`protect END_PROTECTED
