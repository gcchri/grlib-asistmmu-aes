`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wj9C/wvPHQNxlX1dZScv0xHs4vj4hOtAq5A8anfYxSWxrXLc0xxScWuSFwubli4J
a49fZ5GJ4xou/abnrRLUv3K6o1DvE6Y/RG8i9wa8/JgCTCIw2FHA3TmaEWY2PP8w
EELsQHe9KUL5N+KR0hWsoGI2pFtE0V5dD9o1pM/erXPFqOhM8KxWVrGS4KjgQS89
tBC9iX6S7bF7qxImDusQsf6xfMlfUcuOKM6yIWLTAEbj5cTc5pxAQ52oRETM6tx0
IkRR7j9eK/8mWwDkt7VmpNX1Obs51hRbrhCW+jr8XDYpsMH4zkxT752tmLq7lxwe
jki8ghP9qOs6Tsu12H1ojUgyrZwqU3wKIri2EHhfrU+yw8G/qhfRDwfwYPmxS2X2
3SvJ/a73X+cYE4lv9mpELDMS4USD7i2/PCtdLrerIjmPUJJaYvhMBjBr7CzUIDwY
m+S2hz3gMIRoUaHQZ8VecDOpBk93u2JF9CaykWdjUANcpxh/MFDB6WyWdftfaAO7
Hr+U9P50s6Y2MPV7skgSoQJ0mBdwpS59KD/rty7zD26cS520C0sWRBzN/ElX6/4l
VVygU+JGXFSdeiOPVsqQYIlxkXuo6B6ptHnuGgDtAIG9ilcIE/jn2zFAv5r56W02
HEDVjvPdjiEhMpw4zMceV0zUWs4dI8SRUFrTg2JJ6UaT6zNC27aaashlpDiTH/kz
+BNQMu5vAi0VfrBQ8Ss6BWT/uYAbn33s48wQUW5Jh7avMplQg6W0UVsJ2kDHGcIi
4XeXhGVqfM60OVN1BY15gIsCML5jIJnO8jSoDpBt+/y1FqHltuf2fTh7tSNTnMEW
cGgxUZcDQ5dDt/I71Q2+7R0/DlfZqfMeozAzS24B05HNQpHr/o1ypnhgEnvVta9F
HELucG/8JxJqjpUkmaZHijIbzCPwIcQtTWos0tDMwRLGDXXTDNg6xY6BobPZDOpV
8BLwVHyC09sTyn8iefiG71fa0JRxJbG+bBJUfSbLfG0O9MH9QYi+2ELB6eVRG6in
yhaUkNHjvjQ2J2v7pfMrMY8BKhTnSZhvwiC4ZyimzpQQW9HBlQauPjMa46Hs+qc4
mM1rYpjGPQVOZYyNHNzrVnpyqWL/Bs3X8MSOw4Wd4Px86Vi3bmEGI6MHe2OBks0C
BUBMy8fXRYThyDX17S0cxddZsZXafIbw1T0bXeHkZ4ICuKfvHk1rYEc7hTpxT0rP
AwOyvMFDdw5a6Fw9svma6bjIGF0Im2CazyVMgh5E3lya9kZV65lJj9FgVZfbm/IQ
l5lq7qYyUThPBVe+pD6CmciGe0GNMpFqlgpIo/LcnY3ipjhGBj1ieFqIo+/Pl4mT
fB3Gu+608IzXSQTUeveRqNMIQJtXFDUCpXKZov3p3bm0Jnji7sG03ZhPTug1KNQk
RLa28yV0W1WvR/MbmBzUfS3hg2kCj8Wf+fKbBaXjG2LwRU6ePb6x6evPufH/blM+
QHUwJz1fawMOnKeHBuq4iCzgcAWGOZeksytwOCYrn8hP/RFF1K8HtAEARmXi+bz6
mOUwOLuMo/eK3PSlHafkv9eDy6MrifoPW+0osSh+nfTkbvHUW3B42hJ6DtYy/L8L
+M6rZK4Y1Z51uQw3K7m5pLRoHAs7k5Z/JT92GAS4QKbcC6+Qdna7q/E6jQum/zPl
EuncjQpoBk8KY6Arka+a52LG6NrqtIF66cdCzXTd0a35ou57exwjSe9SIkCBkxRs
ZkQKS6IIdM2BI6zEQIr1Wm+jns6WF1ZZAcOzQ7Dm8jghEGFZrXPM8xznoI8QVhXZ
KwFAXsnH0hB3F8fBdO8APbWy480s65IDWcJcIovDHUCcQUAbmtSxCMDRc4ct8HWp
9Q3tqG8yZnFFhFIdm1OKhc9dDJkdRJtN7B3WO09Dwd3SyG8bEaawEvK4L7NH5q7s
dKd27ilMwEJO5IhujzyZssPiqncIyxEudzmHc1iJBuJfVNiuHR51KkQm9LkZDYXx
N9PBIjdFbDVzkIG2/5jppVEx9YGKxYU+S1rSes2UEGupEOOtvHwfdNxmfRH/GdCF
HKep4LMOzUwP665Yo3605z0zayQOBFXYqIZcoYRqX87GuZqPjBJ6rC2BK0xSJA17
2odgRfX2v1FjxdUOOIuatL3zS7chPhnr68zsCydNde2t0SBazWQm9r0bDFsqB5yq
hQrvZzT4WmZnVQJMCLopRHag3OwcUFeoFDtWN79xMWYRm0/DzDgb99AUxSAMUDhX
MiaerwcVcPrMZx8nQlZKFPJMES9vnflg+scH4WqjrpcVTkD+I6egTH4So6mfx1En
zioOtEMMLTpUxgBylRdS8IEduhxHgKPAUoLse0zJTcCytZboeLg4F3V9b8fPLnCd
Em2BQQGRCvOMIEq/35oOd6jzzllpKkCQRamzp4BcZtzSCi1HoOiMg/kgKFjAWsy4
ezzaeW7PJOFAsIFr7DBieABnEBq0fZhbJ2jQcMeN2W73i2F6h+giNzSdi9xBX1E5
q1xBNChiqpgvubazSUJ4eTJcG1EZn1ErWExr+R0w74C7IAIP0HfUCAdxe+ECvM9a
sPZOxp6/mw6oRPiNpdCpwJoOqEri0Kt6jSdzuafLD3bO6wRrfmIL2WHUfORGE6S5
xnxF4gWEWQXnXp+N2iGXOcu3H2YVXc7yko3m3LgHDh6+x9YdGt5Ep+0gN9vYuHW3
oxCiVT/i9au+wYBI8RQkCLOYzJV1w0EXzKqnomTqJMRxSKTFYsyEwXKH2c0ptKup
tAMVK3kBil2gdVlZ2CU222yNHJySA33Ko7UZ7z5stUsfQiOZdlFcbwHes3VXXbOw
drcZOtRdhgVbWUPRGaUwL7qTeCnhu2zTNqlsEPdltzdxWzQq8BAMJ07i8H9lUe4/
o/HLCbSHdi5p62U/mzogb/ZRmL/HGiWRtU2wEOO1ijiyqZhbytiZqu81sZVkFSeK
TcJWR9Pwoc+DBKHa4ccgzij6TYgfzC0J5jyuNJdreHnDARCuCaMFTHB4x95FZwKH
nodMpbWNnyrB6n2ReOobI9BZEZMeqq6cGVXBRyRUe0LpWVq1spbCxA8xSRRcJBE/
NkQJhdhmWMuDmH0QqoBK3Fr4Y4qEgfN+7b8MWJ7tCB3MlJs4bdqXaLtkUIA16oI+
bN5uRLx5UsP1F/HzPkyVpmHUwwN5VXOUfRArxkD2T21xhm8L3VVASdugCenE9kq5
Rscah/NR4s4qtCNi/MfO6fds57slioVpS7YOlZD1xOHJK84Ln8+j3OibMDCcmQ8c
X0hr7hCY9JeE0LVFWTYC7bzQxlGc61bQeBORuDyLHnY9e/UaEWjtHngFjZUXRozd
FU/Tb0Jti9G5BQZHd70/dA8RVHtCVG/U0pc7FPB9hi/huVv8v4x+l4HD3gbjglcF
M6TU5B/f56Gr3C8F9n3dwYThWcqMdCDuYJCegu+0D4GiUcLHVpLNzuBFe1l7h+Mj
Va7WlwIuVtdrY0RxI67T969KDa+DX/BJyTtWnzvWTN8=
`protect END_PROTECTED
