`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g+hYAkzUkhZi35kLOorHSBm1hItXqzd3Nb2qQ4cfVUOi9PXUXrmFn2rnsggtdGFZ
XWvNA/Rw1W4tOBEgizmspsmpXvUcsuavlWGAPxjKfoaePWxI4L4ChcVSkWB4ZczC
nZ8dEEhwWUH+cSt6Y/F5JqU4TFOJtYtvAeh3eZMWYJzBhf7sgDkby2su8IKxF3Zy
ZI8A5lLTPP0el+lrQ4sYglLA+utur1cuCJKIQMlJh1V3zUAj2OGIhUUcGtvUrZAC
yeXVhiwRODSxOcbChuugPR3tk5a+U+qMP4Iz+w258eGthaASVLXoJ9gGF55wuxa7
NKf3EWTi0lbL77IPtKxvZw==
`protect END_PROTECTED
