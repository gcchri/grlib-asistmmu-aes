`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v4k8nafyPeMiVcDuEHcLmk17iVoaoeNBwFO2eymtwSR4M2emdZdrtgyBZUaqe/3T
AH2riGHzvu1RgsQohQZJvvWFFGzmCiinL8PZMHG5lZS3z1hocgOCTb7zkYZjYTok
HfwvJdS2F7DqSUPyb4kEd1NyD941FRNh2RCP6o7tY7Ch52R7XzIOvmvOM0S3fbUO
AMko0MxRSd5X8Zhx2gs/Pef/k+slediBP94BKhydBFdlqLgyvx3QPc0aX7YRyLoh
2mmJWqs7d+jYvoBMfpMTbwPVXkCdfIwNaL0PNBEQKcUHsZAsa1IM7gRJxUnqcQyg
Sp/+9fGu1AVnU19/JuTOYCssAANguzxvf3T8F0iflomj6Wd0vHT4VP67H5cbPvCh
jnwD4Z2MmyFgps5+MAMHqnW5ybGhSx6jo+n6ueNl+f0GCEZzPme6fUJBn/vnzOlM
IcZbh74uH9YFLHTPcSEumW7OX2aRsDM3yV3msx2//VWcQBgBLV4vu1kO1Orfosrw
WWk0TShWoN1E4PRdzgELAbzA/WbxzRZnRGuupl2YgHhKO+CVPDb7utQYRiQKiQ5z
6NSQmMCFiq+957JeZj2DcMmoLakSqVJC8o/kWgEnOdOr+lm9ExmMsvEsgdcCRRZW
47rcztL5eMX7UWyr94G+c+wp1OPj4RcciyCp6HgRjswXl982EcDvfll+FnSOJNWv
ayduzyKdk8ziZqXR05XRKjlvzuqEFjuUBr2k0FFLOXk214c6/G98blWp1J6liGMt
KwrV/HYmJvp7LB8jMHGBsDjeP5YsqgA1/VzXWSck0SOb7PylvoWqr7UyqBKKtAR9
Zp/T79KMPOUFc+3cu4V/txQcgenzSVEO9AG+wDGJATNs12vlRAEMouFtL/TXCW7H
fW/856PyVfHE/FyHIlbLFMoqt6dp4m/UjtOwLc3e/1ENLy8ZluJV9ZOgR0QcDo8G
R9AFU945eehlbg16FZygxIXMkT8Py3z+WQYyBEK08aheBdgEM9bpPMyvAmBY3jRz
urIakiUaQzbp8uS2sNUYJrH72wp99Wx9YeK4JfE8DBrCsF1e9pN54KsPc7FImDkK
01uzP0KJEcPwNe8wVx9EEIyATy+7A3GIYWpu1Q4d/XfNasY+xA9q58jTa9KwMGk/
q8wSiRVMipdMqhtXmD8Ow60Ua9tZ/0AcXp0vngRqDnVl2Rhdk6INTj6SMAdjbz/8
JIsEGjUmULJhdQTHfMpm7cXhvMYZB9VX9iaU8amKtWAMYxHTu5ZRW8V/nUFVUwGH
v7jOFIFTqlM3Gyf/bk9OvUeVlkeGI5g4Mo0q0Qtpr1UD77Dv8NVBoabM+Khi1HLn
2luE6LU48iqyYvX3p2LUWDxyOExPR+eENBdEvzqIk/fz9iuE1LajmjjEZPoy2tBp
Bj9tjQNyRZWpcDmbPvllQYBicdojlfQ3d458aK1+sk/adx3YfwTqORYDxRjlSX40
DcFm/tVUsXP10OE7qx1kUx4Wvzm9RQZ6uFK3IZhA8QbcTNF5XKyJy1ApHzMjaE8/
tzRUTwWOL7SkuxQTziLNA9UMfYhf3KXiru8tCzoU3zviP1nlBJLaGjNMuqShJ96v
j9Rd0emeXvQYIuDWIkyJA1vPuzM2Is6VXu3jNvzzyANnJvLp8mbK9Jdozsoql1mn
9xgFOZZgpquBX1LjahvZunFxy1yqkLJ0RdiToQ76xCaBtPU18nDNTkzTTGwoN6J4
Mkp0geTbw/5VPUYMmODSkuD8Rn3Fd6gdhk9kn2kJcFIWV0nrJ5p/aFbzg4wXsOel
AM6u5JPJIN1Pfdc35fkQJvmAUmiVpWn8/v0JKhb9sCSHfFQlP96WyuzuH/PwsmFs
adeRT02XD+bsZz4YXlnSuwBFxTrG9Vp2OKBYF/7YS9UvMcd9pUV84/hZ+q0Us9ER
Qpe1Edf4k6/5Waf1Ydf7E+Hofye4J8BWOhSNEpU68+zPAOfa6UiRgH9xwxuWHezk
UQb/PCwiakErZMQeWcNnAuODGNQLFDP/Wzl+ibJ106Ly6yHxh6jsx4PN0AOLr531
3LgsoQu2/x0sE4pbnZuz4IGhxwMpohKMh+qCSPJPq/oES1qO/ZGrjiNCVyIvGtvh
t0HbsKcHq+Tj39LqREifml2v/dPrqsEw028NLri2y4Uxjo4JZYVHLfJQ5531CH/X
0VAVIAi0ro3ut5bbCKs8hvKmCUs0E8A6HHezySnRwS/vGm6UZV/lY1lVpZghzAlL
Wo84BobZ/gficglrHwDAVAk2tZ3mxbAvOPfJdmYR6T893N7Ne7Kyc6A1WjuSXytp
y1KaBI73HiNiVJQvL1tRD2kDQrB5e9vB8fwj8Z07e+LT178n0ezthm6/Ecbjk842
rHWCHt9a2QD1zQlZxD+UH5O/KCrQhM0rAlh2yWX58b2Nk86kv5hs46e7fJXv5TFP
g6nEc98o64FqpV7C6LQ4d76Wb46MlxjimBfiqX8mdrvoO03QI0wu3BYHTe1/USc2
hsPabpFywqEqn1j3X2tLukxhAAwClKaVT+tcM5NzrCXyZhjS/oKq5354gecYQqpj
Kl6dYmD6sB0iFCbJ91pxFwiXEYwihqtjEoJQHyqCK4KOeB2NcfcCd7YASKEjUjkK
PRKIwb3ommZ7HECUFgpLkjL8dXZ3kxdSgD+QjFo41zbFltUfGP4a/ybRNKDUfXl9
7S0kqPaNxnjGBnp24mcVJ+3xauFSALTLSnH+HFE84DXfd2D+BXzrvMWrZx+1nn8c
Etl2GvjBpco2qJsFNdf6GT0HFO/PxeGZW9hOts/GxEQ/dAJtnUV0Q36+1u0SGImO
TdhAmEytI+sYISC7peLz8txFRzZrusFAiMAO5/VMOUE4Cs23The6vEKcBI7lg81Q
5yFe9n2DdH3Qh32KYFs2zMieeCqKZ74WCU53Prfi+9Y3IIoXXQQdPeEX33FuVgbj
9HBXUvFE6QQ656jfdUoojFvbYbp4olmcrPZwINvH/PcEFtCR33ZWb5lPLAoMT7R9
YNu9yqvUs3SaGFJ0Vm9IfEsarRo0AQQwuBLwKPKN1XOyqfQgkt9F/GOOl8wxX9kn
IXqv2GbuwkkHLWk1AUzCfFkfcJGZn7+g6ByQVjQl0Y8MBvxILF1K/1ovb31xB+HP
C7WBBwr+w8p4MCeHNPQuyqcMJOnMbeUzGL3LIjLyFqNSm4dv8M7L1HFq7MJtCMBP
UrQPPDkpGAiUZWaZ/NjBoOj+Mq31u0wauMCBc84Ql9TPNvsyq84h4vdHxphxksET
SMV3QNXC3joq5afcBZpnKAFqSTcAEqIWFdkshx0oE9IOXnRByIxQ82MfU3XaRx/J
Y4DVOXM2EiT6yGsSFA2foT++Efer0rCfXC3NSqXYtvLX5Nz5c/0dyJv5bU8fJN/l
Nc8kUMiXQpnni47KkFVOnS7TQE6OvW/3o9DRiWJvB1FARnAlwqb9Lvt6JTOX6W9c
pwxMHJLmJEaHYSS8aTw6gU1sRC8TgvZEKmd7lzKwwVDdafNgrXLWERlPaGxAgFWu
LrRrAT4e1T7ePDzPUVO/TA/GbZ3G9TgA+4kP2TdvF2O43NH1J/pJyv+9cUUBe+3n
2y8waqrSIMfwTsF+YkwRopXmAK8EaW59mLty35dFMQVUTxx5M8pwpZXKrQKLHFvj
q/ocmpmJ4EzoOXmVDbTiCuoyuNATrhnUSE/DVLLt/zjh03svxjnFtM/QMojvDEwe
LBQY8iKhaKYBRRuurMYAxvWHPWrR9D9ijS59FSzUDaWl4iDt4QIBQv+mDftPl912
J+01T8XASiw5KekbMJQEBG3t0lc9OuPwj3M0UsdEv2eSUgTizpdfrzNeSF+qHo9z
IQtX/b491od4/6kDnGTj5Ho/DlJH4MRQY1jJBlioes9YuJUQDAltmTru4bIoCbLY
zA7SrpdWs3GQ+FpmsfoK+0//M4Z8/dwhPJp+1CuFH5gBqfb1ePjgz+3He6hPnd6t
/uFoS7ZhWFBDCu2UenvKk28vdGMjIp1sOGUA0NExtGK3WknR9NMnext+8/91/eBY
aBaZh2KniKAY7e2f9q3gvru0tx50qtBUMvglGtxWsZLwya7L5XfpOMOLHOoSBz5/
bqQh8TLHZGeEsTyVDpU2mMVBkqDYq/9HGRJaAJ/KSU4tpDC+e5A7cwJOGtP085+w
6POBsWwG2qfBhV1U/Lb9ezulR5xkZF1TX5O/DUTvrI98Ev7EtTkHZkIV7S1J4Jip
NwTWFmg5evVUT6kbX59YHIeVznSrNpArnwttM+brB9R5D0fcZ+txt+RlYeON9P2k
dAV1fyLCkedxLMTXuNfC6QoK3b3AMj2HSMsFO5qplv5qtrKlTMNnVwTHBkbVo072
euqe6BQnRQEprgtu6/r6GPd7OiPmLZynu8Jv3JHiw+MAPb7uUAPJDeudj6rsDvB7
nFzSgmUkuJ3BddTFBqpynDgb0TThUfH2FahpO7KbOT/uWyPxQXBgXNL9HCAc7jQ/
kitjZsMxbawFJs5Whj7hwpSFuCaR7qg1xv4btaLyp1mCWR5CE3espNZGQzhxgnQS
cix6Fm5BIAAF0HIrRAudO/D47asseZFwi/7VN9aZkuPd5EbmKXFcGjavhOfR1eow
rkKXKnVOwURKnkRV+fLxKm6sieqaR1PgfemmtuqEiEhxl4USj+9t9pL5qlrKePYA
PC81WnBWZuJSSQzcivCQp8O/vyU0ghyjoNQe974mZNE9KGQJEiC++f00X6fjn+06
HRaBYvDV4MxmhvKyqK/Un/TfOpLFznTVpTBzyh0kXVUO/zcKrt9+sfCFw3dWHCxs
yFkRBNxttcahKpiDG5Y5+ioSmKwOKinekY+OsSOJVJctt8OzawCjE9wBBrzdkGvb
XUHC6dSPlwfGeib7teBwOHyzencLF/pwD/vtCZJ8WqhXnUH/ii6ISjQFaj4DJo9w
pe2/N3n2aH7yb5VY9g58DYiHj65tUQlaoM2QN8SzYoLY2acRGAAdpw4hfvWbBPmv
VoSccNe0OP/jTMolfVgwXZnn34+Wxs4pguGJMa2Ibfui3R1iSDaBWAojfeBdHMp1
nVvgWD/RICmVT0kIeYKOMEfFXEWbRFZwwOcCU4iPf0Se8V3CRePfSdxucm9NdaVl
M644ceMOuOpKxtyQ5TuYl7w7loThy5RegewKPLWjRY4gKKZxUC4HZi3wL6ZinHve
mqTYwcqv7m2DY37eDk39/6SlCRNbaHEVm7wgCMtFP/5PHl2aQp03F2yi0SDdjBpW
mPIB+vE0ypiMZANW72jXpVeH9xpftpM1Pew/cuHhOeNkJSJoRAyEx7CzAB/i0PPx
z9zaZqyO+gV4d7y/mG43KlaOwsxI0NmdMCGwJCeZvkd4TO/4H1Dzw3bQ2YbUhQuI
sn5cPBF40SlUrP1TRZ6dnhvf2GUFjyvRPeYRg50LD7Qr8TOryaIryQNyzU+i6ASH
9W3UtrzXamYq0tBz7WvblNfv+tORM5RkMZkPqUyOVNGRW+ksiuINA53e1KknRXXs
T4FyAMXHQGVMMdoI7gxMIJlleH2nUk/cNzDnEN09ZHFAZhAOtLusmZy0mEJcl1LS
uVjs+eRK3EIVRpC8RKpZEKg1d0Z92szcN/a4W3GqJuyJxxkStVvDUq2yx8rfB7H6
PAhKAHe7v2Em0j0xpbyR49CLXEf7S6ndh7d4wDYoULfg914AXGELfJHWcgOwdXSX
EW3mBxOf+y61FtWhUKJNwnGXSwD49PrHk+0/zt6y1cOrVABN3hKFe8wRTd7bNMp7
RHnXBmVKQi1DHocn6KmurXumMgRKHbYgoOV60CJJWBsYSI3nQr4RwWsxBoyrG5Mg
WflAvmhaIvMVULghyl/LzF6hBIuUQjmrxNDUezRsx1RBPBL7F67cbQvblGlHgfxc
ueZ16ZEGDwF2j1NEcIy00Xvl6Afl01dzDxyE5RpdAbk8bNe+vvbXS6dDTDNYK/cy
sBf/oBNUl29fQkeajzsN42MNhoEea3lnuh5evcfMxAsssN03/+HgvBknSp8r0xTE
WB42vNA/+/y7xUiAIKe/UfCRdlvP2YZB9Ufq2jxmM+XXGjhZEXsMXl4AFKyfxSSk
qd0PJA+rvR+RhrpFB6hHqVzn6CUhZ8Y/V0sDHaKZepFrXSiDVLiFUv5N3WrYxiir
ztv5JvDSe0T1ia47FIXyOjoLvKs+3/ic+0D5NISFGDV8rzf7RFB7MzSzC6336HjV
RBxANwL8Nv1eCpPua4JzqtTXxROPMVpOZ78MXtAfHWe0JAl8e1QxVj8pKidkzt2t
DyvUYi11g1CNkZFFjWKcy0BgzN3JzhEg6dmWk0QdoXgjao/n7eciJapvtlPqC83p
5eZwoEAvFFkYTwRX8KMNKc/rzQEzgFBnaLZg81ncd9YVPSSV4vJayZSm9uqH+A1U
wy7RKZPWoSOxCVQC/kD9SGF0MC+cTYqpa9b1HpOHIhZpafDxKQLWC5+JQRbU5HvB
Gp1yqXQVGMJgiRz70FwlzX2JCSw4AxbAnqsEYTS283VXbLzl6M/OrO9WtkqwmenG
hsbjs8WbpCGcZcL/oSGwaXiIhy0GZJVsxScI4zicdoQ+YABVKGkPDu7Ve86p9N3l
lULeKcf8x/or4t4c0rgBWwj5QzeB/0AtAwWdUx48GNgNd+jZgN0nWbxESfbjAAms
x+6ydLGDn6vfIDv/6hE2Oug8K42Q7IVhmW9cKfh43NlOR+nO0BKVkna5atINOmdB
NTTRTy7aMgYSkl7Z+1fWVVQNgaHYhfo220+oQryLEpLrNIEMBQsxFOOxdMAsOzFu
Lf/V2TAGIup+HnS1R0x2wk6MckKfqDkeXlpSW6HhivhOc3IOFs2MPyc7cS7QpGqJ
axkjPEBke9vkbNlX/4JBO+ljc8guQZDDSUTSAxI6ux0XhNqcdaD/mFtEMm+YSO/F
2ZYVA9IZ/UkFswnW7xuc2R1OQsWlw9zVlpBu8Xtp7KWyjp0vqDrODDvFw8V79o5y
XLCQgaxW/q8cNLTkUMl/5i8idOjYv76czVTdWYONOacZS7/OAHajJ21uJ0whWcO7
zSz3QEv1L/RMN4eEwJWdFfHrdr0D81EvmDG3YO1DFhTy0m264T+jm0dtwV/H48ei
kSb7BPsjzKNhREjYtiytQe2Q6rQKB9YYPe7xlYlWqbxCrhlPGwWN+qMo9a3qQjij
jW4CRV8VFX00jCqpVAIstiXHUCPxiUwlT1nrD1YYWj6VdE4qyB0CNp00ZZQ495w8
yVeByf4pUj7yAli56gNTtXxK3RO33ETVH6/BwE4CmdB9ub0Ca4GMN40gSYbMA6j9
2wksA5YIhWKBpoMX/JJo1aHlUbgBWX8zOwlFdFU7Oc98BBOtceJCaw3YqiLQLmLX
1PPywuPsRnHexriQREfbx31ICqzhsf+R2GNtzUvNzgRqEJ/dSclD7q1SDAf0QByq
qsi39/1iVOTcSRDo7DVIFLpyijCfp/9h0bwshF7Ue84WgeT17706E4XCDMQ+lpKF
jJXuTr6CDCBql0g3Z9COXafEoWpfAU2RTTBmkvNjWVb3ikH3ds7z+uix19apIsIc
0Td90E44luUYpqq1v+k+V+mOH6uYgyVIsJJ7Ywvxdls9TBTn3wV6DcNma+jR1Gai
2I5oLl8qSbL1Fcv2SUz67bO+ikAoLwPFPI5EVdp6682MWobBPZoah9yzWy2Z46l2
bUGpMl1nfcMJadILB574llHId92qnz8wfuwpjiHL/AzwMf30Wvdeo5peEp3CE3xp
tfa3cvz7Ye83vmEeYCZxYW0PgWIULpbTIsY1M75to5uy2PCtf4HTiNEz8ikAEH8P
8Sm2zm/T3noQgKZfBkhiBhYW1B5zSFpX/9NbKtPt+3jEQxnXIHFHK9p+s2iu6A6E
9BSnR4jbEf2QDWTB8tXtNPSCFv/NUNh146trO8l/qCL5pmVI2zWZ/GGO+Sr0kB4A
RSMbyRgAjA+RNnWJ3t1xD/C1agurnVTcpIU70MBztZ6BwEGgtcd6QcdXXzosB3Xr
SwFVN1q16oDOj9vvzu9fQhYoaVlXlJ34xDL3adaZ+9YYLEkuvyE/USaDa6SNAJwY
9LEagGv7HbUw0t5MNEyQBSIS6tG3ohYyJTSwkEJOxCKOBQDX+9Fft6DrCsp857B7
5/XuNy3iXGuoxyyse767ODm6kfPhZd+f7dRAHD5REzhE9EhbNsx8DmU/00w0CGKl
eUTQCJDsh5JnNMAqQrqt6iFQariTcCTQvWymtWR53TW1gqv5prPqz1+AQUVLb7kx
iO4dbOBxyqvaZrqyJ69+zneeHCmDfSWio7lUw75Q6WmIR3edehJ3rbd7k5o6ZhLH
M+ZNEptCkftBVjVmpx2mXmGW60RnLUHrCuB4lloeboM4Hx0ELP+bqFS7nc4TzlsI
7XQvrgiNr5/83Z9wfegrqWIzzokNe9DDTOTbnDLOlYtSnSUFxqlq+X/TJyFX6Zoo
dUKE3tMjvBvE5m446m9icmbU7WvnCpc76ooJA7cdZ0HokTepe7O55UTMFWXU8mc1
mskzLGLs8m8bEiWnZiYZe3QSp2bzGU0ehUe20L18Dhll9V9cmBpWOB9M8tRTHRKQ
wKWlFcL94dxLWwk+ugCcBzY/gHfey/+v4F7+A9LdBCM3jrgYcYUmFSBUGHgBQkgs
uInk2Go2w3QepVMes2XlCMPN7n9/QeoSP2pbQEvJ13HK0HvAg8od6H8YaBIwU+wi
aqVBUcAmVjQbObUTgEhpUy1CW3w3Ouw9DMUFYRUDpO18uMWX9jjDEwcM6taZb/gq
ZZElyKmqE6/o5gWeICYxt67Sf5+ZoWvo4VNfdOEjAHNvMWgpX7AuHUArh/CPOQva
6d0d9XCDGpbmCTMeKTQVvO8R2+Xr685mkOwBoeC6LeaQ//BGUdqQkWyOmiftzvvn
DtXWx0Vx36EE3eNcrYfnG0Mq/66OlIhBHxrq+zzbxe7DTczFHjUIxjBHadj8ZXyq
+u36oEDaZjb1uxF/auaxFO2uk0d0dYMBfLkglQ2ijDFvmAlhiHmwEQFWyrRYMYEF
/lfW8kO3NSwZv3rD4VcE5vQ747dbhxsdj39TkL9VRf1UUd1zEmRdNtHHh02dqEwu
wCaNb6skBDtdc+6Cy0Bg2DTzPJWhJmKHuXFjRkyKcEs6w1DN/XA2C2ihUB4msRBN
Z8gf8yL+Gzy/P5OzJfH2qf3siYiekvneuNFYo/qvf5a7iZ5jO2r4BkFCAAHGJY39
LCzg3p48i6umcyyyJgr/7sbyrJwuWEwEt8n6r6q5ZXWJO96IEm+saW2shA8bPJ5k
sQXtEnZEc7RjOm/oQ4WTAru6DDxeJRTTUu8fyFVHGDQWqEwDk7WLsy6jl+DUMdSB
R6E3QjHhiuGWblV/oyvS+eFnhhfV2QEhfnw/Y7cB6Qs=
`protect END_PROTECTED
