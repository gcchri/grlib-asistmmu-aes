`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ymNuIhu76kTmvVDzTiqyVxq1nbZTzX8mZpSB2yihi7CI8HsHPFCOY3LwZh2fETMs
dPeI+btcfEr7oTlbgc6LG+ryNqwo8m78Cbeej4nophx+vw1XCyvU2pWiNq2NPYZa
9QT5slRBMvmmVE49LaNsTYmqXJeHvGl+04krWZYafhh5SebOTvyGLvSUqatQ3V95
04KnXZu5pXVZfh0eRu2ibuEZWPzeNF94A0bNfc9ZdOZ+Oukhrc1vR2zYJKATKvb5
9SDsbaUcCb8kuXPtUnB58pgZLXJHseATvAKiT3jVzPY=
`protect END_PROTECTED
