`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z6fErBJ0bKqRFPW2DfzerHAF5v1hRfPGg7EN9DBFI7yT/GJYtkPAwUx89l0KQtu+
DCUgQXUdvzJnrYXMf3s1rdPo0THaH2NJnO2wYna556Iykb0aYuHkHyqn3XkNsKjp
smtmwh1dF9lSUWAtRPH1JjuC3TCBulG3q1qWIdWq5KGWe72gKrmHmamjZFVpyUQT
v26WHmIJFf+2xIv+rSUc4q3WRqD+y0/G3rFKJtWnU1sebdj/7pXDzYDn/x/dgeXc
oe4YmuGKPnfRRVQVQI9DcqBC30nZNsRitB6JxVyrWlYp4X28EUIeyJKBXNkewyYH
XZjtYdSTVZG+AN/zhXWwgH0/mOWmZEdXnA/L6qWlpWxctvVTu+mIsdOR9qammp2S
ZCT1ebUC2fFkJKXGgY+IIRxHNqdfa4iExoo0hqLqKCVt/gD7dxwjmc3bIVrAwvnZ
W6seaCYM6cf1B19C6YSPgYgrYchLR5rvqCi60UEfT/f7UiCu7KrEIQPTCC/4GHpM
bb09SmmFDehx/2eiYGFyCuBlOULYftrpM1iNTSNbsBlfWfDK5bJ23ooX+wIUavpp
qMKazz+o0KigozbRlLtiQdl/G47HdhjElDkhHQXb21efr7cwpv/XzVhwVOEINxM1
Z6KzpM6Q8KX5RthFjRvM8LAR6XeNbsPrBxi6OC1T6+s=
`protect END_PROTECTED
