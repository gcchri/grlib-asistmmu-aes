`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E6HepwyP4uVIkSqRel59wlJAUKLAQS8bOXuAsRiQfp+XIYKBzseDe0uXWSXtTcJA
cLbU5RaO+uFZA35Wq0IklsyZ2PWcwaAUcMiClCOJfAa5CXgk24KJQJnFtKj1BVKp
LLzKMUbZM/hOv9Jfnaq5TWLlLSdyVjbll1wY+JqD9ztqKzu70Egl0MwQ7QCinaXQ
L+r1QondFn7b4iyiCWDC2233UNV+EkhBwU8S1Hd0K6iEAMMECFPjhWw+D3VDdDXo
2l1L22QmwEHQ92NBGkV3mAjIsIZiffA/huOzpMj2nEdQ3YgKMKDV+ES7Coyb1aDI
p6KTEHdqgFC4xbnGrlq5BwXmJhvwzTO4z+Ci0VhLSovaUC8dzgx7b6Ptt461dlwj
odVL0JvFEKiKU35b0BVcvb8szePQxUWldmGUhMNMDh3ArNHc9te352yxqZ9s0SDV
MbAxeUgwstI6tLKvmB+8KGaioYurerzjfmu1nJOfneUWQVN9NDF2kFqotlNc/dL4
`protect END_PROTECTED
