`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8XRIzXxBdEWl0MedHNlJMRRCPIMUtzTTsScCuUzIfaUhkbsmZjur2BpLbamW2Zku
dubwt4UYQ0mTy0gneQ1mkoNcy7XwqfML/WO0INsS8foYP37AgGWy8zPKpJ6z/4sf
V+NVNyrYvyAaI3B/mYi6dIHVZNWUqUAm9A78ZvMNWyvV8PDTqJsU4ZhlCxREPUnQ
gQ0heCek+buiACkWfKW8RJ6rux5bBU78taHYPeu4P98SFhS+4s7zk81mRiUBqGHe
8b/A/kQaHMgdTugLd+Ghbt25ArEEAcf8DEzBGmi/UFCG2ElAjMbdx0D6LLbNQTaH
oHeHU47ueh94kBE+lfvK5G+G9kyqhPMv25NjUim0G/TERTo7vVZYq+KEhgu/NH4Z
ENZriZzvM0rXSe368yww+ukK/eXBsr1d4xkTiS0zn5Y/vePHVavcj/Te2JbpnEpP
IFQG1oz4NoTUo/497fjE5gELG2MJF1ac42QxWSA8awU=
`protect END_PROTECTED
