`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RKu6x5CTN37dFRiKZfH2BMfoaL1PKN9YXpZWo4L4PV1BpdPHqvHGl9rmMFBcTE/u
tYeKeWRbXO00Km/5Kl9dvEN0/9lllYwthYC8XwHp1N5LnBNcJXhItKRcUaSYpf6i
40BrafJbgYLIgL+MgnJfq+snqckyNdoZ5sxXqYz6Xs/xWt71QErHHwWD79e/iHPJ
N6wfkSvkpGXJXZs1DoJ80m1b34cVLhTTmHgALBsSdiojA6CJb7jADSLYvOWLv7Oc
ZbbsbvwuZXWJiMzZQubNLGSjwL63kBe9NweJoNq8753i+MZrgtjvzosDX9wr5A01
1X2CSq7fm+OGzP4A0TGkEJ9UrOILF5hT4+mwfYHOBTCgUG8tAm301lcB8OBtN9Fk
kqthUpZGs1o34naNA9erur3njfUpXgOD+LmEKqdXjS3hRBXd3xH/Cd9rnAwVZ30O
i2jI6HeuPccgtgXNuy9+dTHiZSXBkLFX2OP+e1PxKE/p4VKAaKlkRu8E75KV/QhH
`protect END_PROTECTED
