`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KoIPQQj3/m3T+JyL8RXdZ4SRw5R+C6olTnURXDMvg5BpJu+UtgWIDwMVSNdnUwF5
EuctkH6nuFKmbYcalhedabSwBbo2eyOSZBz+Hg2lNcsNV1o0PaThHy3zku1KJm/V
a/R5oHUIguUcrsyoxdANg4hAcvhzaSfd2pUYk/ij1SNZ2BPWfLCNEluKy/cNo36k
H2Q5TK3LTRpfdwO3eZAPIpTjSFoZMzWGpTXj2iYFpez56xbbvscRItWsb9ITHgL2
OEqRjI4VYMsl6TCPvEO9GrDDb6HQde8yJ1Aqoxb59EwYzPNzmmrvkT2/q513gfbm
A1z96wDZgjSYnr1KLBCPQ+gvCZakrxEaN7Ckzy948dNJIt616qbSqTYnVuIMFFlg
AyvlGgAPUaw6D5feE2BEt/Cl06eTt3gTjW00V2jTbvM=
`protect END_PROTECTED
