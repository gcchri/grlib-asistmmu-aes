`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ym4n5gG/t1sSYu/JatgxPgtwse9CfACm2pQHhELbaVR9Z2jun8CuNHqrUgZSKF2g
NFMpoKa9WFwOE+gUblE95ON8USIg7TjmvvnMPtLLMQ7cedKPOvef8L+UoCOOYT2J
/ZhYLcnjhFQwVCGQ8NKdHcSgVVBpabuUXqm3vsKdrPxCstTPgmUq91GNMpcDBwMG
a3zGfYE4XHxYlk1S6rAe8ZZb9xE3fquY3sYNRtYn+poku//TsGGKiKfy2LVX5XXI
7VnvRnQ3mQ/pwL6rFqzbVoZ7z0HfQzHq4T6ExYnDiPN0WWC7ljHNn8r8ivnVzic5
CU31Dd8tQ1BM3pxPwv9IQBKwj1ibcFgAx65VziIklPka36xxwf5rksivOw4EMuVe
YxNaZJbM6GLH2FRsDdwAOtEAMTiB3XDbR/iAEdiig1QeHhFY4c4Fm5vJJv+2qgbr
`protect END_PROTECTED
