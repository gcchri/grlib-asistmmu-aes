`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zALeUY+I9ts1U/KEL60OfXS6N3bo/lbotNCWGIFT36PooKj/g29FNBYS7O3/SBTb
/F6ptx3IglUVWAvFyi/GlFBGl/TziotTsg4MVPtfoyQkM0J4Fn7te1qJzJ/QYp2W
aTky4fktkSnKCOQjww+nD/lmXCj2y9xpwj+bNwSQFObptk1bJlY4+Z3UgdYcUYVw
CBSVR9mngXy7cYqiRSXNIo+4dstucs3HxPVPAiMm8ESTyEwikcmMWhLt0nrDqyCy
E3sjeIobI4+eKivA6zbAeYFb3vmIC4Ey8ATmGcLJ69fRAAbYTTyT7ZcvQOhTPiIK
oltJIT2NOVjY0EHi7ZEvOZH0CwkttREBl/Itjq/dLbuHiWoxZfK33REX1Xy4U5Ld
AetEJppHLjaJUbDxs5T50hPmCe0DnS92ryLySwelJOeZUsIzAXX7gE2pvLGNaY4W
AIrEPfW6ONMSAgWraIvgAv7Bje6wnkzE/MmGl5LIf+RbKVjaqplyTkQkY2psJoPP
+XU1/F0KOmXFtiTBo9kYiUL6STSa59zu8llDKsaCJpGwOTYeW7Z2a0lgjn2E/59R
9XwxeC46OQSVbjRoj5Rv1dNuUQQqj2yVxiq12UXIFOdvbuW/1Gi3s6bBi6+1mI6V
j/iYtl9U8Nsr89p7oQtDbGmsT5tAZ5bO16gsqeGtkDR0AKd+oiXKA/xYEg9TYkCZ
MLWKwKf3+WYFU0xVgfqiwnxiVWKMXdkoku9MWhlsVX46eZNvegLeUAkvcxbkEFsL
KvAk8XINYXM5elaIh03/3sXwpfFFBygtwPU1+l9TYUYC/rw9Nt2EIK90n5a50EF0
35mqMlmQt0lN3xJE7h+8UAjIuNiSO3kTRpoCR/Zu/cIK9WYb59NI9Ktjd5R3KOsE
RjmVA1jAjAd3iYhb2cWcOhgL3DpbP9gZtekHcYvdchRgdAFn9uEhLpjhVmXIiUb/
Mv+ZRKGcS6w9swACzuQyZYiCqX7bT9jJdmhFa2VB69BT5ASt0VN9fUu+DxkS4gMx
dVSgMuj1NIjK+q4N+nKxf/s6OPPCNVyBh5qjT3stqUmKFO/5oVcoA5IoM687iEtK
WNqD4gbpYhr2Gcu4e3LquthWqmxNl3UfJtaihICWKnuyaGsY2YEew3wfDQQqwIVt
KbvVX+AIlwhWK+QA8N3FOKAKoJaHQuNNth/hrHS1+mu9cJ8KU+9De5silf+jdAIe
S/Q+Zbie17d46sHW/mpDOijgTFD1z4muw2hOGXPTd/iiDbz7oX6WnrVjLS8NOAhi
WNn+NxdoFQ/ZPQPWz/JmUoDeTM0DFIikww6CZM6dNTlx/mnh6/IyyLIr4g/qXtkN
uLobb8+LKoddrjnZykCXwUpUX9qjeh49PS4w6pLbyL7ywVjLBwKQDMwX3fXq1Xml
uUvZQYcHnIJ7RdzYXYq884YKQw8CJdR724xcUbTJ+yHy73yB9n6dSSXzVUYsul/D
nsAXv78TXzKJC+5J4j4ME3O1qgkDSXdJ+X5o/F3yTR1rJSMYQcEseiL+Rr9nXxAb
VVGc9tTrg8bn3gkNAGYOpQslMJd55iXDZ0D/o37RFXMudVQ9i7OL5ha8rpu1UEZH
cYX36/G5xro/8ygTdumd37bofKSnxBxRDSLU3DhNUplR7FZjUBW65V/xuc9mR1eW
Z+UdPaxHH2lD8an3Fh7BMaFO8DBZDNWUxq64QNqNNyu98lhCp+LFDur0i4FR5QCf
tYEFlNJJu9teOYIxgpBEMRdMc06CAgEqEDR9LZoOuq0us47dBrr6E1/bkqraYWz8
dwQ+BBV4+ZStIvWpXwWIDr4vuBE2mbseaazId7EMSslxooSRlF/BzMmifTspdOB0
SFvHm9Z1mMoiRP0vBeLxFFRi0hxOE/0bacTc05u/vp1MwVgTdOG7eezzC2f6nmGt
jF9uoOkvipPXIuijfxb4TA/20SC4sqYrl7UKCAJne7mDJG0n64hUwHnW9XTonYPi
QEGB5fDQI1okBxfHUMybZp53qedp40XDq4j/Ehx2mzej34y/aEbkDZ0dJkARNlvf
C0G0ZqUxLZmvFDEvSwXdSQPM3Ait2BfX8VuCKWIbPDRBYwH3BOEffA/lND06cTMt
Rf6GvodJe4uEUr/yIFXAw7GeaYseeJIKhgdBrJQD/0rnAp6J9Khf5Qo9e9I6WdJw
sg8hCxvOH4TDyY2W2UBnbCUh0Fb3ZywBuXL1NNisFPB5dIEP6ypd7UHiue6XTj1k
ftZp7yTah1p5jra99IAMG4dbgP9XOutcoVtqwtBBKyHAVbHF/SeuQnjpPDdHIyEy
qTKFHFI5BRgJEh4soKwAeQmKUNIXNYHUhIRNS64oKoT34U/YxleHdNcVrr2BknCT
fQGTI0Ia97RS4bG0fpdCte8GmnwQOZxeWGex8guzTAA+/C6LHV6OEYi5Kho0Dv/T
NZvCxuCe5rxxAUO7UuynVe1AavETWGHDsVzVGdbxjCmpNUYdPi853l9gSIjaTnIT
KQkiIIy2uEfJQj8VNVtk+IzhJhB7ovMtMpNzzCG/nL0qmiOPmN4nS2GkFlmd7kPf
ZJGjIylvC8H24DW0fnG/Akw0Bp5uJERBmVEKOVUrRUJJd33ksl3O/F98OgHTXQ23
0M9qjMdxEZ3OQ/NdaWE5cygNKYgdK493Bxi0tKVYcTx2hnXWl6eRDyjsL8dXghZz
fdaFcw1wcTp7kUJUrZlEfBPtsrgggJtemd3mTBf0qSp9kwwO4akZnwMmmwsTyLVm
CEhRlneVFmOub14wRtRRB2hC1LBSkKkxYB1rmqddrbVTyRav5SiAtcwcjmCv7l/J
SckIBRlI7hfXQ9BS+3tpYYGT9eh67G5DXtvfE3q3PEDmccRTdqyJqO7vwvrG+Scs
q++SqH/qEEnW8m1F5pAap9yXcKZijFZ5muCtNGlhzv4w0saXGnUMWNHtRp5nly0m
`protect END_PROTECTED
