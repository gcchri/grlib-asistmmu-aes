`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1X74QH/3ZsYSJE1LdmgkFMPezeNUmxHAhsGXnqjL8PhxydU+qXZAPQvAicqrIWM9
SXYohERmA+y8cacGf3men7l6mvzpZ3GSmdfeYruE53cfDJa2jERBIcoBa3AmykH9
ppMWPRwvxB96hUaqITUPfApd1EWn4eKSZiv0iyUNbJPBFeBFQqNhgq+ZMVBUc/aK
Jf/gU+Ne4dbJbcSfzqEiTq2RKs8Cp/OTavrgdtbIi8dSetZnhZIVwPdWVprnAhvi
3gu54YmKymlrcP/3TQCvZHWEs4JjrgK6GRbEzFTeIZjvGfN6qJsUlht6NklxdW08
Lp3Krj3a7Lvu2kUKK/2gPZjyxu3geNdBNNbIRKv839uaNQh00fmQmEjaSLsaUa4S
ng7LSJpVgiqbvx54H3gFFgAYEBP/dMvU6ZjYk6Fpr0KwQRjLncFXDG2d0AZXRETV
KlGMbgQTD4KP3n933sN/ScipDRRNSjIXH5wQO1X2cMTFBAFc3RUF7Ta6VetBE2cN
Jgxg/lyPuSbsyyXn+gzzCw0LZHnQKlaTSPE5kJOoOWgSRzf7ghbX2c5/eUJ/pk62
Zzf4qQ+sMf0pmg30lb+iphW9Gxq0j7ckUS1Lif6UrSP2KxOM+cW8DM/pah+W3GYe
udQ0+cRLEVX5f7adUJkTA6FIPe7GI/ovYS+Cp030LZ2dNjF1QKrF24S3JqmfoV7K
CbPpPFG79zzLFf69mCrBYA==
`protect END_PROTECTED
