`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LF0CwHYXPPIc71jEVkK+hpt+00BpEn4AXC7X3NSv5T/seWxSCBZUU6r6Q+G39t37
tKvhvqmfVc6JV4+AdpQi7C/vBBix4IzGkBfvlhF9ndGZiaMSrFgxPzLYS9AppynN
4rralT+8/jtRRBPzp47jixRPYw96HK1TgWqXUzBQipstJ/f9o2GfHgw1tSmDdL1u
EvoffDF2ZNYyyuByvDmhDWF+z8IWH/9vXnm9KadQAcU9vK6elkl5jootbmfuCmiX
S/m4Rc3lYzR/k+8PIsdGlPEqeQIS/abZq21jj7zKis9zA9G/c3Nr/+tW+On1WEEE
`protect END_PROTECTED
