`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jvCpQl3IS0yDuItaj+tb57zvROFTz0j0z1cOBpUodGzQx4GQ75qa/DHFmy9z98Xm
Z+IMUdkg886B684Kw4eS/JR+ljNbc3LQ3cw2Jssm4lWjfSlEaCgpmpj1PZnwSEk6
HsqXXMApdJePJWjC1ED9D8iUuqzMlYx8ovkrnvIkOctx7qWyK/ojt4bNHfwV+qvj
YfJFgy12upnf6T2AwyM9b16fZ5TovKmxjOtlTMhzdR4lvNbZZsrgRx07+02J2zkZ
As0gyCBFuq+Tv2LnzVcqiMY4TfOvMBVMgCmqcyF3S2kCVWr5IqBUDdvKWxUb3qdf
uaeBGrn1pSBki6YnGFusO+djCc92M/UU23F3UKj9XkD/9iO8NMHjrR8hDOVZqWke
CfTncz+A3xLvbWPZthYPUJsVBUvWfomX1qnmZEIMuJooUbyYFQyy/kGMKocDLCK0
BYg30beGyTjGNa0ltSZ7yB0nBSCrQ7GbsJMeMYOKAucE7SmL3lNSGQaIxVIlA8Gp
MHROu8iIIEp3h/Z832bV3aMzwNBj7ng2npwNj3m5dPpDNPyGn7LSvF/vjt67vc/t
bQe6sxsrwOQ4lq6vqlZo4RiuD5XaYPUM3W/71lJNMaqMtiDBul7/x4a1BClhrkOs
+h1o70Lz6PBgkHhIctdOzOk/SyTPxCwo0hnNJ1ow21fIFY/RuYvWFxlfE4un4ptf
vHTv4s/iQ+KsvEbYOaRjpr/3VGPB5XXrYagUeCO/Ts4xrvbm1tu6ZjWrl4iti+jG
6BnYNm9wrjkHzgD4H7yP7146a+LodNu6d5ClhiXJ0S9jILXiDrvX94EPuJrq2zD9
NiNY/+38nqmVmQxVvSBBAUkEk05w8jyH7aWM6FPN8zpNb8WrDEQ7OGEfNF3aHjZa
f7pNcqZPRpC/NHKQnDszM35K+xPYMlIt6f373591mXl3PbGL6WDvsfOWnUugnq/Z
f/67lhAHBv8JSKh79FXgcdsBaK5yCcxRnCDJXjZOL8hnWBYXHnVRrIUJj2fmjEND
Rn4dvAs6jsnlKiN2NeXvZKx80T8K8IYspnEhuQfjeMpQ6vdOTRhvL2Chhypp2zxj
ZkRWwxWODcQJEMXErdYg1d3P+jcylfRLURTo0XEpCd74M4vxJdJ9wT+UjWpgkKYU
JZlxxTCklt3+FCZTRQnW8JOTDz9K8WtmZvtX4co8b2Mr1v/n33e9NRl0OXPI4VAM
nuI3kxhzxOM2OZ2X6dZJuHPlYH5q6vYIP+h5LAmBN9twGaQuZRsLSKHMbFsxwdoI
S0cYNd3QCu77Yqrru03AB5Fyp8LNEfnrC0YW/BSVeTLgyMfbRYaXollrW4+jM+iE
mNxu6RVFjbrObH4Luxwnj9JbParr+opEoFVrgp/nf0LDxYp48lno/0ieg2cjyiOo
G1pCH2pdRnhCzYrAgntgaXfw7CGto16kTrJw51A0AHmSlVVU0Jja4Hoy70qhRQN7
36OG7ULSLE5MCjzJ/h9mGmuv4G2DZ2ms5vVESnJyGw4aQ5ND50Vn4NPMbgTAZlGc
6VqjhK5kvPQqTHMet3BaJL2xZUvp/B63muuDezIUQ9e+WnHabjhwIZrfD0VcxrYq
Q0m/RDM03644Y8DRhXtYnGN2gAuhCC4tmv34C7qLG0EgjODY91NEXjdcSS2lLZtt
mxcHyMrJaKzYu9T+zYbXlO1vbCUHV+j17biE1U2Hi8cEOv666g9kuvIVuFZnJ6CO
YmtkVI/mru6DyM2TkohReWCeBtu+jbJmOJ5YpsWbjBXejoKFbZmbf8tosnR26tQT
H1bo2lfYGE8WOAFMK8i5aS3VsJfsS/2lE0uRsz2455vcokyosV6haLlYdgMSJ78E
rNZiY3glwT2Y5v8bisLgUHdRp0czc3S635jF7dvrX5e8Q2ttZbzdE+/DzPt/IkEH
yHmpfoOK2T6tjzrHf3UjllEMkL7aMB7SZYn6XMu0uadxwAIbTiAErHF5qti1asUN
D5+V/4llot6ep86633UJHXcJnj1v2+86AObWhvAkmrUdWs1LPeXe9KLoa307OGn+
DU8zIUOL6b3osY1EJw0zBoHX+dQ5ceEJ0wAygKYd2jk/61AxmDUjwqgWGhlhMHQM
qMlUnK2MhBw9UMiF/Fmmu+bLj8aIbFteAclxntrARbeq9pJ2rclW/PyZXJt2Skq1
`protect END_PROTECTED
