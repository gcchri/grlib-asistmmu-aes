`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oe+v9KtXqlghiMeJWgdGF/zXrNv0XD21ni3FepZXGk3nCf4M2npfAit+uy25HSa/
2hH74MOLEzuXCbwWoubAJDsexuoCLyIIq0v0U9R6F541VQ/5SHtywPhBnexkEIYQ
iWNzm2UtzWuPSxzits48tdW8W1bCAWMlBHf6h8ELJEV3XegG23eCkk+rEWnXWrNe
u+UY7HJVPi96TrYlL1G0tVTIY5UKGJdTm6wrcqv89yGb+C9YPgRuHDviiXyxKh1f
2ebtTkHrpWMSwS5EwZH7+BzsjvzPtVC2rdqHlJpRlCsT4Lo79ks7X0Tv7BL9BCcx
O8EPqvBhkbKdJDYlCXxdQTobwIZk/n61KVjW0nM9fpxL0pIeCXoxWAMyi4cVWj6/
5mMB+0tEBpwHxRhRP6XF920misltyTALV6rJeesVM0HSomXBEE3u2PK7Zs5SQyUL
8Yh1m+nutmurA8JaZxd1frZQHDYgBm9g8r4koCJGEMuUr+sdLiuHfsYQ2MXpyn2E
U9MF8eG9hnBIWDNy+MU32h48ne9enNkQ0fHEiqFPZgfy3qcMUfZtMURx3yfr3CFL
gANEnGlTzPcUzhrclWJ9aV+nhieqN9vLwG6Ej9BMicHllHWhQofsylUjP3dDYAMK
6ZOeuStMF2TLqYGmN2H8nHBjRvVuyZLrZ/qxI7dHmhrq0Ij0D+MAXfTkrHIjAUX+
NlKsMfnm2i/UzHAzSbkAY9jRnjZGWls6T1TDfHYfUZ4fkZ/AcT8fiOv72dg7DocZ
fSBgjaAuVI5Mw3f4y2V/6epZjgYs75Lzgvto369v0e+O0FkI5S1YpNUNu2RoRGiN
265+R1+Z98xf6OKZHpcGm9lE5NodWquTJvwhNly73T5P5DiuqWHMumvNXS/K5THr
7zK/BwvArLwXj9jJi45pbpNFtDLi7rnaqjyY7dLo9YvPCDDH6r8WZOPEYUPGW0cP
eBtTw/SIlihliTRRnZsjlPXktFN4aOieToSl4XpFY553IPzQGPFfesMm/pD7iCVw
lhJ3aatKfP+ahCH3aESZ10x5/iyUTBd9d8JHE97J0ew80zk38LdYfusGHxjiv8Ju
UUZReteYB04c/7CIPpbfF1oJkc87JB26cZYMq5jPs9g6LG5OePJahdvVdQRakyYC
vbj9VuvNO6/DgirX1unBAD40kGA9UlpL5vxd6DYWIie+ic5LmeX09I0H6DzPc5eu
vikYky9ZDZRcSxXsWKY+lbnbrJDxq4E8N2imwUo01QXP0roqq5T5t+e26vqZRHwh
`protect END_PROTECTED
