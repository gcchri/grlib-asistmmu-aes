`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
udGQC8ec+jta/kWtn5tMXDi3OC7713V7G70tTUUl+7dOwBabwKci9wpb8dejN5rn
sTLY6AR62JiYDRsO3CfMSUg1PwhMquKknaXTmYsf/ysti/RChgMKlTkhwvu+Su4X
V3RY0os/jOhtMpQWz6cCyj+e0EuLvrf7dcweiuq+hnAKpcps8f8zsjk21n8kH4mQ
68wDKFlVr+8eng+2zRJhjxRyAoJl1/bvBug7/CQbP+B5gb+JGyEBu63wMwNHOMNa
g6D20mu6+XZSWZ6YXJZQmXgoPur3pg2MrN9o4Je18T+UYfF4u7ERONOB19tBVF9p
mBxDSZ4R1eCDDk8alSFCsyPIW7YMq3CATfzLhG9X9B6M1g5frYg72DnGDmNYRyBM
16WQpDnx0XlbMuZUxQ9sgFpETM+WRPMhcE6ACiCHvsYGVhAwqIj7hhFggN8IfrYd
rB43V6+u6X0zYXpw5bvxIoia0POhOLkZmVg6+bN23s8=
`protect END_PROTECTED
