`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KvdGff70UOGuepc/sC61DMumxVAwmm4K3z/aLheMLA2s+EzV37Ulp/YLFfTPZ21E
GOwJCvk+yHpt0TqDJtFBgf+sgp+rvOEtrB6ko/icG2t9DozjUk85boow0aIDlfVB
F30ugpiuqDSPNmHGxFZ1/0LBm36KDTohNYnrVMaCcXhwzWbv9pKVcxL5kOV4x2/w
Kl8zSF4AV62nYoHSvr362vtdmX5lvzfTHjO9rmhYkOVtd8TrcHu8Ha88UfnyjP2x
L/wvvlfqbS44pWOX3h1tLuokrcJCMkgZIXIQvjeByAgZrF7UWO0NHNB8RwViaBQu
Iq9qUqQT5AdsCxNIX4l7DxewzniOB9r9pufT5MZfEzMIgI3HsHufpFZlV1oD0lq3
FMALryjSPpkWkkl0nafl9xzbLyiyulGw6xlveRiv+OG4HuBEMaL67U0GDX26sI7+
jOWA18Nj082QR7MGHwwKX4g6YCtXxl7XKVNVeKe1wL0E/KbLHZLWsjZ9PGbsqWJ2
16Xgo4j5itZjQQ8RM+2c9NKPiUvFanTwaV6CoraSiMi5WdtfYRv4Vhi5DVmmBQn9
pR5MhQJFMLf30yCNTLZktNG4TXcTb8AOg2gyu41l0b6uxtXX84zug7FgoU97AJvc
jKp5dhxrMVAfpVPbkHAHl7y1oDnTj71VvcDG69vn/znCCDOggKod8AM0EGXPOiNn
kymQ66mX2xJDE2H3zt/nRef/BFzUlcB3eyT+jy43KFUL8EnWLfMdOsgibmVo1CF6
ekFYU8Km17L+HHIoSOG1hQfkJ8IvTlR8+SIwgokoo3o5NCc5oHxGwv7lnn9QnWMY
ZjuBHMaK4IgcNPnHCQW4rvRkLy+bFTDQMcZduQFKULAKW3dDzSYsPXQ4qiD8lsbd
XqhmnHf0XRcAKnO/2n/YRcZ3G2lalPNOQw7eqm0KQz4LY38g6ctCWSbXicQeldmJ
bfBoeLI+uj+I5cl1sdt9A5EgNYzGayKpvnXuD1txPhZe2GXdJScIl08EjMR46TQ1
DoXSG055WGp7BhJIdkHlNkEoi4EC/Z7VXXmV4XDOoUs4a3SLdoSbG6HKgX0DUvdx
mLgsvdXeyYzPAjCza7kRdPaHVF0voK+asE0TebjnxwE=
`protect END_PROTECTED
