`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1W8OZeAXvzIPEVqz+dCHJQmmGAvshtJ67LFMeikCZQXypVprsjxduJz0j6wYPUjN
PYDzO/kJI0Pz/ZwD3uHkYsaBzHhBhhMejLgbtp7Zw6DHR9hNcJOrtDB2X8Zi22xf
dyNG4kbYidTfs1JtA93jQc5KxUH+ajIKpSCVgxcbeWAyKXxN11BgQ1tNlGcvB2rc
4FSfjdgZqiO3NjNn37hw2aUHm8uFXk/04plhjIn56LodFsbyefx6vsh3CAuAfEyE
HiLBHm4MW/luaw9utzBdZ1/s02uOk/yAeQOn8bKY5O+ZAg+yC6t4QDNnUDYGwhiM
QmTrbMp2FV8hp2HSBaHHM/YWzJw+FqTrv78oENW6qMBS9d0kH9x7CU8AK+2+WCUD
Psy+oiehap9bMjsl7D/xB2w+NwmXTBbdi9I1kq4v5NDMO8Ftw8txhUUPLoj8A7Wy
Q3idLO0uIigSZm/iM3anACyDQeGWJckfjvwOyjsx6Dbqb3S37iwlem2SKJ1F7Dnt
QuBuqHAgTHMBJp1ps6PhMZhLbHCpSoMkOjSUn+09Tv8Sg6BIN/NpsfQ2MWWQMIud
bs3tmKM7skUX+hEL0kKKO+vRW4oUNxvO9Frwx500cY4VNrH9E+DxnRBd1zmGzTRc
iYKnXxVv3nZPP6geXGJxqD+MBQBKbdzX9GjokbOmaU1aDvbQ18Aj4TmXXE2pWfRO
2ZVTBZoQlKJvHcxLbijisi71EnWxXvdlsfsD4AmFMgiu7PXXaJ6YGyk3drc9QNgd
AAIAKelUy8C9UKAwepvQl6BmuYahg3GPK5eTHJmG5L5aw0p+KhsUwtYy7onqM9KX
0INlrnTMvRZuDySPM9nN5jwryRG7nfvcW2vabSM9360HiKNE7oYCLTziixAzrg2Y
+b1nL+/zfqTpP5aJfn58ZoAqkUHbqKyNu2Etel26xZd6UWP1gHczcobtuscz/dNw
wu4o0N+z6WCn5qPyu5k2fSMbISQQs35Lgt9FgqAoyELlpPfUVtxzb6JT3gse9EsW
8tIkWC+rM8Mz/8XCCWZuQw31IwGcMXlf4oYG0dcAheEdTHVzeh7yUSIKfOj8Eclg
8egEHDAMoPnMLV51LW7vjAD2MZ5BXCafGiaqky4ctxJ24pSqYfkMriN2BGMk/OQr
gzwOlcrbloxc7HSIjagXDl/oEgpd8miZvZPwAyCyvZr1sjlR0ZsCsUOG2AAEjird
pjxnBllk2SFVYMN/WiG19YazijFylrdveLneG0PsOc6VgnvLHbTyCmrJ6yaQlgm9
riqYzbHPRfot4VKcpVThkMmzg14bz8FUGDiswX9i7xgTf7RV3EMDBz9SnnPvLl5j
WHXxWO7/WaNAOmZftrhNdw0URlXs1OEu8H4njZqfya/nfgFcm26IgY41CjUvoZgl
+G7UdX9iV0UgWCMkTp5Pa+eV93Kxln59I+8x0VpVuYbujYKogI0yIZgcAG51lTHF
le2UFe+FgPIlKfRm9XdKydkr9IY5GUWQ164VHt+WQl+65+E9jRa2/6IUuH5iFW69
SPJPtuGqor9RUeJrAYe3yW7uU3GvwM234vRp5dFl2F/qX1MuNV0/axm5Fnr/2hjC
azYD4unsEJCPRbWaZR6WXHidGiFZtUFFf0EQM13Sm9VbTjYSU31Dcxv/V9TRtUI/
j/TvIjmHY0HJc1g8GKXGgHu5DPeqnZtCvgvq1snw735UudqNG1/98xjW2gA85QVq
eG0EVnJvruZbBIH31rvPrc/cso7dDsn/fOLOUQo+TbV3eOmBkq1rol2HDKBxO7Hi
2MP0e9r2M3C506s3NjwPw/ETNG6iBP14L6JrwHc6fvioMzyDBH5sFx4jYCFLQmfl
q3kEX6mPtR9dgKAPKxcec2HadVK+c3Lu26tnbD//WIA0AfF1nrfr6IK+BmxvbgV5
btoWip7lqb8eZp8XfA7cC8GN12beS7CPnJGHTmezLmkfeDZiabp13EurNLEqfCxZ
x37zo4zpMdzVT48OTKXMpSj/MKaJ3OwrXtf0n9zH1NUejEd7v2zxIhd5RhbAzWlC
ZkvjztrAJQqXWT6tuim+2OeBZQx8whFblY/krAH671jtNxg3upp7STvTj2cjv5mt
lbITOxCU2fjP336Oqr2a3BsMeNFITjnmmOUWoMx1JhN2QYB+4kgiepCejFLSbDCL
92MPHn69/Un6x46l7eD+LJe6qPCd4pDs66xDtOLqU/hClUclcq9quRzwtP8rR2C5
xkroOpRpL2ragjHtwV8QysCNzv/mtiofyuBcnR6Aasr865Qevf/OcgNNCMu0jddD
90nzZcX74uEg1yPoruy0pPbwZLMkU4P48TrY3LlYFh1aa3Pn1K0RBW5xm9gyg6Pv
quWYhpLyGq0aAC1Ncwpk6ZZVr/rhiE5AE++/lR76vzUJc0/rzzf5DcAVkQpKC7+a
ML+qoJG1VkstITPglnuVnw3ANPYfQTFp11i2BhTnP4cQFCsRP7VbSflPV17DIbtK
+mgBdb5aJ9jiKuI+KLzpZkvyiA4q0xFg1v09tohoZKJqzIoq73AR08DxD4psyo0W
3kr1ghfSEmXQ81+c4BfuhIg411YYcts7dHZ+V3g83MgVf7VhoRXHKD2gERGYEGGE
bvuN2GRThVt4SUFtYP5LTjRktaV1Oy9iFXIU+GJ8oLTZsw7HbTmA2iCKlBAr3HKm
df186k25gGGmuEou35V2rPCufpo0Nu3VKbnfq59ahgyu75Gwi8kM7ftJU/wbRsp1
B6DIRXGGh5W8LViRxI6AhgK6IMCPkewmMUfGR6+9wkM4s/q9+6jppL1NDRpQeqxn
+S5oqZfghfSXz8hZiRqMekixEP2NDyHuNnxS/p5hrTnLuMy5YLzw1zMj9yfJwHxA
onQNZkX0wDp1GQ11j34iXoniDEpWQZsinhi5Mg3E50e6kSooh2cO4ey1kjIVkYf3
EQC88ZsB0LRZfp9O8N4rljG+PJjlw71jTijHZa82x0/xQ/hAxu/4alivmNA7MqjV
A4WXlR5WhTBiq1D39N2XJrzyU5Bl5pNzhDOqc8UHK7JcDZTF4yCQRlTOQLcysaZY
fOwx6noJH6PbqcwrYik4S/RqYi8x2/iTgKLNMrWm1ejP9jOqb34GDyS9GJluKIuK
GST+S9vAN5BRTKH/kpe1agcv2nWUwHkOw3DeRjJyUhLKq+uyyL+7PBoxqFw8Jutf
tmy21igpbIuiKTsREPn727G1HL/uPfiRbwKWHkfp1LO9jdRzfgm/ea1oFzvhdh4v
AKP7uHqI7lSmagP//lgomZMVugx8Wskk9vXiERyikGZtKsKELzk80F/n1CLwzgba
yL+QKsjempHHnVODyIaPf4kHiyt7xWq77ePnE0A1DtxrIqlkvlQ4+wYq3nh8dK0d
6aNPK54lzmlkGUbPAGdRsU1Y6sDdpgdG3iG19WJwJNfuVZ57pyPKwxhI/AKEsRhK
aTntYJfqUh+NQb2+c3djiTplaVdUwVslrpc/nx4TpdUla4SYueKtEDD7aPy+mL5J
ua/Fsti9lYLTd4O9LJAKzsHvOXIdNd1iBYL1RFPkQa+VoGpdRP5yEfUGhTmm8jvi
24F2WGKK/FiNPkMTU2dZkIUSai4j/Kb8s2j0urXDzG+dkr5A0BVnaIi2xSD3RUgX
0pfr0WACrulzd5EUCNiM0aGKOd8c8yeQvp3tortB/YtYtkfxECG8YB5EGqgBMJHK
wYhizh9YXCfNXO0ps5xssxLNnUpWR5FgFJPldg2wtqeDWA6LgoS8dNQ9JpkA2w0q
J3e2H6OCR8JKx1wckFjxhOjVS7Ke16JSniJtZCViAIujI5vG5BKEsVRxfdqxP1+L
/44+NjBs8mju3TZQgxaETaDKj3kHnMHPRjW0ZQUAWWQt3cXqtf9cMu4Me/ecePaF
d5mo95dXgMdCDOOkysF6GRKKm4l28ryhf2mxLK0b14cwLN1O/ZeH5903Dt95BI7I
PoEiBKebLuTdbCUHBLYBOQhMDBtbHN0RRDX6B9ilrq2+3w934/uFa0y1pePlrVXc
21cuorHHVolwBAuu2D1PnueTz2mPkudbUfFdGlfcHRvf/bbmVbCzt2GRwcRI64HQ
hulS+XI+09jRbgyJWS3vdqlHRPFItwNO0AxWM6IITwyDd7tId2YfeKJLqbQzdevv
dFHssVmZxHIcH6ZJyGiXAUQkAbJvHjujL9sSEGKCLQgDcN3yTC7AJWpgpCFlcCtA
DRfD7m3sHL1nWzUeiaurc31Mz7LJuaIAbQs4v+3r2A/RAVCyP6O4ocstbZPrluLJ
ppNrcXQirtuXZQorqBzMvYDCX1JVeRAgwaI/qmzL/BkpeZFC+BQEbaYUCalrga+0
6zb6BkvVhBXiDd3G3GPQUn0HbEWgEIkUDALGVs9wGBHapJLwEL28kra6/4lQoy8J
xN6PWsTDYpQGooUfgPmuBoEsUUjFXprlczSSC1pvhe4sAWXOntcltouf7L3hZ1d7
SmzrPd0gkMSNNZbyk11vIfT3h6bRbZfASnA9Gx4OzQsQHWw9uIBuEOF3VtjGmYGN
6D74sj1TBDbYI1mz1EsGTo5c+kUIVIPwjIEPA2WLi63bK4yOVXfW0LcwoyqdchfZ
FhiBNBJXZrMu4EZXCgd55pJdrIxpVKF/0lhnfFDGMiDjfRrfBfldgpRioIJCSIQj
yUFaORCr1iPj9QlpHucmoQwwFJKjCWa0BLveSWL3Aekk4MXDQkLJ23KTAu7q4ynj
SN03u3fOUf+3mij6ZQUb0YiL2oj1/54BVAEmrLDrfTTYsQhBuAtYdXdwnpNzeSQs
JR2z5eILIbcLQbEB8lWElQv1lImTaYfMjy+fNxIZEATs9z9kN96s1LQ2cGQ0BShT
M+3HCgUfDlIeF3JuiLY59LGKy81js8WNi5ebBKSQ0PgfK2pUCvEzdlMZtPfM/SMg
rv07Ai4ef149arMUfx0soK5MQcLQEjFSs/Ldw3N9E565HFW/rAn0MRfs2l7SvDQI
9Wj3m2ucnWcFYpX2EZFaQK9C6IkOFjYQulSuICG17sDXqSOWV4s/w9nxNputAbND
UFrFsr/CsU8SacTUu3eU+oKDRmeRdML4ufRnisgJnrIoN5xlJg4QHOfSZBv/ghFC
okJfWBsFATLMsmRfvb5xe0KTS+r/hpDUd9s/MZn4Vl6chyj+EJLWVPohqWshnQ3H
rInPE+aYgD2xpZKD04h8JT/SN5epmf3/qD78w0wAhGwGPuVgVUHPjLZUcKuUeRxs
UAIZRsLe2oeM9Dzu8ASPICGsNlNzUTVpZJA2VoH6sh4mE2IbfjFJI3MLlIUSbFwi
a6WyCL5M6X93PDY73uXD5hyEdA4e22hikqDmUpoY8BNyMTr2P2RdQziYbsKwd4Wt
UuK5oqXY1KR+tTIXt1RFtnRia8OtobGVsvxG0X9e+zlMlKI7o+LUH4q9A/sPjFC5
d+FlyELZ7whN3Y+FWIUiAEpVDn30AmqUQ3HlW1J6mA9Ft3L7p0/EoS9zR/Gwsn7f
IZ/DSMyvM7uXlHwiQopTQP4dirr1WIGfXUUtfvDpnm6ykh72P45y6ZG0mTvOL/Kv
DpdLDtTuBzvwkvIlcAnr8ljRBY+twlXOUcTMMLWg+0pGRItIOU2s1rCHf84cvE0e
F6G1JmjTZU4VQMg2nYgNknFn04J8Heq5CHNMQif9GrhjFxW7bUpau4j5gpPtFdtp
D4kO3aVBE9uoKNCeP7/CdmhOGsPl7mlc1Eru18ZYEAnDzoHG/TkJ9E9IrgTzOF2I
Nu8cfo1fXxD1YpojZd3dyA/GZkTDszgfjewZjn0SgY3NXACuL7MV9x/kRM54QeML
YU5y9iM0kVgPhowUknnPSwe+DRRkTQDkmQXG9HV4Jy+Pvd0rq2QfMW06vhtGvfgO
c7eYu9AeUKlJxN6CsKlE1+9utG4/bhpxgQrU8TCts8J5Ws3T4uyii+HZ9GIhMfD2
8p9m5KZsz+7ALhQz9QWoDxTbGwnfF6esc9A7ibPkw2/jg48qV8NDh5lHPpu/5LSY
JYbGY3LmvuNJfyBRspjhdaGYw4DT9AUvluuvF+h3C5jrnZ82Oo9fkX67FoJlh1ML
SCR9/pEEkPkxcVKbpwZsTDJGwIOwkRgjDgcBtIHhqoxTQSRZuWH8s/TWgzYxFKg7
4ubYXNhmvF5pZ22u7amvarRzC7JG9QPpXRR+/mH00ACoRgtpdlG/+Fpp22AL7IYh
AXLQy0jnSXdaHffj1xCCEL6fqH9zX8ibbvPjM81+63jvbIEEHBeJzZFOf/lE2//C
fw5nuMnXtv6Sbj8qbin1h9l8e5KG5GukL8Lpha2AdYFOmhbICTqruZHaJ91erMHH
2ckpJt5/ojFMblZd6xCz0ue5XPJ/GEZbHzC8JNIeaja/F62wnWQKCMvSUm/gNkhO
/A+7ZRpDx+Do1DS77wump9aS5mOlVscQEgNL0DVE+SbxOep/2Cn9r3KDyv/EA1x/
knLBRIafuQTzc5oTSjZ8FpeRr1VYc+6bgFxuqlmOMPwwbJVeBvS4PoPN0gQMzJA4
CQeDaMa5tfHgdoYaP5iVKYWjKX+0HtNMeaw3OBCGI4PaLfJvX3XzPuPboYAOEQxV
HByXCKdyfJ4b6EqoImpG+KTO0yVJLjvJAK8jZwbqcCUgFFSIZIvZO8YyRDTG4Q9p
nXfbLlQunipr2cK3hU24BRsuj1p6wdqGMSOagf2gVgFP1tmbnjxJlHvTN9KpNgkj
76WswFbuKO38AEIkQTs5GmWOs3dkkjGjYs9D7Ve9Oh3w+WiZkCZmj2sswZLRD5te
zEtyvMBKsplGi90x8xgCu/mntfYbfRjJ35SlpD1+D+398A9niQUu/mFZao2I9ywD
1I2Bpx1Zd2wS9XkEsEI8EeSBSoLWZ51CooEXg7Sg5kAH53G/v6KHOVt7BdbGkDxC
JsacgxfaLJhzPsoB4IrTT/ITKtPgXudsTZX4HcQH873GfLsaDhyC+8Q8bTx5UJ+b
kCHEUOzL8Sciyrh1kijOzch3a+lStSwULa/oYKVW85TOiaLm2QvpT/5OTRFXGW+N
JZ485d+nBwaWs9fRMHWapApnBOV9Vo+LJLp3fQBNsOqaVOcs0sIckxrF4DBhB6ay
u6FuFdP/kCvI+V0r0oNI8WOu/f/im7flA9r0MGd33f1d7jmfbJistJItKAvhFK1K
Ruo/JlH/KBzSQaKWP81oDjqwx/T5Lha4DYhlk+0rA9Z22PRPFY7skoZoJZA59S5E
Qku7Nuwv/FwjcVv/knvq2MfL3Y8pGxr62SkMEQDmnvefXKasvkgocJxNnOWk6LNf
clqJfvKWF5edRg4PnpsEE8nO5oPxt2nlJPRWTcZ56TdUui0wdEBeXq5ey3HlA+3C
xQvyAQgUzoq1MyjDZTH9QoQwdcR23q1BnOpxKEtV8BegJCOi/t/Gi1q7NHWYwNwM
wXtFavWCyW8JTOH3ds+C6htxQs/MaH5iHuIdVfwxr/D8K5XaKSD03ybUmUtXXZJk
5R74Oh5PFNaaNC+RM6XFCWTMvx+VNoEVhLd0X2+EoqnjFzRqsyWEwQx6ArgTwD0M
00+5XjLvlOWc50MNxy5uiFy3iKhwsFhkXtv/TJxQncKWTszHr/MWftDRXOAAELXO
bYlVooOO4Qa4ZNx1JPShlHjgTjmOKUOKIuf55EnG10PcaZ/owFneHcuHX6c+/PbK
ToguGa4G8XmZZj/SdqHMSyc50cC0GbYJCmE/nTBH6f1J8WbgyzT6VVSkoaVli4ce
bMGmHW05lI44BT5d91EeZV//FLJJ3AgM3HReEDW/YDrrJYcU7+wweBDwEapEZJNc
FHIvsM3X86Uu0ETA2ueJdw+WFtUDJyFmc4jXsAgsmPTds2H7ikknMXTs3zQv9Vkw
HoqS/o7qJ7zXCwDKizPwThDiLmlAsM3WwR89XTwz7udFbDehNIMw2dz42tZLVttY
Do0puXz6DDB6pnxGRDCEAMEQDUmUo3OA03GXxNauTs+QOI5cBNeGo9P9cbqEbItx
pr47pXuS+h59y0hmV3qOLvg5rF87EWcK60kSyUk70h9EbqrKplpXZJ+64knIyCuN
uPei+09GSXOZGKfQJoTbUuNLD0mXhU548h3rUuO1Cv8PkvosMu5gjP1xKCH1wotN
pmMoTSzHaZ7z+AD2UodeKz3scrsLRR7WfNOyWwCbCW2OXPulvBlONdqDh1HZbI+V
CPqd65IwlorOk4VOyxjvKtpj1IRTr0uWZHRemTjLo1kL5eYNL14IPHl+YpquWttn
fPrRWtgRAtVk1TmGgm9FcciD6+WWHI2zyUlBli0W4dy+bsGVTUQK9YDYZ9stDta2
u8bBXPcrewooVn50yS+ztIpc+mkMr7twlGVNeiz2hOU1Z/DJd0ZB3lj3TRrqB4k2
c2PPDF8tih8nICa5VGe+9OO1vqq6nRxPNwLOOj7x3HAwc8v2aiGm9jES0l1vtuul
cCfSkbyeFtFNxqZkPm7RSZd1M2gKkjJh8UL0qQlK2gJhLQthlaY9E9ZZKtP2JVv9
BWIN6q/XDvLyiZYDiHQMWEy1YE+NW8Mfk36Bv7FXtQWmyVo57ShRNfAIdtI1ProE
9AcnFTs6/91vMDSPi8hW27S7cqaDVbx2bUaC+9CFhzAPCCekf/uJ4wgiHlwTcWyd
5JtAoEueWifCTJGJFN0xLEfjg4HdUMXSDsvLGp9xams2D801ZL8ZEoPkunM5w85y
+C8BAWwrtc5kIT3kDkNzCoGcVBUr+Se+fWAx4j2efr+KPzPa8peFktbG/UldQxJS
UChktt5ONgRj7e+Q92mkStJztkHZY9pU7aqtjmWB2wrMeYgXXPdv6hlXIHXVtiIv
V5DAcmxT8cN3qOBfszIpVdE4/GwaAFoIi4HLJLcJjqWmXkGDMgxZR0TWEh1cWCbj
+9pS7CFlaBoUOgnf6JY7CsoL+AxWrwhiGFADnlfLMv8HymFme/HrQ8Ttws3qfIcU
FXizQ4rTWzK8y5OSV2xQjYXeHhTZh4sQ0HPPge6prQF3YYTEo0Md51M2YCbKvhc4
iN5V9LDH7jxLTWc1eLILCWJhaYggZy9Jmvmx0MAArswGHz0/PzUzXr7kRgL5jYpM
hMiN+mlHTCZUf5JYPEXpAqnF+Me0IWdOFv+6e60+90Ikpec4Zh2CW/zxRAAZFSBp
kArd88xOg8XYNDo+ZZobYS2EOCq5njQnvnI/dB28If+ByUFvnfGqbhCEfQFZqwn2
rRd3xMteF6j8lkvJqCho5KR657n4xDhuOqQCU2/m/LekUKNXPjfayAG7M5IVd85h
slyeGAcaJMicK5ulrTGdldGfGGAfs8ivx3SK6kRBytt7BLlQMPNYD8boNSqPF9pn
Q64N9P4GkQ04q2BQoveM47BD/Xc8h2cW/zEpc88KAEnv4XAbXFakzbt5u5WHlNdj
fbFsA/sm3KJOhgaZnQ9VBYtLNYBEFhv2zVPkXrGd0EtV8jkkiQd9JtUAMO79dIHe
08Y9Fw4EoqDVcoJKVt5J4HLQamAPKtaUZ0vuSjiO8sN8LV17o3B2b1pKyYE59Is8
acCyhlZavO8YL1r0MwNVAfKmAzdUvGvPs0CriyS7iqW+Jb/TGQ/wCJZ57EkDr2RF
abTlf89XJT4I2YBFRIxc0+PIN/j2XUqJKz2nT5S6V1LpKfSoLMkn796UamnQqgbF
vh/ltPBD3xKljbkvHhXyUXfyyOtiXSAycoopaF2wI/r4Qnr/OzUp/wsPD252hFP/
iKNque6CEgCp9tJPDDQBmyGqa36w/twBL189R/H7JvxJO1hYAQHzQn/iYgeAEE/x
L/n65pLS+RkUqVmpL2hjK8ZW/Wn9p7+I1vUXNDrCoFIZ3BxxN3I1EKClcETfbLMf
/DAcaKNMysluVTx3UYd4DVxpq6uRBq+5lVfIfRz3AAV7DLGQkKK6eogRXJZSFxZZ
IFIf3k/DGAOUwrT5XECtsBIc875CPikHAki/ywVagc73xJruIkipgc1CiF5LPrFT
8USsiAlD892gchHFsdRTSmccJfal1Q/xtOkNUuY837Fzug6/Whc1+eo0SnpU9k9P
gdypCvYcqa8CQ3To7bQI0Qw+Vg/fUEiTXuPDJjRlyh8S8hRrmdbdCuUc+OQZ8vtP
p4PdsQM+W1DGC1bV+epqN6vFGvw+V0Dz4zntC1M6QrKWRV20urMSHSXKVBaYMHDI
Jyf6hUM7vT8siT1m4r8FQl3t8bykf5brFZEBX+K2eOpJcY7rAu9O2iNNnG0REjpI
nD5oYhNIJt2p5vhFYSxPyAjluYQlMI1xvwd5h0D2c7pz8HEOZQea2cVsjRf5A2qb
h51iP6CsuFnyLDVeroz2lVO0RaN1DlEf6WziWTqkMO/kmGe51bxyhOm6RmLJfkI4
5M4d2841zqfx657bNEV1YydrmDAZnuMJ5y6o0TGyTKswAvGWIWzpZUk/8LofCB3c
lsrfMYfEdNoCQRFm/JE+AZ/qvCZociDlv4YC9ZnFVqQmIr0fu8qe4oPYLG/7yM4c
GBszF43iIY2cGvVpFh3/Y+mNRItN+z/8oE9MKgy//d/RAlShstOhoN2MGi9AsoJo
8LcG6rxGbYtJ43GX95TkQT7YkNqAKy90vdk8Agcv5/IDEl3D34PSBLcrK/bhkG/a
fDiXoSRqWTpNXM6XLf3E93F+W1yW3sCZmOxFP8e+hY68S4NHsRL11hrkUsC+0h3X
0zQJPtoZoIs4gXlkqhZ3//yVfGb5NpTRu7KH3i/Dlvq0XI3eZ0GtscuCnoAPYplt
OPvONFcnn/1lYhxhpPTYLRYgmkcuTXC3FyQu2U1noPYlNvWbhzSvk+qcwlXLZlH+
CtrW1ABXSJ+7Iv4ie57jrX3xR0/cyi+YTdyWfWRB6BbevDBC4uLpn3M5SYLdWN9m
4NXWxkn2GsZ3zbkTPKOArKKRd9Fz35YbjijPATIrFAlodDekIB4IDJ1KLejTiL6A
LpWMXjy6n6+4fE7pV/+82HHuyjtG7Tdswk9qFYTPOcVvAH2Ww0dLUU7G733UgOAf
ASKcsNPH+98BBfSc68ZD1ihelSBDHlKVYmJY8QQEZnnpaaZbwFxt9b19YYYUjXto
kljJCoftbzb3miIM+hstUU5nIZEmWdCgcI6QB4D0Nq3UrKhQRpw984CNqi7DroHa
6KyvPPsh684GbxJ+RaNkXWIzvQlOkfMNMwuwz5UAnOCi19LzF1eigcnMW/YXu0oP
3IDE8P/WWFYtHfrBF7pF1167I7zqeeZy1ryPGPr6Vgpv51FQp4aot2vW668+hyBO
qNKDIWTZfHJBO/lEITXN99m8FcKgOmopUwLA/UUNdLxeNBP6N6qO32MoqbK0hz7J
+4nUFTlTgGI8yyUGgF5kaF0sTHGh2lkgiHdHDcUFo62xByWyD3SzUSVCG/E/sN8l
huW3ePNhR4fVPf5QVLeyZMLwKFzvhPZqL2XUd+WjV6fztCtHwQaXjmGJEaO0EJ6h
tIIYcpRov3f9VFvBluA9l7N3oM+ZColwZecXm5Rcl9VWtGVk+1YaRxuyVJ5ukiZF
foT7v5U3XN1m08jVMCabNiMdMp+svXTa2BcB1rVcEnIx5o7m7Y72NcPpHAtRpQbo
hoYWCvgNpScrtPc0BuxX7UBVjBnANYcHoDRAlwsRl72qY4Ug33ovoopadrbDjV+p
OrPRjzXlwGzAHR8D2lx1XfyTHRbOf9vgGGEmL1y7J/iMU/MaANp0hSWTiQicUGLF
zfUlsWK7tyejxgOmLoP7GEz60w+XkrMwYK3adnBGsckfUlINGWlEirzyPPhYAhGb
IGnE8g48eQpp3429cUjQeJA+S6hdMDC+QDAk0hJgPjGzAgePKT6mFNnGcILYrTnW
IpgaAppJ+KGGFIjlHYlxJKCcgiwfyaPrtWSzVTgQTO/k6CRDfO1ERfIC2q0wjxVN
5YxjbOpw5L+Rbi9HchF/sagsRUnqNULcV9Kjzks79IhCTmJQbQlTRTk2kwgZh10L
MBprPOsDEBLveEc68FACcTkant4dX5oSdx9qRR9QmHJUgFeXW+f3PaWgbjywBSLr
lv6mTQeayfMOp4Z6TUuyhOqyN39/zT2BHOF9hGMcILpvV0S4Gfobp57Z0TkB6FLc
j2G73eZRIlEACAAOEViLM5Dy7jxS7mnXNH0MvCi+MyfAaODOTz3UbwL2R+eDrRSK
zFZnf1GS3vgm1aVnWIqvPJuFGQItUJAVTE9uEAX9P1p/ZDhfchwhjlDo9aVoudtg
9V9YGnZk6tFTilVl4qkp+MVON6GKkUddOLumC3FE6ff4hr6jEQ93Ot/GwFw4rCGZ
kaGPrwUXefsXIpLxpHZdC3kE7Ku55mVVzffWF0rc5jefSwXk8YJTWwtsEvXpjiEP
diJx7MnG/kmEtDp7CIUQ30XSs3GaoyG1yjWNOV2QtldS7eouVxPUs18qN7bc5BWq
fABD4mJcg5KqwR5lLwSHMpW5mCqM2Jf9scG5kbAyVD/S7fGhAF700tN1x2ZHbxIL
w5uwkukQWy/0+AhNStV5qTaBXrAZuNwjRl2yBNmWm4cyigVWZPNspn035Cp2F9ND
e8VBoIhJM9qUGGo0BLcCgeovCPPU6ADhG9nZsQoWFa/itfb/qNHOANuFgujwaAtx
fUmdz8XR7a+Zopu+JAJ1G297emsnQPb4bIxRLQCD/jJ1Abp5csn8ahSbhaKJZKFZ
zSixJmmF+RGQKsX/Tld77yRheAP5VQt5DMS7V9bxhOgZuhqd8M0Ib2p/584/Mi+V
0vvwCxhikmJWyl0A8v7OVp4g4N9SijkYKcFoZTUl5pDHzbstTVzl9Qo+k/p0r8FB
TPt6meX/tFLcl4rih8p3oxTMXGjs9YHqzA0tNcuhkJ4VdYAPQ/Ck1LIH1stIpILh
JcnoUBiLMxXrON3yPU8KVBzfnNBeYIxp0yd/UqrUeZTDO7MBDva/NH4m2kSJO+5a
avLN7sMof4ICc1acxgFZdYy8Q7iks4yFeCky1WhJT84uDiaQxyygOhocLioeZe7f
iMujirUElLgsf/Nh7iFbAbW/B3w+H3smtYWYB2+mZ04QOUe7BXUjvQJOmoMJ6u8d
9O14mCTxJEPgGrX3W8AWVfh9A30Z9x0fKTw5izG2h8f3lA5D5vi3wtudVh8WRI4R
69ryA2+KQrf2TcRtDutJc+OUrbNHbodwK2HFydMD4Tz7DC5ST6Ev88mGL/r8XDYz
7EyJn6j8DVLj0oYa9PDRGh7Y7jJCGGzt7ya4oaiv3w3Vvq1ipm1nyvc2tic2WVRK
4Ub7B2oI9qdB6viTYeXgH+FblCnpYN11N3g9FjXxr0aQQWK5Ji6BJRVvaEOxP+M/
rNi+YjWw9+i3pyw6GDBzRucEYMDftfgIK/bW+eGi42vZJ/M8JA5a5Lg6KwzU8Jzd
nfwKe8Fga8BNHLSggRnBCGaul4Mcltnl8gXkXIChHIrV4fcw4LADcDX1S2T33+/E
bUG20onBZvSbnknIbOARiF/CJ6cNODX/WRW5vKiNjhGoDf8a8ekVe25W4cFML+Q2
cvOb52MjaGIySgN4Bs4cg0HqN8otL8Mr1jNRcuUd2Y/BH0WWtq+ZwXSbU3tQaGoR
FZiVdJr1kCsXWh0rxGYBnpcI354F82pHtHy0mknZaRITyjXNdu/uhaif1nGLD2B/
1Pf3DeuynxVBNHi1i3Cnt1X5ZQGpA5WFG/kLpylVPt/kNjUD3nAOAxVD8UxBi7jh
C0Ety935SrOJ42566J2FbS/KWeK+Rzuo21gfAd6/rtsM7UJrREAZOAXWH/nnfdve
DOKeVLsDfZ2Z9rE+YE2gWoDNcaM4RZxa+Rz6mhCFEAKcctsn6hC1tQoS2SFaZ95S
4CpT+tnNJtRo6JVIT1hqR46BYQ8EHFyLC+sEYcZTNoQddAHOAv46hfoiRdw78dSV
y7tavfvyqV5XvA5ucrBJIYPFfXBZX9HoV4PPANHiMwBIAMW9BBwkezcaKUCTT8aA
fgS1eJOoukxvY21OBY8OBwamEHEYEvQVkJNcr1XhhBSfYMp+T+2uaZ6JVTJI3XOV
JxY6bYh4c8JXsRYdwerXYZnm5nRDudm0e5fFvij1Th1y2bMSUEyEV6ANToU6enR2
o3B+W6f32NIX5RsGggiyhpXia0R5cbd9FOaT/ncCZgd8zzCTEB1H2eYvODz2TftG
i6rPTPZEws7dz1Wzz4PX4M18BaMF0gerAExCKoQlDJoUIH7u+MRyZUtP2R3erJFu
mXBg0rXGc5PWpjoftdlw0ZzHc+BxZhjseybq+7xM6iBLya+ieSrcc/mQP8uPWvKB
Y7MzeN6MiV/jEqqmZ98kEs48xWzRT/Mhg1d2gpUZ2duF06slmwfT7TjTSeeHkBv/
yThNtXY8oyRr6nZtt6o7Hilt1e+3PE42KyyMOoQpH5oW1z4WC8DR7HNs+nhRe5SL
8XijzC/2YoZD9xta7nnEcYCGY1SJItQRwTIITc+wVzr0BVnrC/KVLVFH/ctTTx/A
2tKNV4D3IdaW72kkoZxOdtPKLXRhrNKA/zHBipDfBxTdKZtqgPdb9EYnd/p/jaPA
W9k1mFq+GpK7C0rYDZ0q2PjIdE0ZNrB5jOzn3e7qI9tzYAjiinrEdffSW5idaDzo
yaBTns8aIkuLNEOJw3JFgh+g+1OcYXMIBiVI5pepEbqq5pjAvyjOwpUyMSyfV28L
WIL3uaEVcmeiypHYOlAe7XNunHWmXlbqPe/2hCXAFgVuJuS0hhVkL6URtZBgZ3yy
aXF7mhu/Nsjxv6RSwJqTycXpieQBj3IDPvUSKQzsAqOF6M2EjDJeJGYlQZCAfVVh
jM+8+h6k0gghT54VU5xvX0+0ZLbL6k1GUfF3Iz8Xk1do38pZlF0HocHZ7btIGUcc
bGsmi7D/jXgP3LTvD+/eMYeCwQNHufuJC22hiSeHq7KRMfdmhejCiaHGsYss9bIq
20PeNNVVZQ+DLQ/9NUGDKSOmi2XlAXTRZDwOnX/wbeVn1HToe6OXGFRvzmiKo+iz
ik0CwbLVrjUDbXtPSUFb4zxssRGR3xsP2KJ5l7a/E48o+bqwBx2rphAjBsvhoe+B
OE/TFxZ40W2DNuYCechZeAA3bqemxj/xC4xMDF3BffZyH1bTEMs6JRM3oB2huOGL
S/3vsDtqMXhUru7ntykn8bgUpOqIm4EWDoE5EdknwNBb5X2te6v9Pt+1Oz4HYbH+
5RY4utsdmHXcSx3Plra8dwznxejMbSqxBzt7Ys3KMTCPFDJBxy5+I0fLPkewNuxd
UKibByFiFVhdkWIxq3ikOoVj+55dfbKV0lTfJfD6zeP7JBRQrddnCTmW2t0dzEnB
3ddwMDFIEj2MlK32IJCtSGSEYYSFFfzYWB91l8rnz5urt3W1VdQF5JrP65lcbSfF
L7S8VFtRJfWwiI6uPtE+vW6e7cZ/J+SoDHDvv5aLG801kB3HbbXw2DRsPk4QJn3C
n8hPKJvI5pwYWiwkLqmC0JdpEBwLrxv5BItoRr6AZPWz0lDKYdppjp81DeTPA9zl
HM9pPyIp/BtKNP1v1lWQUvTQDrmi/oX5vWOibaHX3WNmfXxgRCvh/0oRxg4cEqaf
9sfZCNYOpj2iVvJCG5ITaM7XmLH9h1TydeEUjvH74UVb/B+KZeI4Fcy+8tTxeEx3
ZCfrk0WsW3KhFkAlvX27gQLjWU5+jK/YcUl6ahLrsSmrFTcuKUQq2ghx53XhP3Dn
SUIVC5nZLuS4pvaWC7OJNDkJQlgwSsdLshqC7bMldooTbYA0xUmdvBtW+LYbhmrD
lg9te/R/gy7qnYNBrZs24WhuQQNpwnkNuZrFCpx2cTrpDbHcMWQT2fRhGi9P0LaS
dCy+tFoAFEY223p7ZTE8m7ie2U73BKZkyjBpAgoiLMhn2kq/11UT00lEhuDrZ4MO
wXr48LLGO4vZ5RgR7f2kimhzyKK9FZmO13F5L0nlERNGDlbOYZfomug7XF7J1ytp
rnr6NcPw6dk2WXr8ecNnOh8hc604QPG8yfu6RtsqYH3OVD82sJ98cwZio6Z91KSR
Qch3/TXLt0Fb8/rzvD7EgiG86sYJsGFHwerUVPEjSYHSKf/QE9oaHLECphLw4MyN
LmhOmtIJoDHO+AZEUJx78Qs0gM32HIX21/t/dMz0fI9ZpOK4UVMhWfkF5lRmvKbS
d+zBkUYZlrtSElm3Zp0KCr0awB9UsdB8vPfo4Sxs3SonTX71Q92TZqjW9WJ2ITkk
DvmwmiyXcxit0YXq6l30OAv60CH8UpPzBBvApAyrbyPvJid09TGf6hGS7//wS6SV
tR2q6RMnr4QY2aeHSdn0/e45vATULZhWFC5RQpXiHmjoR14XptssNhkwUNI9FRff
hO0sizemHXFDK/lLPr9kTtJljcXrsVAX5Ye0PdZBS9jDD2Fer5HfWDpplv/j5kVO
1xKWYn5+t/8j/74ugX8phDTDKbtNdd7i7DbHgQO8GJLGT/ANmhgFExZHaEVvfzA0
/ZvIAPU2fRDfB5YS32WfjHAL90RyUzkk7u2BHDTxH1Y9nlxHwUIh9YrlDbzzNXQ9
2oSmiZCXDWOW52KAVD9rEhAuCyzE9o5DLOJFH0MdLAsEJQ9t4GjHVqeSJcBsWMTK
wLDsqiLhBl85GE4vnzDDMsS1vDPo9NiW8cXlpiv+rTI5MhwFayzne4PZONV8KLTS
XkEWtatoMPdmQc+Jv+wW4CT6ygdjIDPRlWtOje+y/Cz5bVAJTI/LKlpRaOHWwMIg
87/5WiZ/6/EtAc4pNVtuPC7Lq1u0C04lSvq2za9drWD6jEj663vckSxnfkPqEUT3
sG4+ekEtaNbFF5g7FYbwq7mRY7FCx8jEhlF080Br4pUn0DZPhk8HqOQ+6rSvKfnl
ulyrGafr8/Vr9oN7KuDxQK20Qw9sHS0Ip4x0E5lJts9sowc6LBXzVUFVtl8tOQv8
XHfK5iCflR2NqhM1qqW0SQkQv2mUeKFtC1xcbd7mPGtJViQQNid1p0zZ2UZAU2tU
8gfebGvCnUJ8VYxuWa2DEussAO9xAuPkFqg/s6YivWw=
`protect END_PROTECTED
