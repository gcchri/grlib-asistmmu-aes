`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jdqky0IxWAAnfFC03d8V8ZNyTTAOnWX2LPxAc7XuWI2NxIB1ZA1NRUpaHM+rdwsE
cBfvl4OZKxSV6pry+b5jYS8kwgcZW2PHqLKjPA6q1KdnXCi/ANZV6NCMmQGaO3zI
TLzx4/1dbKpXMSP92ldSSkeS1HW0MuZRGvF+/UEfKH8rWGpz1DE+Hxv1j3L9ttqk
vbB3zAZejOdfjOBMcOCVywc4zTT5WO3QsEkJHf4jAfHHqezOXXhsR9j8jKxEOkO1
2bzIk/kGj0EyJ3FxqQmNXKf1hERz97ETG286t6FdjPP+q11sMJOeXg6PnHpRVwgo
VBaRYbFMhRnRfs5v/746oGOvFgDS4dRa91Ifk2OpaNJ1bkP3fPelpRw6HB18orSl
zIbLO21yt3psKR4lGiT9Lg==
`protect END_PROTECTED
