`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UbVJTg/mzOvuwhyNhkloJdyDI1OWKRKEBDOBFOnyNmRGsoD71maSE+q+ltAlwQaq
Nn283mV8uZjbxxtpo7mhroz1JCmNxJcBsDNOlWQhlfQ2E1uLVp87sut6/RvFSLxX
Z/D30t9c3Vvdc5Fua/9EfKI2MvPyUQtD3JfdxBSAJjhUMgIAnNp/y7tU5LFET6n4
p1wcI1b2yv3EUj8nHQU3QAfFeT6dybM8vHguY/eirdUxlzWqOkb3CUZ10lpGwAqM
1ZKFauX7aCbv3H6qpdwJ+Zc9bvyTDw1sLdArvNigNjRNYIaGvbfG69ISeLEkS/Ck
pTP0hSIVS49/8CuYC2PD6KQsNy9GUYzec1VtEcXW2i26+ctyiR5Y4BHFG4tkkMFv
yNyp6DX+IXGU8HGsXk2GawUsHQXMWmn9MnSNPvlAu6BEAml/ZKvjjgrd7KArDW4j
EGppH2YofwP9qpkDB0whi+yxfP65dl6SWykcsjMrZrMZRQaNBNAtmPEXJ1wf3r09
A37Tv5WFo0n4vUT0MDx1L5e6hZC3FjLj3eZ4pwXktuVjg1TrnrUki5cZ7N1gyzVr
aOp3HJt+XMEf9mlY2xIdUdO08pHKrp0sGjt5Gdq+fHm5aXwU3MTzn+q8Vw5FTRlu
4MYrwjQ1wwJuCmDuc2xVVthXgMw3llkiCwxWFZ7MZeYg+6WKsTXxbYMKKWhQ/NGX
o9Tw5XYqzidpCHrmjaOMszeOn2OrncXtogWVJuKebJ2N4jvStR5ckaz73G3O3TtV
XzgcjdBn6xhbT9JY5fUjQ3cDZ0M8OvFdTBEGpJD+8u54GfpHhJVBSzEyx9MGbFko
0p4LlvBpp64AIuklO/bYLkGjXudTMAdtEasPCgrbDpSp3E3ErRr8+8pRqpDQ8IEX
RDwSDTgZqGHgjab+TNlDRL6hOc2pIMHFSmJC7xfI9C6TFkB0mMHLrhRlie4v9bpC
`protect END_PROTECTED
