`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZhOJlfBarxkQoA0XM49CmFi6diuZyD+0xstrZIlOvhGVFuYti3zOSEzevmW3eIiS
6NVACtRd5Jq/rv94QyddbHoT2s/Py1EorypuKue75gL2mIZLDQiqT/Ey0kdkDCUP
4YJ37p5Gj2Tmkkn2xeigQIOw4Y92wB8UyKq7CopTeDUuZZSwHjC5TrBzm6Oe4FER
uA65UJl7KwmZNxrEBr8mzPyeDpbqwh3HEqBCq542udgm5Srxa7Pr5AVgd4DL/ck8
t8PVuF/9Hb86KZzVLzmAQ/wmFzYWHa3NnG1bCgAI8t5gSSMkaGnEDwtXCG55j2gu
d/RHP4HLg6C1ulwdPEAW/96MOp2Gcqp9bwO5L/eYI8n9O5v0ue25C83dUeQOjZMQ
a+PyfCDYPyADvqgYKGnUAgW0c1+mmzQYHUmgu6gUYPWvwHAi1Wr9T82uTYLNnCBQ
siRhYXV2G0y0EOuZsJxw26j8kktFPZaNFfezWJ4C/eI=
`protect END_PROTECTED
