`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2S1wGTE7TBEDCk0rti5UkF7OC6wREi1KAnIQthnWBf5xItP5/afJ73SrrouqFQzh
Ox2gYdrHoHMNQE7SIT4SGE/SCyJXmBNE/bkVUeDDYVnY9lthwriODfW8+ndsEysD
zeY+VG0/ej9eQDOIskALxtLZ0PzYYTYEWn5zy5ktsS9kHI37jAFK9jk68PpFNWGt
8YQu1c/h+rGUkVt3oCkAyKvv1z+A7cxnxL7XNH8v7u6ucvsyEDzG6CKBYcY5kht6
H6fG2u4pq1iXQIrPTjpA0BIq45aDwKL03++DxVxPB1AMiV+ndlneS08vXdJhko07
hvZncHg6PXUXaMsqIZIBOsLm2wzb5qeTO5CcUK532Iu7aX4xTtexBUn5HTMRm4F3
Bnq1OgaC9n4NKWO/8mxGYlkyXsh6P4OriuNXJzHWR2yEeAywaUkKyLPa5KnNniir
+JNPw1MJG+GtKMym2n0sQsm+J/Pgiae4eOgSrqplIzF43jBr4oXJiORnHOBhshBd
Q5bhqmgldUYZxj/RnjDluivY/qm+5jzBjGaa+Z0EiOvambUyyaXAShmTgFilQjmC
YWnVbIecV94XnYvy4P89SeAk45vDH+rcCyntwoaGv3c=
`protect END_PROTECTED
