`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qtERNh6Qu88pyJMTJeWRlyFNnWqGODaTr6d2sXMlx6q55I4pi+eYVPxzhnLfXQ1v
ZzICn0e14jyeMo5/zVsDn9T+lb96H9caDZnnuf03E8oTHOKLZGffSo3VdVhc0SKk
dF9nHqb5gbBuu4RbBtNPKon1+Y55dSHv14D38UN7h+FnjkFZrdkwY7cgZ0AFfcop
ox/qy85Lbl3mIWaQWrlKQV+J0FZ2v+Xwuci5YqqrH3ucVCOptxXS1PWdDh0ozXmz
CYa5xFMt1T3u33C9VrTLCQiM/6B5IAF4wZH8jVP67jFQQUvQwhcJ1owyYv70Z20t
NmUXlJe+bz4zJoi6KPlriGR2Vt6rM3TZyvSLKmoHmcdpo7gAmtXdZ4hvNDFUlJa4
l8PLxPwzTa/IBAbLsUWA+fBqCOlKnRid1ZmS3hEY3rb6bZRXWoGnXXwvj/tZklsk
BVpcN7fehS65SMhz4phT0657eYLSMhfrIjfQYtgELSF2BB80pGJiqTenBJhTHSJS
`protect END_PROTECTED
