`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W5FS/88Qs5z1l2AANXQ4HCw4djLTzjrDKOzuyYsf1UQRBaFqtVYR7QZXuh3I+zc9
mJUsVwPpUGQ0izSDuWje/WtyqOy/PbUdFQK4A6XBqyFRUzP3swgH2YqsWrhmTQge
ZgYjHA6E+Lo5PXT635FxyvGziHGNNoUMdrvmpabmCA2cS82djFeVZyxZweJMWrXW
IGZVeReIvcjA5myESSfUj08NkuXlcCaFR+Z6b7/1eiuMHZDwEjhdk4T7TWI2fOf8
fYATZO35TFQj/Wf4N3EEQRog9uhnEUaPuGvlDAjDuIfUW2fE1sEsBe1zW2GtCSb0
qIn9q8gQ83eW9els2Hw1jVlzS3WV6PPxUDXb2dNle0cwkZu4bYTbK/u97Uy273LF
vmU+1dtFG7V48tPmT9xk3jozv/jL8YLipqgSa/hhlDV+QtftJhVL8Gb04zBBFWug
J93WcVVzUG75l8Wxw6cCfcy/am46cYgDgxS+8xUzuiOlE0azXoZQG3tCm5IJgrjv
l9moWobphps1frUhuswPF4oaqQH+ADgkScSD9bpRAkUuyRj9yuBtkD362HsxZ00d
FqEMq3lT66lGbfkPjA7ihJfI7K4wYatFg9ZMoVxr5ryVdSWeNssfFL45s3X3YzvO
srOQd5ce6zNQnj+0e4HaB68Ff69lhsghqgi7Squoe7zUUQ2HSptySAzL41DoN6Ix
fxs2cDiJYdMtECOd9Wss8lCU814WYIuqvsOLJAC38naq60aXAKCd1XOvKzFIWxbF
nr6CsTz9ZN15MVtBBI1PnU6TM//mRBqDmS6CeJvjrgvFv5MD6YymfjUyVbwLc4Gt
en87f5vbm8kf9ch91YP3pF/48vkbF1aVdbwofv83CUgxHCWC/UhW+lzEy8gk8N/e
XmrNrskxwLIV/vPisxS9h1mTpRkCeDvN2PJ4+J0Swjxyud2tcrXuvS4zUbsl8Tpq
AgZzNmpPEy+plAYY+F124YDqLJd0r1njrQcKOKrYm4DFds8b9wdrZMZtecvAkj3m
KK5NWL8/vStlAx+clazY4rFmTzsckkVw78PcJBlAYJRQ868TevVdohnJOxZj1IsZ
HuPzFw8bu/zemNfroSSHwOQvUs9dMMzBxLJ9D/SUB18SczpRl/uJy4nDYrFRTRWu
e55zO8neE+eLga2dcWZbh4Us8uObfIkx1KyLhrd2F809ya1Z63h0IGNxCRINl4F/
qQHH9564wtN6Ma+zK5V6n6TxT3YH4YKkcsVCN7rwjg2F7x1gRgIOMzywqthhzXsA
mYJxs1QtXugG1plvLN+0eNP5Rsr2ZsQoAebfkK9uiyTW2Ro2R89v+CuQTRegQZlz
+YFpx/kKQseXPHa9ceKoV01Xb19pLY/uKUfGroEISA4Xz+ePNXQfvHPGmNXCMD5/
Kv5Xl5Krv8TsK5HChvC3NAWsUOkImiTn1VLQsx4nLBY5Yqc8E/nRk0n6MKpPNo/B
M2Q+ArmDOrhx4Fm2Vb2lV2oBAzdQ/x7KG/bYzB8zgTefS/25rJVdL8yK/w2504gu
vSJPXBd1PgnQMULB+vA4eAERHZIQdDO3VI3c7Qh9drLpZx1dVUIMZK6OyDGxfTK1
RVa5CsHe28RJhnDx+ohyqbbmZnfJAIqN91i1muf1ExkQ/3B8Sn3dv9dEU3iOsDBi
lgLcX2BzXznn8gKUEF4+gbwPJhXAAeegBfDBVb4YfRo3BrmJG46aDE/V9XJyR3C3
GATbNRB+hJgFwFR8tVr/AZxMWTIyb2x+tcesnYCyXoFtc91/03QZdpo8L81GTfbu
e32x00gkwX11O1FzNqduK9x8EUkDzovGwWzwETXR8WWdA52KM2LXTKm4eDIv0B7p
xPlnXrGDvJsRzmfckYzMQKPZHWNnfY8Yc8eOHG7VVt0CqTS3mGkBNaZFFEDK+2re
5Ci9xptAd4hQH2yoJVBxloWfL+8//qBWd4r1FvoXOD/OjDbF7Ee26+ZOlRdOqVzQ
bZLLiDgObwI6PKoOZ7c09jZXfFKjdGA9FHGH2je/T+tfvampjIw9tbK+KB+jMsv0
hCjrC6/wLYLxZgpWtZucUdJlwzZDgymVN/Bkbxs/yeaRhRgbjxy1dJJFkJEIq8xV
J1b56QdCU2o4IrKrVQJqw6+WyI4WDSdSjdXpTR9NBDrF3SK/KheJX+93nQzC8XO4
/RrtWVnXMRNO29r8cNEMxwH2dB0H6GnG/jKZTq11G15SL5cobtLtn+XiL028Kv82
ClpPpPWMMtu/NoW7utmjSJgt5ifCME7/qJ9tK9NwtYFzVRqbbS8I8ODdLRPSmz6Q
s2z6yb9m3F82VGZdp4H3POGL+vbMNrZnzvQ9qSf1K4oNWXVD/ldmbbDkYQPki1eu
YvJoEufyOnV3d5w+ezo0EzaLE1w67w1ytE0Z8MGlhX0PkWyS0rM+r+/9o1Ipp+Ut
6BbuAATAEJAtkdhUxXfag70xmE1FKGyQILIHvS5DRJsDBKNOr6xr8QqZqirpOYB8
c1M5o+gDXvM7XtXSiGj8WmiKTuuznOy/XIzQm2RpeORhsis1cENjJVxJu7KsZq0Y
s5TW1MJ9cAVG0FkTpFVqZxF7f465d7dxgzR6fi6+SfzU42UxGp7TCQdVioCLmSoM
TqY2W+a70Fbxk0S3gxNtDOCWY/7oL9TyCJfW5IU70SpiT+q6+OSzpltoxSEjkqaL
YsJrcVLR62BcW7x5Ug3TzaA+JUwnvfHBz+Rl8Bbr9xLTnwUe5rukWwLyL+KICJ1r
C4n0ZnpF7iCs5VbAToQgK94xGL4c+ErAnt9HQHKL+csKtEblhkUOO8jCAKaylF+B
TzPTtU7OpY0Z6Hd+w9AtalCSpfWICIK5aB7F/u/YqNDH3mHa3iI3ID0BMlAEGIW3
kg1a8mREYQzdMafNO8F42nXWVc0WkXFgigHTAkepHRj93vSYEdz5qFpcQnxAV5FI
pVtK2xfvHJ3jW8Hi/8ttVz63UbGSlm+72tTHe2ZKkRc/763yKidI/9X3PqrkiCWm
az9oNv5DV2gmGN+IW4GKzDTyJFckInCmXHfQCo1w9CnaJlqzYH+vC5HfouMUoric
Y89vIP8uayXQ+OC9LzF82eR8hJPuB2mTGm3ZXLt58StJny4rTFDVnisnVEqGmeWP
kuXYDo6sS7EtLFHhSG0LlgNHgdHGMSmXRF6IsiADHnVZq1FoGluniTJ2vM+yb0PA
P3bXUL7fySytde+bDXPH+EU/vq5MUYW5FeWog9YL8PKlsvwZp2PcuCzW/z+CBOZo
kuLo7LHkzYqvUWR8Oe7xoHAVpGaeYzwnnuDgohvyXqvlDEC7zr3bo3kAlAkjT30o
Y0stOn8OZcl8DlWpruVfW7xwaAPBJfLBqpUjcGm8DRnjDrYW5Ag9AJZKfkXHKWGr
KJH1DdkvUV1xrcPrAehR6KSrmG0rT1LN46JhBWQOjOlEYSgd79x9J9jOF3oTzwcr
nmdfLe8GzhbWgWbr8oZWldRgEFVdjskTIqgwO5yD00GdBDGiQtzI9sw3z1ctlALb
NQvEvVwHfGvnW5w1pVM/trOpznHXs4+s0i+tnuOoARfCZGeKYN/UKE0aP/xsgmwv
r78oQG3nqV4L5jrrP3V8VMGkgYp3folLF822lfHtR8J3WVI5nAgOWInPe4CFY52c
7JZl7fd03q61XCI8MHbQEJFxUD4kAKKFGeEKHhCTRzUqXZed3gUwSKiZbOymHUUV
MZuWaySajwPU4QHS16V2yz2S6ammLEVzL9myQ0tE7VW44aQMBub8/WdrES0NQpTy
/p8u3wlH4upYlgbzELFtWykOHT/v+lnFgjkmaawDpCBe507c4z/9e0NKw91kJcuq
bfI7SBED7idKpZz7d7fmHKA/6w5dGvwkqC2z8LTwGELjL/GHAwwOZf1fNYebCxbe
FkrE+SG6LYT27NfpH8vumWo3XGuTxejBjB8AoK1HY+l6Iu3YLTyAs8FoyA/scZYB
DjaXWSyUd4yjSWA+/Ipyob0NXIPis6utKxUZra7sF6sqZjjFfY8HEPYV0kBsS/bR
sG5ourlAnRquixGpkZj/J4PoNprb5kIZ8Qx+PIc8dMCtNua5+owoi/Im7RqDmdOD
vjOQYGkDp4aEuYyIwuyfvyOhs61h1Io70ZxL5y2PmiGRQdMljkJaYVt3P7igh9Rc
NA9s3vX0uQoH8T+NgbAct0A5qfzbafqNDfWEhIfLOGH600v6K/Kei8wdGLJRqC0L
4QeFzyDqekV5e63zsuoKmi0BrcSLiipUXw8S4VpfCJLAwReMIJsZBTBwDyJUhdlf
4W+VH5BE/MHIYwRIYp395oD9acD89GOy4k0e1tLUSovuoq1yKwTGg0IP+Yneiv2z
E0L2vRkg2ozZ9+g4my9g2KUhf5BKY8mGeDSEw/eHpKsk2PUlE4I2ahNlVVT3woMu
a1PVJebCWhx8w35Hp+HDnZeZs873YrDt5eupiY35KgJpbLll8RYLLNFvHgadi76D
81X3in5kgluls4ogTRke/dvS+qBTO+n8C98g6DJilFEtg9d0MJOv5H0QXWeBcuV+
CjYNE+e+XlO+z6t/j7kyRgzfc7Ec6BXxvBUSb07WpE5sipd5OHwuhPr6nvmGcSiG
gxYcX4GqzC8PV6Lb/sbrKdTIYHKuUJ0YFc2UzFTo7KjAdjZaMZhOzCcmz8WjghpW
l9d8P6VLvE10O4Q7lERDtD+a0INPYXSPCrrsP1Sz3BQOrGpAzZNxNLTnKHy2G6P8
t4LYHhs2dVwtRTiqinRGVuEhrN0qyxJAIcNdpzGuo6JXodjEGcYRj5UpODGeOe6x
yfp5lawjRKCkRxL7wy8eNH+84WoVDpc7K6CU8IBF7mkWEpZOGmdl5k7CnxU5ybiK
qgxCBcG11Zefu0U1LLxurwOoLAqAqhLtLmoZAC7CBRF5HwbihH3RjSEL+DDeBJ1z
7iFfzjRy722mlEyMJVLkKpFq/3MTJT3VT3n5YtAlHY8SAhA6ZmHtXgzW6IZdjXfn
D71qsj4kfYELxMZji9Az6TulYguhz3Q9VULsOlxOGqbWwObwSyP2LzxX9RgPh3GH
kJ/ybp1r7WbhOAZOxmDIJTBx6xclKyXqTSLyfUsRlKVuI6gCcs/CPvWg3kTdKU/j
e2s3V33T/hrNKCq3Jxmirw2nyHttYMFyshQZPLHJsynfzLIkkdio2TMMPhepeUed
U/1gJI3xqfzNoCHeqA1+06sn5ixGxpwodX4wOd0c0mJNeJ16Y5BWzCmaW1CYnl+b
9NF7GUsmaB/X5/Qe5q1FAmShUxGeLcEX5AyWygfnJASZY0h6jxeZiCwQuEsJ2lZg
FXstGqTJWAm5dQj/MCmRESw7Uap2KR4YiOVspE+xzJbWRYKSiFmtBrYwFVkCqp0V
bwGt4EH11W4OoALGkjgVWWCu29cbT+szNHiPmDOrX2QABAWJlFHVoHCzxmOn5a9i
FzqGJrrUaJ1fi4MK52N5PCLMMqUIbeIy4Ps/hfsEBSM5S65QkQy4haa4JLq2mh4L
d9nXNbl9Tl3nLyR2J1FoYhevcWkao8GOFi8n0xhpvvjMwNM7ZcUFHpNxVLGY+vGj
ZVwNmysCjN9QWSE++PO59ZUQlcuLjt/0/Oi1UHun65RmZ3zRvmR0pi8FJNaqTtuS
4le8M0T1uDq3wok8qfvD+otoSDX5FL4aKJE75OfS/gEuZCliYp3yd0elC5aq5RPE
En4okXFYnSDn75BMt5KFnmmlWOBg7H4FiyKX/u8ynoZAi/8LAMWxlLQRfyBI9Bnf
qFWHvDhc+EQ9/O86V6+h6A1O0t5lb4rM3bxslxsm9ryy/2m4elQkqfwNSFpnASgr
g2KZFUOpNW/mGRUS/GFDueBuVrop7qqbJnGamVCxh4cyhEkn2+QD/OIYJ3kB9BU4
hivWMB6pEwOjsqOaSPLeuqIhsKMPLd5GI507pTxwSrdjaRPwlyCaO3p7s4SAsWPe
ALoRPEAMA0tdMWOARgtogKsFosA6flwFF8pcR+myAsbJL9lcG8VbUACJyMR8pKBm
W85HOTa67e6wNzTkEZChCLdG/GA/WiamZVwr5YqpxijBt5I2+kVOhKPZ9dA1Z+z6
vTTpMGrpljPXRZNWhZ6q/Yk56r2/kHeun8788evxb7qkD7aoEuUza/7Eekssr/x0
JtB/Ydn9f8fy/gS+rT+IpycPrDHuie0G0FmbfxiOUeClWo+WYXEuQ6E2THyqWXxq
AFMTfAu9ZdFHpgEdlxBrVjPQUwMsvu5RkVvYZSV1OWDG27Zmua1VC+z48A5XAp9j
khnebYDG4msU+ZvzX8MquEE+UDkbukeW6EV+WB3wplilnngwKI31sKkzikCmJPAG
/GMbBIpuAvPX4T993EgsUq1tDjIpIZqKbCib5lB2Bm32PmP9r6BWE0tEO7rZSbbW
11dU/ew9giw+3kU+8E+71heahl4WQQB12I16UPj9NeXbRmrQJeCIVLh4jsFh1XVX
isOhMa2gPnquLBwNzrKHbw07sTA2GeEjxUNu1jkUH7aKsZevpIu0SU8a4J6Jb+Ng
TWcRECF5IgcYDHMwCXAVKsYO5LYPH9t7lzDSfCSeDdp0N5boaxO0pJ9G9qBaqAFz
g097yzt2i483R6vQgcE6XAvuMvoZoyumFj7HZnA+d11MISFe17X2Gn58nVsKDm/C
0AAKuN6LDtzs59O6zigILpP2huc7dyHoLu/19nIgVY8hMTCoLgI7daxy+quXZWI3
hjnjqpeWKgPDv0JD0vKZ4UOLXOrI849kDJ74q4jLcVGx4RRI9JULyEYRlaOhRTJg
banue7e/ZyzIBs0O3Ifa8MHiBoYhn5aoVMB1R7n/eQg49Cntq8wWM4+XuUtLczzE
KNryhhNN2ePU4mSdCwWJcLloQHN8J+3i2sOgSJTIjZQ8+L55lf1FvgFxGC2Rmwfj
cSw9E3YhdFusBQQ5MTnXFEosIPtwv5gOit5CYNBK+uRIEAr81F4Wh0gCNOq+1KR/
XvLrM5MpgZEeEfVMUPMUhhac5xZ31KaY7NTQsGcT3XM98ElUf42rOyYd2ifA8XzZ
SWzEIVA77UJdIkwB/gJUv4AfH2rOkNGRrDYiFsgB+pDaB7f6ds0hC3H+w5lrbWOx
gX2pq+2pJ1QVNuxXDfT0cJ7i6uFPmc2Fca9upCY4J2PKNk1M5fZ8+rCT6d/HAqKv
kevwz2D09Nu4V1ZKQnhRi3Yq6eRGouoV++tyDytsXY+/btP1GadJfWX3DoF/opi+
7u7Enmpuqzoo9ClUB1RsvC4NEpDM4/nywCQjwTwl3UMZt+bFC0ahRTjiwp7ojn2y
hVokJIe3PXF1HQIbGCO01Dcs1Xf8uv8Czm9eYHhH+t+JfE03zlkVq5sdHYLzClk2
F47SbRAbK8xq7PkoY8K5F8KXrb06iVpARYD3jlbl65eWjyHut45hMJ/AO5t/IZ8r
3rBz4vl3V+IG63BCBf8Qyg4zGQVfuGDxqm0hKfEwktbiiChPjm9Lt8WSZCcuzi1d
T3Xp+37QMfWulw41wXJBlPOhmOezb2tIu2rEh369zdCOFyG4TnNt0CykquEJ1dJW
HWDB1MWp8VeBfVx27dWDlQqhmTEpgaQ8USAYL7KxAgwGJJxVPCucdkHxSdGzM9qz
62hRMYIeuPXYDYQ9gnUN14gRBpEqj/7gab16virbxEkfNBzNpKWnsRP0r0mFhs3m
o6UBjFrR5jD0qNMMl7TNXt4Zv05Ewr+rJ4gCK9zHqGg6XQ5QSBg/2zKCVd6HJPy+
iQiwHQkXi7EfzfHRhfALk0J8iqiw4V9w60jktW0ZlS8q1dk/hQwOVdRh/LaMZpRy
BT3bhCFlxSYCFjTGXQuHJ381BIE5SuKSw7HNT4w137h1O7ctIIQ16tu+ctWko8Vj
49PNdUDP4Sr8xioqLRoCa8WIG9o1+AWNhKfLBq957e48u1dxztgUoQbodkPyHjl6
L1gMuSrpcFoPm8FfopKo5TokLaa6Mp4bcsQiRlNoExWYA+dk8/RG7rHitKktjqVq
xKEiHvPmxJlq14jE6hEAQzbIbT246fB4lZIyla5iujAd3EnmceZJcrniq1VKdNv/
4A8oj/X6PmsooUS3riEyTEQKUtKnFRFSa1lDB2rna0WlRFa3XFn5mzOZIGJ+eg36
lYrsalTbMHvALfz33WmMuziEX1L6BO4ju9MqGpwg3a1LVxlmP0Ulfn0ozvketEL6
mW7NuXHq/dA6Odk1ahWG7SY7D/CLMV0Bl9sesNkEMOvGG1hLaq7RPFSmVzVDW3rF
xoToSWI/Rv4nUpu34eAPQNQksbaLtaccgJU7th0AHedHq1t0UzrJTqASuIFB3ESk
ehVYldTLR8dnrTiRvePiXbJSZwdL6HAzd/oJYxOyMJLLbo8XlqWAA36o3Pfuu62r
YlBv9g1dagsUvSfvqULzAVOUtV/Foue6F0cPVOuPKzqjgU2eTcKsUCPtA2RwO6CG
vWqH7jAowRfhcfcACn/PHjlbIbrKq91u6/wwDmMBjB7fzFLTgflZwdD9lHoxyzJg
7O39OpUAkObznfgYOC5HdjkIVdrUwrLPuc7TJWHmEJIzZ5m59yf/0yG4vtMT7Yts
mUBzqJEzhWgF786tPE08Jmq8EZLK0Cln9k84+SUXp3XLlaLWk4fZuhlGaXqBjEa3
FV/A1la3YXobD7rZpaNmyulZlkthrqNl66tbiDYwqdS30FMKUzBdldokmMEnxLSN
7alE59r4LWmMPQc/tKDvV8zkiXc5Qkqki8QPmkOj7QZ4whACDPiSGsitWHSggeB0
XH8HPnK9txP5twC/3IAJb+M+8IbLWi1HoqUpu6ktaDB0883UkzCy04DOrmW2vdyU
O9wLbib3JY6nI0NQV+pkgJfGUMJjxc2ZttzosdDPg+qUnCfhw9h4FAQ4sqBG4l+F
85zDzFZcW9XFyqfVC9TDZNOSFQJxFhvjWJVhYfr5d1jhH9ltDFrHbvrn7roI3ctt
lFrS/PGKYx3vpUnEcdyWKHuvtL3aeQGMupVqVjQllY6grpWYTjF9Xhqhxhyl9Tuj
rU9190/ppFL7Hn6s6nxFXrDA29N9GfYiZ90i4Prv9UO+hFpH89LIeYGkEeXraTCe
0//tTY2A5zo7hC17/qGSu90dc9iB2AkQdAF5gTiKk1GW/e0zHhzKuV50nvc+nHKc
4NDXc6MfBcw9NNRQhgp6DKpGZCO+R5xknA2i+lzmgCUyYWUukTdS5zWzsHdl1fpr
04OJ9r7ORlQR0jvYDtdSs3UvI0g1Gaf33tYcSKZWIaZHGUTKB+RzrqYR07+KneG3
dkhrA2m7C5jAhyZBPtjFCHDlny1h3rZzTLbqgiNSPH7CBDtaPZMkQF147zfaS0LY
HX5/bBex7f7eWl+el8oy24ugS+9y7rPhQWNCXVsUu+FAv9N17i/dWMa8R0wLMiIn
4HeaE0gK80iBIcUZnqTaOEuEwN8xEVmx6rEWX5XxV5T75/VWfqp/U03PbFMOeUrk
AiK2VUHpFYM8noGvOHyzLgYjukgestxelbrVeEYD1o3L3UABkJ4322JFxRoW1d5A
kpYcPzGCa17EUhY9j06S1NkVj/4p8j5265ou0w+b8QOYsuAM1gQ5cWhy+/CgFnOk
zzcyNw77fEKXyS/gxPjLHT6a7opY4BYcnYoviUyUUazcemJtnyPQpUK4SLfzUG+q
zbzaggRlXwmlKs8YRHHAWo74QX2yO+rqDVKSaY+kqEb3aht+B8OeCkHW7f/Jwmju
`protect END_PROTECTED
