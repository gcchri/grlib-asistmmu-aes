`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ykr2A1vEBmdR5NqE22xl84jAclWGwe21OHq6IpKlidhu6u4XoRBI+clb38G5UU50
X9B4rvNsswcAZBtCYQU7C9wqQ31IiNEEcpU7c7w1Hq3CEDVYJpNx+UAK7EDWM/zK
MlIC01onTFtVvbPwS637CYj60ep4IYi2zNdFFh4XUjpNdFG1zRrJd1VOLx5wIndk
FQI3LAJAU5a+I4juo2C04dPZ+NP3q64JR+BpRccZFX/Jptpnqm+9APo4Rwn58pnz
ZvpZcVS+r/Tk0D4YcvzGAK346Y9qUFt5hB1/yISljRs=
`protect END_PROTECTED
