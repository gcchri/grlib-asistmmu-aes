`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C3B7UOdcL87yR1QXsWKUwVXXUzBPnnsccr09lQQsjgW0+z6/7lTxkj5YAqt2v/LY
f0FS/8lWTcG2/3H1uXh3k0yk/MfX3HkpBVWMv2vE3TD5wE8HcppCWCSPiagtUsMX
CUfDl0+Oys7kFDQ3cY/pI/NqgBfDUeLsVytdJ0NkfUXE0mMPUPlPlnxB8gzJOzyH
OG6ODlxiSWBWgl99J4LUwyyf9LBCcDZzukvjEHhZXtHtKyMRhnsJamm+/0vAYAh/
L3aiaUYgYOVQWiNxhRtgwNRjXCaKhDmThLMKaq4aUM9p/+TuGLoifBLkcoL5OWUt
xXNDKeUWaz+QFzkUTodmlr8S2nV0AAYS9h/S5M4d0cxpdWvMEsX06YWNTsL/X+Hh
/CPNFAk/qKDnkbuFaZVMXJy9yVOoXYEOE4UzvphgVeIcskiOeoQRq27MJ9j+h4BD
X+o3oBiO8SSpoEjPCgjdsslecU7SQt0qJEddqYSX1ZhMHfp1FSolu6yRXgRcdC/V
`protect END_PROTECTED
