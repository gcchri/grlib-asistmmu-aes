`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xpAZfTNUc8T0MvCP25xfuSXmVd+mQsic7lZqMILsS7GKYAkS5stkYA+15GLwvxo6
OQTcAB9bLT2UJtMSynnvxleRr8RXnIFzJSW+45+ZvVW1I6MRDdQVN9c7py+IUAsv
5VkkL6OLfFHS4uyvxCt+3xHKLxF9VBA5aWcwd3/H7DQ0nVaMx7az4X/hKBb+b6ke
ZDtlbPevWpHPzszXFLw9UeHzGxGh0vmIFjEC/xjGR6R1w4yXyxk+7Bc1zxgDyrIL
HlqWeNA0Tj3pw+p8GVYDpKWQHrMRVNwUKPZmNlTZrgTEvJ940aJvCthQtVE99ODr
fSxznmRBTOyxrR4Eg5KikhcpE5bkqMy2oo8NuZwxZdidDeFboPb7kgNxxxZ5rzkb
nqAwMZ4A2iUla2XFrvNIm3CRNdji42BbbSPZFBAsjs/3RDFwwmuXbsmAtsdNcMcq
q+iOHNEYzwm5YAVcIpptPPj5u3e73PP6RnuAOImmh/9Sm+nirM+NeleEhyczWk+W
IsbR5WKnou6eRgNhdabvn185iMOuLhTdUGdNMnUf1GlfTv1Z7Wy5cmbOBo4IBO/N
Z7ufTFSSdAAnFZ3JIvLNy8BjG+ttCxAHJpe1PuPdCN/oqxnVbV6QCWWmrvCerfEO
T1jlcP2J+vWHlYjWdegq0+dGpkHI2NOV84eEzJDJb6l+7X71GyKi4wpE+rz8Q6vp
a17j2RZQN+pl2ZFGJx0aO7vi4rgtoSbjC+7E8y3QEJ7OXyzDMCArYIO8wKUsqP1D
Q7fnLs0i1fBcqaIR+xCD52MaLFbEZeBoW24ZKC4uzbwtBGfQXGCxfRtrrmfJl/gy
vpzX/fAA9aLxweYQp/oROR3o+7A/1fbK35RDyHS3D3w13wRZGKPAVCvm1T/ozpI5
VWej8JQ0pHCMXBpf4DIkaNas32P4bJXKOdgKfpMOWNYpdzaOvr9m1Wsa5ZfrdG9U
W4Piix3nlAvH8drpWTWb4vAF7nNSJ4lSQyx9J6+xHG/PYZVTxQRGNb03bUNVoi7b
iHyhtT4dHI89fNDruIDNhDF4sCZTn950AvugNBGNSrNWQdhqjFxuAA4hQWVKroeW
fmKkeWaMZmgIBsoemxbR04JSmqsCD5s8UZivwBcLEhgzXUNyaktMkY1sR/1vs0hf
PcOONk5um4rCah5P8+MCaCyG5s4pQQdqIDs3QIrCQ0s+XXxh41KvhvRbOgOz5dsy
`protect END_PROTECTED
