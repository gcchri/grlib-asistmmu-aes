`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rOKE3isVNJ2eoKIv8htfEiqV769HidEZrsTnp6ww5VBFkSx+9WB6YY0jXbFVQBvx
4HRzUITxtZd9BgHhOK0G6LRmvgMKKLevNlSJULQ0bnhM99T5H26xTw7st2Bpa/a/
1IiZmIca39xtCysl/sh0gQT2ARGQZXGAZW+duiuJqBelfGtW1ai8lOmQQCGet+3B
JJ2eS7XvI3AJEgYPp6JYJs6UB6H3V54l+m6vs9xEUzFf/gmplsHQJ57RZwFM9wCb
mf2/bSL8Iw4/GeU4SFG2zFXeW2P67IvOR7mrBR2yWKNaXWZl9sC6yr+wLNDJjKE8
s7vPPMiXyTgkdQVaMRzLnaQ/cyk7r9NVRmkJn+fae0ESYbJd93INcGLl0boLBcTD
5Xa7lOBwU7xGBuu1R1mqBhkyIM8UqFTkMxRenV1oPlICGG2UF8zC+D0RLeIxdRfd
JBAVvvEIMs9N3m1HcAfasvFIQZFZm5N5HdYDRJpdT5UcIzURmbHdXFLmP1VDQA3P
giX0zQWFpHwXcgBwbwd8wEscUQPTaVTXOPvi2W1TCXg=
`protect END_PROTECTED
