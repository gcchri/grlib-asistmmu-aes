`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mU5XhoVGCXkNJ8PZXfI5NoaWMRS2/dLhDG4LC9EU6G3BPSQKxvOLi6vLPZ0qD36Q
EyBZUoNkIloQae8L7IQVs835pWW8e9Khl0DBCEfAEqSkMbIhKKoLEDLwy6h6/YsI
4NYfIOeMyqVFjuk47KjyxPfbZ0GqImsCmrD9KPuW+44DimpfvVsmAdtxufY99zhJ
Ek6rd4EtgjTngIrqZQFEsw7uitU8anzCe75FQUbTpVYDiu/6d/mBw6yrHdMKvuk5
18MtIrtgG8mD1HrVlSdFhnWW7C5LgKhZV2Fu7oCQrS7ZZyuRPGpjl4Aqy88GV7tT
xR5361qRe19GXZFw37AUXghqEYXJxMd0JDfCWLnOFVATdhObXnPHaNpRnC/+f1NG
j/PLtptTdyehax31HBarWtheYP77XHZJS64j11d0p163ZYGYNtDPI9TXZm5fLDbQ
miYzglQvf7gBLtgm7vmV0xfbOsdnrca4gHGs7l9cKng=
`protect END_PROTECTED
