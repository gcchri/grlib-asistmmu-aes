`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fgz7tqY/H2iFzRklyb/yu2gaiDcAUR3t76znq2Az3SZNEu5h6yMFBzH7ZUnKMQjn
jWfiqWo7wS3jljIjJLBnXHnFm/M+U5IRRCDuA+jgXp3hCc/ftvX3Wg8rRxnJVpmq
nXzcYmFZV5SQQdkWF1eZaDsbDcAmNSz2MY6kHSaaePqgnru18XfNKYWWrBpmYtsw
nNQ5kS5haUuOTGI6ChJ+pXkqx9dqBD0nV7bNitvNZyUpRRFS4ZI9/T6OPqpgLcp1
K6mRiFpJmgzNbjBrIJj9VFtiF1KEFBzG8rQs93quuLtS7mzIMbmuZ76YrMBVcDtp
G5fFtp50j+pEjgKyLn+Dn3jOxMFvBy4nAuzYOpGjFVKzCUxdr66XfaFx5RTZVsEi
qeUTtPjXB48F71Z46RnY7O+4XgRy34FoDdL3Dfuiq6AHHc5arZgE+aTGpFe9XkXc
pjZjj8Bg9iKsXYCTZXiEpO/czpqGpqSZfmfN5Jo+jYBlnLlNMO/VnxruTft35PeA
Bh3qDSPN/68ArSI07unO0a5cy4+wByFmoBhVW8ReFhweup3YHCdijc7QNWKfdWE7
gUeQ9MtQM64fYaI0rVyJFwFbQD9fvLmRHAARgdCggC52DLostVucgk6MbXpIljSM
Txr7rPGQjdaD23DhrrBti4IGCEiubgfbfPOdMqWBYgd75zxSZdtzex5nUWPjKff4
QsmlsGufY6r6MrWMRAXG9RoQybbYu1LF2AZ9Pvc+jOmOf8Jk1Htxzn7V3x5rK2QI
ZlFQWeooWXrY2Mccq62UDsXE0DgTSburFxnKA3Fa/v7oHDXM6OORz22whbC6idg/
pp/UsBOb+FRy32B/JtBsiZQ60W/sl3A644wZn21O4G5j1z0KVaxtNBrqGSxxwhkP
NwS265NETGs2506Q7dO65UK79noJ46VMagiYoRBD5tNderBbms+o7uIAN0va7sWE
HDfPveB2lSkWyVGgrWDlECVq73YLllCQ6AwnvytvuAAxn7KR/PudCulm3/hK9NQH
KClV9oztYk8hR62i1VH0fYBksxUQPYuyrgFRjJwGkKMplTko7odL2Cw7hMVgZgUl
UXSxW1IQBVIrhigF7Fy+I2AV865ODdH8oNCNdYJfagXfZB38k2DQpOgVDMG520EA
K6fr+m6tZr01kgtHKhGA1N9CjvXgOKD+IJvIfSRpeeAhAqWCo0L3Tyt71/N/RTnY
SXTSie21aeVCHm5v0AhpEJ+yOkFGHtzHlg9SsyIKXTswPDYZZ+NsoOxYHbTBc6C3
Jvns29kfP9NkRevPMlr9VaL+1gz635bZAGy1CCxlB73yGY/NQL1r29+5W/XdSxc9
`protect END_PROTECTED
