`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fazctX40hxYsBdzK2jRoCLZ1m2VbdowknpMhCl17nKWTj+WbGrutrBMMnIaU9yxm
kSEyi4TET/M235PW+VQaDB5i9JBNPB3ywC8MPWtRIn1fSoqZtNKxnvzdfD1yA1JA
6E60PKGdRd1vMuC4n+6h3CsVccjn062KY6P8AgG8jqfQQdoi6hn+X/CMoiyKJwQO
BsOOqelYWdB4iX8l6IXZpI+DfcCb9mCmYsmOziDw5nWueZVfeOuMmM4dq9Sw3rlJ
WwecEbVGCEr8HUF+mWp4AKo3amkhjlWcTvBg4Goq/kZ2POMnc30XFYDB4vTZAsos
NQhR7E1/ZK2Sr0LesXpfz8tUwJhAAs0RxGcptyh0Vwdl/UfkTOWV+KZbjaZHCByt
Mt65qOCMSnIVckVnv+sQK8Oue/SMWcxVsiSz2Td7sFJtJ87oUZpBR5dki/xZkYEV
HINZTyvrRvGCi1L3USuP2tNgRspKlY+pe9t/CEzfoUv3noQHTzzl2HD+kzdfoMV6
rbALNtG0O+bzQo9Zx01h9MbeY5prDHtgiBefrgxozYBN+BQbIv6K6rcloiGBGqPX
xZD2QbY12lgv+DJgwrpuPnUNYFFCftCr1JLFRj86Syxzqx/Km4ORzXot90rQzYJm
9GCPSrmtGNsvidtLwtkhCo+n1WjqvzMfCxNdjdDosTk=
`protect END_PROTECTED
