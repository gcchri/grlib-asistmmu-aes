`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IRqpmk7PZb8MupwzLtKBgeMZXbibPAGuVjzjffRtbsVZ+KnokN5xZI9Dkxqyu+t3
aKgLEOgCpTHnQgb08L4hQGZTNRVkH8/s/GIMFlrWV0qnu4iUZGiVvML8EyXjwmr8
wHWMZd1pgXVvgBUutKg+IyTUzJ1qGmGmcDEQuFxw9h4H8bqpNIp4wzMRZHPo4SMT
yn3wFcbpLpW7Vu0iY60hdRfHBTaTR5la89o7gX3zP3DztDh49EwxHKMOACYtl2rA
MAUg3npT7/YG6HuiN0xRMYPv0oT5NmULmfVQzgorwncWK+V5Tlz4FDaxeS2qqNZN
1bYwfUCg1hrPsdxrZY8GeQ==
`protect END_PROTECTED
