`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JpmJNopHJuosmhEZfPcsQcuZ4d3SYKOAUVV+6Oqql7+mIreAK634YV5PCh4co6jj
RROwf6XKlUuO6ZKfdcathnWke7/gfP4ylXM2O7WYyqoZ0/DEjar+UIT9SPbi5zo2
BTpz93BzVnfEAm90irkBPBQWeBww1QpAj7B/cWikGwDK0RLe4Y+ckZHxLcAMn2/d
L7ifolvELCtjp5Mb428zlSxh2NjqFT7T56E9iRGYTl6uMZZ8HY+4jAATjZJM3Ox6
17IlkKUiX7QiWhWQG1VD84vWYGL/4ChQsJ8zI4XfojX7GgmagFXFzdjjP8pq/gCT
iwn0MwW3KFS7HYpddNe/vQeS28FG+bTQVrXpy4Me3NBk3E6OOJmnN9IPgCKYiF+6
UGGeWrm/y/6eS6x+PQEwCsW9qVWUJcWublv9/5uFhtU=
`protect END_PROTECTED
