`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pSi70jcc4sp7SZ/XiuxTPIOQjQbubjezuBkptbxH+sC0pBdYkIs1nk2yM/DGbxdX
k7thOaG9ga32LYUzyd9LMqSqopyqfWIFfjGNvICtg9PB3uclHvbeMEJq5ETE1rk5
+sHHczaXzhKBDXD44a+RkreZGIcrImyCNfZpWdHAN2InHtzIpBKX3uBp18mBoVuE
a5YvV7HhlHhG41/tgFGyj1x7OdNNfsKtKV0nhD0KhluMmcUzBtxF7sgfpF7s4+FV
j+OxIELN8e2skIGNNzp2Pl4QDnHoHjKCLC1+2cqFdG159KviazLrO4iYFlRJqe51
NiS/aVjnV4xbfz7ONkgNSU+USSeBs6QLXkHcYmgNF952DUDzaUd7XLzF4xDaOCsn
DJietXRGbB2WKjcuEOYJl8+EiCEjt5P2XDwnemKPfB9hZ7z4NL4fM3ZvSNzaYJ0Q
FSGX5XkkvoPnlawXdR+0uy1ehF1NNX+HUKSdvj+0HAMQKFOLTUdWGhx0HJWJFqs/
BfPFFuhct0MFy+zjoV7UsmfZy6JmGGVCPT5cnQ7lR/HuhhTSEFOmtuB0zNaT999Z
86u3YLzglioTJYrXXL85++W8giNRbtK8L9FXUAEpil75V61Ua1QlkTq1ClmZsRcg
cyyt70RT99kNGNorj7+QSO3eq+q+06ldXP8vsTexD33+7nE+UHAmHpK6dlZBfIRw
5UiDGbYQww6gLN6sXDSDXBONxrmrODizdUqGLOyllEG4r1mMd2N8JU9KV3gBcIGd
DwJGwPmykZlXoug+OfCWBP3jlv55e+RPz5LYdlWEuZzJXboQ4DDnS2/ubXaHq8jb
Jkha7Y9iTOjltH2sOndaTNVQqZ/Vp3XoSmwG7Ywo3XKMwiL8x5eydRbhfMr1QN+o
G+VImZbaaf4sWYz91xzE5g==
`protect END_PROTECTED
