`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9aNXONxC/64PpRBAuOSB28Wme+gs06ZYjuVQftqmpbdwVe/Usu8kSPSSiU/7jQMi
8eQrf1EtTA+uAdaytFJfNmRtqPx9LBE2Q/mFgztdKawSUgVXIjAAhZYnR4ULIk2J
kT7xVnuDqTBu6GfFIhzwQ1A1X5VCcDfHzMAiGo97EnyrC4/u9+V8r1Vybexeyvlw
BlylejqmQRzfXxTeaP7UI6yqMUqFVRyongVLxpipW2GfGunSfneFDRLqgs777TXo
GTkmnk4zWGjV8HUbVMkNQ+kpZn5v0XjAxIfCJPviKZpK0QHbkJr1C08yYkqCw/cQ
JJSpPsqXlzCkE2fIAouBionGV37oySenIPC/QNN5F8KQtn5EycljIWqkjBz+4HOu
9aG2ZYep8h5U3vlSv6tjX2OggpPX8ex3p6PI/2isMVP50OtkWJiHSehMT+H+CcPT
f0HnGV23VEqbScr1fxUSOFkP4sb5gX7N7LMQBGzw6r6mjsvQqPOcxYW8w6XMIbCo
No0FocRleOR3/RI/qss8jhxYKUHTSdMzrdQuZNTVZz0H8HPQYURJjvRD/5UmlfLi
wsWdID36QynuZ//pe0NOBBLyWZPoP7dzvHUUtOgEG79yLnmsBi2BcOiS6VOmhS/J
nkacSy4ahzb8zkEDu0/+Bg==
`protect END_PROTECTED
