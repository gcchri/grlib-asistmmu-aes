`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xaRac+gLojHzqg8mLvI94xAaDLVbPSfwQ/XzwJa0ItcXeIyH9ww38aU4KIS9DowB
nytuqrQ2MQRFNc6VRrAwBTZ5NN+qRRsyf/DEM3ffsW7/ZoX48+M5H88WmFIxHfeT
0PLhzYdJyFgRD4Pr7thy7MMBVuF9SmBc1T9h3v97zJgb7RPwJ+GMDN/bwkcnW8X/
3eQWO7NonCiWfQAMsjPLBjyyqLNdrTRNjXOVX+odeVNMEjRN29rNhZb2xKffjnE2
KAxpj7DTENzcfKsr/DvzxlQjHpUJZNFILEGwtcl6Bz+7a9XUngHq02kt+v4jPQtJ
/BjSiMRaTPdsVTluHPH/8W9nJf8NDHMzZ/zbQsPapw8kvlFKwxliz4Gx7X98t/DE
xbQ5amfz2iw0z+j5Eph1AiIrEhh+3jW0/+o1+yj/tNz4HQf5y/8jU+oTXhMv8s+i
KDoJd//Yvh03RvjExJzVeUFfd7GP1zjAT4tzWgJNEilbKoU2UEMvFSx/Il6q9YqC
wEQ9z4D65kej0+hA+7UbxD+oKdUsgClyA+Lg6m0wLiSMmhlf9lEaJBUGQxcObgnx
oG4nnT4N8TcRLElbtsuA98gsEk+IUJUnSzeihrhBgYqOpipZSVKhXuiYCB0Bep+x
ZhqAnij4mg28m7u54zipe8lBCXsgHLWKUcdjBGSJcu/VCmyv++zVB42oDWYpIUHA
0l/qyxnjINc958BvJlAydJS2oOjhCE1To8wIuxcBEY5dE322OBaF94f8frDAsRow
jMiJyi4mqjGduWfNSaO1iGLfcmaCLYJKuKN+a2KqaCgS67IxYAwPqCyMbjs/HNEV
ePKYlF/wJVNnwEKp7H7Js5wKsCenxDBNVfFRoFF9WYP3qd0JoYxcN5SUGSJeFGZJ
iO/UaX6/GJlRfkiS1WNMA2YsNzUAeT8m3YQ9sFLm98ZIo94DPGy38zDZisAPPZqV
ksCg1zUEdhNzZiA4DjHSkQeHDvDYuBwkeRBnxgMhsQnjsrnTVb7jRC1yBfUdr3MY
Wrl0r+VST3T7vGPmZGG5hmUoC9rvQ07pWk06v7zzYKs0lIsVkJ3SNbSX0nhUm9xc
6+UcNwxM05zbbY3GWnYjgt1SOBGYIFhsb7KGcBXcKTHFi9ROce6n6CKOo3YYDrD9
wMaSCtYxkEmySGHDAq3SJO88wfBuAe8gofl5YxWN/BytFAolxGEICdnA/OP8GPHu
z/etfaFhyO/qqIJxLdnr9criG0yHs8iUMWX8acskp8BRhBUKvnGhI68ggXnYkaZr
jW5bM2Oa9AWCuva/cbRWnOU8dggRVL+xlllpyiyeIwY/0ujHut4gviTf4+9Xlue2
ofhiLQpmG7o+ELmIqKT2gaXc5IWzdil3rTOre6eVlvVkRyzm6Kp8VXf1NgWUvMkA
mQAi245IqFal3x5acy10+x49CVO8u0UmqWXq1FTwx12FiU4dBmj0O91QMuOAXYTZ
ztk3/9U9MoB6GfOinjgq9xdhIS1GBg5S5O5rvuZCzQCradh2BWRNi7wcSj2dHdAw
PXHxYvglo2Dim904AdS7Ilz9V0stndJ459eku4P5aoqfrAcdO5uVWH/tGU+V+4ag
hLDg0l6xY6GM65NpqZkgB1Oq2SIG1BoNeDV7BZTaPGRS9oNr/uzsckRHJNbHsZEm
nBkwFgXra/lzudVWL4d44+wLHZMvvAY0v/E/ekcuNrEGu0LNa9NQiTr9IqveD3nY
6yMGqb3BcXk38KqwLZA1SsFKg8sDTRe1iJSFJMmLLyffbUVg2NR50iAFILN29UXP
TFTzHksJUvPWYk9B6doRkE8NtrfAhQgeJsgnmgz5OAy06h1yZKtbYTnZCAT07EML
9lsye8iMeTFVB3ihDSvlA9OI2D3DC+JcVWcOYIJMlt/PkaHogu+AlIuZYQaafuha
UYpAKJpwc8hM3AY1xLpJLkK0O+ea/qCUX+146Q8dzHGANR0ixR67BeoyWS39bGfg
p4J8q+c3Rqa0/WXbvrLF9EBIoPRs5q9NLz3Fp1IunmSNp0yk9u8ifhsB2dpVhmRx
opJwMtdajf+z07ke5rgH4PXoifhAwAeeiH4PGLEBrbTzD6PoUcNjvh9lLYNWJkMn
f1sQWC7PPCUPO8pq4t7uExtMG84ntg+7ENMpZZyBF0ZTCzphBHeyVH3NOIzmdGL6
`protect END_PROTECTED
