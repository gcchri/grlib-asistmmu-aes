`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XbOh2sm9B8s70kU6CalBrLJt8r1m3HAl2oAgzFUGHFRXf3VSOXvbhSwEU62rGDRE
x4LRnfejWMEg68W/UmXGnZAMZ4xGnFb6yyZbop4Ncmvvgj8QnMMUNaTTFcaJBEqV
bUX1DuTzczibspO4lE/qTHWLbGFypVi9HWM+EqqEXk0C1rqaQkq9tBqR1fNcsAmL
xOXXyw5Dnd8U48nW/GE3ykuDAwsy73oFcJvNyA+k6lkYBks2wc9eUzGEaGIH/aLt
yeAiXVoG5vhPOYkS+954JDoNjAtzBeHXymff8THWd9HmofKZ8hHsd0a21q3ae35U
24DTnuJe0BziHmLvLkNdStr5McxtqOS0o6ToTLZAGpd0cOqRXOZ12Q0j0/aY6cT7
oAwy0Hfuo1pH5NoVtGyvrEqH1lBFKSBsrNLONLjsIUDbCW9J4/AuyfXQz7wsFBZ5
ix1I4fy1M5I1Zm6HUHyi6np3Xx3rYkgJUPnZu5IOlR6aQ1E64SCXFTi/4H/ACH+j
2SUV8h2/rOrLfbgevl38wPlP48waDdoQ8v9+Xv18BDoTnb7Qp7zO7RCkcfOpmXhy
kAPEPSXiGNDOHJjdu5bwXn6ZfvosAysqXGMtdHVyNGI3Z7iXEfFcOADuGpx7gy7Y
kQWws/VLzteBy+f4lPw0c1oXa1CxZqRL7apTprJghpp+oeU4dHRL52vGxhp3AGgN
0IUpivx8/qsfxv3Za69D9ZifwOAUmXR4GxCZh8801vx3/FrEmmmNDIWL1cGG3/1a
VvTcBuCzygMQtYxloYC4c9UmkQkcwYv64BQ9tNY7MM7pz4dpXNpGUefjtvx+UWVI
nJOjfaaUYpHX2y57tHY2aFmS0XZAFaAKd4qH1N7zKKFkhBCcTt2+wUy2vwXE6mXY
se5SlZn1ebFXEaZu7zb1TeDAYXBKvRipQ01Aibb9wHgwDrKzGmH5k6ObeY4lfVdA
YbRJlshbqnzzul8VOId8HSRrS9rIkkufu3/92lcVpxWJ2qRaN28sHeoC247zCB8T
wt/gpN3ce2yQFsDv9jqgZQqSfRpNwMWFypIxxd8bQs/+zkrtJ4V2hDFvNkA30qdx
KV5aRonANgkkHg78ywpP3dUPXuP/fxG3esdoLPhRuBAq/WEvqaiRGfIOjJid+/gn
CWV5ADFTbJSSfnwaEuJJvqpExkrSQSCR4Q++7w7Emd2MEQht9UQAmfhKJP3Q49er
F7hmmH6tg109fraYYMveld9KYj3sUxWYyitXGR7TlrZE0oLvI9doWvt+hxGyRVN4
i5y7syNu/dizeX+Zj/4uEZV8ciY9O/haLc7Qcy1hivuF/kOuuupzi26glJxCK31P
7SEXE16rwG3zEkSJLZoCLyJnEYqhQKGdapjWLahiKnQGJGjkcCyXdruLb4b/LEfm
iaEcBUMIRyfgqDiEylJOuY+TJ/d3EhlQZcZj+N08Z3STXRfvsLmz52EDmLvBkW8e
wf0WqjelHKemCBc+gryOSz+T0LwFWya4h5MeM7WxnXiFxuNiM99ZrQS+Dcstkmh/
/JxcwrZ+M5V7nNiWSnv0/XAPPNvViLA4HDd67Q30/thLMS3TeYKTBFQd9Ed87NFP
dnMUumRuZOJZYdRGVgDmDCsqhu6KUGfrRC5TSBb6CH0F7gFiDX9J4VW2sbRBdce4
DBj978+vF5Y2HKRRKgp1lKVQ3vx/gNz4VUhVLc4Na63whBGAPTwM2tMt+GpEa5uG
kaqmc036e/XLgu4WIyWcvebZaCO4NNADCgod6gR3WZMDV7nA/E0CzNhNPZfEWG3W
/nZO9rgAQZlP16w6lpqs5C4Rs2CWV3cW/NV+75fE7xH4QMdaNfl5bAQsXG0Rde8h
iGvxvmDZlyumBaSI9POHiLj6SmHg7SojcSPl8fOmZFWuMRaY89dv2i8kBVsQaF4q
GyQDwI2IjJdt+fo7s/Jx8G30RqIgbfDJQNFCQlUpS3XUiirBkPw3/qNOTS8yjgHJ
fMUJZWwZ4bLVDzJkffnVb/5fkNwkhkUFr0lUXGzU42uwVo9pByEjv+FEGLmd7z3p
7pBf5n+dGcwCSbY+xjG8Efk8rER/vogs1wFKuwQY4VoXff64t6yMVNZujJASQUoh
r+JHCuK/pJ025F38lMSpMGKVBVQE/xuiVj0qqoffaHYOGr4iPsyLnZFM26HBVfPV
k0cri9ytKZcVtNJtOxlZ/auGn08Km5DEpBNLmCSpwBugXZymURhJ5hRkriwEWIw3
+N5XHc9V7WdRVu7DQfLd0XrcngqiczHL3c23hVugDcgBigkEodx81kZfNxjgvs9/
ryDyr5UEGilxZsKxmHXi3o4kuTduHI3iIuFmvfMm7dAzDpeNRQ5WpLu1EFQEz/HW
q9Rn+mxwDiwvmoTGFODgirwn9VuQ6bpDcA0pLdxiwXwghw/78brt4oB79w9NvptN
BOwjoVS5kPMIKr5+13N7FRirjFqItNxfBM7Mq4XuueRXo25QNqn+lRnHn8MVhVzy
6NeaiGFHlaMu34w3jmc9MV2252vtrjRr0zSuW0O8kYthewkgL7LcBy3Ip9/KIZWg
wX134cT+HYN+DWYC7RzMN17im8dnUovw7cuAXZCfzoRla4ngDI85GifxM4zywmDs
3wGgtU6RQQPgu0cJQYusyCIaIsIEC6M9NtFf15t9zOZlqWcuhjlIXnOeQNVQy7LB
2mYigeCZHVQghZxr18UgQsCNEyhRIDpzFsp49laU951Fyshf5alJE5U/Pf5OCWiQ
LZ0IRP5up4ivRPl64H8oZb/pXyd0FfnXkMHqMfEnHF8unU5juiUUBrh6DYJCSDbP
bvjkIfod3CwEL+dje0jSCQnVZlVvHlU2L8d1z0LKHBel2btHtY9mMUwSOqPIQ6Uy
gCD05rD66cKbPR0bYXfXu/RSnX/V6+QXyl7LRv3hlbTQbHA+T+gaiIj7ZpLJExDt
1WNvbC4/BuLdAtVsoz9Ho7HAS1/Olr1FYJOpUdXLx2WDIXb9JWh++Jltq2uE7l6i
SHrJpHphh9WPGo+viubZOACbura4HlIyJDfokANJLqYWWLSn5fojGehhQ1gXXwOm
du8msGcSJ+W5Vqp97Y5IjmkDQV1WFbYIblTUYJsHiSKhFV/y7Pz5DwgSvfGbm2Co
ba5GsprL29OIgDMTmtQ34nPk0Fc8sRqqM4YoJKrhxWHwuz6NKgNu2UwflMGH9Yv5
/sL6YHqWgS22RbE0rNFgILlmhP9+jJepNqf56ggOyoWO6tFZQsHiHHYnshxN8NLE
KG4WbNmiwwkkIMgid2nrCdUqN+FDhx6KYRlXicEt8hgCW1QUT3jBeXaGF3fzPwAl
clMM3ha4QIBZl/HveoiOzpF4gTbPgS2jLkQVvJ4PVJthII+xbd0X7JkpN5WBk5dV
zDwWYeRZtRwL8dr9hFF4pQsQa3vqk4l1gzpZlKo8eWDVBPD+2B3DfuDAjNxJqipa
WwbwRTX3jpf1o8W9akosRiHBZp1QLoesumoqr0uEETkAxhjZOnSQtEsjE17stnrb
CvXRcKPNJksmSQktY7PfQekZbHSt3u/EB3hBASumw799yhw597k1uGB1RHqYi4Ih
NYSIGVUIXd302g4WqSSGgrGJWofWdlwyx/NK8EFDOY4t68n01oNaZaiqhuOO4IYb
TfbnFSZ9LSb/h2fGM1b7tv0FWpI80fosY3xf9XQ/XNAw4UeXccs6uQVknyWD6L/T
As2QZzoa7fx6hBOmchEpN3oujeed8TXJQBNo5LCYIVU5LwKADrr00blFEy4XqTPP
a/kbxXgIxaQKHpmZCeRN4yqrNUAuJE+xlKsjy87OFmAzGV5D2vRLniFJfk+e9cck
szmHzGUwdjNBXNzS5jbDPDNQpd11YXErWZc8jQkYzNavhmh5zBc/eosm3/BdyZDu
PpwnKt8Jn/D2x/eLMBypfYKO8rTIDHmyOBlPbyUlldEiRExvPBlJgiIwlB+aQUot
o+7vfl9ZxFq1TJ2xCQedw+h66bVdxK1zXSyw0LJKsMRpzMLQDnfIq2uKyuA1bbGq
CZPmVgb+mWU6MwfRX9aPn7xIlxg9CMlvBR2qEIReyilVmYKKcs1Z4RuA/lmmMcJl
zGhLeaP16Tm32PxVVIztDFO71akYUDWw/xqCcfGyWDstPbWvi/PD9pWqdhAl0oAi
XBpkyD0pW9qM6PM9sO7MmQLScN+3DCx381vaQBZfq9ZI7dV8bOXMdlV1Mxolx72S
pZQqxCKraILBxz+1MYC7gUrbrZOCf+IeLQt/34YdYHCzFfEkL8aRpZ9/6JQY+JoH
gDt0pba9Hv1BqXSTYsBqlQ9j66yhPeiuztjamWrMbnpX71dOv7tOVQ6Bzk+DXxeF
U6Cm8deoQzJh5TIDTWDKvGuOG5c6ud5Aly8l7Fcqt++/A3twoSVUQkTQO7pKKOoD
niPPUn6J4LtEe2fYnao5k8NckBH6GZQ0lY/e30sbYnGVbZI8kZr7CeMRaoayruV+
ddOhSVjK0NVW7Yca0d9QSsw/XKTa0vfOMOzS2o/XypyeKK11vbP94uDYD9m2/zZ/
6XZ5Se511UkUxLyt0OYiOY3mkr3avcC0poP3V3g4opycV5r0mQ+z/t4dAiNp2pW/
6N03Mj4kznpd0O6//oxe6nKw/KaCoP2GMgQQolz9UwPSoYrMqBE76UwDanwB01C/
dtwuz6mDyvS+t9UR33PKUo+Q6UZkUqyitGDlem02Hc9eBMWKFKuQ2OfEMDU0URml
4B8o8k99yi47PQ7wEC03cfWVjO3MYNvHM3A0pTZM41aXQ6h609NzzgCAq+1rCJ9X
txomoYZ5zvRGIicE/RE3akmcyvl79GQ7jVbz/bsIgY2uPFsR8j04KH8c2cu2XKjo
cxlm9ABukM7GlbpU28aXDoFARN+GFVfZyobD2PPDu++kR/nZJ6j2Qkr9lujzy//K
NSX8HZRnke5a52aFe+v3v6A+DYMU56mXLk6OQWKz4LrN/7/z54FxHz1e7m47jbj9
0pewiHmLXAetUahjDqaNcFc+ynBiptPV7tWGrQn+JS0SwfIAxJIcmVMWNCFqleLc
H89X8yTv8LD/K+u7LCsJz95DTXk4cA94UuFtbkZiwzuJXFTAikRWealzmY04bkcJ
wBGgEDsy2nQ+s2ivUzneMXy6O7vyJxKRaSU5ES/qxnP4EE9LsqyC+FWa4bBqxFoR
tLa1VJNc2pkTfTaUZHOB3/0tU5q8mrohxybnZ1E2d8C/IqIICg97+ZSz+Oqx1nsV
FoOeiXaaSS90W0Yzfxp2ChGz0ENnlHDxshpmNl9bpQPxD57E/V9r/Q8COuOTrBIh
/J9b5y6SZ8wzPLvxL3XYSMwX5pS/l11Cuf/qxxTNwBEhc9teaSuE3a1Y/NF/nSLf
GwmrhFEbmUPT05SB0FF5/WkBgLkDHRw7q1lq2hSlQd/haJj8X3J+Z6xhqZiV14mL
LqRrxoXzEy9OOCwrZLqNK/KByYysBuPS+MG+Twm7rwUhtrPTu+eHiwfEO247S9Xb
5LgUf0Z8y3vNoitHBpmSDG63trV/KN1I+BRhtjNeEJPRani4szUtsjVmujKrrycg
Y3X24A0BMt3LUglSd/kIQIlvwz2XdB2wiLrh4nzziV/DLF+Zz3s2zMBkOW7sBS6c
Hj9EOGJO2xgLM6ZMwbo30WxeopjlIOGuReM/Ww2Vt8f5Cf49XxIlpux4wdA528Qs
ms1a0WQStlhUqcsYCIPHfEHmNE2Q4rdMXuO04Kyg1vl/+ftCD3dpG6R8t2VvLMm4
VcAHDa1aBIStyMopztccLgostYotGZ+YWlLMZr/oJGNTHg3xaRsnjUBjHFwZmNTT
+skmAEjhgPMYm9xFhoeh3hCygN7NyFl5ox2/0ilgAENhiDGr22XDiHeGE/tc2KcE
CYj9EPXGAuUyGHFzt1xYBvlct7TmsBh5T2JGs2sk0dP7VxhdBtKwSgZ74P6PQRxW
rkl8iEoxe8ivV8++1e5813hNQFHsSdrj8YqAHsnSv4kwJvqmTwVOYSHXSvUYVUVG
k7oEMZd2kR4LPXgqBDYWMX8Q4gFW6EY4SSG30wI2m9DD/z5DyqQ2uGjPmXyw221K
HHpKXrQ8yCb8Z2nYpWYK3SE/NM1TCfNibQWlyjPwY5KT1MQ5jXsExig+2/ryatQE
VCwHls4WJoAHSl8sxcxalyAIWIsbhKfwgczOFLYiWT2xBEK1fM0sqDbYw5CCRd36
G03I/MR4gfOL322JypbSApzgfnDGLqt7Uxl87kVGaEpYDzqTEG5G++4KR3hxu4kc
NS5oz2Y75tS4Kl9ePEGxJ5SDIwWBlHVu9u6v0iYvyMUdmG3V9u9nUFCdCP8harnV
+lSz+wgcnSoMng8S4xfJGl//xdnbi4o8hwxmbhMGam6aNzfBmvcFdR+3xIslgwpm
Lize1gj+EtYMEgf6ZwGI2HLxgFjTfNW4MWngc6KIVp69HGSqj8MeUsXAGm4F5g47
cewcA93rML5Hq1leJUmEdAO2SrgIOFis+03kpYwlKRtOdmMKxDP3U4AZZyXFuH3f
Ufc0TwI91uHsHxOCUgmSc7RVI9e27J6nWjYMkjGuSXpyog/CWF4bGdYNJ8rcw7OY
V7p17/eepB8cSJtHY7YK4hYdrrwU+B6yjuCThstVeX3E1NmYADQx6Nqr7fGLCcid
3GbtgNTBqWdjDOkb5lwYGcH3s6bnJDBz1etBoS+QHvG+f+ctcyXFY8m7CqFu3N6k
NJ+qYPo22il6Z7AKlnyWXgR8okuCJU/+d5P5MuVraISq0zwXIy108ItgScsDn86q
b/iKH6zl3uqsKQ0TBcVvn4MF1uFvN/UPmMZ9izGGQSHMz1R9+z3o6MFlyK2Sh+G6
ivYs8kHMxQTah6xj3zkSA86Mp5qWheo3pc0nptlSaeaZzrcXbjEua7m4hY2Arshd
EDM0LaKKwHRHlRvQkBsthr2TMPgRbmZjDmvz6ymsVUN8jdGoHlDq535SGo4pfNwB
BY4rj0Fiv2ebBgF4dSR9bRGxK5iefaNG7/EPSQzyItwi9h6/dJBgCiaQ4/+TpeOJ
zPzXiqON2T92HAqXN2205y2FXyzeEU2xiqsXgeZeGJNTE9tFrGI0A7ZJtw833fBZ
GAQUrB7DxDPpdy3bYPO0eZK6ZOFZEKrMHB6qhTl5/G4KqPIB7mquf4JwyshnL/n1
rSGTfJO/3Tjd5YvIkYI2eAPFRJGzVNhPpRLkTc7rf/ysyp2O3Tqx+bCUK+3Qe2dX
ODCBZGAD8ypmaSgXnRAfc+8Xt2T9Su2sRx7usXP8sL/ZUtvD0AH85VOfi06FtCRu
3+bUwOoviaUtmn9PfLldaimeYJIapVj4HpGR7jhIYFQVpKccsiiVKjFyYfeiv3Rl
hPpMKiNWbo250meUPoktZACFZqSqE51kgQhZTzxBZwbV89koDHd4vh9YNjKSFpAg
JVJEbK9s7Bf7sgcB5BzBn1Lz1jnmHT7ZaY8JihCOubapcSxjLGUORkVKLxMxp4iF
QhZilZKIYkidIvlLc81QkhgTMFPv/Seh1VsP37L7BL4FxuUwjzdfv46BAUxhtWCh
baAJKTAjM+cNNwaZ0p9WWQdTvsrq/8t03lUhpZ+qDRt/Q8fF35JiwYEQCybXqHxC
NPBEaGstLB2ZHkzTyz2JQCU5V5sE1f6E9+EWz5+KYJGUU36+6Vf4cbflo6Y4ql8u
GHlgNFI4wanHTuD734wThC2xTt6HJO+706RPqhmled6V9rvQEgKXSO5SgbJNR13S
TtayH8H8KOR9gg+HgzPB67oOFgVQdOxfvDBLKTvvtqcjyAC2dw7Q1//hqQ468N6c
nywQKdJqiz7EMiZOcX2ng6o36B6K8h6Sn5kEV/QkEZZkr0T/ZUx90fJv/cOo09Ao
qb01JBJ7Ygo6DNAwKf/39Y7xgG6IEOV+PxD5xcGJQzoPg6RabTdDB+RtjqUea1Ya
1Ale8yEFpbsGhdBRO60J3QBHLmbQuNyst0KIMyARdeiHdt2u2lNVx1xTbDrMsqNM
Nu2vPQFpnWjapgsTqvDHm1VdWGvbkPUBIR5G6jvhgeqwjfZ0VbGj/An2i3JNhcdO
kdYAG2D7R5lYCp8sPoEClEYNVU8QP91YktiSI5IhgJydcz9S7gkqfeKQqHlcrViq
SgEIjGE/LuESnjWh1kcTPBGDOwF2lyDhgFjd/Kmm3NMBIesiWnJtaVAC+bJBnE0c
Q7l05pFLChLEPMmMbe8bCdZ6gi2x5qGj+eWpVUi0LzmMQVzBfumM9DugQZqtHtP4
793NxK7m8cA3jgMb9GkMZiexhQtZiylarEdQCBr5jSyScP99G0ANRaJb2OKgmseh
CvLTvDc39isByPQSkr5CMLBG28jOYqcj0jZ1uuzbEudQdJG5G8hQSUELIZ5eRB7i
iR+RTD8i+5sySWgJivSaZp5FO/izivzbBQeUD5XTUEmq1QW9U0p/Jn8jWvbfL/OU
M/fki37p3TerDDehLEK4brzM7gGkmbQZ50o//qAezxokSihPhxJWgsINSy/ej8s7
r1r4+xNP09bXoqdeqhuTd/vBFsR32x87/1UZ9j5cAmpkGArTJfUkuAfBwaa6kkrF
WQC1bHdZlj0qNa4m9kA242SbYvzrC762mxnSo2scqx4eD3mE0ygfnZBLwk0kvNrh
BcXTlFqgMxk6cNJhkC6WQJKnTSNP6tGn9Tjz+sbiXBhouz1liKnkntFgqX88enqx
Djd8Ub3VZS4COVI5qr9PCZHMCBrRYTrxd++KMCdkts/G+hfGzVKzttODO9FK5MjA
rIjlD9uTlopqtzl1YgBAShubHDWZi9RpDj/5bUA0tuNx7xpTEIQyfnJ5/vLUwBOi
tg5zjBfXch86AFFFrSJfcFVSuydZHJZSt6+eE5KjUma0vqetOa0Yl4pMbTEW08vc
5kcKrWosnL1M5K8lMjacY5QwI80JhpYaT0jMbE2Wx18FdFJhD5ph1snew5dHCLPo
V6FBlblAXKSxb7gx0uMG75xc74joW/QLma3L/HDf6jnjjy5ExR2Z+JUQvptLqdaz
H3vgpGeV3II169ex96ETd36OfuQeVervGAA2W9GlKypubKRRaAplUGAaK7nbiijt
tqwLdWFGe23QBeENbbDruMdIbhHcJieHIQKgCetCwHh6q8nMWeBOsgNkUtCpuk+V
TF7SwldgDpaeP7EsEHsUIesPyXYGXA1Dnr7rt4aoTNSD85Fgb4fJeC/Gh3W8pXcn
yDi0+9HbpoxNuIS1scx7YcEF3r8WFEWaxnq8x39XdY3rLWiF7ZgNvUZSdi2xrrdq
AjEjnvnxweo+tU9gGhWsVV5y5TN6bD3yZ2H7S6D4Hg6CI8CD4vpOLrF0GGuNZyUc
wrSOAtuHVbnZ21/0fk7/m55ubyDYRz5lU72Xh8dY+XDsXTPv0S2kraNffUvO9Y18
BVo8/W/QlMtxbs9zt8jPgBVxNaYECzC1BJ3sFQbbc81fUH9Ki3jiDGFv+ivOGRnW
WQmuSR9Q4lpVehGg+aYJqd3ik++NbSYBSVGvDRXbv1ZI86SiPwXpTXSFN9PPbhb/
DDJpJOX6xslc+Tz5qM+9rU+C+PBc3eAOokaRVN5N9CK8F4dGaor9j0nuD1GAraQC
f4ncRBNfQ/a7iDlpNoifccXlWIWYCZoxPhSQzpnB97A7d/8iobZ+w5egZYXa0zBS
DrkIxkEAvX7JwjsrdM0PibxD9RdoOVr+eZaKbcjyyUo0if5jj3rQX+i0m7UvY0je
WBCDdx5qGL3TVoC/JvoeX8erOgUsZSRIdelAu4u1+XR+5nc8OKgj1TS3bcejTHRC
OFWK9PNozJSgLw3DyCiyRapW6StTkfomX/wNT9gV0WFyKHrdSavSe2CDhkXoK1L5
AWrFuKdkaCGXu0Eaa4KFpYI6qfA5sPqRT6Ffp78e9lmRBXV16ph2ZB2kUk2hjTfQ
Ob42jbYNoYDrVwi/uWNVG+ObmYZij1EfpDiFqflfsqf4riAfEEMHZ7We7CyDIFHE
eL99kx1jISiffVpWNxwt8RtiAgaJwLLxoKnNCGDAIm42lsjyai2MYxpifvwQMdSt
ps4o4dDk+sOUMIBxIrUXYycSZWvRIbVLBWeLUZN1xGGxW7UtgEtqMlCpmotLIpAs
oQWw1rqh+QYy/X8UFLx85iesrsf9CY9Dxx2Q5S6z5xvKLLvB9v/zZFWcX8uwJ7wf
3Kv7NmM5t+rxklkRA1BpvAbFzJMBa1N3uUb0n1FoLNJQ4yv5oRffTVUIdVJDhUJj
oib6oW5/tJfOgUVZ19XFz/SuWLnrZ+fJbUThDai0VVrX2Uz3flWUbi5dMe230frt
zZrimEMdGHdBRX0uptqkQqncQN8BI0k8gne3TPbS468nnxrGkohYYFpPsEYUmL5A
LPHy68morkQ964AlMWgY6CzmLNxLVgs32CTc3WIG9xtOCtJBwpcaPfCglcbB9Rk1
VkZ2WMHjazLtNx+HfZJi/JCF2aIbi6lf6FRgOSNrwFTOkx4mQxP/+/CxFvansoKb
RSkw6DIlO+tyN3IOrMTafVz/Zm3tn8BobY45izQt1di1qcw6ukqfuERGcoRNos9P
fyFYvCm9W4YIhhTOpfhGGEaXQ9CzLYPNBHJSWMXN+txqD6qyhiAxv55Vi7Yuuh+g
6ZDerJKf7F5aL42SmeaWoVkCURiwNw05VS+r52Tq11vkA8vluD6p3EPHFeP5MiwE
X6gkTLqrTRGrpexQQoKFljaJZ/vac9prEJ4ssgTg5wshuHpXJhFJsjZFawuTJpoZ
DV00XvfUBcVgWH5S9gGrl/V9VUsP3U5IrAZFe3D5AG8x7vuNNaDmEplpZdBMW0Dh
maqot9Ofus4Fm2k8B1PggR8hhsDMIcaDy4YozGSsWda8f1PQsR/nhTggrucDtlx5
yjyedBmEeZzVSnQhBSx6Ck+L+cxgXgS8LO4z6wlKWO3u3xmlBLAMOgXY0maGoL93
cboLWhMyRDQeFRxpw+NQVsVjnhYWMD/IDgakj/ReU77Lpc80jqvK2zDRc5F60lS+
EfKVZWF7u5KFy4zqArWZM9p9H4qxsyHMbcncJUuL52FQNCS21FA1g/WEH2x0fxIY
5YHQDml8P2QnD+w3mhRv81kwpr6+t3yLztTBSTJILJjqOFApQfYph2zgADvIDVLW
v1boOwq7K4iQCIbdTtCTxOIKLef8ylHvmKRz++lmWUZ5ZX9OTxx7qGQIsBIi2sKt
IeL+G/jYAITUDFoCE5ZuvVhCQ20nm3xj3bzO9WHquFKudv01YZUi6L0T8oyyc5hL
vKPAaY3TZQQZktdrNORGMVFIz4qlhp3o8ZwITorF48nEcKtZUsTxRMqAQ23Ug01u
gIEHN3WMaPCAYhmuvxd38eXXA7Z5ovvv2x9/cDnAGjk3hjCtlZ86Yd7A1zLsasPt
K6M5Phd9FoM/4zvdctNMt8kW/Wz/655pcpT1XBzZ7rK5P5MNSQK4UyqL2iiL8Pqr
7ENKxi0VbOe3g4HleeRMY7hcKFbHwwt8buSvEpa1CrWjf8433J+yw5tgjCfuogK9
5KoaxvpXS+h61GQ6TpCE4U+xbbXMCQIo6yerVKTrIft9cX2vNqa5BrGWjapxo76c
JXqhkaew7kZQ2fb91JAztiZ6Y0Z2V2+cboFU9VXNBKSyFz59UlcxTsZ1aIuGr2bQ
T6JovfcgLyYng2pZizavyjuHSoEqdNc3L3lg0ZKs8XRRIp0jGtTAHAR56S3wj6sV
rFvxrtj9aRZCu4T/OF8QaIaGp8S6Yrnf4MsbwtqaJX9NhXfLKbbWgsUChdGLmthr
kAHSBHUR8pZ3x3vjplts2S6NdgPBiVDZ3S5qvFJoL96lN8GMCk5+ElR+WYTKXLfw
o9egaG+gQLs85OBlv3QHHw+nN2vixemz0mWcAvFScZrPKBbwT98doPRHIttUufSt
J493/TxJQpOfAB1VwmlF+CUbLfvgBfl4zGTJii86R+R9fUfL9SuDtnYqHKhu/bj4
ozcqjDXIKcWollB5L7tuRv85HR3TwCppyn93eRBz95//9w9Jqy8+hCUAUxL/sZpO
qFR8awnUuZkQqyF1gRz9xieYZ8dxD9iWgcKa/VXG7Nrss+H/MVcLWQHPPv6j8dUM
1G5iOeI8/6YaPAVuY59kH9NQKzi8G3n9Lrd75IldFt00GP7nufMBGsTpslHg7n0V
fiH5uSmAn1N/klwXFU+Qfj0l1/2+4gCT4n8Wm8aEQpvr1H/hnQQXvntuSbdcxzUA
1AOAC+DM8HgQImltJQsXRea4jWl6loq+m7mKetQW7VK+XCq/40AXT1U0yal43l4S
KcUyzdrrHA7aRitOr4vEq/HFwcaCZfWxIp/Um+4HUFBLLFHI6rrtt3fZnMSMuT1V
rXvvQ5BQOlBbGm7XjSTI0rba44+sbbreYObzpVnVBTjLg3FkjnqXXva1La0NfUAM
Ob/RCCn+MNPkzGxaa0PqURC0/gJq8mR2cCtDumSzdhxJ+na+O1UQLlYG+ziuheCl
8J2ALfEe5zO1w8yaJk1Gj6boM7bSc/cEGGwagM+s+TwN+x/WRjuVvO9gA5SuVi2B
Zo39oeZ7oUguVXdLCarQZ+32bBXs36TWYc3GYe8tRvqVr4eDnLnPGwtBdnM9cYye
Nf/0N/AsNdOn1c9IrAW0fBCRuOmZ1zWnh6iCQnn6tYrmlvnXIBe3P5wnKjcM+qSX
Kdc4lWOLE/qNKsJN1n8Z1/SMz/npfgAo5WUw1dzZoJpywg34mf+mKhoY+qBko5r4
tC89eF8axLN9mbzCF2d6/8pW3s67gQvOfACTaVZHAUW2G8lxfw1UbGx4ZURLigSc
OubuF0JcNCWfz3/rokAvjRy3zr6bAyUb3A/kKciaCYabtDgN4M8CoxiA2GcrjDZ0
WsPZZE3wOdfbvPxo3ykfjtRZhqYA5ktThMwrD3AO+Nwb2fK+vseXZSJLxR0g43Ri
dNRuGtxGTciXGxnbAx9fQzY76srWiBl1oPgoo3m2cvN05aCbciEwt+mL3K6wtXPw
Fe/pY1/YXeT1LyqeW9Sf0VI+BpQg/NDbZA6ytFu5gCjO7mJgLeDaGtPRKOBG6vdc
WmPhwiswDxDY+RlPc39okYZxH5iivz+HrOreo6FkRFXpHUq1+zpaZL6Vwxf+TF1Q
AiRNs2Veb/uyLTAKvgmIJYzwlPnaNQR3tInnA+nn9B98u/XKhMdyAPUmGCgP6018
xRadzb6b0YqY4jaKSjpiQz1kRQL5a1hOAIiMuiOZRDcCkYi8xTUgVc5riP1r2FMF
cL+XxXdcyMM/+uKHSGwMSP6tHZlMx9y9qypiSv8CQWH5fVFlIg8RFdsAbqg1xtzS
44BsyGuo3sq1JEZareTbWlAnwA1O0UxNs5FP+8UdAK7emjAdrL3vf+f/2PXYL+8D
bgquCQ5wbMYJwzLrvyuF4CRAGAHmJ+izITImT9YK3lq3GkeMN5O+FULw01stL1JB
h/cbyH6Y3nh7E7c8m9T7XXd01m7Br37+a6TwQe7aEET4cwmnOj+JNKKTpL5tHrOD
G/645zu4khsROKjTMiFD5aNbd/FHK+P6RazGGP9xOInL3XDlEHdQG1mA5XuoEBU0
1KWoz6Q8efh5aQ9/pnqqIMIaCqw9R9eKQRkKm1tyBqhzf0QGcyukXbB9ydK2eUHJ
B9LuKUrIVZrG680F1bFUDy+ZoegTZMGhqZOkCH23BBhYET7o7/ZexRvg6rQEcGnZ
a3CvXQqlR+T5NS9S1qcHoja/YLUcR8V6dA3On1dABpIdDzAHkyiYSzF4D2pW60O6
rt84naABW4QCDfYsfpNDAwdqwgcWJg+8gz8t+f8skOfQ1WwZwRXs27xmciaedXyz
LVAPYYI0GEqu0ZPrFWfpzfqkyv/nGXUSDvp4j9mDRtiFIIPzI/6zDYejr4Ay8fxA
0yTMRS5zXpIWsegNrlGMHPE3GU4mq2znQpQ1tvM1vC/IuL+6SNA3lOE3u7G/SJvG
KsnvTEFWLRWFOuJ/S6mRsmphbeLSrwgjNvLE7za+K+Yr3LC+FGEIKKWNkBjw/nGK
Wr5OJtqUA5cDyyDoW1P7J8Zu7Ph48D2LK5r74fvCJJ+OJIx/ctQS9HaP2vhKI+SP
uTFvC4IKFo1WT6QY4iwt+xlpdfveLmDuk45Vi7cudC+afX/b4qOcuEQRQl7wrLLC
1D92kUVgzipPwRZq1kAdP7Bj40QgmYWpbR5O5WNekfnGMungxZkW40b0ZBVOx0H8
PnjSzc1dhKLYEiGsszelYcmDFcqrIOyqQQ/H35UDc8//wbX6YTXQ8Rma3yuR47Gl
HWBqIxHGzouLWzjF/gHxM5O8Hep2L3fdLsL6mO542Ez8nB0nuApJkX+pl/eTx312
3h+MCh1CbpGW0m64VQyiiq45OkF59LAEorPUyWQxiM7wZMrUcoMgWw9SzezigH+U
t8yIxHu+ue9RfuDMQ5grb18bt4wLQnI0R9QgBr9ZOIfQhu2lgCkvgnLPboc2UgNj
3B9A+08k46+bDCfhFIB2suo+qN6plG3AYGykjbiCnlFt3NAPM9uf0KFcZiDBj75t
yOvysjlQ8n/LUq8TfU+oXW0OXwe+pQ0HLn4KdleYHfeln8OBHvmbt/ZRMleE6qzS
L1wiZ+N29kye3J7xeaxT9a8yY79czc0qNBA1qhXYrUG6l6ymyii5B4fU4hUxivpi
9+OxPD76UeDdZmEWnveSvRhDlpObmxybutI477T7BxOUl+DTVIBkovR4CevO06M4
juxXND5zXc4o8QD9EoSdLejgB7qwnj88zex1KN7pD1PiQjRJs8vB1FFPaMRe3oee
yDa4Tr4f4VYMJQaFSxAONrmBWsU/ga3jabQsUKVkXqE67OlGAXijCrXI9E4meSSJ
nj+6EhN40HYUxbdCb164PsIxB+nVvcTkxwY798hAokdrN3Y2RcUJrBMTAYKNchb2
pfkXfF9uSavpsTwdYKSkg/SyDHYU50umXQvsQ/j/GIdd5dY0FAAQrmGUh5vDyNVD
NEmZLRIiPEqC3pARZJ8jZPYG+JnWCydwpDiPXLB/g0yjsnv0tJ+B4g1MF6JqjFud
sYURNgNwiehEFWDQHyQaKalfvuHiHH0iZjSCy8vJ/hVf+GW6GH8epUi3Ykvtouln
IZJxpWduVxpxvTV1wEXwi+GqIEa/+3xOfIGMKJqGHUmk3Avc0iQp/TQu1HieBJKY
Azw+F9cUW/JY57qbUDe6pZeFt8WTr/FACDDkq71lVqAH9p91FVSmwqQPAOEj8A/s
GPiKL+7V+glAckcj1wL8QydabwxgkpFpkmp65kOE9vO9yOBVoIc+fy42aZUUTN2c
LMEaXz4xjO3/8Yx5w1jY/1kvp8Ym/lHLjx+uKTyK8U5d9BxIdH59UXMgOmvUKi0v
n4n2L1nCBuw6rbLDK7GNdw2xX2dsK6B4p4FcEkxjMAoQhXZDT99AaSrICv7Cs2Li
R04JtVeOoimV/MHXkn+6duXwdtU7qVY+MXz6+utqfRtdUWjJ/1hxDARjlNThg/x5
itQg275G/4K20hv8kKdvmZw8x4tTn+gIgWZOVvjydlTW8IPkCmv15Y6ckl9VOjJl
/nbLQd1zdghX2A+Wza82zrq238bd+zfw2qNvf3KN4UhVwnJjxoif2cTbhgzLpIfl
5ti0bZ51N/Wa5Q08uPr703PbtZWECGouqh4bfw2fcldE9Gpp0f2b1KFXID33HMqW
2RxnrIrfAP56vxDx/I422YLwWdI8wSZJjHzvsSpnbKrIH+bU399kGAx15jbrsxCv
HdWzQ09jxHY3/BkvVoDZnH+ioMNwEAQz+Dq8bZI7Qqc5fNmxExJHotdd0zAx+whQ
q5Z8CpUhYZ1YoiXBcNn9A78Tnb6o7kYAj+vooRZPOIzmnrHFQYtWMiieCWozYArU
dlPhoZ3AiIgkRl/q4Cf579eaJml/tOCCvLewUZHhhNrLvkiCoreb8Ib7l1NDxSOr
AHTAV2x4abl2ozldsahacOr8Z07AqSCt0c6yrW9TZkFRfCRgFW3KuheJUEBZWi/u
oV+2M9lZ7cDl/oXUMrGmoKrGvykcI8GjBVjPwDYaQUygqPqJSimvDKFrDRLDMCrL
z8Mh/sWu2bqApvwOx/uPKiP9eFRvMbHYxCNIC5/072Hgif68iS0yupUebvzchfnQ
FthQ2CB6IAAmYVYowp2K1g24DarMa8NtNm0/QCeopXazEqvvEPMsTreB2JYmjf3S
iYTvCjpiiL3Tqn/NT1M4m4mbCilA3WcG5WgZEtq9YIet3TA1aqS29Ie2uADE3jNS
7QNXI8PWfcqFXOkyQ1soknc6iiW8RHtgFaD3pAUQM0pOOXUFq0YDJmEs7wEuMa9z
i42p5pZgJEm90ZSTQ+H5lyCvUPYdzLMbPr5sK+VCKk/6s0i8wC3xESYAZ8o2nBGh
bVt3HxCpTa54aSLqPid3k0//XN/eeRSFv0piglv3EF/O4NAYOZaAHd2xEkqyo75H
81qKdzI5TfXjnQYG7FWQwouak5Ulzz1c7tp1mriocStUDbQxR/1UusPylp8WbGFz
EJV92m8MFRypQBQaNulh+JS2wfOaH4N1b4oiMvVNiJ/DErOvmt2uj2paZafT9C4g
FhPQoaE8D7MtSxHPGnMyW2/v6KKnnsPk4HTkCKKjEFuFkrbxVi42LteOlFiEElrD
3BMMgPWh9gn9XipSrsx9YhhHlsJfJra4NhjwZrh/KlSf3eaZ2idkv1tuNws2ZiqR
pZvhE6iXo3gbDZnQCjVQUDU6DwXMkb5M5/2vdBVHxZoZlwyh1FP1vT00hD3OsrW4
XAQRfnvUcKcHabUbP3kdLBCpd/z3eJ4Ih2ZNpCW8qnp0JO63hjSUCQioPGAY8eKf
g15g9g+44ihfra8xtwGUDNsxXiZwUORr4R5EY2gR4NhT/m40CEDngJqRQuXPYwYE
7mIA3krjUt97RcWaKsngPdlwcrawe6sJH5kiUymCUJEyg7LL9BB8qLzpGZMPNgjh
gaxClsTyogkW/XhbhGDS5iBszoq7UFhkKAHxcSEW2UeTXnmZTamgpJEeBp2T2lq0
3nSsKknJcEQ/h8o6zhIONOMYPHL8yIgdH5yWhzDIqFLgl6w8DIRvlZ0ibM+2l+E0
071sEnoklO8JmoUu5oAOxF/FhY4agR93f+IxiO2PAl36LyTom0BknitXzfkvx3c2
sMI46nJoq2JUz49yViom3Ez9P0h57+QXyO5PAFtQPER9apt7LcM7n3J1Fr4mBbwr
RzeKC1MjUaLUhYOI1dMFgKTh5nve0k7+WJJIxY3hbM5FXWR1CcdSr8DlYxZ9lbmg
LaBu4/R0Ipp4/Nb5aI9q3ZlxQ8umww45fVWOCabbe/nwJ0NLGqlf79FkVSl7wI2K
QKLEZDN5zVEMZyhBZVG/iiSMn/Md4n973VZaGTvVExP1OGIKlbVIONwrynUj4Rrz
xS8685QnJkrAM5iq3tMgh7p3TbArBScYZc67UxO+EYrJ33OSZXUGTFhtCw39wWQ/
5UtP9evZams1nVyvns98117v25oEBNqxcVJlqBoZPYNWlxrZxjgZ8+1KJg6kML/2
ihh9BrMsu1FYVbCgEXUdauJdoBYLpIgM+tCp6fvIGnGqNUPkQYnoLBLYM6bSaIGi
vm6uKU3Xa9CE80k7lh02x/Qjza31kRHCQEZBPATWHhSSGWeeBGMLqwN+5z3ZrQdA
wZ5u7jUbTRff4gjb9yg43VvIUPUQ+8EarT3xlIp4Ce8eN8TbeAX/o76F9zh3N10U
taox8F3vTsAbutN7kOHJthi3PBT6K1aaVk8+MoM3uzv7jUFXsAda8/rwrWnLWoUP
GwtispcG7xoyS8JplRHDSaaTfdYk5vdSl5OCqvMkdYJ5xcxcHbqR2P2OkgJlCYo5
NaDtttMlUU3Bb1t71p9wMQryiG6+SuZeLZWyfWAkMSOXSxS8kI+dtOYv8zP25Lj0
iXScgp+FjZ3gfJrjWKE05/RHi+rh7I4m2AvLKEmPFM0rDysAazdqxjLQwGniL94b
Z8TLt9YYI8afsoopdSxtw6atB+mxk3el8Yh70GYq/mZUyfZOJIbDMvrMpL2mnmTn
DZYHYPZ/nlt91KnICXTmK8YwoOgOncdMjO3uRUW8ldtzwdjFiDjCgEhMC8s7jcMs
tOXZekjnWKdmDQGPhaiBt7OApV2HnuyLpam+Rbzl2WEJoS3xdKtbzPLpwJTzJYrQ
ro1usyHYjX5rkYeZOWIVyqn/g+XBJNit5kTc0h/ZIxGzGpg+8HMOyBEM4u/RTiMk
mIRPuRUxG5hNDoaNmFd4GDn9HDuSvwOI19kAe7R1nw0S3FqKTUksDs9yQegpqVJQ
BCksv4Q0iphmbPu7QjYwqIdZu08bGhrX+DkCoOJ9ahs8G+a+KLblLJAlNYqgCk2G
CLBAnA6Nar+fXbn/RTahYg5n0S69feT2l5zB4SihEmIE/abNHl6WVua9tdHorpOK
Le2giaw6Hf4kXFbnHUTKhp5h0J0/PXoaHa7UdvekE8mDdoCsT8eSOoYLADOqwR6j
NFgNNnC8GRcJYmcDEXlPreUPbZ7KiAKqPQDJLgatkhlXXbcHtYgoKCYfGW4ABOy4
Iax3Tu3QZK0cIwSuigC25o35q8eRPumxiwHLWZEyVSmv+9zprVzMACgdU27ZCiNs
f7Fb6b74i3dt/sRDFQkRcfX/Qve57Wa6HnXAukX4vFvxOSAkvLcHTgySOlpBP5ZX
uCzLW2ZyOL6Zdht9Lrg7ghFd9nqaShS0RGO0A1FuqsdFFIHVs47IuIMQ41JxHM/q
RzY/BOC2oHpYsTqNVcWg4uG+u8MnYFc6aqUQ2JzItVB7yyFL7BcVX9T3zVtz34UU
+iXp5M/AcQTZdxJDR9rNZmw3dFIr6M0/JQzIBod/tUBkHlmv2eJQDv/r7qVrhno3
ZQKl29qToTydyBl2eN04Hbl6lqH12VW+K0AYXxS9MWXyeoepN+xNg8c1hCgA1TjO
zgzrgZCfz2xSVMlY8Z+D60gbn70zmqDbk6zg/HKdoLaxcm1FC8X/NawQdF3BWju0
jhcWTE4nff0fh/2bW6/s4ZWjkh0MPY4oeXhXYn6HBXmAOl3xSjK4ewXItoijYILZ
oU+JyZacBvNPq5r006UzB+IcMCwXzICoO2+ouEMV0ImaHSi82MF+mWzzv7yB9NyG
s2cwVd6Xi9QE8jIIntBwXMUQqmxi77lJEJPGv06GQKfpN98jrWJK8lLV+Zq5Ymsu
US7Zvhhgof/gvazSeUaXXXxceRcQKIj0nxZWB/fQ1a7kA+cGt/3j09+VAgI+HZQX
t7FyNN2rGUfbyviZZ4vycBxKY6hyngzHTaUbIGQCl7vaRNlMIHGtKghTOlASeCAe
YVk/o5KUYBJlY9v7E1Ya0El9vwiggJHRmZEG2YIa4jgc8QBkoi5DdicsDT3YTSMu
Gvw5/xircgBSrlcpvXJtmvft0Z9RoGYgs9V/85dH97D7p9VpMkcfESQcrtol+hoG
c+yWZXgfwfsUjp1i26Z8+14mWregEkQTDlivAZhnJB0E9wqQWMNxAcEvP2YR2/TY
/h0fRf+sEcl7yeKASWP+5mmJ232w/dwDdIrWs+Nza4ekOwd0CxoGSqIHCTkEZLvA
zymSbqCKjNnLUJdkMfPMlNKjavG2tXJVulT52bOh+KMkIxJrCIzjjcmlgiLTScZG
AeBs/4g2OsRj3vyDjs4vscU8BVwJ/eDHjsK2H1Ah7+fih6hAW8UJVHWCzU4xQAjo
j79DQsnxNyhVe/8f4PE8TTdRjEc3qm1nDSt7mP+R1x7t07ke+czKBZZQV4lgZWcS
1p9Hy6jh6cUDK+dm+RqHdok6IWWnv85D5S78l9Yzr19z3ZuahNk7haslE10Tq+H0
v0OeFgLxr8qnkqdg4ENU8HuXlNLYB/7D5dZr0WWzdL1wz78xcHLdoqfinx7E9yRy
lXjsVrBQOrAxr93z9qoY08SvzIEGROYnuZs8588S/U8EI2hyDKhbBKVbBO81cmGU
zcxHbFDqB+EEYUfqJgrfZ5obaQelzPln4x1ojeuMK7v1fykYLNkp10EfXeNN8Dwy
8IFBa7q5pzcP6ZC541Hq7kcwIjfwZxo35Jh/0LkSFidcv3ET4MjFCjAtTcCdGltK
WPMEyrYuusa09PJXz94qgb0Z0binnvDawKs8PVqDCMfXYu/6GEf60nXoiCiBbfsL
+Ch6HNMy/t603k82gUBcRA2zRhEKSc6cGDq3QFmuVap89CD3r3nPCrEVMeW/4vuG
AlDnLpvMVih/IfXTPl7dxUnr24roCSvvKeLtP7S+cremL6Tn9Kqtgqjnu6BBaFLL
IcOo7Nj1zwt1MwLQI82ototLH+EOCCH1PC4chu6JwhlCt87koDPNwzPBH1SeLOwm
dSSLxJcYIbYckjSZakDD9f8X7gMBZTSDuzegjJHLTwdNi20L3CXCTnKLWvGx+jrg
YC4plPRIoKtwwcIXcdLiM66STUp07coT4S/cwPbrjbbnkG18pxLiE4qZbtmlwLeC
H4we5uOFMsY69CpmxSZ8bOrwMU6gKx18Q4xHvyqEo+OLYpcOVtnqdnRHFQBRF7hS
zXy+zg4abMHj7ZoBb6lQR+6bvt/59Oau7rl7wO0o5gYZuGshJE9x5zRbnYYwnckX
afqkwwEROn+9u/jk59Mbelgtg9n5BHR2D+SKKczFuweNfbBGr4QCFU1Ba32i0bXA
YYicgNXMHCLCFjsd4LBy7767n8N0OTVFzsOTTlPUOkE4n5A6nVETeNN/Z0veFsHY
X5EZetxj88TIwF+Rv78wohP2Nb6pKOwpL1pDuTaqir59G0MQhW84Kmcy7zGjmZuG
DVH37aTdbpC7++eUhIi5K4qLcIA6cD+h6PG8JtFQqxVhKyKJRWAXcj6r0v3izWfL
i7RPF6ene4tN1apBXbaBQfPPmFvjlnUQsBexAGRTnh9Dp8esqxe65l7+rFyxnd/U
df4AyZdeVv1MWWVjZg7ZTVl9OFOX+2qb1kiSUP7FJ5c3K+VrUspz5D+UeG8PUvYQ
fyXVS9jqhs+gVQ8K/KuLG2Ae9Ina5pY2NYg0kodc+Zpo8YCS7snzyT0Ct2Dq7sPR
ptrrMiVEJM7+XjogoXnXfSVvzEsehtLw0ZX1sGC3sfZbOLpfff5WYRdZB3V3IlA1
IEUe5Wjv745BE66oejYqT2/787yF5L/FxO6aercImw1rxyJVdPLNKaHryFYmqEnO
W5HMF3TKpzXulkzHQBak6QFY4qz0px0J+lYOITh8VUlehOa/rMD6dDkKSkf7oucJ
jlHmaVApm/7G1vJyT97L51ge6jeXLBBqv5TA7IXCPiKcEP8pY4gkYPOpF/Q3Qv46
D5CNLyGrT390iOWq9xUgBrMlBwJvmIc+eaxzEuk7ax587tLu/7WNDAtvqV/y7Tjt
jXrZ84j09oKjGzb9+1IVi6JPkfZ3u+NW/R0Jhf82mc0d7xtrmYeCFFbRGxhZIeAb
L5jzg4LImtsBY47KLO28L5rlEfqfZIZ/hlxaSeU3oMwHtfvhjUDCkN1o0qLQ+5EE
BUAlwqfjRcjoQS0zOPPveBmLHkUihC9jevGV2sjF/Zh/AVqH5+/7QrYng31008m1
Lf8PRj4Tlz5pN7sMVg+DZEoczObr8QkbhNPIgCw+lyDLqAfUGlC4ouBPDe0bkyfm
vkSujlJJtetLoqsczk1Ptu/D8i9R1NZUYah+XyI9nIedEFMAXCqF7BmKHyk0r+uR
0xhRIiZQkEQwl57KGKqbG2SPW1Hje8ObOK87KUa1mdb+T9rUvenu/fWwHCxPIqcE
U3mb86/scYmEuJNsPr4nCW8e7r7eJ91fle9F9gXudGUoNugBjF/OzYuzBNHd9C6r
/gxxVWS8fwilcH3AWnPJG5IL9cey56iWzQyaGfDTNbvfZh1Q3BrHGZnd+xeVTKk8
lGz2o2jLOIseuhLDod9iraKuS0NSP/eV3pwAZTRuQaxGU4aqguENycHUbKUJRMoq
i7aIRfVIHCc7M2YIOO0Bz/drx+PlhlbngsEMq4vYo2tp07LDhyZDJEkWsK07Qsy5
KtaOV3OVmVC+jIfGuAgn271xNoKML3VX9+gOM2MVRAi4ja85T1JaABEpIfAQDPoZ
hibiDu2vpPtFq2kmAw9CRRI0siD+g/Sl8fGHpp272xm+3JCMra10zjCyO/286Ie2
PI+p4iSiQMlWv5nSwI3XNf7/MabB+Zi3YEO3UK/9v/tUXXgOld1RoXYqWRD8n6eW
9UH2hhQfLdHjojAREx9fK8B1uPH9IjBkBVrEbKJerlg0gdf8Z9BfbzyJsaDJmFdH
LTkb23ql232DaK7y0zxt9vPzkKc8bXXtwzrVpZh86aNhqO6Y51qtJ8+yA23MRVxq
ClVJBrfykunzamiDx8QLTBIxeU5tHIyaFF7UKqkn3cwfR2xg/sE0g00XlsMUMnOj
7j4Ue4P9FphS277v4vJsTP80cmJnvK4Ng602YsOuQeSsve9D2ODmoU+sew2+GNnv
LB6X7u8bwS8mPhFXn7DwbFj/+hqZzzZJdb3pixJex6hUIKYUMB+xbwVdQ5zr3nDE
E7yb3HgQJDd/Et0X/EcSI5bSt6oDwaZ0iRrKiDlM7HgEL2C/m5AJgs08XVCXeoL/
t3xzsO81u5/n/7wdrsunkX5kB4RV0l8Mj0wx5kvPCXHcIxJv0uAOZv+dTI/p6Lo3
JmjTcfTP5wERLu8UEADRhFaqsnxENzAdGFTIbh6TXWz/8QMc6U1Vgj1Yk4GWo8eF
7i+XrXa83thjn91wHRcstmGZ3O0o1SuWbZ1Mjyj2P1u924L+O1eQiuWPB9YAWByS
BKwKlrHAThQpIAbcLw+UR1vR+paWSMUdDriXbBqJVv8PbUTyx2gHGtKfsPVuia1t
zASmucEi+LGrEiPj6dj4EazzLFo2tQnL2FSRHDmNVJw1O2kdZEDuXTyKLnXtvSSr
zEklcOz9bx6892sREqXChN8hJXfiwhiW5gA9Sfauv5dxn8MdrcnLNRDlYStKzDho
TzqiLtFbdAZRoE9rLi5tjDEOh45y3HL7rf2RuCSWaSqhehToDQAOPT4ZQlHeWky2
V8bxkLEWm3u0NEOFzLX0u3VCQ08LLwsSRuwBM1Kv3sIwuJLypr5Z/xLYwvkEws6H
xUtJT1n86zFZ6yd8ZbngWmxorIoQ45dCAB078Zmw8JjcZTsccZPsf+e+Dgi+M05A
dfE1bHuUoQRzqr2o+LF623Ty8nk/za0pkaHBQ9RZGOLFpv+7O+TCyNrhKqbKFK9r
+9n1DS7Khglw8/luZJD4KyxWnaeYQrRzPubYUZSQWACge9RUBHBazYMc0LsAEkAB
bTO0VBZgs51L1LHB26idyT/kYPSdubUQ8MS9ZKpZ2sBn9LvwPgxLGJBUnsLTQ/P6
jGdu4qXn2KFDmsBfu2+ILl2sFETEslYJWZ7TlLrfGcUKmrqaJsWdJsORcT2nEIM5
a9w+VaZDjF2d4eDdM58DRncx50BY+C2hxeSg86o1AGYTB8DAsIJidab0eRsdEb5Z
rmaMTG0IJqnBDXU+B4alyR68735LFTuXK1zThyqm/aDIbt3kFWLbWOBWJw5aSrLO
MrOxz7momnJbVPrAwt/LNkqvEl1E2xrESomSmkkglgqqmmfJ7TrWY6WjYJk7NiqP
vyEIJtOHyZKBMqTykpzO/F+g0T4T06Y+yOSWrPJVXahU46CbNBT3mFtwO07dXTGl
hh8AZgQg0CNrQXJfoFNzi2bQurpm+VINwuZtitdI240FdYjqqM/LVQu4ocyZeEBA
FuUIbic0JfxVjTlMtZk2Uv/1YLiiAJy6AblGoG8eq1kKH3VMf5R1V0mJXbDmtsRt
iz/IC/x5Be2KRGiiInyIkhHHwSS2KDdVOOzekUoCX4aTFp3AATM8wVMB17gsgF4i
Dur99PXEt15Wj5znfWqcp8XwuRqCbEAWqbNccNIgvCyd/D3DqPPDaRsuqYFnl77w
f3z4cpxdK090tVTGktS6xOdZPCLBSs6u8bTgExXA7QVUb+gGAoOeOMsuVCojnvrp
yoHdMtK1TBxFim1o1q3AKhFSSOHgfU1LLydDIbs087dc92F+eOPbXFTTGNCOG35I
eZCQHCTz0Axi4Va5nlJr4T1bKz2LW+Gpw3hx3TUjInB1gsqQmCSeMgecGOt6+uCJ
khMP1lGnTmdhQx75FewwTuyGJX4KENPI2tJtR8VclkRS1r1Br1yEoiSHAdARSKK8
PHDvJ1oN8UUB960C6wRt2FiUeej2fitCiFa62b1HKD5DWc1n9iie8Cfo9I5765zY
MOxXVQMMjbwfqk6bb+4P0cHpxns2+A6rGRBGtkdhZGNE2COh6x0qzO3uLU83rMo4
YhMNGI+O6paDNmT6uPiosDesDnz3oH4NlccB5U5wKQ7Tp2a87qFdM8fQfybbOPln
A6FeEp3AJBY4Dc4oAa0+1aVm2i3X7Cxf+YYqJQKdKlu+5SjLS0q4K+E1NS+xYFSy
UqTwuO46H5w5QWyZL0tbGefo6Uqsz3fHt4C/W7qUsrwI/8fVoDMqYji95Ayr5DNd
nvDwSEBC2bK4vTHFFDUWUzpuHFTSZ79iuIweBiJNIl04XCKw/9mFEXYHI4e68bTA
LHCAzCU1o4xtL+s/FSMyGj32PhPaHuSHN0W+PNmj5omxm02elzwcNo5fjEJ7neGC
fhYYtO0y/oYFVVor3v/aIE7IaF4wOPWtuCEXMVK151gq+r4MxCh6aVcVL+NxtjKI
L/fPU6OeF/rL8pwkpPRCZaZIbz4thM4IP8JlHeI4amN9JOU0xVFbwyYq/sGHXpLk
eFB+T4xIZjsT8RsUS6vMOaaTF3Wb5Hhe+JvRxvaAIxOAODUfp8DPo0AHsFvvuZEr
zBQifdXw1P9qi/rc3WOOVLG1j0Qx+JNKZp4jmKVynvNV49gV/EFfQAjfZrIQrKyi
C0vGZWZs6qwpKqi3u+z/pMTqpiE3KEJoxx4MYi/8wJQm9OiBLMnL7VnNZDBH1Nui
V9XYIbwPwyUxGS/5C0BlDDi5V0RClVj05p3+1xhoaKlWbYHIbJnWJUbyFanTWgl0
AtrWvXJYC7KkCqaoYypOes2zJV+akgnCA/5kMPF2AIeO7XT+hgP6lBmbLhmP//bc
NebBbf51ehEJh3l98AE4QpXZ5bDgFQKYbgAFRu4CoWNi8bIX60U9+jRoN/dYSo3k
S/Th469b3V45StPYPl3Z9H/a7HnVKLZqR0x/o6SXMJXFYZ+6vgY9iIy+ZfKU5Pif
1LAn/sh3oFgHNvhx/WnyNqrBo1WzrfFqZ6zPv1hUsNz7wdDGsA0Bc3CMfGv2albj
FWsoz2mNullEDBiCDinzbp+HDiUYJMLiU0C+oLQLi6ApjY1cAaerff6f11NFMQq3
l7qNfw9roSut0e4rLXjdsUfhtorISUPdCdvSru9RKATfjuGM2Ow8QrJ5ZxAnSl0h
Tqqy54xg9kmqD/UpSQW8ejGXN7O1wbYl9wzIqzpvYRsVRjcpvlgRkzUx7NL5yJeZ
R9RmF0DUuYQkdWLKbZ6IY1yn493qU8kgxNJbRl0vgLZnezz9boVeJVzLY1eHpQaw
lOVV1G6ke7YFrLIcsqnP3Q2C0YzRTFlSo+VjavrXH0ZTQ3oOe8H9xT1aFKWkNNrS
PwB/ohb8j8SdgFID87V0NghmPqHKWVlYvQpQ9BmcWqw6uOEuSnmlteOnVKsVeF0W
SNKGc0PVVgew8LIcXOeGuIyVVMt3kEQZsp8+WYw1vOawjN2FXVMr0Rzdl8dU8Z0G
EI05bff93rvwo5M9JQAZvQZH55HuN6sNTUfaSoEHJt23uP1mNVo7ltrokgj+Umua
Rutd8bfzG5lx8MrQCwqeWQ12XsrpBLIhy2cF/VjxsqO+8RUlPB3uKVJZQS9vrpTn
103F+g63mpAwbhZkv7ObjsPgZxXRRtlugqlsaGr2FQsfW7AQuesNubmh1LPvUp3N
8SiiyuZxJdNvDUbydynMeUaMgzrh0wm3DNP4VBRHf0JzBW5JkRdk6UaePRnV1uSG
p2l5lUCMq5F5rx2ZUB1mkDHsHsV928ycXDv7OhnO1W+K7jhgk9Qf5tnB7dcizTeG
Ae78BEIPljBv4Oc8U/5afO/kjiksyGK+76x2aaGorz1gzS4ePjpyuLwePnamRVKS
glWYz5LdM7fNnq36RRvXcjBIel4b0wf/WFjNolck73bFqidzyVfVGLUtMty4Ljja
Ewl7k/csERVxgFzhm8tBopR8Ao6VXhU03JSw8xJ7NoklkMvH7ZpnRMmo76eeBMgB
CI9KQIwRjptKdsCUYXl5s4wPIcqCRO4hyN27FYkdWyIn180lAu3sWXBO7nJHYCXk
rc+vPZt0RjJRuKpx0Gc9pRXn0dLeR+lNduB5qyd9cSw9ljeiM/4gXcP/B+hN4piS
TG8PpM9D+Qi/ASvfx7ZZSXhmWeyaNSudKeF7UtkHlGORYXe2tyPNNlkxhCtAxAcr
FYhvUzuCY83IY2ffym+1+k6OuviYI6fNCcZqeFotvNXRjsZQ/Z1RwuAAa2BmVuNk
TlgTnFz6viCPy/SV1YMD71ByKBQU+FYDEY0ZHKmFREiHOiJRzvS6y+3YdHay9UVR
f+HAg/0QBXrWrj/Ta6DT7oYpjmycVbfMHah1JhvY5DdggJWka5x7UaR9bFJS6Ql/
0x5KfD4/zUq3BnKE895WDqJp0qF3ysGfneoNlKLDpWuHiHrTtP4yqSlsBlVIIUWD
PP3gKD7V2isMBj548Qz07MUioW11Pkjb7UcESFgwkPST3w3HKknUUuoZTuew5ioz
dBchA1G8YNF7Rffz2lplj0q/iIvuXBxA7yzWnf8bin0M84kWqzF57aWkmSV+pVW6
k0gq/YLhaRa+NvPodzl0Bc09paDMiI7fQI32W24cbUFmvfLMGJTeq2EF7TWue6ED
rf4fTdByboKU62k6sin6A5olUlgbkqnvq1H7l1JlQCDKohYnU1Ly9nAE196e6Gpl
nKomYIWmlK7usv8aWce929FI8Nj3LWbOKWS7JbFodhSblyfYJB+9uvgUTrbm32/d
vwET3Ybwr8tNMqz0w1PTAnnEPPa1G8fb1vkLwbpCkRHwW8COuK8KH5BWNxUyHsly
Y6h4RdvZVsgv7huF1yAJKDy8zoovCu3BXFyFSF3cSTIChXGCoqPJL5IU5eP3B1ts
kywYq4rTJkJAfVSJg6SfPgBrEv/M7zfAoVt1vBKmU065nJLfTf6x30RQQpHHl6Hh
q4uiG2YlfADvD6NhHh6SoReDP/qQHJg1rXMgfUCmND1QGWIZsiDbIpmHnNlEIeBh
2Sk2rIqGRFwEQrMxPz78107/b60IbbB+P/7FRQy2/C5hue4ckXquV46yv5oo9KvG
XaW3nrj0rgZ1pg7nQ1El0Hued0Ho2KwkLCH4VVDwixhPbO4KkyFSd1qeum6zQnhL
nUgSTG7ZNPyJplraEFT7/Ay0py2ts9b5BF7CFn1kUl/DOUXCpwrtxEvu+UIbTlk+
kF2Thpm58oU9hyk8vtMAO6L0RDXMce2Rw7yr2slj7BMM9VYCUSEqDvwwvzbrN87W
Jm7oAwbw7epd2TwT7fiUjukmGtEZTmE07ujchzpFSHZSscNT43f2rv/mYJRl75e8
QRhK4C2Hip9Ep2xTuZ0/NgE+c0tr7DR4biMTqG6rRsXmCg6QojbvXjzy1oPH7iaO
oIANC4pf2y0ptHMgSSARmERKnxboOsygVy0zwYbYvntJuLn/35gd07hhXEnQT1ua
N4K8o1POU4nW94MyPrZkYZryWrZU7Ie3qxTwLFUm2DHwnam9kjGfyxYQymwZDzWW
F6Wb0BWIv+JdXnaA+EY35Dp1+M/sUagGLiuVm7DGw5wkX8oyM7TEeVa+ePZ+xENS
JKzlWAf9pjk7T7W0DCAMdBrYWGAhc7SahgoPImzy8eiEFi8qR3UqeJmwk4WXRfOF
HzDhWQylj1AN0LQ9qfUPxSvL/EtzTStnn0ZQ1Fs2WiDS5pE1pXyYMpKgWk0tjlkz
zGzQhbOMtHB+/aM7xmfD9B7DcmswVhVHxy+UR4qEa0NoiohghPx6XdABJvDJbrBl
RJuKGPnbn11Cm9lPiAJ0IyCnykQEIjF4bqo0UT2zCoelUHt/ePHtt8tLhmyK8IHn
sZgaJ2l8uQMHFtQUvcFVHPx5vzLo0V3gqBEl/I34EQ6PmqKJd5bWDzhrkgwxZhn9
lmheBjcpnOnp1OucKbUPRpy8ngUDin+AhClZjXkJyQ76cJ6wiI6GMjdkFf387mht
zwz1wIHZsUT627Xre3/q5T+D1W/DSFzjM1PLjSuVFQKdnH3Yp37ODny4m4TZiWUg
2KfkSqlY7gTB78KpJ2PYzif/52DbH27STUoNhoU4tY+J7Oqbq9nthTAGPsG49AWj
MyEVOjN3nGQV1rBodJapxBx9nAN9OlW1Fo26uomX4Bfc6pLbIC3yg3iRG3Y2u/ZW
TmQfBW6AES5xywPSHa+s+4FlYAlcSQYun8dCdwzibnXcL6IaDrvxRN6cNGv/Av/8
dWqTmlwPy9gBabnVN1GyDaFOSTTUSFaCShIOHQWoXrX05ozEtKCePsenrPiChzHN
/KbnYjTNOHEPT+felZEXtdN6mSbY3kulRJ51jcMpQ7GPvisNI0VgAzDOb8rh8GUk
o8GceHpdoH8Di1aqhbFuQLQnTCsj1t9SYq4IVcNWGJ9uTFjno0hO1is4jVsiS4qJ
SrjPYgqHuTRcRK16LkQ+4UP82rmj/S+4tyeKdFDn6AKVO50HMXBa1OqL3+F115oy
d5GArRz9RQ4uU/VTwCj/O/Gyk1s+iRUzU/jNmqd9gbTYAQG7kKYKjqwsAI4E55Q8
aUJycKwSzGqxhL61Arc6pHHaZWVazExk75xDlfAFFi5PhrquGTV/gLne9n68N08k
YUtRg/78gnRtBpqV02dRg5cq4HG/+g3XTnYwtimaH7dB+1gY+9kNWWW4UxtgyrDs
KGdb7H60pd0nHK53XwgbONud1TLaR/p220QZLJ5mk+89Jqsrrap/BbvPpbMn3EmB
VVMTzC8UF6fyj0el26UVh64XlU5u9ZLb83DhgILGIlEwFmtDsY14Mi8Styf4GGvk
24W5YMMd/3rUnxhlqNZqx6oYD6Mn+0og/feo27yTqTfHjJgWuv2SOPNO5YiUOPzs
LIojhiaKlHpoPEH0OR5oVISEoT1Upb76SL8aqAYvtSNPN+bARwszQJPXQFwlSgr3
JoUYBo/wdhu1HGLykK2NB4USB65lmDA+bVeyJtGU6ZLbBLDGpx9bARajkyMdIEbn
TxU0bfZDX3KdpTnA9Vo9qoGNI3kvkmSikuB6r3EwwnMY4L20VB9MeyKavPPRu7Tp
MaykN17hnCyv8qcusfrz9i42nkvnghnQDkGUfh5IkEahm7AbbWffp1rkCVUMI6RF
IQ4MTP0UEiEofo7LaZEerD+n+sTBAofE0DfOXFwgQ+o0Lx7aO6+5q5DJE1JVuWvE
+FHVceAcn/87bQaUvaEbj5tktkChZnAS2bHE7s/kvoLPV5YrUvCxbsTAtffn1xqU
c4Gv4ih9GlIOgLqfCgK6abNsjFmwFRJHkurmoBp5yDr4XIDCePWI2x39LNEwxrEl
DqkLfch+uKi5BysWYEyEv+a12V8ZY6jTrtvZwfLgrc2FScXUAeTGxpk4gTwAWh9h
+XeM02Bk5hijBuEMaCHsKCVWeMcTxXyIrvOjwCaJ3glUS8OcRN64xFvVa8tq/zgq
sLnyIesH5b2hK3HLjn4GTDfkVLnMKTribVepV7mEBgGcbOn56C8mV8tTH9hWLvVR
lgJbcVIMwiVn/eRZ8pXgRlUMF/8nRmVEG8/wXu+4WslVLn5NYKM3pDNRng3zBwW9
lvb2Bd8dx/pMTU0ZvOCo255NUT2C7UDLafF4mIPnHft04fwOaB/D+Dfze2eW3a3D
Nb6V7QPyaKZJ0x5XpBUWASQ2YdYgXUj9LPfAOXpPlN5aZCbNXby6VUCe7K0nGMoS
gzuc/GGsfQvMacvoL45g1tYyfnvJEUde0g2YtukZBz8oLPMCQWt3njvJx7SJsvZA
KelDxduNTwLdfUschC4Iiv6St1U/CUIYc0YIFX9wPwS5M2zctAtl8QI5Mq/Ss/3Z
BMc75A+vM7KAR5qeT/ZUSvU2uCIbZ6yesQWa1qjCauFoNYHQr8etAOCdNZma7Vv2
S0N71KOgZmJ3L00hHYqhse4vEmEy6d1ly4erJMj6XV/Jvu2Cn4/w/1xUpD08qtLE
7oVzmHcid/MUFi9w+/Xa2ycLqJWWT4LSzuRPsJa6bBIOhardijXQCvkyBGlInFnG
NLu2b8U7uJ+pJsPYDOP9RbOQ9EK1hR9AZ/WBjNyMNlAvHb+WN2SmF1pR3YiUYfHM
2L9d1IfxeUL8JIj6iZEzIJCSGNO0e3Eg+gC25ul3cSR+GO2RLF8mdizRmD++rJ/Y
hMR1bOtLXLJVqx7jA+sZ6iPQeKpPh6PklFo0X3PwcjISQYigmFvfA9iOpuEWB6e5
7jPJa3j1hgnVVzHjmq8j3h68bQMAYqlRcjPogoM3CKfwbHJAdtxAeSFvd3ZuRhz8
3IRqwZkDG1Dyce5+09CELRt9oFAXQpGwJ4XoBR3qX/4QOdVu20p8/a9KV/Fy1/mr
Oq57tujM5mQMNyAPk56ebe8adUkyaDHwRNl6RBm9RLbjxvHN4y57dXU1crKDK6ks
dE77xPw9qU00oesGx4nL/IhUmOGttK9Cp7WSl6PsC5wEv4j2vx7gNN8r/LxDtbMa
UIg04Xp9HtanDU+VSWniPYTIZz6B1JN+9DP8ozSwRBHSQgOIBxkievYUgvqmfxai
vOjOF/UvVj+LsUI9wUBZiLgug/MF+Kweq1jHTooWT2H5xvHHu94ZdcGoM80WxCXB
+ptVYdjHEfKwUM3+Ib+6UhKebbUm6Nh2N8nwB68LX5rnLRcYuosILbrISVphXljt
zuHBF3BoVPiWb8HyCuGGwUbrAPuX8slk4wIkug6BfxjwjiqxOgyDubNSl5SKcaOM
c6C2h2n+WUd7NddSjONYJY0NCzUk+t5bWQUiEcEfVekgAf7wM4sAT5VvcCmqVDBl
+kU1MEomcOx30SHHlpdn3e19+RuKgU9f6r6mcT6KiU69XkcWXIGF+Xwbp+QxJS1e
7sMKcJwsoUfioJaaWWYXGT8Rl8LaxTl1h1YmRLwmcGCmi/wZhsYmvpATzPvUCqGr
Vchi2Sy6wLKwevQVr6GlR6z/kvhzLpYRqOpJwKG/dSG6zTjL9ZjbPJXlNeKxhVI0
ucZZxA0s6kzxnW6+IdVr7nCZGJh3tuze0b10q5d95GnedPgGEMwHqw0ztZtFfXC2
+WFu9G9jqznep1wp/YYnoATD/aIQUhrfv2hweciZNZeNiUomaOrKnFbSN1YpJ6DO
+gLtbQQoXo4LRVCSUirLTIMqdK36mBP31u00E+yhjwZYgOzjHNGHNcKKSIHyXOJ3
ZzIiXanTDi7NECG0ONa8edGvmfpxHIRp6GXCSFo0GjS1YnYotQdIvaQgyHvZYWAt
+0fx+V7aXt5QFMHBIt8W7axUE4wnte07378+CWkdTZICkCaL7Zon2xBWWuNpQNhN
tCIQd1JutFL/qIl6I1+tmVCdnJdQjB5fzRJ8ZlXabIZFan1UtCDOPL8h8ePiSrvr
/+thydHlqIdHm36U437/sZvNoM+3951sSnGWca0lZOtEDBMD56S9Rgq0/xMQToW1
uxi0/kkweVNqlM9v/2GthgaoxXiXJPJ8L/2rv//tfhxRpKb4UYdLoVNIWMPlpl5s
HWV33wVRDzgXF9PsNxusD5P4bD6oORnKhQe3IRuJkKpVbzk1Kfe4CA+v5FCfPdL9
f8Y7pF/+CUInqYspHQXaXYVHGWZuHi34xXslRQj9tYs8X5x8TUu7BHgHMh2GZP3c
qcRTLaI79US+L95AzVxybxDN3Jbn8xzZ9JB9W9mHrC9WAW5S2DmRWxBNnpboipG7
eKQLqzRHXkF2CRfY8w57ScH6zPpoWMlkB0E+IJHs8i/D40FZhEvFcOHLs0bd8kzb
cfRFaZQ9XngNinQnj/fXgNqJf/TgncRbW0mNxe1Dy6XA39Vs04jnM2QrorjjVd7e
ovzJPus5fwFCj7NGcmYGkZiItuhWV9lLsOXOZCCIrUxsDTTzKWDRApvKDQ4vdndW
fY+aGowb8/Kpla47RRekCCcYT9f0t471UPUTQWGqYPLi1k6GKt5Tx9dcS+E7ZTGt
gTQVQeCdHEViDvAFN0Y9jbfc6jkoTzL8foaEqAe650R2loJjrd/iqvviUXe3WObS
Xb7oMDk/QgeSjdqoK9SVEyBYj9y2L3XaVKCbBLRuW/XAH30rPe5JqMYBW5+6LHYi
fbXMX+un7Rm8iezpye8bkX8Kw5DQsDsvxO1p5wZG/kW1WjhnTAuchTYN49NJd+9h
395nAV2ZUX7GPBI0a+bUejOtTE12n/m8srxGxl+umGc+fsztO3wi0CQy4ixFJIjH
BEmTBn7tzpXSR0n/GPWHX+rKiddvyC2XxxUjRuBuJt2RxBW/3sHpx3gItldf4wai
20cp5Z/CB+EWTx/AYRkBBC4f41WW+g32krAxI3UEO7xd2EpZnP6QIM2NE8+k7i7O
+fbKUuzY1ZwioRJPZ8oPgvZja+GdTYYao4Lx9ri3ptIHctuCjSwkjpBNU/xu4fr7
FMtNXtdxxQhh4LEUbvRj41DONv7u9noEVG92S727z53c+34HA6OFqiEQDJWLxb2p
wHyuEmAx1dO3QzDRtvP0z3IxLoYIJm1Q6Ba9Qjjxh1xvnMqMVSRVkzJZIqzY5YQc
t5x+gyaAGhMPcjr8daSbZj4Bgggb9JgkvxO1SC3UAdO84e/kVooZOf+a9ZoZYLaV
ai18UN30OmvEvGo5hTofklfu9HpwuV/h1aKw+ok7/HTzNcktK3hoV6vueIUIMoqD
ohTGt41ywVmUEGIJNZRgmMDH+icAFb1g2xny8gquPDmxULea8r5lR0wBthBstyJ7
rVNhOpVJNjvLNWFbMNbsBTvI7gs7Xnv6wtQxFc3lNrBnFyAugUX4jrwKw7Z3oBP8
hh3eBwtck8fnCe57hTPA8dk63ksu+onG7zP/bMUz3ieOya8wyhKvX5Uk1VRSvcnS
jb1Qbb9OYXTxvJ9mOYPt8AL6t7DP9JqOyXqvmhiN8XV+juIhJyGnlv3OE4aDG+fV
91dAtfpWGBzyEt+iZujzRJwXHcd3Je2inWUDshhh6JBnZkUj7nbUia1/Dt9JlF7B
On0q4edsubDmwm67GV06ZzM36cTZ/IF9UpMek72Ld6WVlS2wiyAbxsoU5HCy4jLH
VMrinN27XU/fm3DNHmeLjg+lH95OOXgOGTixM4vH5ciSpb3mkFMe1p8wX679gaaR
ON0kcYk3/EM5QP3qx9dCjWz4dSRtlCz1CzmaG7sPNU3uXeDs14KTQ/uCLpo8dSRG
mtHyLQxgQ5eWrjaO0EGvmlhwrJ4EJPJKVx8XRvzQGucmGHMXJB4u3t0I30ZvzGq+
ROxVNOUNPB9BKEAk/VoZ/tuJWphuS2gWobQH8XxJqX0tgjjimMS97xT/SakZhTwx
/8hmk+yppPvdrJEF8nWpP7XjT3zMicZRH8GwRcgC1A0ijMC6vhiB+o3bbcEk6dSM
UgFXU1xhtIxNruiWybhlNv3hcHkPjApRPV71n815nqtnfJeWv8CHqOGFiKsuKHxc
fne2KR7MRZcUS40U3VnvHecCrTJofhfhKrtTASwB4H7xefl+GszsmyX3Tl6jnNn/
hhADIrMY+6QIR+W9WsfkT9ItQV0AJCtOHOHHoYIh8NLO9KsDMIIKvk7lm6ypk1xr
2t59+DQASMMe3JIqTLWoFBgueKuZYBmA8LzPg2KuLzQz6OwbhidsFTGL/ehq9t/3
xLOCQMWmUUsSdI1P46gFUVqb0lkYVio0bgF6RHVEY++5MgoiVrvSh+CZhU5+HBM4
d54asRyYA30G9nWPysD1bofl2QgDZkXPCznaXhqMHhxya6pYyCNgPlJwaRoxozRr
I+CaMqjj676+GHKf38OVlLtDE5/oJ2Wis79uC85WPSqUV05NF94Gc/3Pf/CNspKc
9NIIlVrv2FEt+fBolZg9nIcRaEVIWSmiCptH9Xr0b2z2/M7Htnhn6xPQvzj4qSZN
0kOq9M+IHw0ZBD4XJ2hny2vhc1tX6CwA3T28kjv9ulApEQje6tISTATPFctUJuSa
IkarDi9OMgL7FDW7cjWXHc09DF5xQDCcOoiBcObjqT06iqOeB1DBq0ZYUKzKwd8N
V3yVjzvkchIZtKPixf2+wqoXwZ+lMrD2Eiwb36YRvnxzImY64158fmbwVSG/v7z1
bztsBLVBpC/gADIlHS17ZanPM6E4lQ0nlZkhQMQ9Q8v6RHliZrEW3qE2Ocvw9cBe
oU+c5eSS2IaYpVvzA/Y46v5uuffIvYLssf30/D66MM1+A8rgTeg8mC7WQ/VhjIe9
dQqudrixhb2CBkjlLpcRCpZfGMANNtOZSwq6oPTqKERCXJkMsCPs3h7tWTUzgdiF
tGaNw9dWrXIjUdqowqV/wjxa9bJR+74ga80W473okXrDvYMW3vlKyWjMw+bVw5cd
GpLNenpDNYh8Tnx3Cw3kaP5twT9z5fz5Iy0c67DhtSE6iRkQr0da/4AVoQlpEi9v
z8DUskS4ziNZLaK8PuBhAuq8ZVPTQ79G0AOoOippX8FMx4suL82/ViXreIj0gfOd
H0tGIdSuQukNGTADfCVrzbXwc/A2UhnksKknxqCjdadp/Hk25yLOHID0qbU3i26Z
Qwqa8lBVMIROYq6aoEGx6DWzEGwPmDIT4fM5tN7xcpR0Dft2XSg4QBQMRYLyY9PZ
bM6DyZL2C+KI2nXsdLDL5hSEVjmNqI6MYJbQyeU5ZChDXk3eBf9hjuT9373CySgv
zy9vhmkp7i2ASWczPOYNpp4RqmBxAs/27/x2tKLUTF5fEERZvNaqC/SYmvZKsNQB
iV7/0hcm37brQeFphUsSh5hcdIE9GD6XYMUDtXATGixq72zNRUoAGfoq2fLLtzTD
A7kbS0EfNs9b/TPCimdKY6FCgqbUDwqL188pnibS1F3GmKMJkM7d47P7D7IqJKdl
OyyboWvlZ1bJZs3/W9GT/lJmzQb7PgJzDtukhp4nx0HqFwZ8m3lnIT9NAe6p7aG8
HsIXWmAgpg/8J3w8yUX1t5TYtyIVrg/HKuY4MVjXXvzPdXxxduvlywdP5hM6ZeGi
PtheAzub/mI6Br1bQ55kqRMnvb3PGG84sxH9QC85wi/TDuSwefAUDS18EMC+irgW
K4kGJ4zpbegtEx9wgZp3IxyUWq5KYZvkGES5SfdfWNHuJE9D2/YDu6rPxTjWu/TG
yXFr9BLBumMm1i17vKPJNlC4upfAP++ySoZs+4tHrC7KZrnrzJQDOz7GeYku7kak
1DT3BYqLA1qHrJ2PteaUSvFqtxEJ99DzTjFHXuEZTdbysLzYJsiVlCU0ES4/+idS
HdTqUY8sNgf2Oof8AdxODfzFu3K4ZM+ekT3hRHijSMImat+W56PG+xIZ7KgAWpSh
JMAz7xUU9XIqaqK+R+edac5KscyZEHsqzt9eYORFIv/+tFt3HjPf++zwVXKR8iQT
pnZLu+Qq89ke1UZSqYhqssRWtJe1PswwEM8+ONJhgWac0elqbrXs+/oJUrsGPZh7
baVbcMNBVCeXemufC6e4ExNnDUImV8D01WKOwE7o5JNPoNmF6dDAZmyQwKGB7aVU
inW9jPcAqpmRKwEliMy+UPtOSsjMSTUoBslV8Dbww2UqAk5M+w9sxzYS+JwaUyjC
aKp/P8S/00h8qBZSD3q48dhzaLW5dIXssJoO7GZ5L1y0shbHcTne0GijRSQIhAsD
9pskWcsUCFCT11E+yjn9jT6qb2jYghMaPhlwGTFvkR/yW651chHrHjmwv+kAla+I
27wnokvMs3FH9PIgYbRbt2OQeAY+trz417bI104TZbm4oqDClX+hbhCbGqLeEtAC
Q/7E2cPFUSlZeew6rBAWi56FEIwczLWKTu56qS+bj+pvwZwZ7RaUDOzhjL2AEAKr
TPY37RJCFMLOLc19M+JfM/0yZp8RE3vOgIxHwZtPdstzl/ZTtb6aSIuk6pXWxIco
WFJfypyVFj2nwlk0lmOPLpX5hbSORaz1IlWBKLQkbkmIxHDwjjbI80OETRFCZbQU
eIshBV/dbIZhf5+kTQHo6ZVewuoq3PT7rtQPRE94h+EHdR9HoKzKlAqkPMnLU/NT
XGIAFqUm3XNJuCukGYSDD7wxeT0j6Lxj2X5gqdwvvnBssCZIU0KvBwBmhtKmNdn7
4BmEZVnHfPmFA15uW6TCzQ6SpK6xFPbstSQWOqGUq9mytX5OQsebRy2KCgBppzK0
EznAMq2DdJfKStQH60IhPwmu0CN0J14YOqIprqLGaFNzTmvHPLLA9u8hnNycjmE1
R98xIUnAE217+n4yzZyVoRt+damx7MBeLasHwhEc6ot/PLq421/7FJI5EFeWpKs8
hf3n6ZLxGO9B6ChXfDCH4SyuFtPTu3NGo3O0NWenSS1r3q0kBDZONf7WXr145Str
KuxneBDCAdBpsxsu5QFA3mO3fHsBS/Pv3Q/Qejamz6qbGbh+xMko7gXl2BOGHiud
OQ8ZuUGigvUQEbqVODrdYPedv00UqaEizapLWvTKiOuEnLERdIqjT1yFth1mrb7V
cBuGUmkSI98hAL5i/LmCLhnOWY0LMFJBDWbiQStmr/LE6V7GxnmjP9hNHX7Jb6gl
QtX/EKxgV/wBGD1lxmqYZ6QYjnk5CrjRYOCdQVZvKGXg5aLP1wyMDQi6mRpil0OB
zEc7MC3qlrZazu3JnKAlyzhgADsk5OQDtKSUZCKD2a7sYIPt5uRfSluSeKu0igT9
zqnJClOFyHla7ynGCMF3M9LQKLZSceRgSsCqErpo7eCUdcs6++errcRaVfpZPmd9
OVL03o8g+o6vs1DIEfDYEQ0dL83Klp8+1Qx+7BEsvmXRO69ve9KLjMJv5f5qrLDu
s/3MTAOUSnIan6JhsRPf+Ry1aysFdNBmVDhmeZY20ycFEK/mgMSYpmAWXYNVfTu3
XwHqV1TlsG8aI/VddNTKS4WBHq8M9aQf0ziY93v8EZc98nvDm0QChz/pCgWwcCQn
6/zpz8iMNxUXZMHs/lOWAlYtlXrtFw+VpAJoE03wXzym77OIeQmv0rK1QwchnKjQ
/24t5SFktkgDJRcaYppV3mNv3R7+wNtYzkKGHzPF4ZjWZEMswYnaTxelXPn9Ipf/
ylng/CAltR8ZRqUTS8nys6dqUM5hOo2MK1TQddBthC5GAq+A6K+FUZ2VZ80mb52i
fCgGs1MtvoUbfvUawSbhyaZ4Ao8ogq+qA8e+HQt+WbuEA5koQCnO9N8g/gL+m/Bl
yI39rMeaxq0B8wPjpREkrbdWH/qCZeAitFUmn2zknqM70COilZ1bDKQmRgbYzkkE
sx15uilukce77CJxv1PdOfdPuFybk7geHJ0BqAq5ffTVSKyVod76hS4PJe2hssJL
PWJVJs25vMttBsfDzG834psJ33docKc4fXYXHofOkbOHDfXaoc2oGfwCrOIfj+MS
fW4tBhxuNZlcLYtGBgmg4DxMqr3B5dLEMqJUESkXnK9Mg7AZ1n/gzZNfZb4Bs+Hz
on0I+rfZu/bbHHxWQ5wenZ8TUSPnenSxTh7+kOqLZz2ZmddLmUevdSdH9FNl3GLo
M5bybNGj53R7YHBgGgpQrdXiJh5Hm7g+FrytVqrVqWOTPoqcQXES70NW+ilZV3vb
ybMzB/tc07LPvW6r4HG3kfdxDxfL2p24ZtgXoMLMSjW9LnpaA7kJERONUpysWGXw
83pp+7NYNi7WG9r0sPIi+SGXXjKZJP2btnqhcQZBmjsD5wRV6UK8L/4S61yAn+bg
78f+oEH+Hs6Z0qvgQ19j6CUeaUQsy1Bz1/k5eG+C5Piyx/P8EhxhMzg24/eLBz6w
a9l8d2UUNQQHurAYyOFgAJZjMkMg0qJdovljAn/2OqG/IpP9WuBeQNybTFtf9UHL
O6EYQxqyg2/BYJUbU5hKzISpho07zwBenY/VMWUOuK7r4iewf1WZngo5I0/LNrFk
QyZSW5aSiOvQD4IIib/IhHhKt0CdwoU7CfwIdDbR/UJuB9/fIJaK8gPMaXcvjOvb
gZ4ia+fZmVLYObvnKDrTnJ7FSIVzMV5shBFhJ5uTQ9nGsLOQDVRQg/Q1EuV9FJiG
BZItLogBxMQ+fBdyy+Ro8P1yce2WAQrhE8/O7nJ55R9N823Rc9myZfYDR7w/C0mO
LMnY7uWCzNeQu0jMmx+WoH1sLB5xvnrcjeoNMniU/G8eJhxrfDHEMJGnzelUtk+C
jUh+9IeUVc6OMmL8dF6U4xASDV2S0wmphby0FyDh6lTbEbqZCTynZ9JzlsiTwgLO
8jK99frZzYRtCQ7EbOYNzqS+nn1x/SDIrmKZLMRSq0sfbhXFyRcF2FJ8hm+7NjI+
6INbDclH8ic3KhJ58uw5RPqCkqSZetAMXX/Q2YQpKXKbCSfXRoNKL83T6PIWSFBm
zx61fLeVA7FqRk9lKW/0mEqGyiQhV1srV9vk1Y9qXlZU3jVRjC5cX6kY9Bcl9EL7
OU1VKhjetWJ/JWXNLa+PH6rGuUGHGpKFrG9w7hEIeJjirABXWTOLFClCSy5P9642
txD380ZGrGhaYVno7kN/huOhCQGHguhoYMXFVd/pkkBLtfTswEuMC3twpIUP3J8R
1aprVdO1Ky45dkrpCZJn/y6HCwN99+DgZB/NXU5fdtfwy+Jrke+t0ySf4YLBhrUk
6xLMD/uXQjojizJpawwLnPbuxQ+Ex6IieJ10Nid5bMkLsGMg51Zmcs+hrRV1Rnyn
bHJN72ye9gCxBodvjZ1RsDPvvqwakSWFu0kEtEljJLROsJsmNCxxK7EwkLF+Wf+x
6ezgrCZVgkTTDCYbydCdTfmZCGqDDbUXDCDJK/L14fdLJ7AFEFXocVkyedl0NJTd
/o2uk/7imdOazYc2o44LP9cfYMYZauxNPNFUrXMcHFn3uvwu6pKYtAsVgDDot4D0
SXgkBplvGIJ3FKwMK/ihTRXMNz9H0pa3VpppG8uQ77fBeEMud6jTXE3UmGwtsf/b
vL/d4msT5Zpx8ZrS2SeJrQcFE5HFwGRxyJ/iN2Ql/oXMDmbvGMUa/SF2KSGkdqld
S/gxgVdUm8KgZvuaiyUDkkQ/u2iNQhcpXjWWussKzjRO+DxAVQNiC3EDK5JHPh6K
bXhsCbRIqQQVl/MysgxrXQ9VZJcQlh7vTIZvsqSuQR9RNEPeAKyoKrv1LP3pw358
JY+bgCwmSEtXxNVRbk/KtZByJdIv/eo9b76e5ibpkXkPf19E4dKZ69L9oPbbojiX
eSNCTQ1pp+bNtiPZWD928S3se0/x95FtCupyNFIWDcinbpkMKnKT3/NwG4ybM7oZ
sHEUmwTXU3id8esLwbb4qHAvq9l1GxYI6QwdeW0E5GuTsacisnISYg7Sd2AoGi4J
BgnfJo+MfRuPDLkU439KOhNcKn9Galo4IbMZKWhqAIyVIWU8574SMUGJjvL5i69F
THlKz+WqbYq4cGzkuNVmNHpHfVl2z5jugKZmx3Ny4k6NXEp6o14MTKjkVHG/kh4k
w8D5/VFGoAOtY9JCmCWQ9bbsj/x1aVMkHNSVCAgq35ynmZXDmlacgC4meEiPM43U
5SIj3lnnXVcPNyM6nXN8HnQJFpdKpGS0aVEdAhpEWvkJPiu041yQp6FLs7MI0aES
2sc4hQLa3kypHRgqp/ZBH6wvdf2XDejpAxsbWdkiuDMx4yuYqAjDyPLqHiBqAgRE
tv0iz+BtVJa7eKuDAXbvyE00opdMisDJq7/BkXgIr48CYERQSMSytNw14wnEioUp
vgek8QOVStI8ABkjhi2Sucec11FxfbJQgULBhRpEaX9OGFlcNxR2TtdPOrzQ61cH
vc2JfuMpYjxBcO/GIDJXqWUsEB4ZXIAESSHKIEg7lrAqRPFDGyH5QtKFN3D9yNnT
c9IuNp1/WmOHRTk4AIn7o/65sWTEAmgCwrtZnB5+xMTyrK0ATgS2bYdxTJGkrWFi
/V4o5nFSpWDQjCVz771ZJauXOSc96j5SQxNEmN2UvIbf3fwbAtyb4o8RAFMCua8z
74/aKrAgkBj9f+a7/jXqr4Hj/aR5gC/pFENh+bPHhaRR0xYpZ8Ag1prhEfkIqoYc
MOBL7wTImhgkmjJF8way5nLr+ddqqyq+TbP6EdATpixvoNhJPDpHXe0hDzMx66Qu
VGVWDgCCj/TsiaaIcPO9nQHv5cx8Z2i5gSoV+FlXpAWMjHTfHZtcYJNNYdv9nXLG
iZ1lJDlARGZW+AJN/nktwcO8csi5X1io91oMBbC4i0owNw7K5BFXwuHJN1KAWebC
+KMXNB8pOJNyRDrZXplXx7trCfQRzoF/q3lGHtBxYGUzNpVFc6FLTm4yEh6iZI7y
n6boED/KjCvXTeQlUosoT1SLcyxJkfsEMB+d1oNTTKdA5cXPi4dPSDcuJs2FEDsJ
n6NWjSXyP0y+l4WEq7ch76DNHEGZOUku/l7oXIajRZGToOe1lkGfTZwzbf8ONKVL
x1R5RVjla2Lt4Nzdy++9MPtl3Bjopb7ijMt3fsFe3l+v/JlBenR+BYiw4vfVs1AO
zYjpeBGS5jVkx1Rw/esyXE0mJmuNLtKvroG8IsTrFgdSIWL3Hl3rxGoYhRsyVQ7n
Mbpr8FMZAJUNh7nSdvQKdqf0BCPETqY9zrN85jkIhNITd+xpbFf1ZirWGsojbdSv
49tr41aZFJfz7RdW2jI9UWAA33GEukMz8gviPSfMKcFu/QGLbfGJf3ns2cSaOgSo
7pNb6ClO8Tx2r8k23d+XoZ5S57pRJa9+0xpaIx+8NveU3X6aVu32MulXiUrQ/v+D
/nvhBI61gaFvA0Aadcn1biiq43wYE6Rzc5WDtxxfxT8GDOzv3+AO8jpr72/YO5mJ
B2Y/r3XvoQm31kx+/NgmV5sGOor/lxdjKXQa1hnKrH3w6P+pQlaThtzqL/HJKt/R
vEkB1WivJscW89a9cYqz5LpqSzI6Zsjb8LT4WTB6gTaeaQO9LFhE8BqS+vsjMnDz
n1sjhlnP0Sk6uxkEK0BQvBtXSdhWrkChjl/Gwog8bQc0umCkoeBxj9zg8IXETsKP
XobAi61rT1Y9ojD740ylrS7ZHr036atNAxsXNvthrX+Qr6wt6D76iL1jL0kB6SCA
HHwHrMsjSSSpIvlB3/Zbkgfkp9e/z6oJ1qj9SfCo1DEwOR+Tx+MGG9MKQiS3K+m1
7Fi51Xb1K+LuGczBlC5NtW5vsKWc+N3Unehf0GVBeCszV87wbYZyOUniPlM5IlOw
YEjei1MGIuhWbATH02dOVux2QzxhIJuISOA3afjsnm02KwGlINd85Ht0pj8AJeZs
KeRRKb2BJbnVOZMkLdltYEbuZMPY/1/YHOmqtF/rbEw8bcKmvwVIFeUOmEbq9THf
NmYZsUllePg1u+HHc+X3W/PC6AleLI4hlh6CBlFL6GTm2QTUN2Dqf7E5IGREkOP1
6wRsVpZ3ANOn6Wu54ev+69IjlVAQoz2OfbXJSj4mEXFjwXowGDYTAZOczqv9sm4u
NGoLl6Li3fw0MGlCrY0kxsT9kUDQF/nfR6hWgWg4cZkAkFGWHvcVNuxzqeP4mukk
bjwwsiI+ySBX8o/+ArWy4NZky2SvzRxVQq9BH+t+i8v9LvpWMWPqNxAZFolBq06d
RlUZkP8G0rBmSGe5k2oxW1mbOR+twQLrJTYbolyu9g4mOtK/rNcC4V8YpAA2KS6V
SFfqOsGJKte+aWeppwQPLoA+Fb3NpPpSVJJY50zrZQd6jm1W/TY9zD9e/gOX5q9u
CvpLBIrqmkppdTRkmBoLMmZp8O6E2qAcDb0Bex9BVxt+NATg/YTHhoqgyuqapo0J
1HoiYz95oqBUsKGEZkbtox6/gJRWWh0/Pj0Qanec3DiDVixA0km+x9FQMiVwOD+n
+5dRPLVIkcp8yYwhDoINs2Pkl/OX6zO574yVRIb2qSERcyQnoFY84MDtMAAINJBx
MVpboYDYz2fyGIuAeXp+a733mUyf8wiiKYYW69eDsEndmKNlIZ92k5cK9ZjOY/t5
0nCPdamTOZxQ/dmIaMYPn79sgwiMpWyABl3DbTyrfW+2wSvT1/uQJ30VNamfQ+wM
HwgcGNuBfY6/GM/X9nTg/TrSAgoULR+hSnb8q2UpJY6TtJGkn5IiYVEZTeaGMXoo
/dnKcTPDeeGqRQIUmUCCwAEhe7DuoISzi86sboCwYDtHEy8euG0NOCdySoOO0HoS
TDCSShH8/55VWW2wwEEiLWRnAKNvcLMICjsb91w4qDAdUXVmy8yMuJgDr8ptGRLu
ym/RQR9HBn8DHYItUKaU2UnfeOSmXixjIzj5FhTQseDbk4tCx6N3kJDaKRbOaOXt
vlrYUMAQ2z+jgCQpnBf41Z2dbHuvfpuFuFErhlbo63cXuZL/7uDhTT3TtsevJXTt
+Y0TPgReKxBwCFlf/3Nn6Wb05um435uMgJOME9+96Vr8+/Rr7slOoL2dYYnBbovS
2H+4WxYJylv5KmN1pIgOXAIrWuPTzg9i1vX9igoIzchuLl/Dw4jWJdmt2lvHbSre
OzW8Mfe+kXPAfH7mHxNntRfqbAwB/xSropdy/GBEt6DM4cpg3dcyOwrnedBqTWCM
HCSC5A0NuTGKxeSCjzoaLbSQY6JijAQ2qwOhCvOAhA9ArqT90KM/xgAIK/0z7Mme
PfGn/MubTRYM/rD3dzhfMMq7p8vlt7UfH2YMqvShK+GBtHF4CNl9eCBP8pfLiZ6r
eHHotdw1iStzNgyNklR4pgj7czeKlweHth6yzJuN170kGVtKA0UsWdrB2OMzYjgr
EvefE6mVJVO8PPYBaHKPgs8rCIj60O8RTcqdnXxS08TAXb8pxkhYS5v50Rc/Zk6d
lL53KUHmQlnTGr6cntdW7Hz9NqQCakqBjU9mAlzHeY8FmtPJE5E45v2nJJNEkC1Q
zBdK2rLAsVJfVr+5q3cmWBOVafFNd2mT8BgWavcmA0uxKM4gTA5/8fqnlzfMmiPK
SI+Qxiw4zZyeH664bzoKfKF6tDHU3WEeodPCIwP04yduZsIj6Dn6nduoySMB50qA
9l4X8f/FHF44bY0bT+LbtZxRcPY1mpkjdmFXK2YD6y2suMK6zXSbRuxc2gFGqFUi
ezyJYnNGqs3DV8V33rEInSCDPP8n86uJtSFX5hJlsz3bHK/AmiecHPyfrFefZPwe
QlEmoiePNCs8u1KYCwX+iSwx4yHDM975cSXAiX9SB2fFYmZ2FKdzZVTEGtyboIi3
onzcMzhJeXfHbSybE2pKMEmCf88EVq6obaqhRlEslhE34O2L1+C09R5zUvFqZvM4
YSQt7PJzM8jL2YYnxlkhoC3FKcDuA0v5zp++CbRATbwL1Pc03YSfl19u7685YL2H
+w2aJQWt4kN68n1wexhjWyIqhUxaZa19lcWTKOF92f53VeWuEtEvB2LSknD5VKW5
nGDw7NH1zw0XP+L8f9qJJ4lbz1yi0MioqLqUm/3onN7OcE97rAGznnetlNeBDG+k
PHZ6APQBpZ5bb+ojxZN3Uy2YkqO3GhZlMtavs0od7Wxr1bgvhd3LXZg3T7qYTyJg
nqRtjAtu54P80c6vgC0ErR8EAs8LhLjOpYXOjhJ0YVGpyL/JAq1/f9fZ3osCCWzi
HMwtLmA22WT6WiEpHjyYOQE/orRebGi1DomNE7ZQHMuDhfFY0SgfhEU8V7PBsnmJ
l1wMgvMww6vpgUokAgvUsUnoS8T6qIHzd3KUXcVZWES38Dp8XNJhn/ZxGtD8+KaW
OvGaeLido1XMeD/VQuzi1Prd6hpUvxIxBILpy3m/Q5FtEUKnMJ16PCiMiM3PKnh6
TqvNgcvWOWpOsM3oxrrJQ/0kLY6Iq3tLvaEnne5SnqFooPIcgWK/L9nfPCnb56oT
Ck5oQpKVtse2alrdpq5xycNlRGjrAN4QPWzZGFuUCnTNigSLQqE6Z2PtfAcsADpa
fBI4QlCzwy06VTn0xGyvr2WmHkBBgmrs5l0q95gxytkm0z0gVt+X978DcDByF57I
+xi6VeG/h98NpnR02TkZQGt/dfICLm1ENrIeMcsK4bL2w/N4tm0o3z2N652E4u1o
q2snzM78q/gBjxaf01IiFVwdUQ5+AA0EwEBvFNL3Hh0i/N87ZhjNdod5joCe4cuz
0OrkMmwBn9JyYhWJWYaog0+vbvPr7I2M69e3tDNf7SZsv1auu+xRVl7To8ryaM/R
SIa+n3xiYUg62UA8fjzc5dc0CcgZQPoiWz70CRZ7XWxEXhoTCsa5n/bFyBFI0u+2
J2FwDKTXuJD6G20u6OAdMwcomZUFnAq6O/0iiMV+oACl+VRGoeiRnACk8GTcQAwk
CD0OEX2RX4TUGKpq8C7LdhNsPcLhpTPRqDeJ1nkw8HC0nuXY3hji+icBjkxzGNJ3
ulpIB7s+Pzx19cHlieR80eAhoXE7NDM6Y5hrDKvGtyeSOgN+cJDgcuRWyqXdfddG
LTbUmor1GVQw4QrqOihNYyPd5/JbkznvJBXwlEfrPTH4KExCILYtvT3QVJ4YM2ti
tpStls1BJgMmW39hlo9ItT1/GaTTbYOzxmEreW2Rnq8DC7MBIntmXejrSRXzD+Ln
zrPYkqjJKxYELm3YTQjLzBcJhNJjB7iYtym1xDKVJMaEWJrbjX5+eCpiBvf52xqk
cCFyBSIRZGxyS8GQuR3OvfGgjiMEDUi30fj7Tp40gFdCipjlcP8lr6ij2kec6c+N
rNb7A2XwPX+vj8LN22p6bb2ue7Jwu9qW8YZ8iHZymHqDXjEF2wfukkViUwRCdJ5J
QcURX7VV6wB+nsCOpJ7nPSEQ2LcTuhKe0/+ObAcHymP1La6K3au2jdifWeYaXYi2
6G1RNDPdKj4Mnq3i1GzWZcvf0k0EpSks/FGz8hKi4+q1i+k0RfeDjXDq1OsJo6xO
1TYFXcJ88aDXg7V1bAzOUR1ffrvXZ3d7+7s8f/ikjypthZVo9q4C8qfBcumy9Wy2
UvL6QeMN/koNmbRu7cTeAOr28uTKMk6GYxovnnCegqr++lRM5SrDNDSCrgJwTKDn
l+IR3JNDcpaJLuGULZ3S507cSthN6kqyp/JbOm8l35UVWuwBt6QeIxuW1iRevIH4
MyiezJ20m90DfFd5AuI28Yp1jKg8a/qtVpdymkXSrbEg8wfOGNifPrwWMbZMhanE
k3hxtRR3rWEZWcv6ug1dYpgxa+OW2lu/42OvtDsPcHA3be6bz2WzdhF8limxMz8m
+yVFxk+C1kFKILYxPjgz11kA0TaGXbM6vwt3KTr/bDfjpBitShypiktY99TEXneS
/1DQTZNav5XSgM0ShyGeFxK1kjmzCyKxyO64QctxJlMECBKrWw14Cv3f7mvIpN4u
VGPR5C0IvjGgB/69Vdcztkr7ez2qdrK+f/EfhiX0P0tNuHUO53DrJsMRPTJQjXee
MKRj+L2esYxzmrGxHNp2pejGKhRnHMD4e7WgcDup04RT1jORkfaKj2qSz+EzxvoC
LNw0p6RylR3C8jMPH752DeHO2ZDIaccoKNb8af+JJoUQ1EDWIZngp4XQJZzmNz18
QNrRPt6/45Q08FPcSHW6tks4H5TTmPAZENv5hpu2WYMQpp2l79BuOJBiM9epno87
xoh9mxqhxsM3WYCm6Bv+ldP4vMyzujI0T7yTvqnt+YMW5XpKE0J2hwyjYjMkCrF9
uAUXvX97wHgKV5szCfhwls9U2OsB8E8ib8zLZmSEaU3PMujjpthYsMBkdf3FMpu3
UL+tnMr9yTMI0RM5jTMJYk/f8JYR9LoQM0G66uHDY3bm2uE2bKCwA8eT8Hg6S50B
RYBSI3HcpFld9e501w6fxOljQASsAoCQMnS45y/Cnwa77SVYjkRlegQ3LRiDgWK1
e8FjXyz/H/t6tFb/xCoSsL2pQV/aeSxMnuyO0QvkJUliCD8RctlavJhb/YTEPI7K
zX7JaRo49eweBNf7k8fNpnaLOCfkFspfVSRBmAqsQGw5WWjyUF/PwuId+F81B+9o
cwbfR5IbJ1wE4N5ecr7FlmRD8kLTEl5r8QA9fS8fsxRXF5dJ+bsdexAh2Pr0sN8P
IR6WpqB3/+6Qgbdl5p8WlI3SHl2Kh4sYe2BpUXrxhUULV4Dit1OkuIhwq8geMBUS
ziSNkGuDLq6puO93+wrwtnge5zV+XhZEiFoa/awvuZCDQ4dZf+XY4TBqlA+dYI9S
t8MVsGOElWrb9KWmiDJYIOHeoRc1hJ1X5qzNZNp1y3+perkla1stFmyaap91dr1q
3wiI04bXC0DX+aXXCMP0RLRWyJuJ6tEYY+dS5XTKnDcO87g9wUBjVsc3FQGYGbos
xiu/+IR9SlOun/H5UdlernZWfddzqEoFkkroPP4PdifwYtf9VRToakgmgcZh44mO
j96A+7O+tM6kLh+A2oB5oQywC0bzZyLxOC0TAVKUIZF1ezpatQ7IeEUru2Bleqg7
2A/7u5SWyJRmTgwGWUQRmd4JGoydstT7XwI8gaMBu5NitKBObFuc2/GKEbwDhDxh
jp6I89ueCelIZFfTJ8oTbi4sfpAWtXMaykwMJuf5me/NCS05PfrJ+t1OZILOIBrN
Rc9MnAh36pPkWfiu1/oY9ReityfNUHhbbH9YhJ71N/1xlRtwkOlBsniP7RNP0h52
qb8BZBdylAQnf2LdcPZuBG/OwcmotBVYZsP2wva32Lin976ho60+WX7mDXP0GOFy
MGSEsZI78KdUMy8E/nZVow+OGNIYPdmQQLr3y1eIOVx9M0l7eyMUd/EJtrN92mqv
MdU/QTs7H4OyS9GM74I8eu4hY3ViSa0DHerw2yzzpDzOPBznmUJkkaaXk9ozUTbW
yglRjIIjLQw57MtGWselPJR4WIr1ZCz2DEKwqUwPhkD1uI5Jymf2mD1RhaU9Zeea
ur2d2JDTFMyEdf34h/6vonkErtVzlOEVx6NWs7/0TP5smAQqagiwa3dn+EjnYz0B
j9jFJ5UgVggwj+eobe29BjttsAHLRwtMixn46adnr7wj7U1Z1Q8rvE9S+O9mhazl
8KZiWgnswjNXI6zPbXMyK+wchhzUE5w1LROkjLo4u4/TQ4dumTeblCa2ppJZ/Ngn
wv/F/UWoW41jOH3L2GZSIlkP4j/fmY5c7vhkz0LzWh5Dj6AVeoPosomTLaWZfAsV
NenF0kEaZEKQoLR3hi/7KYegUeOFDcOz+bw8QbBP9JNPWUZ0jqvYVvjuEUajdcNT
jqpeTQmGr/8t7Rx9NCtbM605CvxdudMUYU2PUOx4JZjIfhZozjUDkBNKwejqTY6f
TWJV+zgXc+GhKnQk5XmcIIg9y9zNV/0zF+KzfjQySfTcddMbK7kiDctjvO5zWNo4
L1I5yZW0oL7hIswoVU1A67SNZ8LqA+GSl9Vg/tXpaK3iLp/MVNT+iFXzBi3+0xWh
wOaI3PUzhSVX3CoBnvCFBHDK6P+UvGL45LB6l536DkxHnncJh1wrjua+Kid/VGVy
rOJBQyi4T8v4sBLWxnc/ekuwbMHSVtAQgtAURkyukW/g1TsMjWtrDalvVCyWZiCF
L01efyVWZFvzbk/lAzlhLxA6XKq9IRVbFCgIl4hBLHbIDfzDWrk6wIplWWAUx2BH
DbnsRmE1T9PexjQpIvI0M4VBsEZG2LShsrw3LxyFEvWEsEZ0wyGIuLsE59J3zzTl
Cm8t6TX5nVZn5eKo7FA2sUF2K9zeB4+vpSKnKeuW4DJy3BKJqvgKPcXFn27nxC+0
ZKDww8dApBrnMIdNRqprFpi+OY2N+Kg7BR6MGm9+gX5vmlIDS5SpRvk0JRc1UOaX
uAvJoFk5jo0e0UnkbR26PCe9Rn7e1MuNxa3O3CVvwV11ESLSZwOSUr7M2uDOKNI3
ulHi4BXL/QO9k5pYT7apss1ZcQV9HerxpBgzwB1a3aByixUzk5C0h1AsGUF2BU3v
OXIH38ibrKSgJOh0QeXIlmmITMd59zrBTEQlcZciyX4/8tGRK3cnQEq8NT3zETrL
I7hyfWhYZ+vqKMUaXNgEHumwYWX6KGenxAl8SCjYfAZOF0Ssold7tf7A0aZUE0fV
l+gr4m2R2FEGWl5qtOwqlkC1SBcsE49tlS1n6rdHbXX3zWrpb5qOR22yJdieSqZH
EZatp4lf4nOlpFJoHX6qteADhtaJUHSUWY9PxudVE6vUS1NlVUM8ntptEslGi/nO
JygbVJPOcAwOKKiGDshsJfUjN/dFYWw8MY8485a+DUAVNhblXF6TmpftKoDbAGkz
OdYBWOoBCLWLKt2ksQ7E9XmWpp4mU7UTn/+bBlqnHidEWUBNGlTRDnH7wIpl5Ouw
9RqFh+W8MkSSoa6uKPo3IO74TNLS96y6fx8DZo0w6WO7DAySxlVhAxKRK1miVa38
RDoQOq0rqxMrNQcoq+d95nSOPtHjUgK2u891zFBiRgxn+YaQx/iqZ1Iyn41FGlMW
CWf+6/3FdO3IVc/T8i/92K8Gv4AhfgLmPyRW2AcotmLVmXTyYqPgoXGCoiP+DCB4
4Zrga3fySKLGfFPyz5BGdjAztfxXr2XnbmFs7INFRTVtjlAfAd1AFZI8C542qFaY
nENaB7T4E6KJkOev61RdrdUJfHmizS2D4XRB338mDkbQYaTJX79/3qJen6REcxw7
tuVjUDtKdfB/jr1jOQbuSyOcUYMwEpCa2ujxANNW2Fc0lPP6bRUmpqso7iFWvAbF
WRC/Tkolod7c2LivHHkJ4QFrx/wtcuQvR1ikBTMP/KaUHA/7/6Oj4Weu0D1PAGru
xIkE3nuSnTmdU2fNRanlxXehX/YbV4UzNBED1Abi788vv9bAR52EVwDn5xx3RDs/
NKjlKoBUmuTJFh9dToqFeRBu4YY2ZxrLJJ2I9snP7N7eyyYIP/8aTb+4ODml7yhh
zg9+/zlyA0hZsG/k6WhXPbuVOP1MBB9tZeoH4vjG0qV1kJn5N+pfA6G/tqpbpJ1w
Vv3gP2yDzVOhIKT/mJr429mIDrEsYSzMt8AxP/II/O0IOokAvH+0FbwoluMdaftV
qwZDmx+beZSKSZZKjxUPnayiXNq7wPkrYnIainkTfscxHv6AMKnhH6CyVFmNwZzf
ObtdJ0eTrchTDiDuqiI1pzZZ2qyrw6612WqYUhK6F0JGJ/pBagZteDRYb23zU11F
jK3lvzfDdMf7HjCPSlY2Vf+tCSxk+AbAbqYht4SH3TssSHCU2AEBL/nspK90uDHb
IWYuTDfA4FL9AxIZ0E3YXbVMn9aQ/c0iDRMuqrxLvRt6RDDzFKwZwopR7/w/mceC
MHZQ5rGF2xK0DcojpnQ4fvFy3d6H/S++5MssR0gvLW8S7OQ4qBfnLgj8Ok067pn8
koIMoLgO6ZOvaOGKnDvZFhIKGxisExmbW9C/wpXStKaEjJVjFy3UqipzUHv+Iy01
YaK4XRlOeKZzcVgsACEp2RNiWXKMc7PtdzhA3tU7Z8+9QQOu0y3DI9Kp9sP2J/QN
izrME+KI2g7B48SMVO71NSOV94jhXHuXh0QXrZppgmJ4oFCMFf0bS2Qb1AotzdAV
7g+WO7Iuyq7/ODJgDJAyOsicJrAlreceJoAnfDvzkF8QbDuDawgg1BWXDjqOZ0wx
xwxmSGaY2m5L5E9puteEx2wbfgknsVt3euKBXzYRBssy7Z53rgTXWmFhsEB7vuFS
CU7iPqyBZ6rcGgCo1+g8aXnopja9cAdBO09ryoXboLW3ghXkZRtOYEYICM7nhKy+
CCFC4guLDxPmZEJ4B81xF+k0yZTWHO9NzAn/h1pttmx/DJEruiBMpsnp3hG+FvxC
kUT2kL0n+k3KHPp9DVB9wqjQqRgzGZ1vzt4nxQGXXpbdmx8nlWScXlv5qccyZWQJ
BY0HZQPGV47bNwJWBuJyP9fv8Ho42jC0evBK/UHuoniStkt8B3HQX01GEj9E5vP9
eBhu3kfc+QQzUCVOziIEtCI6ivxGDW4FqpHwc4X3ysIbqaAzEERTrNPQA/b200Sf
mgHu+ktp1KS2YMMwjEmAqiXABb/1s3odqkN2leJ/qtdZKwBgLOTMGdfhQ281cZrZ
Cf8JAzAm8OrGZE8Gy4YA5FsALng+nrDAhsWKuLAJZjOQyJVdUYmvf+Xm9quX6bVx
msW39CCv73ZZG/xi4SKatM/YEBGN/NapTl0UeT4TYYEVE9qn3YrfSpJmhQzQQ98f
hkuwBQzMyeYQya+/HZfdosMV79Wrkky98wzB0kkoTp/cfE1M144bRgkMjwRsIwwB
t1DzUMMHHHPtD646M4iQ3lkI8GeafTqFCaVX4Gj8PgNTNsLFbbdtM7E8d0rZkcNr
QaiRCq12f/VJxjbhr3TyLdorIWsnN8SEbQGuNVF17opvbl9zDDvf0VWxWiyKFsVN
RANJcTuCsr9OZjuDDPxMUfOmNCbJctWhXPJGpETRM4/ueVG5Nyn+Ws1V5etOQ6Un
mRC9+fuwQYVbYV57A77aalnrAaRXQWAFlaAul3+vXUJSXE4s1TiXB/7dFV5xAZZG
dwBdcokxv4EHQ+cTmq+1Ht6mHXR/Bn/sT3J64DUhELNQ+56dgmhJx4GUNf3EoI1g
LD4O0SQrzueR+dBwoAMDg0dmOBjMjaCVYjJh0VZeMn29KJ48xzZgvjEtVEuAvdUj
Q2GpEQKkr0qzO0ki/M4JEmVlFHS0ZXOilJtV13fvgGiNQH2bPO2tZv4+xMhUrKsE
C858jj6JpwNUgpT0lP2jtVNoEdD6giSyNOvuonOMt9qRlCfnNjEPExCQY7hOmrW2
exdnvjko39SqYsm+ZL/PY4wuawW8Uf2MmsZLCUnQA0IYRZSr3PWHCb7y0UAhDGXl
zC1DIHy8ZQC7dqBnKdpbEil4h3egXF3mczzrd0MzWKXSJPiE/klNRgTV4IY5Ii+F
8uJa+yiCr34cJ8pJ6GdEFgx9mzGsTdQbthueHXy1bJJsp7TnXhxE3ZGt5wcsMbqs
7/96WO4jODpz3+OnVrsU/NyWGmrUVDW9JuCCgKqPt3pWkG6n6paocaZ/F8vrTzbP
jqI0jPvdmT4PrwwfjO27bu1GhjPRIh2CiMaMI14hcjz6kj45xoPlWavvHXlif6Nc
VQF7S5El7zHEMJVVL8BT8cvoYicz3xkP1EeQeQtkXBDP8gy/yX3f7/mXsVUKF4Jt
g3rdHVmr8hoyDCvu2aOqRjho4Xv3XEjT+1ebOUb1sn84L8pFPWDmWt4qhevB40A9
+Bl5u5mP5xKi+eSZD3GMs75BleKEjOI7okjtmFEL8hxaYx2Vz50iUrDnfjS0LhaV
+cCeyQoNRmGoudVOt+UZ1mDS395VIzcz/9zzhznVOd0QzikiHe08J39sLJNKp02X
NzT5m459CIkMsUVFzZFu0+0/EjNhZo32CnclCGyGILOwbZaSgmpa1zbSXn4rTN8x
5d6zcJKa88XcqL5eAeHkciRCysJRh9fCXJ1Gmr7PSrVVBiVVm2wrXG9TnFYoAJO+
Ee36VXz7vv4CWhhUobovacpQZa2sxg323e2oimsPRilgVWPmdvn27XzSKe42AjUi
rXi4GTmthc9wwMT6MwS23IRP23oZOJp1OjZVuRqZfuOLAF6tBrDVD6+7OqXduZ7e
OPur9QfpOIh9kjU4A8Iv2fdHNFhkGIEiD1R0cQ5kJa+cohwLr5XhgpzUiP34ieIa
tc6vvoSSYYFgq8b7xJHYIS7bYDl3AFMoiJsg3Psp33Gxo54axg5salERNMkzWuIn
uNAIM/9V7St8gu7Su874hxaZBZHhkHx++O4YsjrNNAKlytBVHlQDxHmZPsmWfceg
G0/2WQ0udG0/U2prFodku7Q6JJjsmj4YfMdm7rP9yfcCTS+c0cKrn31xFKRTo4EZ
Cr6ozenlNlYIaXnDDwLuwLPuQZ1S9riIFT20cUBDCDXqHTKGuiSbHbBrZJc12L/j
YOZum24KgpAECWXAjsnXC5oapXs8N15AyhPX1Ck6LZASxAGaZ6oMz03d4a0E5Iyx
DFvT4BPsKsSMzkicwn3BDJbVnbkMaJT7nVIfuO1ZKPOFpV7RCwjycf+/017Jyv5M
kVOW86qCSOAs34FupXtlOT7gnqG40sxXrhfiVOhrqx7BYI0i+kXckJM8xz85Gr2y
64qQ8y9fESFWs6W1gDimwZ/3HaFK9UJXDeChfcjpdJx2sjULXijqPPoq+/xHvy25
/uN6uLjPhhNWgxvEis0TfJ+hEgjqs59buDVpTbOvEwn8SxcZ8w8yXlGFLIgghKu2
RVPfRj/48yEp5x9Eqr53JnH6BRJweM9ZjRBIgAp95hPLO4DxDY8qySWUx4c18bHl
YLPnlJYUD1U2LUEFzob/RrqoYaBT14hRNT5Kcpe58TVWns6Id9b+xZbEAIgmAvS6
hYo8L8OJCJ6KfMidUtSvVEC7686zE0hAiq5XTPe1HezLQybL1dWy2xeiuJYokrbX
OEL/TsUdKBnOQv8VYwrIZ+y0jNpkWzEkyssuXTKVh3NW0g0q3S0fQoByBkWFDt7F
DKXQRac5Js7D79UwrCqXWZbqaekqAUa9ss/93i78vn4HdgK/7PW3WCPbpAi9Q6LV
UOdLNg0cVPXTrVNhUgn2Q6Kwqe8MF1TSbuzNPxNWpFg9aM395KrArWFeBa2WOd2E
RoschdwQrRHMxZfpQas1nzIAw2w/6wxCJr5fMTZS2mv6DmgMUib7jGHrX4yF4rRJ
fLQd9zNmAJEMU9X4PU0W0GCnv1qqxnOS9ZPPiWY3WpcPpVdWm9Z9qgq2GJLC+ss8
CUhbiEZRB5xdKcfiV5JPFN9V528OIpkdqMSEiPUhpDLQ++dIl7hU7N2nFgIKM0VN
wH7VvzGNqfo045jpnCuydk5ud33Ssqk3x0xpRccP2RsPGm1Qer5LIxhH3ZBt6u+F
/mmcTYKwZrvmDd1kb4wMxktK+rI6JqwVVqwfMjossEtL99TXKW/hmPjmGTx5n3EC
TPwNXKF8yAK545ber1XUqvT3NtGl6OT5FI3ues507eqNGH68NcGBWpPFf6LrXUog
sRng5b7CXuHOjy36/nM0a3ElqFpLdH2cBqoX7ssDbXnJtjMRQcSr9ugzQTCXJUg+
kXrAOBM3uL1DP69OVf5U7DT8tgtXzsfj6KI9QtOwS2WkPSwAK7g8Qye/XMhsltI/
tcJqWyfd1TTuzgeV0C3I5df5tzSEJmzUp7RVX2qtJWS9fZjQ4FpklA078+W8wUnq
wTRh9OZQMwAzOu4OGkSRPd56fGZcnS6TnH4PvSfE+dA/2g25cmuPEplATVkLSB/7
VVYmwI0x+npSdkx8o6DvPFfFujb5VZKd9HNr0DSK9KwQCtGwgTBRxjTXLQP9FAhy
yUdieLS8nyBBy5nRT8HI9TRNeXcmagP+j8+tu/Xj8+ejSuhG7WPRxT9/IFSr0ycz
Z0as1sGJbGfLsUv3H1WX5TosHNjCFhcyTJJ4wX6/gYfViDjYhoNjxy9AIEuhg5m3
qZKMDYeOeDq6esV40i+Pjse3KUArO3JleNVC1r5CHwWDymQUfVTjyVUqEq6edKCo
3SgdErdLuYx68hBxb03mhWrXNu4hdlbild6f/Z08+3d50KpAKh2J+ecdZ4tAtQuB
F4BFYzucNPnz8mrMZhX4xQDHZMNCIwsoT6gbMK9uGnufoKkjE0KmSzm6TbHteHNp
/TrARemq/VpDuc0wA2OPuL7V/UKk/e653pm9feqs2gBxjqJKppFfbPMAPv7BgHaY
+xXgpZrTCjpVsc/QgO52z6wzjoUNSO5nd9IBDxtRLsQdhlVapzRnBjNfPCr7Am3Q
Is+AUBM4T+EQkfwxWCcZozczZXU+FEaTrCeW4QntB/HnQ0MPFG3gk3NDFZvBcGTN
9WnZCPBIi0wWJ8uQ+9/Lz3sDrz2gn/AHg5zAWS1MY2ZMaOCYMlrxcDVSrgwEtd74
uZyUsBL/bSMKe8PzjSxXOEgw/kMJPBFRdeGHzv/wCMXFPWgJU69OLuGhOHBfxhT9
SpVh417vovNez+k8QfTgcja1gjIJksL7DFIuUc3ghG3ONfwhuKlj2llykAw2py6a
smUxU24hgy1loA0RjMy7Lz5ngiPBZRWwRr8I/MuAxn+pgDqG5fmFeIaEniLpz4RT
nKDbixOKB0dLtKu9gJlk8haVAXUKDq4RzUz5Os6EQQn3Jk0wOTTXMbRUW0/itA6p
sgrSwEMTdPhPplpw3EUAgfj76QPqf5yTjs7CMcqrW/7pYnkn5A7wn+Dv6n47K8sq
1tOeDVP33B7ey4S0Hizb2ef9bnjD/8BeuObBj2fjk0OeMlDHjqNm+a4n4Yw7ANCc
hfQKWSijf6JvpCuQ0Lm40GE+gOZSeMArhK/Vz4dCnwmIYnDt3jPemWgBkG0nIrvB
hdFyrHpLby2ApbBLPxlXhvniw9uc1jxp6u4Td9WoRa8xS7sNl5USreKL87smL817
lXCIk48Vq58uIMAsWbWQxCltJg0e2oBfd0pLH2GNheIvoLbDLNEmSjdLs3iQ/uF9
JKcMUlfhhb917jW99NT4fiE3nTkILIIvVD6/auB9s9Rpffr0G3ELCydJqXRJOuGR
rwrcyQPglUG9tkj9LkJ+ReMiAsZZBnyeN1ndcLrD0Un/KqLOu92cXwa+FEzXkNpN
JMCMw3sR4e7HugSeDZOZilRI5kXlWhqe9segGGu8mUSIDqZHi9agtuBoRfxShtSq
Ttqp96hNYZD+f8gb/pgA1iav22qCgb+rKpjoCdnk7bFVmPC/+AFk7LPcrlHySH4P
1seXxTnptbOcK7ahhiLphtnUq7n26peMzkMjy0165mAROVwivOSOEd2xnXyK9pMx
VpHivnrfXvlR3w19MqX60Fy9xB3FEIc9eYZcTj42WzKlK1hxWeONdatNjT2GAKHn
fc6pdh3HiQEz9MREjrLt1bNkTq3HHVoJEDkiWOTUePgTboGbMxBoKI9f4XOU47x0
4rpdwCoWH/KI6pzwYSSChek61ZJCod+fMcs7tStBRzEfInNPNKUHkzYRj2EJRXwz
AKWdPN/zsAAU+lJRFImGfIMWA8X+GTZ1ayWFmP2veZCWKE3XH518pzXyR09CHBVv
+9H/xR5lGpnYtFO0gkI2Lcd5uXxCfKxY55VMG9uNBVSwoBN3NS87QyEtSDL8lg3u
rMxJF9w0o0i4VrIkE15Z52cKCs2xoLVjk/f8G4NyhOnS7C0hMINaxoBIf1/ROj3j
Ed+C5xRIdMc8mVw8+/rnfwCcdZ4FPzl+Obd+ii5s6lskWeB4UDCL2Xcs/p5vrSSa
udPTtnv1aqieVBb9Fe7tfIk7G+urdVnON7B/CqiiwqCA0gfeRnviBjCbRiFowZLt
9OjWUEYNOCj9OY0Ueuwiq5MJpxfPfkgjL8ySPMzq93nykdATv8z6TIvThnonebYu
yi2ky7sPj6EFGggt2qgKkPcPEC7jHNy4e3x8A9nAa6KfqcbQTzJeO4jKeSSc7V+a
G3fUAra7MUVXWiu71P5ryrKN6fjmphzyfD3iZLLLxoqV5ejwp5RwYeVxqeEZZHeD
uh2Ttkt5K1WNcpIO/fp+TbIoGHvn3c4TZX60NmrURu/EBv3SpF+UqU04GQrByKXF
REsHUSZGidKu/0AqBA8Zni2B/bVE8Sd0SwzgWehR/COSONwN5zViClzuOCulN8/Y
t/DE84vc0SXJQJWHl6ZHZKFuEC+DAMvigFHIQc4INJR3CIZhJUh9GuHUW+Mw4K/Z
OiUfdWWYfM6NHKhwR2tIPc26s6k1EljXuzUIlNSiHS8UxdZT2xjdL3aMBSoV6QYt
2KVYcp/LdtIt//Myr134ZaZ3tI9H8ORhN3lbSONdFpAPMjL9Bh5GMryf647DaMEU
q5d/0e1gUoT9c9V0Uj9uUCwcy2lWumGbr5Zb/AVFV1fNeoDWB7tNnGVhkEEqz5tq
JqWfOL1I1pz+llCRnq69Pmo0gSkqyCVgz4fA6PgykVePtrLq+DcUj931QEki4kdJ
NgYfzjohoQM3fZ5fu7+Fs+u8IFN4rtqKKQ5x7TMK84I/G7NRs64HxOeC3KMWD91T
NsXSdIODp8B6Po5DTZ8YDydAA6zlVLOl/VBmN4tMzXdY4gmz6FDBm8E2S+aAm15X
uJBnnKlCpURz+acNfcdUHNXS+jfA7jkWOylIRGmqh1pH0Bs5WIY4PqvA1sbYEcH0
UovWRz2Qh8bJ76WQMLmhMAgt4SBvgQbaHjFNiPMsJml3UtWKHcJLmFlDdEKT7c8l
3JeOonyWeWabNwV5xhFWCER5aM2zyjA6nSNfRirARDupkR8CtkLB3VWBcbTACHH6
21QHkTy7Tbccspm+Va+EZTR0zE1sw7Dm3X9NS4x1kWz9j84EkSQnE2DSeKOufSYW
D3vWnbNREXSfJkaYa4V8Ix2DFTsZyl93+me2ETu/I5diEFjap+3lefOM9/PdGDrn
iu7k5iCL561EaQVcxslm0D7Or3CUezqhm6RHoIAZD74KTwkjUNy5a77U60WWTFPY
DFc6pXGuBRRwY3/1H7VeQg9PljrqWIdbXyTIKyngL+55EdkNBxRZuqd7QuXqbmUB
1YDEjyWLbOd13T8raf4KDhXYy9UpHDAhp6HwShAqhWldmT2KCe+vvdPx6IqvhQPO
wBn4u1Ttvas7r/Jgl6PWz5EqEuA14Pcl616Ahu1fb9yaarR6ZhNVjhg1lMxUbRby
hIQbSCgNQ0LiFDvP3Ffn07SnDqBYpiEfMwp44inrpP0/p3RkCZBGuXH2zA4qQUJ4
OlN305LbH2qAFvlpZaHX84l1aSLcvnDoI/toVtTafTWVsOoOZNynTlcSOi9rTRBh
vgLVqe2xFNhhTnAuLqUaUREMORENw+ibPs5290aLMglX5MwAr43KoidRVUIoS2QR
rsV3Dj+pKwTKMMN0PVCZfaz1Q6Fu4Vf7jBiH3MVLcyhXkvYTiLnQzAfNWHnxOUx4
BPJA0M6uFwtd0nJr3UDkFJHxGHMsAoGtC5Zwyp3cvwOrK44ZKG71+8KxoV397YAx
oBBwKM57HTldKunH3CX+uq4k/hf0wURTVz0uk6la2hvqfM4C2rpXDQCAl33xNNgz
eI9uLOSRI0TxW3t7f2l8geItMAxiUgtqt8vtXXwPQKdA4zrKDMb/IK9Cs1OnOKOO
oR00lWeJDHabHHHx22gw8Zb8eSjE57xZc7yIwp9NNg5TqJ2SRlxUyWBh25974Vnv
N3/j2hF5sG4NZpX7mT47VQDGKlbu4QH8RCIRmtbYB79A4C8z5HamIyb7epflnQ24
aAyzaUjdHQYQhyQQEj+zMdaiFykzTN9Tcw+YOjBT6g7vnmY0NLxhxUmDPu9Qo/fh
qXBHrAC6Jtp6w/HjIUM9a5Tft8HBi4HbJioyHOx8JUL/kXqOUmiRsQNTLesTp42S
zGxaGzksf3Yk+5GU7B47nnmF4QepTPoUCd7NG9lHaMyEkhyhrLwZyDqV5Hgla7uO
1xTW3y9hFC+/Re3EPEHaf9aQs9tdpXHpcBhDjx82UaSY+uss7D0/fh/GgUShrLCX
jca48aYuKfF+JPAMPoro4h7k0By4W0BIJkDYfGAvg3K/u77SwFdbKkxsC9/bSzer
3zFP8tylLzwz2hVxpTbkDIZKdMnHRBGBjX9KJc04zj584joXBoExfsANKUcVrc8G
WjsumgAA+6T/Uo1+VXlrY4Vcr+JNNmbWaHuYjUKxUc5B6dFK9ajAX0jzkD86MiMh
Qu+yga/++xx3GHYgS0s9N/S1ekf6Z6d9Xipc8xqPsTXM+X0iQzEniJMFhdqADB96
i2KaBdEufoWroKmfSRNjysJaEA01bQA6Bq+UAqboL+5T/02r+senYXv3duBcX41y
Xa5zregGJQEEBUZSa3iZ3LNKpdBPp37o3wAGWKzmlSh5rW0Yvrvu2e6FYxT/mx/A
l6m8smRxDv26NCCgUxE9s984NJ5rs91NydYukZQ+vnNfclM416eDmVT82g9C9l3q
PxXXtTTelVMocL/7u1dKWYbX04nWgNn9Pl83U6Q5EMYBIex0a/yWaWAx+b+VbkCu
hU9g07zqmTYyMnssNbZL6B6jSMui+wiS6R2Y7+rt8PeLRSqaigmYwBu3ot7l6pJC
ulVSfmDZR77ihR4dkxd1/P2AHh4gpAIBzLGdzx5uE/ITJbjDhoggfmFNZp+MEVfD
yJBPT+JK5O6LmJej3yz5JNloZDrTdPBzToKLdxdqYPQXlvFPbaOxrKxy26mBU4fZ
spRcq+6jnKYKT7MvcmA7RwxIRQoorAY5K3yC5ct1xpaoG0JxLYIUejzwSsKvnwQH
VtCmj3hzc3tnzUqOfgLtlS5gpCVKjdho50344tAw7d5rny5TtQt8b+h/STN2gjPi
+ScO9WL2ZLFRt1Z25ZPj6LWzOLQNOiUvHDTfZVxZlOny5pTz0hQgA82sCiWKQ1IU
/ZTUifJaXsluHuZVeRSwBTRxVPGI5WSBXhziqntuWOEyZyN9MbUqVVNab7aK3Sj7
qqarzlz52huLmLzidWTN0Y9k7hJZud7HY7WFg2/XB48VTNfQILSZ6IBY/XuE38Wn
f42IF5PZI6t2sdNl8xhaUFoIh11d1h/GTYixuyYBc6bSe1QI2gLf+B6M+VVicUtY
aJP+ZhsHVEx/OH8WtWuzQtwlEV6yEuFnHQhmzJLgyXpW228hiWz8vI+E7MY+tnjt
67T2IXY7vDbFt3qG1oAuZjXEFs0rxLztOFhdY0W4gYpN3EHPFaluCE5OIj4jS2H5
UXrGZPPByWWq9N1fAFKzy7K4tRieCVl/QepYf02l64lIg2z5k5j/IUNQL61LBNw3
fih1/PkAb1pQTNM9emv+qxUPOQI9WMPANyzDA9le4d9eAL6z/u7Z1vV4V+T3DdVS
dSRSPPhmiDRvBkZaSnzWvLptI6BFLkCdXQcJBQuRkDCk74RRvkgxdnTXliInqb2K
Rst6SgyJmv1XG3mf6zgGEx44G9KVLwjs2hrkW5mQQhiEz54UfN04Xn0FDEme56Ww
2P0+dEVeLzJ7b3ZDd07ZahnaV7DufrExNbbJaVjjZSilDJsc2QUnoK3CX1yDU2lF
C8ub9XMsXfOmmHUwECcq+5zcx10M8UScJRjj3xuEKpSTW85syUdEuZNK2BB5TEXB
KPMtYf28EMW54e0npiD5LjLwkiuYmtikXbPeblIsqT/xfJjiFaaRBlq/sFtZEJVz
2YAETNhNLp+vhsvjnBlI0f06QAIQJdzjPPn8j4jHY9T0r8QqsfiR10jej2JIPQnO
696adnp7JYfzKJ35j4eiFUIugrtoaxMhXJqwEhcnrN4S7IBJp2I1mnL924lYr741
S/QZaphUGMrPXrtUdlChITlGh5BAbiuVuTF8I5+uuvExbpbMs3KwrameJLfWAy+g
cokEg3wQydD1yLYeUruCVwo0SNNG4gZb5YKp/T0H09/7iPO9ns17/cfsuebdjrPG
UXWTyULgdx9YmfZOh3uKEskC0MTyVKJVSx0mlmA6D9MT4kaSiFIK9uonLIJJt4Vs
yR2UEdcIHNlUnOMMTjkmPWYR1nuDCPpihAKWjmK8zDMGQmBetuUGrV5uoMKtidDh
e13rJv3ele7DNsfUhco6efUzMxPVkIfEtTet7mH0nHUu0GALdINnP7zO02nvFdM0
e3HxI1760QiOxlATdHgDEQENrU7W/5bq/SbieqpfsQcNmEoOEZXeqFkbvOzRrbbm
Li/Amf3LLlQXiUbdai+pTsvbiD+Eaqv+fRCpBJM/FJ8RDCSEbx+HRbXRdn5Rc9e0
uzLMrDyIc51NGRN0CWxc6thO5fmpKpcy10t4swtzp3/w8brgH/wKumy0nzb/xZGm
6wqBDwUKLTuwqOEy9rMh+LOcPFVEVJbG3CYVAHku3qR+gbdCJ/UyRRt0o7mQHerP
bMLYc3Bry0Ku4kyuOiWGoYV0z/ZIEYjXdtjlfr1bx87WLCT7zGtgL3N3HtxBc2T4
tXe5UtmGTkPHeqZX0mqhj4BB3O9xIkjWr371zBi7Bk6f6H7hIfxF48ui5Dj0ypHz
VNHofZHL6VJHliqOH4zNbT6O+yE0sb1WsT9xu7s2DynOZ6NpQy2UHn6bG8eNe92g
GiVbWvSZ/DpXEcdTrAOaeFN4XO2p8wq17t7Yow5LEGh1vmK1d+QAAjzKN8imS6bc
ArnAmtaHk9r+Gasb/CYhpNQNIdsu2NHF4IIYeQO+H9chyeuBB9dpLnMFa9x5EnIM
zzreEnQPOue+UIyXnOvzvWB252hHTZMOAsvxfI9ckHXsX3zr4jckVAKGpuPJml3p
WwJrB4WoYiXE0I1XRyIPLC/dWAvb9JXZ4sG+WcziywK8gSNLC0lSTntZb7vB0r3P
d+vSdQFYZtHda2y4uYehpR529gU0hpSC/TOhq86ZUh1AxxLajUXcQ0NW1gsMfxxM
5ndIA8wV8gz8WZN0hNojVJ+PBbmpVIfcw7Np1n9y97q0WMXYP17/lGdpaZ8duHpb
0d/dRiT99/a07+Cfwa66hMd+R9FqDzxcDKRlX/CLqiPkx+BLLWJ+Kwmzhze7Vz+U
YXI2CY1L6lPzJNz1Kp1iRmYwkUC+AdMaDtIGqCfMjUECMyTGzTnv4H/axHPznWC6
v8vgwzG4+QUiENT+L/wdd0qpmZclwzQgdnp3KX/m9DzwvccgpZT/hhcpxCUD0cX9
Y9HxcN+gWDkAJ8QN+nZzOSLwV7rpUC7b9brjXL6p9sVz2s1z24sL7T962EYByG7L
Ue/uNyNPg9bI5Oi5oJZpaUYa1t3dvUO/fjPU1/dlC8U90xazvUZCAo4o4lcNqW/9
/2dMOt2gF7w8RZRVI5xP1cJ5f80UG6L2qkLU9VQHfBepZPHLQKD/3jXxUbAIDsML
QAlGo9z/wVtf0WCdW0AU8I6eexgD3TDsEJmyPEDWocB/VDa6cdTLUkexSCnmYuBB
T1QbW8iiw/AGS2fK196IhK6q69FbfOZg/8QoZDN1sT5Q4jJ6p/CBo0btDKJyv/AR
D32y/ei0Fi6lu6bAGd1cjZN/ncWCSbrTT8JoNZPrcxPV2DvBQAbqnIESxvK7r4V+
wdIjIUa7i2lWYkzDqQxxN1h+lwiMYjAa3aedlQy28O5cFYrvyCXFRmbdCP8lYCZC
MTJHsBJYDmHciLrQPJCE7cvhsmlsDh0unotcK2PlZS0Jcbbay0CdAyyq9eP//aCQ
bciibWK4eLOBL/MYnKXeyXGSCeGK6a8JFeppUsMN37glI3i3g7Iwoi78MQdpLnhX
0zwXo48QIknvoicQCAho2VyKMctQNTjUbkdTby0DRopJ5CuUx2jk12W167jD3soW
zOWlZEcpGaaV8rbES57ZTI5VU0Om8eBl9KxwkOq6aGOiKhnfYbMl9mA53oYIAh6E
hmzY8sf636cEGgpgymhgNY+rg0kKahd/Ad+p4LHXXbIOVxwBUnSvUpC9j+OQeW4T
jtbsmXRcJXqSUE8Kx1WDZVUwUn6VXj6vkRhzlQM7E2wM57UAZyc10SxpD1I6jntS
Px4t3TKi92Y43jv+k+gyXg0vvGtmfQjgeHQrt2eS0+7MDBCvYOMkZxZ+08cMiLDa
rOSOphASswxEk4qxS6FrXRSv75fmV87gywD92TmZrFqiRrBgqsPnEQiJ71ZC/3Tc
mTeOe02tRDmLBqsbn2IWR3dUFa+pr9l4E5YnygiC1NNbDWiwyx/8JBY6cWXKHNI0
icRfJYEbJfb9mHWgpvOApLdx0fkWF3o7dZh1kgTH84h/RmxaBN6l3gTtwt0RQucj
2fGe2XmM4DZk7lDLh4EU5hMKwz+PbRtGCcbSY5PJg/U5QKNMLGKly92WRXm2zh1h
OrO9q0bfmw7d6acFdNTseGO052+8eBpNMduw6npAQV+GjlTBKpa89pIoNEL2DI4D
Crn5xCX/W6/E3rIzVsMgkCCykiO+llqhg1Ob5uYEtDieRPZuCdlX0yzzyuSLko2F
aEcY/TrAoh/4T1uVDEFGOyUxQ99pjHHA250u4vjLlpBR6YIivZ00AkG8MYPa2Aup
M3syhMMCN5tPeZSaycvMPXFOFxZVOhx3wm8iBC4IAM7PmuCbTeXlcFrNB35WbkYe
1HHj5s7S8O5G6ImDsLpSFQQjSj00b5mg1ABM3Bbqtn+rGZcUAWKcjJWxazRkRPg7
iZJ6aajECUgkaE1nO9wfVqAZI0fWJ78x5/dgix5H5cfeubB99J5qjoz5mqkMwqWV
FwlNDY6eUT/xAGol1jwmDWx3LP4r2UbizHwBkT3TkLxnnBaK9xrmHV9PvnrFQds2
3l2z81BiOuqJNon6LQJ+S15QvOXunAu3oGXFX8S+yLoZJVBwENNO8uvemKa4RWqu
lEzJf7Y8SsBDUdtPfnGT6ZcV4jG274FSAZLnDlS7g28KXUzreEOITz/d58gHcn8Z
0GG9EfiN6smnwI5pAZzs+CMDMYSxGUvcIqaEkDYbmVqBOl13qy0j2s3cjLjN8DVJ
lKSm8Au1wPugBQsZpA6IYy6ionU8TqZwnM9zMPAMcg5Syiz8+IfN/JFmumHl4csd
eDibXWZJDxqM9J75wgRmMfJfkyzaDCvcIEoBlepHxOcZWarE+9R/xxY9TVj5Hm6v
wTUqgEcM41W2gipwwyfmuU/UWdrVBALTOuQvenbosQk2x3ntFSgXSR6vesQzxaQ8
USTmk60rba49+99faK63WYLrareyZyyy8qtwQ83i+EF39X3oLOwEMSTT4jVfzuNj
56+RjVlymG/SGOBZo5j1WhZJo2S+Qj+MS97LrV6KgXsHOE6g5OXG2up8beQLMAcv
OYZhNyD1lA4JDD171aFEAtNu1Ab345M7RD51DfhEJJueah1pBNnuj8QoFovvW7Uy
4YagLXLCZ02YtT+KwalCDVdgWd72u3X5NPh/lZkX/m/017zZAkYTlPKvX9u6POvO
XPpjEj494n77bK9E1/79He6RY0hTdvrCZ2Bsfca2tQJs5Vr0bSbAHsXPeH/3Ztb4
sSga28DUhG9V0xJpb8O2Tv3yjyjW2OaJln+qoY/xFIGtd70FeIlhk4a1kaHOtKpz
nPsv/RmWGpWchkgZ4sC6eAvl1WozHT3kpTqYyCzKxEarvYrUN+6Ln+uv0wuNles3
eL9bi8chdGKzMsryLSIAGZC8QvCIbXVRhv2FnHiKBIoGW41YjduzxMQy4FgGeS8N
PNXxKKrOZl0lQuBdSDCCvrhkYg7u7TB+Fps5xo5r7g4=
`protect END_PROTECTED
