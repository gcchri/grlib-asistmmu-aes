`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YlGtj3GG3raA6StAYLcN6npZx73zt44ZtuJ/TGJBzusldpVqxV0lsLodbw2Rzua0
DdklQJ7oXJqzMKsHCD6Xas7ASKoQ1D4kcTLz/q0hHD+AjZelHPM0cvEDbuc69x2Q
dcEIJadycutMHkFDXZZAchMJjapQO4DzjK9wE+gvqgwRFoQrKHTo0iSpzYZ7lCpV
fO56YBjbqtu0b2SQf2vfbg+L2oUhfcyeOwA3L7cw2lh9m6Wi/2st+9XMIoDa+0BW
WbiDqvN6+4jtYdN+d3f4AH1RlLcgmN4yehF7eIaAbJpeMFOSLEthy7p9DVs++q0a
cpnU9WoRB9/KmCwP7cYgaXpCjYmpF/3oP6fKA0eCMtV3Ka9noNVCx37FbpA31MXJ
QyfwQtX5TOMOIA2KLSpo070UYa0G4aJHCiEMsk6J6fM3WF/9VUqvlvyrJonaBA6F
KCpy6vSP1k1bbZAqI+iwxG/SU2rPgK/22DRDtvOByU5BO9DaL7CbSszp6qleIZle
YAJvx6+VCeRA1Psv1XsuOxTymjNJ7WVnHf0685qUh3X5CffKzaB3b/Nsb04/wlFf
1CjKQaZmrQHlwBlb4KrCVIdGD4fhhyJlLLiOnh1x6iFSrPEvN270SrWMjnhgG2g6
Z2sXYaiaqggbloFCcnADBLaO3WhpO1ImFKKMkhvQs5QovY/5Ordhbm2XBvQsslp8
e3411Zy9XlbcQneHFXDqvmmeCQ1EVs89Wt3GFzWy+eG2QWytmyvwjtbLSMEWOqnw
C1HTQQjGTT2H5aFQVevHvH35PflDAm22LlsLe78CxZhhXoCn1WaCxJ1IXCPz4Dgm
qz0L8tfz0AKUxj7r18HgzordHzNHTOIeJpPFtN8sg3+OTigzdSSn93BdMu0G4VDm
8YAL4AtIZB8qnUvbmLfDTDKPBDhLquF9J+xOWzQJifhMfbl0oTtehKBUdyZtDoEM
EcXLWqW35X40I4zrjOzkXCLkvY1x9XubBLNgWuUpNbMn7PW7aDXjWmPyyw7TEyQ7
4gOgr6b9ErA85bXwE6DGXim9Te/Y/hhNZ877cnHt6iooSB2x/wyqAJL3A7nM2U++
Teswaj9JkhnNDDnt9WW2L1zhY/H9JaKpB4q3xfNLjlWctBKyvCHbHn7VkxrsUgy6
MnLWMz1IYKS+KqkrSU3Ut8iFq0kSskCms51ZxKIXoofnl+L1rFwPWUf0Eh4YQU5h
S513ZKp2iLOM7jDu0rRq0wLx9w+/rajdRkqTOSMN3gBFDakyQDQgIbZ6xx6OW20p
VVXZTxBV/pE1M+cywSWQDAnuIZrlOd2JFBHZM05WOQv8CuBau4onvVrYGZ1f0+YX
EKbjItzcBPglZqgv9+iLZeRjspVhvVkNzGffonwSCIPiugA2TvvKYda0Zkr6dIiU
gCtaMXc2TeCzGrAYjoxOiw==
`protect END_PROTECTED
