`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xj4XCTukudiLv/I9jtnS4AbVEbEIbCB+H5MFpUQyRxwp/MIg/VCrmfXhFyptszn0
s7jBSmEfVZGstNL/P82QkxXGDKTbmsupA5iuD6sZ3uW9ev+D0IkRzHS3R9WJhaJg
96vNinWRTu7gud72/CUYnzy77KIXrzGhgvMUwBD+SyEzURH91TUBLLLrfPIhorvT
bdsDgiFrhFuzDmrD6fo2fC7cMVPdmEhQtzdtGl7fEIYGHRhyifiZJsRThs7gJFIy
e8JPpHmrnOnF0FFFcz1vOjUT8HhIXXZEXHDe4VVK2Qg3K/FmzCtdYm8Hit4+Rah+
92tyeHiLQg2s2a5W+DKF3wS0yuNmeYL1eSC0Z28GF39p+46wFHNxHq5EYp6CTi1A
Ql2Hk+6xSrl0SzpnSB6Z9sz3ZO6si+LntMOBeJHNwLRBrdFtAMZX7Hs8b3ehusYX
9UY8M8LtB6ZLzn8PoBBMFR7Htrs/jj8qJnTp9VIbYJP3pwaM7wYA1gqgeW5nQcSo
`protect END_PROTECTED
