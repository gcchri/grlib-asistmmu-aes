`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1scVkLCOOT6AfFFPbcAfc2rl8Zt8915erKL/6DSmrVXdESEH1qvGjwTSl65YGD5l
r1jeTZ/wImW0lC+0RAGOF9ZDzGM7QvRBF9hwwf49HOWrlJvjpxIXiMoIKXEKCUnx
aLWUvlBB63hp9GgoNGldTnHseUGe7g3a6PCGMeOokrD5vPmGjkoVOWmqyJV5C9n5
e5994LXAVdzr0HsO3QvCnIo5fHiOHlDiSGmywlt7nTpM7uZ/diyAW1E02AEO7InQ
UxVW7YPhk2bKcSHiOZHxsRRvJCsK/jCCBMtPBX4ovoZXgB8dlAp6OLb0y9Pcr21l
m9uP0mdqTY7hNDGvZk8LBgs01yA7RAEScFdNOS+SroSuGf1ti8PV6EAgyNjnCSmw
`protect END_PROTECTED
