`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vx7OlLJ95DaTG+VP1O5DoWDa5AOiyPW2bJFfJaBsR/WPKg8neKqmf4Fnhu2dhAmf
xLqI1IRewHHYMVEregdQ05QPsJBh2Uf0Pms998HYuo2skbeQ/y96A5LaMH/KDQA0
M0lCC/JqUL2c5ZquqXvf8H78AfubTy4ON0keiVSVfujWas1MnYmtRSM/Mzfgg7gC
ZMdZtLRaMWFWhFtONivMogdNt+beU8xwm6F7Z38eO2chzNZ2GR0HDY2e4lCFwOlL
Ax7kgvexuoVYmxIM5BNzDQubbiHGSxdcsYWWfLaaOhk=
`protect END_PROTECTED
