`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UGmFH26EbQDYsnJAVY6ymSmyXQ+jK92jBTsOuswIO5ErdULkc7wshZqz5lAelCqG
LwRAbXs5Jejmbtx0W7CkgRbt++nzuP6k4aqSmOLoJh4Q7rYOhfJCeWCN8h6n5xdL
balVgUaixpoQaPYuvBq8htIZw+qVa+/Za2dByI/KEOYisMH9BaudKpcB8M74KyIw
z/ICtlRQEh5dq/Ys48dg+p3PpG8no89zijZ5PwKzATr3QoeeAA+IDdejGAnen4mc
xq40tWqmAXc153SZXP38aXpTGBzfq4dV3qVa+sgXpmsuCT2yaid0f8UMt5pi75Nv
UfAd7zoh/LfSEz4l6R0lLsh0cSVaMhmeEm6Q0m6z8QWikgsL2kYOjz84iPZPJeIM
VFyF/enJKiNUY0qDOFEOHw==
`protect END_PROTECTED
