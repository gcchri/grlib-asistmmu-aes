`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r2rq/BVYqyZN49jDlzGnPnrYrvFXkq43KwxdF0o2rvieJfS5zREz179ytIrFiZwZ
B11ByT6ZllovmgvwlmguEuDxc2aBdt3Te2QG9zWuK98HUUfc9J0f3DlDKhESXAXd
Fydw7oa5pt9F85eyFElL1nGg94jCMfKrq+OoEHI5jdvDGcB4LvrnVFIRS2v6EkkE
oNJpxwoSS0e6RmiqemUzyQ9GB4w3iMzWh9bVnOOEsJByyr7ivSRkb+XOn9p0beKu
S6M92tMhzhTPWgA15roPdQZW2mw1l7BdvScCdKNmrqOF+iKmWrpTlCC8b6HXcsvq
2f7bOhzHq+pcsPGxcVZpS5j75Kn8nzpsuwC8k0WMM42PAUp9zSzeaX0OdGLSvvcn
ETPO6F97eK7iAIoq1sZd0g==
`protect END_PROTECTED
