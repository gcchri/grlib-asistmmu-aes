`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f+1VvHCL+IsuVJyxVK2XBJdBN4fgoxwhpzRrzDjOZYyZrCRElbrSd30BwCPrX0S+
EbO69W4OJiiYXZfkS4zfDCReT6NkujtSf0t8C2Ay40zHJmcjqaVTl2MpfO8H4VfC
9Qr5Tky2HWFJgWi4/clqyHOJjEhUsRL+eMAtWDDRYkzp3s/SmwyXHqDqOJ7ixzED
LK3+8grUtcdUZI4851Ce4t9UaDxiHCFBO3mCNX7BE+xlBP9scHk0uBcaYQzL/aji
7xhQ0RJQjXx4fS8PXEei12U1YUr9Vptam+AWSdCdcSaXM5BVSDD/SlPA3G0yYXNI
a4E08SVWq6F1wArgS/P4DLDyT1ntYXkruuzc7izGvsfYC+3xCj5MKhVt3r5DeqkP
p0E/MoJShuEOrC3nyOVidg==
`protect END_PROTECTED
