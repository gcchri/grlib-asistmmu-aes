`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D/ejEy7p0KDxHEqPLSqdgKNdaYSR4QuJmMR8hR/RpMetYhfY+mRmpYU7gTEGooQi
L6gk3Jp/6grAue7vAwn6rhzS1B/mYx5o48ERSb8BSjG+VlAXsDqnauGM8KrMc2qB
EKnMbTh6xt1QwCLji0b43Z19uX/TUsNjNCwGT8DMM5zFQYkZoeWxKdClnTtaStUo
HRTf/0l7hFucfyDx0uuIIUBwPrLlBUVeWOEbxjY52o1G+STPA8PpFmGakpntQvHJ
dZ1flCqw8nQAfziixzwbaA==
`protect END_PROTECTED
