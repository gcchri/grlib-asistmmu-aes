`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DXmU+HKZQXCT87EseWcUj5mPdSgexQHugm8gcTVd8vYVOh0GHyNxfHvqUhBx/i2V
a7j3hyf/C16i63YbZr5tjIYj8ZaA03CcKjz+Ll36eU16PsQMncDlM5UJAIkK2Quu
iBkg4QmferK6ePl6qpEyHpPYl6Hsv1nu/PcxwXpZFNBck7o689wZUKKwM1Gh9NY8
n+PnxO8PZ7Ag4WCASTuFQ6y6QQKjFSHs5RNxRNc23D6AkW0g3SUh9ShktUoss3J0
lOIaKohnopvINldGvr2dcBg9xRI63ryfStz8wI2pDSl71wqMyoN1n9b7Dc2Uerka
6Dm0Ki1PRNQmqQ3ww66RvqZp8dMt0JudkDJaFct5WPTw2vV5bz3MVCeg/dJml4Kd
dY71FdYFcnIoETOjoFVzWjw2Vm72FTEQ3Kjl1Lx8ApYRDAjsR7MFdZPOLGT3eeoy
`protect END_PROTECTED
