`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tv8mUUWQlSm2WqPqKylipWtsU1GqWxYga0ezn2vklAvdMygNzGWaLzMF4RPmsr8J
ReWTbFMf59whF2lZlBZ/KyM6Ibtx5wa3e1Yd+u+QTa/js7XX5GjDyV42AaL/rFrz
Bor8ZJf47VRQQAaG1CVfDyGh491eRdwpDs5xBNyec/EsSmkR0kiIJEWZSVz48DnK
/zwABoXWZd5X/m8cLIzj3WQhHhZO46NYAvxNc2BAqQEytkF8Az8KJumilamZnGUB
qvaWpZK7DRTxAj3QNvCYVm2pRc2+BynMPqM5F8CD04/9+YGSxmwEb5aLwogB1uOK
dLjBn4CHgtPggHRkLZWBZ+Qbb/xq+sTIvzwVw6+YpJPjNxMYpjpZ8OyNtjpTmkKu
b7FWDnPGIBrG6wYF45h7EWRiuuYlnQzVQuu3nVg5dfZdsWQrdkXo4r1DBgBqDNEK
A6MadPvKn1RhLtEhqTdUWwt5MP+Y7ub3dd8MjxDg4UMX7PYBa4y5COeaA8sxba4y
l1cjZXtf79hzNOXiiUiceWVMdPoY8zUeyr6pbIWj1WxxLaohpuvuYku2Jb7n+TT1
N8H46bgsHA2AiVqx+DJ2iw==
`protect END_PROTECTED
