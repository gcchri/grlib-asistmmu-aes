`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H7P3nrLkl90qw0LpLmiqHxp4XOvQuwMhdryql/JQqXj3RiDDmNLPGnjGcwhGWc6c
emsTvj4iHkQpQoAjz2+YUAyXuDSu0wysRaBQVjru1KIlNVtfyWc4Zd8N7r5EI/Dq
fmMZy6QaYJiqCAwpL2KX3q54DDAxwXS3uyUSibhk8WBCOS1PUTXDZBqNOv13Rl0e
9ekW27B4nshvUt6keuustT+Eed08NFBpN0zLTkf87JEEP1ppkV4j2GgDOx7j8wwr
pMTmIr34Z46xuKPiPlbcmTQLLyafcpcIYcSgMgpyUY7cmabJUrUWA1SB3Av/3hWI
9FOaIZcY7EHvnYqJE0k+wSNwVisQfqny+237YfwivhhZ699cGU6GBL4KL4/aDmKf
PJI63oeu0zJs/zy+bh9kZQ==
`protect END_PROTECTED
