`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t/wonZNezGhPfgOIf7vdEhMjiCBhtoXpBADllN9y6Mqv5YIorxXeJbvbheSyKrmz
hQ3PqATdVLqXstUL7mgrTAYkTR8s3h9/gOKPUFgvpoXIW4Uxm4Z9uB18lcyJ+vOV
1br+8E9uyq31I4ozMDZjoXdHtrtrbcQuBKMxohfP7WeOztFSwGuU1FYRl3ykpBPU
2ccSESvoxWM/7m4BPOVfnveAs4eoti5XXmzkxuvMyq/taIWLRoZTRAPu4Na/7nzM
ohWAtqoJEEFJurj65mq49KUw+WuR/kVDBd+7G+2JK2K7vcelLtTiz/NpGkisX/oX
7/F1/gCeulI0jKS7JfM764ZekYcoKDgi1NF5sxI1+AYl4i92RatoNI9sH/3T2nlN
IrvUNVx4/sZESa+RiXjtmELRPMsoGGD+Opt++eXZIKkceVsmSn9XebR2kUO0G5ZC
lLxtG1bah34kzY/+4RsL/y6/v4XgKdpb9iYDsL8LNbQ=
`protect END_PROTECTED
