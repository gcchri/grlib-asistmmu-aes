`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WEkq9TQR02qOrFCo0810Ib40WeaGlr2Mb4SZ1+xnq+3+hW1+gmBQKfMGRTdVMS9Y
oWaZvel+L+U3Z1dbpW6UTjXD03EA2jefQ8upfJNUqAzRTIKPDpoAhOOhLnamFmGM
nSBHPLZXFFr4n8Sz1KTzfosbQ1KtPzktIt9rL2l/uctjdLYu2TL4jv72q4X+kgRQ
vVb6aOBScIAdtxmYHKI3ELwX+6QTFsHNycQJnewZAb5sW9s3UiEx68PhWA7mZY8a
aVMDV8EK+We6qmSCCapWE0+Lp9YfnNKE3aox+E7Y8/sgCis2IhyqWlPmo0x0BuAI
7yAY1/Aomq6+i7P5i7VIHL8z2KZv07rGduS+YS2quKL1gXO9FaSLGBIJcYgDr1PC
X6RKwMDKEnay2gHGu6fULEEvr6v5RVHf29vsGqYyT+c=
`protect END_PROTECTED
