`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O41ANlCvi0uNkbtg8Jnhp8KoX44N2sL+fs0X+esKjJPgK38Zl2lTIuF8mZY+fTqI
lIzn1aJX/IE69W/sEQ0LetpW8c0o3zcU/unHtLwu9CNbmcd9CITxJmb/ys9l9Hc6
uLFMqJCMd5b3YP9bRTA7kSAyfF5rSDjPYIRzCmpt6SKv1lklW/OtLhW4EiDEPeHx
wwJoUHLndJSqJABSlAt8yPD6CW5NkblYD73JQKALCO26+Uxm0oDS4ML/dI7fBM/h
1V6j1oogKsbtsNrBwLOr+kSf0/oslW/8IqmjLVaD3kQPKD5mho8iTsg9VI0IfaWT
/k6Zy+tidfu9zYPSQhz9whXh+xsTScYDNT0RViowJJ3UfXFnZzPGcCEIgYZqla0I
AvH7WKdKljq3wylG5SbSz9gqAM8VrK5SCgnTFoEKhXOVE6YZ62dcarpbU//xPMEe
uehjcHlInqiERsVpld0xvd0wVdII/2K41dCsgRa8SnmPEr5UMSBWLQlvwXBVoiDw
E+AtAfEFNU6qY/O4fYMk//0o6zDqHYF6E4WUe9LGAcFMzTGAte4P3DtJDfpflrPJ
0tnfmbcSydi7zMGPNMQwTq2ZVaQ3pqrw+SiYMUr9qG7cq1tp/UJj+4gbUfzirY5e
LLRMCjXsrdZ3Ym69hr8n1AUYd13yEkf5RH5YPJcExVWHna9wd2aBldqgRgeTr+6R
N2u8QuU+F8ohl9P0SevyfGeq1bfJ5tywm6M+1r9IXxcGIMd5+B/PucpHcAENWbGU
WKKbz+z/LS5mwvb92Mn6X7EnhMA1gZRB7X7B4+NUqDeAFcn8R4ZpV3Hef2Ey7yA0
CRUfnCC+YLEs4goC5dG+TX3AdDL7VpLCBGCNWXniP2xvWrBkqQBPLzDh7nBXEK1K
aabejRf887Ms5gUDso83BMtk3QskEegxh28cXFo3GO70Leu+Chz6m6hlAAK8Xpu+
dxikH+IEh4RHsSyy3FDvH+5vpcYmYlGA1N1J0jiIbfnYt3IqIP0c+XrqCMHJdbXu
79S6xSGHdaj1RggQFkGlvPq27wBvKwjrt56QgFyhVTe1bH6+lytOuH+iEIxpuB1y
VkoGiQKrb+mq8Rz8txjPRIzAdX3wCRBhdB8kvyqp3rBS+8O1Zwxbf+2m6tt7RgNB
BezoMPxFVXvl5lA2awscV5U0idjZAQVUB5ow6EmZRO3oYjJ4zU9fjTqcuCpOcwpC
z9mdfQiI3zAOm/1UcubqYODRAAwRua1fhFjxPFt6DskuM5Z2IexA/BfyDi1F7wfH
x4MgTimt7BG8Z/JZVOs7u5nHRUHA/UzGPYpTqds4B5jOTozL32vWhi+S/odJQQB5
PfRj+QD6CU3E9+Wcbo+n5X981atY/cV9mE6W+UyMGiRe3pixnBu+OoKgOBJTFtuZ
tG6osNKkxonugjnkYmBgNIvBKGybTn5JEWPp92jqu3vTvp6BaFFarx91dxLjwviM
L6z/tJDvv/MuraELkN2gbIi/vFZi3MDsVrNRPpynjw+euI6RTjt8NaHFLqTQ26Z1
HwbSAjec2mjlMOmTS96ZvxseXa46kLmZNvY6X8Jygm5k3n2Gvhp+Kr3/YywLU6G0
a94r+ns2uXj/6dstWI/PxgzYIhwAJiiLNCZETuJoI5gH6/9BZBLiXFkpmglX8Afh
85m64Ir+sGwpjSknyxO9XDmce7Kgp8vQEbFPY4pi7+0Rc3xAOzha07luLhY3MF5c
DHi3RgZixlIl2R8sDM854973OrT89QH3in2dKm9qW36IzOtx9/YCGAQQ9I0Dn9G1
DbdpWy2ZKxMSShBWGa9xlb+YIUH6DjxGlhcKI6YnF7b53zLhoVXXKHYoxQ/yZHmf
4RUogQ/nvMB+d1L7VjVhdVdULt1xnLabjAb+RLT89bM2qW6cz/YAESJIpjISefGC
cVwQMGMqg7/PogpveBq9CxFl8l8rEjN5zz33bBGX9vFYfWfFycDktX8n/K+q86qS
D8ITZj61jNykSNrYkJhACtFtYCSVWe7ROySpmk03EdOLP0dvGck2TlQDg/XEGxul
/zjAz4aSj53118B+xjilDpGT/SGC2gwt0u7GkxjrcpXIf98rydJJVmgl4VoxMwDf
ntMn1JK3h/MPbl8uArUnVX0x0UM9um0Uoe8fAJWC7nqVG6NGGKQoroqyA0m86X9V
BkvW+SYsL7ZLOLhNfXYvwi1h6pz1rWqzAi3jsXqjzmyPjsp/04IgaGaBwVwxY5IB
y/k0qUOkk2PS8PZmRXoVwEEWuywvoABKwCwHYH9Fdnm9D3viuVfulkp1k/Skr0Ma
w75Y1NdwJaX2NBLCbrHO09MIGEzX9Net8hQwXS0RWjuQiEGjhVPwCeaeAuzbCVPV
J1XUC83Tv7EMj++o6IGtRmc7/8V/EAJmlgVYRNESVZ52UdKPGwg8+piOTsIuLgsQ
e2D4lTUI9qiudSohIYaf3UOuB6jwJow9Q3jKHwwCR1QqvwtEcaU8N7OaivsP4DfT
sdFlonfjQDsXF0QanAgm/6bArr8frA+cZXoesRQNXRTcAdploTyYVGQJT977sVfa
8exqrGMpOLZ7Zc9eENWtgbGrGp9oLOu/vI1ic212z6T765VxWw20r7XR6lJoE25r
Gm6DscmMIBFpRjBMY1iS+2JS9gzqOcqiZtkELfYGSMkbjnVuisqF7lhsHiP8WALz
sXu02G50e6uASx0i7pI2taqEhICOQvu2gKK9rCrZlr28fgOiNoclRZRssM8MHZP5
5WrunH5e6Uq2Xh5vY1eyo0zJyRjFy/02aLuBARdngQQdBqwfNGZXuqZLzCnpjGzh
9tUq87iK6fYMhOs2UliwR5oxt2MqF/HkaCbenV7LXrDmvHndiUqyKGhRWAvH7GSB
8QKxU+JE3Gwbostvw2dxNIptEY3ODnyJnJIiehFTrBpIQzDPuvQHDa2AnWn+DHpy
mv/A6XrmTtK5flDfTSi8Ifqf8HAp9c41h6KW126xUVwO4E33yo/AxwcmF/fzlPb+
usCb7u8pls/JAabkuPB2gya4f3EzAAQV62x8lw7xIWbKhak3KDqz8q7uOqUF+UkX
mL9Ivhab7eHkmRZXLFGd4X//Re4bGXgN8AvAmmRCREzZ7egKvvS3uMBcn39ULBex
1gdYFUvSXTHM5445m/nLaM0nDD6Hv3th1UsqusASdXcy3C5HbEgRASXym6ee/Kgu
jKZ7KSxpixkRU6tknogZyhT3L45PP153SHtP5xmahhIITI8ekhDStVHu2XuZr8wS
vQBe2NlryJIys7y2k6lveXACXcIdwAZCMcSSNwHHdyq5b2cCXsIWEoYtYhRhc2xy
e9lLnVzPrgHXxxXn56g9xnjuFh9ukK+q7e8f+O3cl+oOcfODHMAXCQQ2kvx/dbYz
JaBLPknv8Qzbjf+b9zRTq0Lz96QZXZ2rtt37uLf0LHWq72RzNgXqLOtLdlll/XKi
ruZXq47+QG0eXD5ASLHjk5IJfG35N7RxaUUxFD3uW9l/0xXyDACQqlLdGAQIhAQD
wOGQKgExSaDHCd2kBASMOKs5ULKFdkOddqvk6Mq18+CADFMgsk5maFM1IAQJ05EC
N0aD4aFhEQLouutPljhXez6EpBkctaaDT7H/a2JFuDYNy2+v9zpmD0s6h0jx4n4N
dQGJSHNfBXtGYwJgkJmX27Z7Hh7zYeIbU3rD+TItG9aLeZEX5yUOgCW2LdgJUh3N
BWKlyPnLEPi8vDRU4hURYmKdHPkprJpW/uSrxeKseksvoTUyLut1S56XTM6GNY4q
rui4F2FX9tNWwpKr77LLkXNQEvc58YQZjPbuXEnD0tD8uK6dWc0CcBEJif4xMQXA
vTVyF/P/HQMOO6sdqcw7bxShfYIJN0Prtiy9CaX1Mt7CcGDDC70EUFXZTW0puGMm
v8weufPH776aSjeiNoH82UAjT8Id/axJaWmILfMvN8KZLCbiChPfFJK1n7OMH/PI
ZIZV9+TNFmOFgQzQVYV5XeHw1yT6qqbxxDpxhfkllnrpEA8cZ59v/10k5GO3m6Kt
a8loO91CyRb5+kme4Me7aVoYr4lRzKvJTUlu5/y37adpmL4ha3zUnp5dGNVwA7PK
T68b6a7AuoElcDHX5N9ifh+kxzZJ6HAyj+3MQCCk3gx7+s59+4KxqH5P3CK4V7H/
5FaEe7mZwwkyhNNEzORmLs/q/B1RrazKMl8z3lQf63u8E6cPVOWakifV45In4Uul
q+rTTkt+hgFt5yhVI1lDfrTdjOxijOM8uKtuWnUBI21xQrd9tOS1TarV62XqNBzg
e46Kn1e8npV5k5hFXkJgU38SKKrhGpq26ZxRWzbAl1VQ6ox0tjT1B0TgaED1lULB
Q+LHcAT45q9Zm0OVCE5YDx3hIp0XXIwW+v64CixeIWkjrRA7el46CXXIP3/VKtpv
6qABm9lcZ3mvbqzJTDqPZb8eWrXA+Q1gOpsnFC8aa0/l7FReKGUQIxzIpTg+00sU
60Xe722O5NSga/nQ/jSUcY93F7K+Id33RaIEG34uBjBX3rHX6o+PiiuS2qknNWH1
wLVWVtKltwbJr+iteearV/MJRcxW3NnT5p1Ufo0z4d8qlsDfjpeM3TRRfsoQTOVx
OrL/cNltYG6wQVnvwbrvWuXvoOjqF5TDVgGMYHPpTrfKW41jxAX6RpVWK9nDyWEk
gXqQUIkrVZHqGqYmP2C8YhoKWuH+asrgKTZjrDypIbWSazIky3Jb2mFao4L1Hiac
l8cEBHr9KKg7jax2xhdgPoTJvA1Au9Jq8GwZRX4FSNiionQt2+YNuBau6QJLKeRO
ctyLsPlAr3ARiC9hEClvn9B9jCygJ1tNKORXWoKFCLSxFBJ7s+JyjQAmj8Afst/4
1fGpWeSPOsC3V7QoEhrtJkxaIqcVOg988yQ+m5wrawSLhT7Fq7//Regty6M2RWRK
dP3+5r6/A7ROSWJ3kocertWe8h8Nh+AHAx/3UkDSvBVaY8PeM1wak1hEu2Q0kye1
YryVvoLGUkGN1wLbNU/iGUH5QKF6prIgVmUBdQR729F7AdvNaD6ShEbe5OL5MPRN
NZgWAv885/WJShbnKysZuJ2oG+g4ROgXQeVGaLgGFTEgJcJQ0XbUaThtJTjrxmWw
4mA9BCfBNj+VjFbG8yToNrdQQOxcJ5FYwxyjMJxEZ77YpGXvDCfzE6iqmckwEG+x
a5ISLRQhK9lIl6Iy+kHV0m4fe4jyEZzZoREBRMPJUwmS6mzDkOUaEmy5V9pcZj/6
B5Ft2v8YSRTilIFIYU6EInE1H7oQE20ysYKZBCOlL9lrDdTL4oWhcittZmJn1rid
3Wjxngnu8lJNKUrsaGVLpDizJva4H7qeSLwW0t/UTNfrjaWbH/m3TCbrOxxMGpOv
ViuDe0vCz3yprqTjQ1PU7RfxzqogT+GD2zwmJu1jkXRoJT5n44AAErmPR4k3uq+R
FBWkPNTYNUvQIFCMgVtJmVA4GeDoqmSn9CCoV/aRs32oH1oHrMVnw2/eu1XrP42S
9ycA/RgNOKfYFBnz/JgU2M5hJa3B6qzxCfzqfi7oXSylblDOmcaDWHclnW64NVJs
1VFnPTOzfqfZe0SRKB42jQ8jEXsM+lLMMZ1ayX/eveHNA4OgzDFgH4XhJLUrlmjD
RevkttzHXaAwD+D12Kxz2EAQqeB3NfCnsWG+RJUXYK+XHSdTIXm5HLtC2a8VtEez
tfaeLZMU4qgGw8zgZDRmBQEimGiOU3MwWy1CVJCn/RD13jpYjF+F7MLoGJ/K3IXG
GADxi1EdZ+wdPlMNRaXqZOVT7i5fjSa/ovbViA448GG2u3Kx8TrD++Rz7bQF8lmI
G3RUz9zeALNpfUKVBfTKin+iS/HRxZB11iXGlXRWGQm2XaYB/UV5pJ9nww5BX3tm
zysH2ZCWlh6baYoqr7tvDxkcIlqdg5p/KRKphz2Gv3IGfqNYHw9k9Dpw/TGToqlT
PIeW6sCGy7FTFsEOxaNNH27Yzt5wwhwgeDJav6X5WURjNbZkaWxOvhx/Em+/OcqV
K7XlqUFIVsC6pMqeV8ilzj0xBmicF2WwvF4aEhVH2qVqpxgzgUX/a+EtrDg55lKf
lNeIMCPpzbJg1RT1jq3a1xQC313auLqrWTI+r970n50eXa5E8mkDErjJtteBmM1q
k0rqhQIwK7Shgp+4QiW1CjhydfL4MLIW6/xMpvxeklp9P2yuoUcW1i/r/1JLvHng
BErvs0etKntaeWysoZ5SxWg5jByENq7EwXybkKPve8LAkEYmBqrN6AUSxP4O4Sc9
Er6FKB0W4ZrfEyEGnT0lBp/hz3w6CIBO8nFJJURDkFCfIDIIwFTNHrQZrISwrstm
tm5EaTlJQJJAqJ4mqf09/5FGWilXiXafIrqrANXcHq+TdPdBgI/tgQVayDp5j+UW
cHxrXalGqVAisiWc/O+/zPezLkJgv9nmh+5D0ap+pOVM6DLynt8tZLAWNZ/TgHv8
WwD6zdPNIP0e2nqbe6oVEQIROWMS90k2voosZZXOLa6RE0yRqqbiW7Bl2jLWglJX
FgcqTmtk1ppVzutIxJqt/C1iWHwJF26Y/JJP/5OvITgQ69oggyBg95xIwy5j2IYz
EPln9fE1ETvz7rQcRPuzq8+BEMGo/NkMYKlseWJikzTKRIK5q/unzlyuguTvtxd/
pEZv2/fUIgyWoyI8JsytXO07LCLyHiOiIBSRRI4xtnTFdThXJZLq1IYv1A1vrdsW
A3leQaA3S6MM6bVI8U9tmpN8TkSzazY++JLn2xqpNHWI8EYEuJt3EDvPP/pFCSmK
h7AHEMtIA4viMJaHYkkGM+e076isdYNBNyp19pE/C37gbk9cTihdBN8+lTQFHeYX
8t9ugr+IARV4umVxa1ksYDfPF2suG04qhzHpbOFLqDsqFluFbM4lypy525qgVj21
PseV65zmEyxxfQx+YiIY4f2ZqC8amZdzjMuIYVzBYY41nyXmsqdEfzW3bup67xlF
WkMRYHcDSdSgXdEL0E3ZuoJWQjHtIVmHwEqCW8AMRjJA6M1E/QdQO+rjnyAailKU
5zLDT8jgL7CJyOcbk8ZNYuKvkwpG/Ma+I7SvCzkWTwqk4/akzOgae+M0Gg3aTykD
L6R7U12aXcFSb+mnELY4noo9J4xfQfJcjL8EZ7EgCyVpeZOnuz1yp8rqcIVi+8wU
TxQDFiItQsbyLVQ9NEBpXWubvyb5G02IxmfkuGlpTyZw1ex/26DXYDmAVzpkQxQz
Itm8i/VsWOybB2zTsHFdvHSOSQVyypJOdBT9CWlNmxCUHCM6Qfw9TdDVwZIpTA12
kQP0u7U9Nwwn89Q1/WVRuXj/CgrPBxhiDn4LSzyEnU7Ww0bR4E/vfS19HmLyBrZ1
MbhkPuHTKT+9ZVDSSH+4LKfcNLHuveWKN4iWvhXgH0JH7JSlhrZwJo+fG7/nqn0Y
NU2JHSJvkIj56IKNUP87bBf6acAk7nAzR8lrnbqcsP0MdEHdVI731Ghw0hS9oquI
4Qe2xzDhU3eOrUYpdgRKMLSUm4/yWxSWWLqoWfiXiAT7SB2cBhysI5LDuPk/6K4M
mDkWh+seC9qDMRfVqmlaiNqlAsWIOKFQi3Maw94Z9HTJ2orgoYlPC7YOQJ6OEpbq
Y1w0fAYz1pWtGB5HM1c2IpeImDTnQXa3TlGeuY7xH4xp9YnjHHfn+hpUWs1f4EQP
5p80nvwxinqsA8HPluhL2rblMjoZbCo4CcpjyonD7cNCxcrWWDlC+YhzJTBTDzn2
SP7gJdONNzj/eIml+eBz7ie9GE/E2sIWTU2I9Z10xdIICFFaQlIC82fOH1EU1Crj
Cee5dA6UVcfUDxOKlnkz28Imhm+4cr5/MhGJtkF7yRQs6iJjKJQiAwuKXbSYXxeo
gGSWaIRgl99dVrAlQbc4Nnns+rHZU4rBDi8XMfeqnMo0+dzDvs1+A8opaFSsLUjj
yIcmZffsJ/WKbPVjw6eLK0LeOjeuJAVEG/CTihg6Z/R/NhbQiGxUp7P+EaL1WA0R
5OjBnBMPPvyHxlfTxUokfaJkLEq+lK9CKyjw96CgkBKNCI3nmIDcpJ4rCjVC8lOE
fnIsASbhzRWHkmAFEj6QCxxA0lZaP8VbfumH/WZdmLisgWqeeFaN3nWaGa6WzVV9
Uzhub0nTgWTpVSxIq3KggyFAzLSiEGBdaTiocSEbFX/n5pcxO4ok6x9sjYqDDSQu
fLKQJJnOl1gWK+j13V0xGmqZ4DpW+57FjQnX/cD2PwWyRIZdIvU9QM9SA+e8c/bW
41QyzBNT1BOQ7ofFk5A6m+1eYKdgSnBV+0+0dTHiyh860QxN+xBlS0oJaDwoHmJ0
Tysb484guhhhH917KGBbXR2mmTZQSQlMnG/I9IdWzAimuhiZE/gbwDRafdm7gKSD
UOZvMwNttZKTJsitWFXNe38+b4YPbJfSWh5auIeZFBqqskwEsnrjnrVIU16ytJHS
nBzmH0nKFdAL0i8ieBbG4Ri9Qgj1f5RuFnVa1PyaeIGN99EF9/nGcGhLSe/0RlZd
ONg8YGbPp0VqLzmNwzBR8L2GiwDe5Lr4lNGOr+ZW21TjhhdeDJkSqd8cRc5au/SF
QAXlnagYw3OJ/u7RkNwuGMKkmnbYkap1tiH3wz643LeRMuuZKkJltySSJeApl+Uj
kbtB3XYrRofyyn4riepqCQMpi/VUuMkxgWMEoUX4y1NMRoetX3qBxJEYQayE9a0N
z/ZYao5Zx9ewB+AtqE3DMS1Loas9aKOFkoEwYrygOOVqwXNvDDzncf1YI90iTaQR
dHj5MBdM9dbHWPgfJou1ROdDXis9m3DVicbJCJWaE8Wwt473ymrgLwEX8zOu9igZ
BFmYScycqzp+fB5PHjc5xdlsw1siOrXPfVqwY//gXtNpv3atw0kb2TwqJ3KBQvGL
mF5JQZmfAbZhYdmDrcUundbxAKtQ72t+0H5VNMNTZmsTse+A2ztRRmeLyQXIoxud
bvT0ilCodQqfNq5sywIjzBZw7Fp6LkEeO6qoE4SaIYA/jPyrHsfLTZd7X9Gbj9Xn
TXdKydQXv1++70d1JGVXMSu7GrwLgw5D7zM4N0ICUeKEfsF05scwOeoU1LeNFYXQ
rXNmMKeOYJ9YVfewtMcW6wRHcPSLWZFLgLnuvzrUOOEoqL8DhyCJ6h3lNd5Q9tO6
UJ7dNTfhr4wXoCKsAVGfZ7RSMU6CqEzrtBolUkSNpiCC7cXEeF83lLEBIz1BBEg2
W+JWSq33IafBi6gFovaqp7Yi3EAmhPKKT3EbyjW5d7GQJA2M2KJJ1rys+Kbrh1Hc
P5O9cJyzodpmCno5G//ppnRfuj8YIczijSvDP8eXlVGHYLSA4sUOnglQyADUJIGY
pBtMxwut4LOv4FWV0UPmjDQQPYw75kPN+WVzi8MD1ueWWf4gTb7lzLQ4/26j07BK
Dx96oRlnL2RoZBTpLX6StX4/xWmF3ldQhPvce4I5pwYGE/i2nayuyrZZ57HJZuPx
3n6xK5NbyDD2iqb4hdkowsnUq4JexrtnnESZyIhHCBm5KY9uspMr3HeJ5nbmu0Zf
5XYzxmjPFmqVt1kaPSLIwGKz39/Gx6tRqBHHlf5Xx5yvVDGYtVJI9pKMwhKyul9d
u2MnUL0rvbJRlfqbAUx7DTqfmc6wBMLV/7hbwU9BPG3KhWIhbMs9D+IgohGdTpgS
qr9/P1QPQjAd7K0y2UgHgoSKLAO+yDbnqAYjxzoxtUEBuCp/pWNZiYRiml+R0mEB
B6FKqYLVyOUhuNUFH1D2IfBwzdnpsyjf3OTbXpF/z5muv7oovP/zLu5NXGq+51qs
ppMJSt9TGZ8uzKGt5FaY1QDeZ0rM+jeuIHu3glS+RaPkzUc5PtRyv1nPNqhWUkXD
DP0K+8Tu3DAhfLNSYPkHITkGdTl/9vj/8zDEeu3OMb9BhNut/RrE9cxoKP3vbc0z
TaEe67A5yF+DGtoRw0Idp7/mgUWL86CG7TIp2BDwC/cmZMPPhxBOZMYzSpNXrwdg
0yj+YxpL7Ef3NAe9VSzYgaghqBm/n6dZrhjexAjB08VCgvmb2hnOBQgeKqZRXUJR
+/YvskNVBk6YF6dYjn6IGqnlYjDNijASeESaDQ1ELByT/m7dIHTx+cVGUghLHOgE
/702ctQXF1/raJ4txwfh7KkQdVSy9daO2Ogz6rWWGDr7vq6b5zx+wYMQ8TqnaTRN
SQsHjnVMSIbctbcZjqv8vR5SKFrwUg3Kwend+HkqiJIZlguu2SkTH89fjklCwViw
HRDP/yvS7+/cEKT1sYbAzUJ/LIhItyYfKm1m5kAzNe+bDtBncdsia29jUrXroKiY
FdnkRl6jS2c8Qs4DLgiOaamDqfDBDpxVP2ft16+TfONS4ENYpo7xd382O4tTU4HV
DOA5/OuPCxDPGOOms9yovCUsWvwFkxCgsEL1K026M14+05UlTbWnjxqDNEpbuSvU
zWOIXwg4hFeyR96r/B3dSRrBoCStEGaOwtZz4ipNdXGau65MDdFvtlF8CW6Yslav
u2bJ4zzRi72RW7IyJduP0jJybUzYbuFtj4ZWUfUQ7IugVeOWhk8B/0Rkr/0Lgoqk
KJ7Vy3QI/9qHl1bjbs7KDEqfCDUxbw5m9C9gVDQONB9tJvem/YvpibeKCe/jbllk
E2vYpxCmQ4jD7UBbtiqtGl358oVM8H22Da/HmnKUR3bEuqkBansgtFcTdEyJ2tt0
rtB35k+BN2U4iZUqeo0EXkKBwS/l7zxkmZyxMz+ZmkFG6fogLYogvPOVZ3EJcqIG
EDrwn0sHtfXmgIhLYaIiuPJChWPnS6huPM81Mci70a0Agi3QP45yzx+cAbBYlHpK
mHdo/TH8TNx4mjVfWykksPLxnnswsdRObqOKm1srfIndlk0WRYM2c9013DQcr3EO
pWrloFsUrfb02VGSXbn7/M3l2IQXRaaEQYO26YX0WnINY+dKXemvm+JfKq0Sn3/m
yEP21JxAGaYUoVo/38Y27tej66+IOWlQ62dQ1CQjWNCpNetzBVI40kKlegi0aEjv
j6sxBjMkcafp7/ZZZh+7fpKyBQfc7qDKQGz+8OHbUahraaoJNF3mfly+hfvQvJGP
yy4E2pnc5AIG/uxb04O15WXiiOa0m7/9dKdGOn+qWJ4qRBSxcyc8aeibNQIv1WCP
OzUHkXsoHKAl5EiPgmfLJbEl/AC6015IAxMoLk6ea3uhANBAaiREau+KjUwBlBsO
Rp4ymyXpcCf6EuPgmBsR7tfGXRTn21Pw1MkN8U90lwSl2zDPgSDH5r53X4Mz1wGm
vwLAiQ2tuKUUK2xhEHgZDkoo5ojkttaGLdlAmo3AOdrHH/SObjADLAiITL78iRFV
VW5tnrNreIplG97JrpHFHiGL8d1wLX4mXkuc0h4xuq935y6uTN3/9dC8xs0WD3vR
L2vvVDPDLG4n8ZEM6RAf8kR0hirtGJZpsmk32WCqnnDBgeVbJJVdKSdGlbRAWzHP
f/qG7RMKTy6iU9eiFvKR5udVS50tcRe9peAmUlIdky9W5ecdY1sV9FEpVCD2I3KC
QpoVJwMhxeFar43CuJkvmFtWXvDE1F+iXecpyXM7roByoRmsgJZMObVe/YKxyRIf
WKulJCHWuSN+qVKuVKoUW+oxGikSA0JMQQ7IdFiigcHh203XYzhfWtKrFLiqZxpS
9oMvZZTcCyCDrkXqhvzyT7nXtWudx7i1t1Ez2PiriEUaa85x6h51wdNJBxpNszcA
y5Xu8/YB7RQZbMTZWFO9KwTMTdiMNOCNtbCW8HKavP4YH+bfPeLzzEUDjpil3tQQ
`protect END_PROTECTED
