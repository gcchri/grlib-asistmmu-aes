`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KA+97H1c4bjW9kXGpPdnBJrpjfhqkxzhovEphIZk0dmlKyl2JvzypeJ2++sazOP/
2RePZTGBrK2lJ6OgC6Uh3Sji4tbXTI4VZLfjJjzYxgRe6ASPB9K7jpAfd5dxjEzS
30H1fNjbFOExxTuVtBtvFaGDZOKk4zXEPulE5EhS5YwiXupunn1sTMy/S2on6KxA
K6a38nVyzOOjx+YBoQgVEx7WYQcDRPqe4SZHB6pCUgVdJ2iDymitJXKU1jzJ3tbY
wtkkLjzSecN8iQcE30pJqfTVZOaxz6IIjCmn/I5u7W0cKRmRQkjHRsy42cO8X4Nd
eO5xbyM/5QGKO9Bizn2CD5/o2qURLdyGRO2uy7R7Sn4og7HrCBKb8jvoGKbstpB5
t3uQ2Y+LXN8Y0CUlHMPnMw==
`protect END_PROTECTED
