`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IfedtPQIaXMPcnzl804/WnV6YyIsgf8UeZAJtQRHthZZT6266UkSkofI1w4h00yt
XUZRDEvbdBWexj2o3YGOsoIHWhmwgp+UMP6J6zQqvLly0SgQGNKmaZfs/23wphmO
t7/8jcZr53UFcrYVzvzDP6jPK5adPMJrc6U2EK4YuTtOVg66c0kADjVMqPTY7toB
ehC37lnhYo0bdfqyoTI0qybfP3nOd9SvEO0pqDo9r+Zq2DByI9tmaPTOX9zzWp3N
UGJDTmarcWDghG/H+1yn/d6QGhLAoyJpqRzV+9hrRQPU2SfX4yONtYzX0L43fthJ
jktM4bULV9qs63psvNVSwn+0URSBeFb0h5xNMcaZvQR6RXHztyDs1N8vT7hECoV/
5P0l45WlsQPsovHlGGDWb7zUDtDFvyvfoXgb7NxCBM24oko+0EMmgRgYcfP/RyRA
wlkDmVJ1+qL5Prczi+g8r+sWvtJq/eSzsIoXNTUZo5d1Bl3a0ZyEiatsx/CqBxxH
QtbsYh+n93M/uHgCz2eypQdrQ5FKquaOjG0VW1J06i/jQsl4Lk0b7cWPMyzEmluh
FKPPii1t6/gc9AQPlA/eNcBLt2ijYahZd+Nd7PiAQ+GEMi//GseSBic7N7XZelcn
N2t4/uCepCXMz0fYDwQ8Qml8OLhAb0C5jJh0pTgJHUc=
`protect END_PROTECTED
