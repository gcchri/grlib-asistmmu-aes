`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PPCqbDw0ozI5JAtTmYr3b5OjvyoX8A2Z9we1wt5+CgvjXJ3r/Jc2MZAPbQM5pljM
8Lcb014XwZgjwQoovBBW7dsdXveap8ebowI5FUpnYFndtcEO9D54GoJ01BGJ1vX4
WZHrcW10OAlIYCR8yPZGdIy55MAYKRKzEyZr5J6y3kR0NLop7lOcM+Fw8nuEM2vC
W2REsH7NhzLTut8CsBKEoGIjgrpACKzD8jdWJcGJTSwWJPNNXQV3iOvyqlK25eJz
MFm46QXKhtOj2F1vm1LEt3zgxraMdvOBy0BTZcgzgVAQSUFkSfT3iWZ3o8cPbqAI
Ih0YbxMELn0CrrOvOPNTKCwPDRBA+UHAwDRhkBMV4DCsqMkXN3U7Ak7SlfzCFoR2
psX+lUDgwGsZY0gqya0D8HPb68Jd+JMPbaISX9whne7e/jahSUcg7uOugz9v+QHJ
AWPufU/odrGgjb62A6e0MVQLe0fPlB2/TqlrkpwX+44=
`protect END_PROTECTED
