`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ORwQxtlMzJOBmYBqGKwdj+PyFQR6dt0+qkZ80ti5J0FOyI7D6v3F10+Vn8olYKme
D9ENQvvgu5cWhLm/cjpc58K9KTog9yOF8tCu93wFnYnEtgaytIMInIdWQFy42vh/
XUoGNsbyMR4ded+ju0FGW7bHP8/ADefFs9gCak6i1g3c6v9iik86YZSpKBIS1S/6
VI7ybRv+0bnozkh+Q5qU6qXVSSJN7P5BZ/GbnhpFSGYFnUWp0VqDyfsGYkQbC03X
J2WelDFIHhoZOCejZaCMd8RpXcSknVx3F1udEDFXdQF9Mh7mkfOWE0pZQ7kZrtxL
Xy/ozflAWanV0WMSIZULYCaO5AqV/XFxz86XUwJogp6qfrXedXJ/25Q3KTO/PtTH
`protect END_PROTECTED
