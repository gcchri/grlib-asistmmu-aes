`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OYURacOSkMrlPo1cSQiSUHcB/eoIXh0kj8EIncGJF/4nATaV7cpELuVZrxj56g77
do4owsezLyvKIJIdviI2CyoFHKQAjhFFSU9/YnYzboUvPr2cROazB0XxAoZUDe4Q
DZNs27MmSJ7cStWYaJqfMgEwNF+e3omE5iTHvFZ1qHSCPniqJQlh66mWhYvRPdPb
YN8KSdFuddi5sHn1HTdaRdlCzF57mjK0aP8906TiseDG7K7Soq2THauKpc4uQNPi
36f6e3A941mgLuA2Hx4osb/DjHMOGMzk1IFOTNQmeeA3ZcWROq2hemtWlUM04es+
jjGHFLvA+oxfKBn985Q3jhiVEfppxutF1PEBNTZyCb/9rrK5EdyExejoreSkSgGn
6EYY8Re9+MbDgD0lBh4dP7K/xr/V8y1HO2HWKiYzrhsagUMq/WjM9tBn2w0TOkXM
Wbo5+xKxTv3IYvx22xdAewBC01iRXDRQjNVE7PN0Bn+eFalqFjA9Fi6sXbOWEP7E
xt+WcK6J8srldVTfc6xBaMAfrmu97VdbM+m3iUTYqiT7srIlpYdFIgc5z75yyMak
`protect END_PROTECTED
