`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+7qqvgjWehLmO803iciz3A0rLYshPQiCnTH93VFvzZZdiHTFMdB9nq3FTkiIYtVS
fw+fg+QBVYXxQjk1HI6xylvhprJ1CXWPWpC4WY9x+uUrlCGOFRaOgtMTsuQ/qEDH
aL3Lmz7vZj/EFhvQYOxkr8ML70J22Gakv3cv9WLfHU93wCw1ahb0OmpywEQmVJbQ
icC70FKHzwAeKr0/PH0S+7SRieFg++uQsWcuFV+kSsZn7kXyJFlao4vS0h+CeBWb
vEjsFipXrzwRWP46k/vHvQ==
`protect END_PROTECTED
