`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fSrkps0KsYKIw6QBJ1mMLHA5Pw2uXpCX3mUv2t2i6dnUbYCZN6ieBr5Z1U3wYNLL
meV2/KlYSqbks1EEzkhN/0d41rExrSikuoxV/bIy9ecMmgnTBKeYkmsjBPEPLUcH
7YhPcz8T61rckKw6QMQekaNHKfhg7HgcibRrmtJJJ4C9gVFRLgb8mQgWgYKsNcZe
BRwlmytOsB0FEYV2gzjS5kzsTtsA/rQ81ZDuej3G1iJT6h3EziQAdEQ/uVLHtY4n
wJP2BNmK2aBwpQi6H1EXPyjjaPui8bHG6VP1/1DDcULwL126uZ4IE0fP5qdbMcyo
lnK9pyAkkT4AX5PZakSZ8jE5tZXQF2pgDOjN2+6YYTvHrv34jHpaTHB99IrGbyu0
Y19LL9/7oRLGlmRDYkHzBznF4sGvklb86Tb5llyl5onQo8yaOE5uSpi7A+tFi+kz
6KKQRT8Ie6Bm5LOfwk3aN8Og9mZ7nH4N635552B35lmTlXt/JA/SNIvHLjyF7cCI
zySy/uUEjXdIew4CzvCLu6Junf3IiwNF4a+yoflq99ubCT0RNR1RfO29uk8BO9Kf
a/WRRwnjrVmqzT8VYsW+4gUP0AkWb0ZxSQvBQeBZloV8X9mr1GJ6q6Gt/t8WV+X7
Q1tErf793/rfbBNxLhFP4lgsi7JGaALl0MgJJK4o57ubMq9KYTuydGZFDbwa5fES
O8AEvKWfBaOL9zur2bR1c96UD/b89pFL8w4xMzBVtIxQO3SqbDE6UqwjtzidCCC5
+AOMfOF7iE/D4jHVs18ZTsrvOKisVOCt1I0UiU/cvDeSst65lX+5zBtjO+ce7vqt
xXHMLIi7e6TnmpMooumOvoKGxCLMob+TSQewGnLAn7n0iZA7h2SC2ES/yga30qn0
zLLEW9NthB6sdtEHx7h/orsjxLfnx3a7oHXSfR6Hq9rbn+ynRqIRLiArgCCilvMw
ye4Ab7rv8at1aPA29wcHpijI72TZMiI8j4cD2WYs9X4KQfAUwynSZF83fJAoY0L8
LMxPMO3yVVzl6tQ0CZy6oblk9+I7AKOb9wjC7pwkz2DMlMes2/WPdWSGN1TZ+hgp
eignW6mbMwOx9+vQRsP5RqCxx5A3i7R8TJxfzhmfNd8ts1r1xiWOLQ+uiBXTJFN8
uW3V2bL/v9UCgkCDIqS0Zh4w/xZka2+3C3aQbu2BltIwFKa54jhH5nnV3fCV/7Uv
3b0z6JJsHHjHJQbd4NRBGIbbZMxfN/nNjZXofPmGwmz96N0jNu0FVc/R9vVuaocN
aRvkotoJH6OkgpKtvdOSkNOQ/KCLAzHgyTBVWBlwvDTHkRr3Pp+SWw+ocDZsjUbe
DzQS3nLE9vsic3phFgZr0hWrPF9IFq9JHKFO94iLgNx3jkM3eaX79u5g5T2FUFQ1
s0pmmDXQXwquqeUKrjcUNLWElSTbPrENVIrv/FiWmXf80kdC92Zmjsb0n/ypblJB
sY4YwufYt1MnsV5Ko5FrdOAzPcGFg9nHWh3GIlXA23bL6ohm3lG9/ha2gVanY8GX
VQJxxU8eVImw6RwDnWyuvktV2RFE8I1alH/mBZLCTu11s6BgQhNaU2g1tYKddDRx
nnpn6KYRsu39nS7W5NRztC2zfrCDhxT0jd2xD0SU3SJcc9puyd/gd133VQQSWdMM
LU48h1CWB0HdYIQ3+GJN9KSbuD31LXHTIGaSjXiBJl+71a2BigLOJ8t+SDstF92t
SX8ohnfjNgB7Jh1t94q2rke9WgPmrAgg/8orXYPvX6zacSEHwfvVM7VSkV6bjDyx
mJwU1o2oXKP7EEgD2YCuVp5NZHCT3AM07jT+e+pNtI0DjG+p+lsMGaA1dhi7cUTL
o6fwaUoaiXWtxYxzpateAtBN0cuMsd9PmSdgpcTk887rMkfH1sPUgm59PsOmA8bN
PHnRwK01oWAEuwBf/6a5CyPqIgej9oT4abSzbaej10aBPtRRWwv3DXmuj/dMbhFt
SVFXCcoQnrdlbULZd+i8zB6C1AU3FvkZLk8W7uZ6pquqb88kx1qjyr8/wlkWcPY9
Y9eup9sThC9BDfyaL32h9+hTlhetg/HdtU1S+TVs3V1b9pedYjmdZGzvsIwkv3ki
RicsxMHRM0CU8HsjC41N0nvTgoM2arzR8dmUJ8F/LKUtYJ3rG8c4mMTApcRQyA43
Mk6YrARNJXcAvQ46AOxhTzVC3jo6lGPvAvTIJ1K8j6P7GkjiuH9yKL1Mc0ZAWssi
rr05o6JL+7M8sZwzaHYVPo29xo4T6dJBv4AmMYPUTat/s+o/Q5D0FqJcaNfvqCSe
/yPeFLvMfh8va830lU0pzZKg31HDQfqQzDHW6FXOMNENp9emm6wOJFHfPHBRdFLI
7PZo2DxJAlBmofBh2HmoCVmQEl0BfLCoYncxdXyKI/LOGymuKDmIGVXSRJowRYRj
RxRViLKqIZIu8rCPIEZtshxrxdjSrubRavBvdgtu3XohJVKd9HZamsOuTpg71dll
Reg7DdWfn+5siCcdzeDoYNqKWvJ4IS52lzeoUGP7HoQchaDTHofsZgs6HcqIhvLR
TE+w4AifwZpWBuNJM9FxxrCPqqxvRNn76UWFvg3oFPTfTDpSorR7Vy5GIVEKfdBf
OBE7RvyyNFq7jhAqgdvFA6EwpwaViZudHJ7ePfmuh8PJ4wYV+93ow1h0gB2e4B64
C4W9AwMgcA1JtWmSwrIuihNB0+JYRAdWDhARHbZRE47A22liptGym6pE5q+L4H4S
Vxv3MQ/SJZ7HTLmCNpsQReAVexNtAdv+qMscbRVkMJ7iv2MRkK/p3KQBjGV5PWqY
GeSCo177QLQ6FA0TyYFAQNWE7W7Edheq8r/XsOcDklX2pe+7t/UHrcp/AvbbD22k
XriDD9T/Ix+KSpJ8tRfyVQE/XKXecuGVlyGGusYMWx0uazTjtjBBpCu/Ucpi2/9E
VJR+gADt6G60y/ditdHRXwYitnNVHBfX6KZkDRR+Re/V00AV+tMb2eZIoE+GRNE1
Gu+fDbb7mDs7HThXZqP/T3CralJHquYHMjUtjhIdR4gs9ijU+GxQa8pdBUS6iUTJ
PeEfwbIAPFNvMgcgkoMI8mmklYCqOqE/pShrzvCrgusWgHkRRSPQjrPLuvkrvSwr
UW53Uh0ZKsn42bNo4Z+oD1H+0bhklzLT6ldQCHO94srs0SFn/jJjMaIYwMRq+Z7e
VkSgEV7fLYzPVxcrHa6hTnuhyvDlq0e7c+shtwBbnvsbtMqR+WlBJfNE2m8n4lMJ
3xC3n/8eDiRkILemBf26wQ==
`protect END_PROTECTED
