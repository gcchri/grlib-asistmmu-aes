`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TSf/we70NSC3jZImGPi7oonfJW5q3xeTeCeKxp+2vmtZ1fM1OKbXSgStm3lDpjxj
E72aNhJ6toy81urcmugiUIadC9KzpRlWROYNVYbtXd7yWn7PXnUndlapwR8CqQWD
yg4pHIxP03QPTW5SJqYgKKUAIppYK9otr400iM/suLTUUavAri2rPiqo3hnCLsqI
NrdDT+vnFwfK/Q/6i6KVk+kdtcgpUzOtQzH0+ZtFVCCfXB6VdKDRnKdrXMiMj4yn
vW44RqafndsdE40+d2iR0D1xLvEws8VVU4kMlVQ0beiYQhBjpkc9Gows9ukvpggG
oXZk5qV04KISoeSfniCRNRTVHhv1j3TVK8X/HOreQwCjOGiGeghFcBD0hWsGZ5br
1BHZqRlNE9X3E2fbdgPWZt+m7G5zYTj7XuHi1McWHpY=
`protect END_PROTECTED
