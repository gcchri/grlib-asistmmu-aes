`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8XsDcStHc0WYvlkU6IkTEN4szz+RnT8g6plnjGVkAD6FqcUs3gcOHFqPsyiJ7KrU
L1JbVWCdCRX5USpRGTtTBjXGS/+8pIISViOfrbx5yzJAi8fMUVpv9g9GVHE3e4df
o6X4AdHm4w1Cm5vQqejon0CkreJgoNUstnxihSp/lgfuVc9nruRM0rKrfD5Tl9OR
RAAoB4xb7+Lat8DWzDc9o5C60KZ3gKofmsvV1Sslb4igJYfHFUXfIymQYSmb3Jsh
HqqI66WHq7ohpS1jD3dZjv51Z44STBwG/QE85xH7Mzxwx1C1XazLJRp+NZRP5yei
X7m9ZuowACDpzn9MoC/ZVniqvtScxqnTAiaTlS/KwbaADz6B0SmAqFDOlZl55/LR
Xb2dEkxsNoSZY3QzwCYilTEJ7//MdmNf8oAApCvK4OxNs0QH93Q0B0hqxrnCQfd/
Zf24w4/yuEjpIA3+Kct9vXqzXRCnpggRoIf7D8T/fp/xNpXWx/gL1RstxXKtYa73
`protect END_PROTECTED
