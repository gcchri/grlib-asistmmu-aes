`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m9Wh4BPSlgvurLdMybSwQnisymmCw31WCDF63sAIPQ3KfNY1mgoUCjKwckhySXCv
SaAC76OPsw2AD0N993NzTpCsEwULwfIwFwxcieZp3Z3e3Uea3w0YR3SYrf6NKAWk
W8bIOjTm3CoiL+/Wb3qcgbhQPXY3cDP9xIkqz0CgWeqJ+gfNEpEZteDsVEkTxt0Z
s2OSBGAi3s7LOQvmVLP875/Yg9AdMi8bB6rdUmPBkNEg/lB6qYmSe57lE21WZ0eY
PRTXJTumxMz/dcvCawC25C2di42hzQ34Hzu3N1iQNUdpf7c+N8D7OdC+OLLaeV1z
SvnFftyq7z2C1urcaU7e3kt+Fvz2+HE7rJv80TJvlqJFw8yegiBAKkRtu3RD8No8
bSyFFIAueRZ1/p0gcRJyPP6J9K19LAYbmFyJJF2EBOkc+9NqkmjkdBtqrhLJ53sJ
IrpVrmORdpFAOCss7iZO6HxtvqpjdCB5YHz8AmP4+3dqwq8RGy4ZfVUzhGsYqTuB
yQTFU5GK4Hs+TFimgyz3CX1TW1mQfLbgO7IcrUcPJTmW0sUHTV4Cxrtp6sYF+CcY
KyNKtzoGCeVbl5cg52pEtRHw47P7+dliTghSyt+UUeszhtQivW8vGq7Cj6cxTJLc
4wswJKG/eU+8Kqoa52p5A2LqblLZQzh0lXHEqMqH+VMgICXASBFsFYTmoZeBNArB
yfhsqO8lmVMDcDN7Qajd0Hha+mufBOrDcEKPtfx9ah1G1Y5QNd7koXIwRfxCymX6
v6xzwlG26sHXOPiLBcpfmLqtnGtykOI6HPj4gYR56CSAzX9k9qbYHBOGEihSd4iD
LFe2BE6mti5HZNb+KZiarop6ZT6iUmgW9umtGxmCKVUusB5iyhg41LwceyUEdrZC
9YXT8YQd3VWOjwozJhA/d/8J81caeljf0/laT+EzVEjWGeaYHyri0B58mh77aiHo
WqvFjW/PSncAMRGRAt8vSQjQM9nZAZ+UWJS2Muubq+Zw0mRnmwVwE3UMtSm/Sk1j
luf//QB14ghC9pPenwuF3ihzPz7er3v4J+cWu2VaZ1+HLNWsEjhaKrteAztARA5o
1nBJDh22i0BkTifOUybKgxmVYPseCYhg+QLDANqwZ+hhPKEmrijD2UK+nhGkdvEw
aVaVTck6t1ZSwqIcejroXpIxkluSZttEib55d0IvE7lCJvqKC0XNlhtAXMXOGZoK
CNhTptikjRGxeM9FbVreHt3bnhT7ul++ghOB+MLLaiA7/66o4m5W4YF7rMC4yd5t
tSnZ7j7c1kvUuITWuwq0m60H0MARDDJHQY1pc+GsIU9tE2s9i5VrbnHpNRmvUoIg
GZYiLjTJA77b5Eam6otZ27RRS7fcGFyD2VoCjjM3+VyhbervrhR/U60C7at0BnM/
WlOWl7BUqjgDxXi11dbMohrvRq/YpkZE6LBgL1HyZvsFNoLtgzVX7eviEDqvszFF
PtUyE24saoZpybq77V9wRQ/5nI1k7lGkBSbxR/oJ/R08FNe1ibRLYKwJu+fbnEj7
tw/dg83NGV/U23TdbTBB772qNi8ag4RlXf6fi1tqrAdijW3UZKXftwXVTt3+Kjfj
`protect END_PROTECTED
