`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WwvC98HVhsLa1+h0zdnrVB9pr/crKBqHeq7WPhTLnSV+5eC5JJTvBzfCgd4s8bUA
L+02t1k/RROmIs+i64ja2Qh4fDnp1Y4hmGaB6Uy9tK6Qtl2HuZKa8oievpffkXHN
g/eeEtksusOghsA+1RCkB9bm8DUsQmjexlHmy7kblRNJ5TpbiZ7l8mR1HOVtYEmA
amTXu/DiFFcJHwFsjn1y9qSUH7/QqosgnVtXV5CRqetHYfIv4fK3HXYfrC2v6ksV
pbHh68Z30s2xw7PRjvAwc4U9C6DATw9v34QM0GQpcKcM/scUaGKEMHHNp7PWNkm6
bGx2ASTXHHc5f8Jsxn7+TbRO7Tr3edaUjLrLTfMv67eVPjtAny2g1o7IT2VTP+z3
jmJLiFCSLPha7BKNA0K1jOh2zauq3PC/+ANBiF5AS7F5EM84t2BFBbiL5ZQyMzk2
p33Na8W/+E45maq9Gqb7j/kXrevS4BbyqXOgD6Huu3pmkLjjsB9c4eKA095sVg8n
3D4IkQaSUjnb+RojXmNvLsS2x/M64EHKc2RhlMHYA7AXBtPTRRIm7k/7oc9NYxWx
F1siE6m+lR7VlUb6+xL2yj/lceThaEyCy0MoJ7ZZHxH6CDaVMl/SK571gi8w7nh/
WqW8TvBv3ZFBpdmWtb7UD8wgx4y1pBaZSFcZLBE19YIjMXXMcO24mkJ7tyei9HGq
Q4ck52dxKFZUHpsPcqN4314XBlIArOmP/qi31198IhmT9X9peKhorM5MNLm8657O
hj2jtByyUdMD9EsJS2hFRDAp6EX27mrwVlUvb38Rm5Nup46KM3T5e8kI6JUo5aq+
BG2ISnPIBOq4ntK4WP0VzMxV3tAsHJ4VJv/YRFxkKHEkM8sY9tcOcMCkw7SbRtLA
QHj99eEPOiFoBjNk74F96HEKBfq1RkpyzEJLG2bFuqD9pYVm3DaPTXfeHqaoa3fo
U9lNOvE6z+QHcdd53gOAtK5RiapSSEE0PZIpUm+Hygcvao/Vn7ahs0hPT7BbztTi
RDTtOA8UN2LhXgnCqjB3WV+4A1VrR7u8NREZnZYitYIp7rD4exC4zTb6Yc/4Y1YV
9TVId+Jk8izhCEVtPEardgHDOJHaHWc+zDEUUD0TyQcvrLT0lfTKHYuJUHFgPymR
pShH9VZgTBGve3hjnwF8tVo4SqiSOYU9iYNLb2+/qcmNI0+YBmD6eILbBTs1BhjX
59YGQAWq0QHXo9AaW2TcHgPJnELE1nykTXFclLNI96fCVZnU3nLcMUguZ9BVmcbC
czdup0lAisTAyqdIgtMNROTmLKI0bfx1K52P9ekMOgIkzdPPWxx2hewg/XqF+iHe
z+tec2bcki5+9lgnu0uFSqim/ZQRW5VO8mPaA/9LLJkMDxCJQO73UxQt7JGkqwc2
rPAmpckROzJnEJ3RAgjyeQjF2EsiPYiommnscMA/fTleDURRr6HbaGM9Ybmkfc1N
MvceaKHIAnOM3lUXFBhuXdvbVTUDXRVwjyStb8Q848hna4Vz472bXhNLNU28Onlx
41Xjb00GZ+qy+BUXfF5sT6pByeaEzdTQe2zpx/ARWJeYiciMpvrSppXyf3OqzCye
GyHGcSix+L52HyarBg3KbQ8AQkBT/tFBoMGTyt+DZzqgeD6WrPlhtqoEJIlyMj1Z
yOCuANq2IautE0vp/JzuyUPcXG4+FIJugbdkesNsERE=
`protect END_PROTECTED
