`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s0wK2ak5yWnpZMFgfl1IiZAJQ6wEQuqt/+ZS1w/bD/y1UQYJ3/BXWzXZ/6MOfzUw
7C8bjd9iSduNLg0FaWa9D9fQfQ6nytX8t6MHxpE/52hiT1N/lIVlKV5E4p/fmD2m
oDz+jNB1BEnmRktC3O5bPDWozivaAoq+J2LC+Qp0mmggM64TcZ/ZKVRDQ1dDBrF2
1vJI+RRaF5gCxg9dQrUdN8ijGT1iw37VXNnbxiblYWFMasPx1PVedZWcAap0FF35
8a03rnMifQQ7VSl9J1s0o1+T/p2BneEUvyBAACNBCPS0dC73nzwuNxiM7EK9Oj82
N8OBBSppYIjC/NxQfJmEiQ4BdO5X0V+IQkfh7+vWs0/ZKOrlu1Mp659qV/6BiBl8
jRgzYdcyQy+KCvZMfsRPnwPe6tJYH4OkC00USxYlpevOC187w2X8dynoHKG8M0OS
5F8gTRt/AGgVc2b0hwONuAJt1cmKhxDG6jk5qAZ4NLwf9qFWD5G6GtfzJ3t+4N/v
upnr5WqW+JZ+JMH6JTk2PjtY7qQjD5hg5Kwa5XiecqbVdKYk8fweMfHCvJwsIgbj
2VCA9Y9sH/ZvK+wN5p3ty7gyYMG/A5B0yKiJo0dRI8s0pK4PuiSBgfdK1iWeI5Ek
wzkhoAwBgXcKsB6p3rod7zYNCbqdd/aQs5brVCk9+UJwDLRP8wxIqZXcIdNmpaZL
rLTga4kuDiWQRAgLX0/yyuIQ32bgcJgDb2ioskIrA2b0hcDf4Tt1HXLBsD9tZ/pH
cAANERPFKAjO1ZYALpHK8LXFk/LSL5Q+zzJPQTuYIaHaN59xIMXrabjP8+Py1ae5
j6s4MgEZr+cu4ceWzQHfmGKVKBf/YVdIvTwJD5y00xjLZft0DjiQFTsuoUieT5Bg
HNmoqTBStS2q11M3cIWTrYXyJJpzRe0M2Wp0nkI28BlQH/4NVBrOq0AnAbSkEmUr
9Mwdgv9ak5IjAh8C6LhyPXlG2B0s8fiRw2PfVAvSPGSajb4s1G5/HxSYZ/NWx2CJ
tpLaiPtWsbs7owsyjTEPYY211Hh/aNOr8b9RXjMRhlm9LwSnItz/vLPGayZyDEkm
fkfqvovDlnEsGLXoS/n6mltiRC3tzEKC4BtcJbXYgt8sVTmJCEn8OlLcdvWTrkhb
sqXOSS/TmcrHZ98/hGe4Mg==
`protect END_PROTECTED
