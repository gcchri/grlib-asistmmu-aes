`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fBpfdTfi/Rj/BlQmvczCZVgz8cm6EI+FFbbyi4ffDiNbV0XelVRATsL5qApBEdxq
M7rK8fUBgX6HNxVfZPmTcOqwHBPJZiTmAdRdd+kbkP8N8vHDxuETz1fZXw7uxYqs
WOzTQTV7Oo6p7LfbhaQnXqZx7q+65ISHVNjDcnlSDMWmgwUhjfhFwss1uD5Z8pIp
50yucAS8yDMmwxyOjSoQ4Tb+1KrVFV9hp8Rs0Ol3ZnHRw+f/wID1kz4mNjcDBzY7
gHHJ+mfnQrgzLnNA2G55VIqVBJ6XIL1yC/3Gf63gCpFdm2Wi2VU1z/ncuLOT56lA
ISm3fpax9GcRlxGd4iUbh1nnyvh9NozAf1LqPzkPX+HivgfL+RVKXq0ST82iLo6T
SNZi3nLxTyaJdYU6NC+GhpVB6N/XS7kGrfD6+EyxHADgmcHBK07xKrkAJMEq/4Z9
iVpjniriuVRo5HAKe0OIFcTV5/8hz4/e6ht2oO+ttgvWvHwkTHSr0Gqmua6VkLM9
amMs7NAVtgRq6yA/fQm9Cw==
`protect END_PROTECTED
