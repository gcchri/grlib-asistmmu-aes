`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sobb3EGnrXptpmhOBqS9TuBiSKm0JUJ5pni16sLMXqBEIFzKCHj/NydZOBzzWeRN
Unlp01vstIzV1UMbaMqVq/D9uiJMHpSp2g8ThdEt4k96AB6ZGH6brX34DuFKWxF+
T33iLyHWNuwCeeARfNgK/0GLMkFZYhoiYLrhA4lpzbzZ++1v6l8VSNZmkHI90ff8
RcG2r78GTGu3KvfsgeM09BlGoOoFFRrOYaqxThbOFCwBnw0Dy6eULuAxBiKTuyFg
3ns13CtHrQZVqrSSpWxmd+rUDtgF5A3jdMw/MK7hm6i9v1YIHsnoe71w2dbfpq/k
CDcWBXy85lZvRy6/Lqb9XA==
`protect END_PROTECTED
