`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rm+eXAAG2ZbYh12z10We9calDjK+Uptyy6iurTJoSnZ6n3AbhZQLCx9I12SCQcCh
wbXKpn1NChrvmmaBNGxtKqHPfL+hKG7E69+xAwYF3ObkIQJlFTx4VSJjd2mGFlQ3
uznIQViVKV736Ce5SU+jqaESZgZ82YSD4Gd3fpH6hZCDO2zG2lk8Q5fjevLENzK8
rOWwoKZwUNs4hmKlxznYnw7x8Re+xruI//gHNZ+lAuKYe3NnCWjGOmgLZ0hUFIJA
A4VfYu4ekjDSL10jR0mQd1l+9+5x9R09GM5wyf50JV3FoxQ1tfUfjYlNtVx4O14G
2szkoxIxmWUJxK+GBxQl2PwJDcrzt9adMdewBbqQtOqlZ21llU52j3NnfiiwuY1a
x/zRKYr8AB61XvVpyIZgBhx47sZqFv/gP1aKL5yPErRvGWEBz8fOk+10n+QmE0WQ
i/AkBHq9BfTLvF8n4SOKTVDy0/vwiIZncaMJUnUxhnc+GN4zd1WdTl1jVjsudiLh
7D2xtXExlSM+ht3LwnFD2xMn0hUvqGRmaZToy4I80j/efqxQ5I5ulUmho+3ng79u
xII6aUsjihAWoRsO2CHRP+Nnje84cS9APdOHKRzr5NiIrj1W+KpRU4sv/PygV7AK
skMDS/GeZRnYJdc9q+eJZf7JmAWF0G4gOmJIP0JqLNtfPkCYw+EbTlC9jBqTVVcU
zDD4dFln5MfIj809hPkSZzuextY+0ty/AbuV1n/1eploN/s+HlXUyUwdABI4Saru
dkGiOsOERmNdBKBY6t7LKSaZBmMVUvR54+pJIZ16lyQ=
`protect END_PROTECTED
