`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
im8rTlkOhRSJ7Vw+a6qg4eaYyyOWimAbT28R4cKFX8u+guoovwsP4GWnpNdIjUKo
aIWgFhmm9NY8KGCd8LepfnmouDcwRhLgodsdlPVSN/gzHGLSaQHG/F0A10xb4Pd/
1HD7ASg+KntvLh6p8yNQViJZTen+vGyKCzwPpTiRpIO3OYkZRASpT5MeQGmp1a8/
PD+lohDe1WKs+/kgIuGZMOetkQsp0yByCF/Tukc+euM1BOyxyu2T05UcATCG8uqh
jaiRiravFUdFrYBJ1CTTS4k6ejyI5HEb3R145G+4gtnhMAoF88bkfXrrrQjAP63T
ZxWSJ0H0K6QMJk8WY/mFUcTtLiviBx8P7yunj1Yy3jh0cYwEz5qLAOa0shXWT8bj
meIy2uPloG9ooHQsityfLGHoQUI3DsY3ed6W5LhSLcCNBpEq17Yu3o2loRPOKRXr
CreHNXxFAx2wDOcrTax7d7da8CJJM1VPrQFezDlQd0BU9Km0YTjcEnbkhjzAQ47A
SeJKet/Y1+2JDPhJi2LOOaBqV2QoxqOD/8fePU6Lh4TZ6IHZt0adh3R1eu8k8m1O
D5dML0s8Wc7ZnZ6L/O1hXg==
`protect END_PROTECTED
