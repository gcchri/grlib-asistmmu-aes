`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FFsSLfYQZn2gA/BqBlfNSj4xylSO6u7RzZKdXLQN8tZqfRmWNKzbMk4hAWX19U8r
cjsxVZQdc53BdFW1kF6x1gJHwvkU3Kjdy3L2hnZlKGpLZ5TdHL7NFf8ymi8/XT/D
4Y+gNj+QKh5WciOY124FWofLafUJCJaJunkLZt35Bo6FWhlnVloLWSNI6hk0rLXi
RditmlJzqILZS6xIgWLQnkY/rxJNeSd9AEOIT6b4RYHpKG0n5DaygrKVeh9r9Szf
kCK3qF1cK9vfiOJ3cYIxJ8mIsSlwUzh73rC2ziNRYMl3ctVzOK07rmP6Xoh1LAiM
uWDybgGK9yPLNZOn3aU0+PguIoe9+GmZ8ZhrS2yReEGeyrayBPXIzgq+cAFlMX/z
xCIJc7AwvuTOxH+QvfZPkg==
`protect END_PROTECTED
