`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JjQA0+4xXkvIIsGj60MNSS538fnFRR9V41JVCcVaq2qDhbEgw9XsZjbE2NDsmtnW
hW8iRPZv/c5oJ2AEOhnNeKB6Sirhpsq57JLeGpTpRAS92bL3CvGupMuPgkfyDIx5
9PR7ZACXnh9WaN+ZqxvFCopgjMcZ7UUD2X7pMZ/NetX33FO5KBfeHvLq/i4sY5wu
nWdZGVBTKM10VuC4tGv1Wxs1eQ6IxGrngsguJwIamQ7saZ+MVpxkrZiVRzi+v46S
rqdikA7RD3JeEyj7rgD6SRu5QOMwUGhxNEcORHpx6PxAtNdX6vBSTCHWaKeDq+48
5S70my3t2NCszumpckVKDB9ciBzM1ezLJ8n6xZM+E4Pf6eTerq5AwrzxCRtBnnfW
N7ISvLKh3QNUFLMawB2MxSEvELv/sMvlNgPoeeFO8FWHZWwY+tWc3ny9kueVl9lx
kHpFhXKXyodNHu4J4ht072zgc0GX2PQUuoHWuGBAoKsk8j4fEPnfDMRncUcL9nkj
vxlxcFinSrXNPQC9Q7zgEUI7l+Ira6m9eXMNQstVX8jXqppe2brXWsSHzKCNiNIP
9bBECe8zS8SDvCv/WqpLVWvlQzVUJXXsol0UL4qWlKNl8XipDyr8NNSx+G/xeNkQ
VU/49XD24UuYa4sqfoidxkZ3+JJvloCGUPAyKFGw1yXe0Co+nOyTCOgIj+CoLCZm
nyVD3RxEFuPMXDAUdxukY/MDyKVy0P6ky1j6XyAeCqO0/1qIDNw0iyMDH3HbIPbd
hcZVbd53pYMgIMnY8L08XslfJqeDwsFV4bjFa9BVkXvL00DClQJiXw2FZZcOV5U/
MMx0L0ro7ViAfDu6V4y765S3amJE74k/8TTXbzOodP34B8X0F7BiUDkQf1JY03sK
I6qRI7DEFgi1lQQZYLRyZrMuaaaNnjzAuzplrvtmeqMMAWvOtNfCXeXimYYGDHuQ
mfQClFN6V0KEmHS2pQMYTUaS3zdvHZWQhXwMLbKolHgr/3hzKl66uXPjgLo/mbYW
glpDoKGGPLwW80fZJBR72xKMj/Gab09avypHPhbAkGxPdLUbPgJCwUIs+r9RVq1u
GLKTFaRohopf2KV5zBylYCrGDFSX4TC1bRQpRZPibFVE3CdSpupbu793OhJjIBtj
751pdhzDg8xce7+GwgRliKmw8mzwK81bZPI7lzcv66Go+HYRCCLedf8j6s816cMG
qNBswbI12av3FxW+/IXgj1CQb9uABswg+1lL0hYjcIhMnz72XHzApCBkCo/EyYH0
tnc44PIBHuUuX5BZEg1sg/bTpvQVafpaMXCCtS1nZBtG0X4NDr6+4km8qiFfiKVr
Oogu06soNNxXqi2pLL5kDwZyc6sArYst16YsJ0YLimtl/XdPix22YVMaAlMA9q4e
JmmAB9XSYZfllSVz+HGyWFRqvIcSes4DDkEAz28qAv6sjZhYqdsysyfqO9KElYAf
DAjl0qD7Q1HR7HP6i+d0yuXjkLSYeuB+R1tPpQ4N2aS6d416c0ATAaDs+9trpgyM
Z/XTex4FG9z0UG+l6Lkj9I4AguJee7wu2YbLJkw0fdsTgKruV9UFW8SEcm5QZ5v1
7NcXSqtmvBARIqlwx9eUjYLgBLqmBjYRdcMGR8wMdDwH3e5iDljfctAxanGLJYbi
mvTzuBBAepIVukjjBS0dzd8pqutYQok4YwKkp7+u+B1vrtLH90O+rD5ueb0W60zv
uvz8LMpirs1sCZcdLyyEk1WPKcEH6NFTYWipSERjSOxH6DAmPUA5K4K41LnRbovp
LWhNulKzsP0zto3cWtSYSYL+HtA0rB/pF4vqPmuibrMCeGSNLMZLzi7Zek87bxv5
Ef48A/V1HbWdWJ6yL+3GzfUfoNk9oJDm38ahRXCs7Ibau8LEFvTu+12DzR2Gc0PI
RittNlrzvZFL8LloUSrRGloyqOrC8/mWFO1BaicjAEwPnCq1q7HGYOsvh5TORncZ
x5P3PCeW54OrDaE8+OwJQ+EjI/HQy00/Dv2Cs7UApjIh0+GCxvVlED5eBbA3le/K
iSSY89UrwlbEqsJ9xy1tcMQ7CtQKBQctxazxZbqoN1VCf+A9JlqIVr36LxZZ6KRo
sBm77M5YW4fdcwfwo1bRFH977fAjuAPG8ZQPAhJfh44j3h7Ps2gGPkTMtl7BvV1M
b9Kje6oLr3cKE2ZsMUIShUL5/zXuM8nqlrgQ2V/AjIuhZtpHsHIy5zU+hGgUblQp
iju/psQUwVGqDpjSy7/+yQD4yXs3be0kFmjEx/S4ncnGeLujBxdGLs8IlNVuacla
tsGKrdni2pH6FiMCyiH5Gu0ZLqdCFlWaAMMIevoHglcRPfVq+xWktSCgC4CK7BZy
m9Y3aqGeiszcQwMdOZ6Lbb/eir/d8qY99g6HOcBFxZieVaVX9T708izONnOdlIzR
GtmSMUZw6XJZA8lK+C0NUXKM21apCRoWC0d0DOCMTdOjQjDM60WWgfcn+PAxwoZC
siFqSrCuvczFZucMTnGWC2Vw0hPiVKM1aSc72Un72i+KUQgcZj26Cf+zRFCmnGvD
5hmHc2xq/76/t2azYI6G5pESyqfon+OHKs1mEGDASQvBs7Bp4cvOYc/vYF5kqy4b
o2mg6iai2jGLMxZW4dUGdGjYNTBSbHcUg/NsXSfOEoW0jzIzIZg6xbiyPHczDxwL
jn1uAu70EB/6x/X7ZY7m5VTm+xl+ldgSBuuepynCry/E4KjDGaiu+IhxOsL5NMMl
yqwuAQ7XLWXxtYa8QJBvgFZQXX/7Y8DPM8lqufH1a5qc3BDTsZcTXDIfjb8Tr/W6
atqsybN7DCCMvJrZvwZ+X5PGakbhwvri+pWSy/BOhIDYy4xq/GUDtflKOzxgxLeX
SX3FW9+IuI6lZWxBvwdC7FnrvBdxLL8XRpzFiOHsO02X4DKCFdZPrTxdgloKUScI
q/fhiAno0dBGBVN0pIylXJwNdQ86/cXX9M/FnXxhNrPquHALw7W4hxbu4qRzQFrA
vuD/z6naANtAPowDGDcOmgBcm3/DQwEM9iWk3OhrGa4imNOX7XRrKWhgj0xLA/S9
ZG0iXFmtXrPoYdAKN9zkoBSxebW7b4pi3uLy7+RgknJT+I/m+++oekZcGwYOi2t1
n3xBIQ57kNHHe3rPjOgnkXSwZGcwZNdoNEMwI82APjZTlltpqPV574dgyNoZVgdl
dCh0tXQzYU+lTeBOdIl0TixU3S4NKKP2Kky2tZOfxU4QOcmdINfPxD9tAO3P0K4T
+wAGqKO3s8X+25BBl/6XYOBweMR25e3tE57L5p5PdXJ/zGrG+Dcucz7EduMaotg/
LNE/uLhzQFHK74GFeswmos/fHAkTMd2NgeLecp1nHTynEwCRLGN4zSud5qz1rGES
lPkn06nD+uNvnPyFcrF50uVctGbiQSXGOU6ItbLoxL3b+B3Pu9B4yOJFOaGROHs8
7w0v5qMIqJtrW7KRDRXxhW0KUp00wC0EOCHqcLQkbvrykEGzGsCLXHAIVbxxVPzt
LKfYhBg87qv23gJipkUVhPs1x3A58DChFpnx1GEtC1ouvmYObXXLlk6H0pXc1OTp
kr0gDL9TEEkGz7R9JQTp2T8I+HBRT7nbcD5qZSjCQ+/VUMroy1r08qlwahDcaaH2
PIjpOft9FY+4g1utmfBQBgR43qfBXcVXuSo/QLq+1VGfzyGDD28TiNeAmX9PyA6E
EZYRAgeEcvA1XuJRf3/xPafFr4dRhK/rnThqwAA73RzPuo+QIU25FWOLhv7F9E8z
/z9XnOPya9rCrQsNt72WZ/orKSVFMW/IzKlP9fUJaar0cGHav74MhugRtmEqGBfm
evGQ9ifHg7NkBX26c90w/aJvUjxO2Y9yY4s03B41S6RHTxtyLxF1r1YypOjVw5EN
2LQO86zrCKPZfCv7YuQhecqKI6mIIV5r97mBZ5SIio8/eZUqE5Ane/htydD0p9GZ
im9MG87Otm2FglKMlndbgtF1ZRkJfhM9x2bIl7dRCh17UTnD01zY79c0HzhA66WC
ZLAxyKVnReYJVYmojiIbbKONjO6syO4DL+v+LXxq1C5xjzrcf3Jft75+QpqhyvSC
YgDaxk61qyafceRE4dGgBnCnx8k2cAfD4tvrofPE7XcrPsyTITfuI02t7f19lcy+
pdld+GXYEcSlK0vyvYelgRw4rzON8RKcYeH94D+UwGYgmOnGPYhUFGVu2WnHl6QR
kZSIdGfPY6IxwaCii25krrL5/2au3Zp8sMuiXPY9f32BX+UFKq44I885C1pBh7Zm
QHAphZmhNRBs8JZCsALp6mCmkHqYywnS5vfG1uNS9D/fgIlFRX94tiNRIEcfbxsR
57knFRsFcCTuEgIGaqgit0TeE8bgiWKf2fQa7W6iq/EV7az1O9AgG/qKH+3+HPvW
TRku5mZ5UYq2k/dClwYlFNnpj/yXq6r9LpgfrbaSLELP4SRCmMmsnQMdEQXWZjIi
WgFOjkATwjSc/SB775KWb3PFjAeQ5lMlTcoMUxPFTMJ7Ud3YvtTtUU376z3O1BVG
mXI2hsVEle8dMRMGr2viVLTTOeCWPq2QRLWM6aeaVK+o/x/SSk41HatMiVlJqZvD
HswhfMEgO63sKVwZDKH4IRHdU7Ij0ErdMoTsopapCvjin4hcX0Ax9ukfpewg8usg
0nO6I3w8kWnPsH5yckSXyCBOLYTheahd7U+dOX8SkmF2LwN/79ORhdk6tH7hQIGW
Lp1YaGuDlPhEyFWZ+e6YyhiEKPzUt7sQVrWc7OQIGtiXa/BGmJpnE6mF8ev9/xYi
dcFp+x5nVMnOx8AC/+q1bsmir63U//v2aGLUMiQmaJfbMm4RPhBh4wd/cCbBn3kp
BPOuCDDdAetOlyYF69P3Y5BDZPJJ60Gdg56pW7CiNfQLW/7i4sdK05Gl20V3JezG
ZpC03lmhvbSK097WZjPjluz3xfiutcfloeiQgg4LecDFgabv6fS5IfNUT+UNK0/9
ng2Pmnl0rwn2Hp6j1t71YUfC60oumdI+QotCXlNfX3k3uzP3KhU5mmimpfzznRYY
qqXo0QC98e08psHrRtOpLzL5ms5bdSgemlGk0CNPwXQC5sO5b4z0GYzUVGiVk87q
QdnMHAmdq1GoFpjXg42V2zvFlWcCZfBx6vTmCsZje9uq3/XNWlDqW+9c6GmSHnBK
vPGTNoWiqR2qErTUbTdC2g30e3ugr55g4zegXvPTnUK+qbiy+P/idKWJ1g2r2WqK
sSbGzH8cRI9n7S6nLdMVSdgVt+fLCKHEtTLhtrCJAnWbLtsBBFq+6wN6+EzPCHx4
wkCsYbCaRvpAx1CY3ZbNosBQ3ki4a95pfP6qCFortK1XPaKD+zlXHDb4jfS12yyy
dEFWtcY2/31O/e4RuvuWmVfL82EX4TgRKJm9rEu7FsJbSY0N7fvil5EP48rfDa2I
KOqZTxZnxIHUHXVJ778IexQdkn2E/pvNfaViGp9KGyVEQyr2rZXMajmS9h7aCeRJ
VvxApSnOrU8kmwbZpnCoyPjumgcvIVn9RF4Qyq5TW7BY9jdlHpYeNEVNrj2ZXGQg
K4rwevdEhwuJOQFhZ0z8T/4cmH3N39vGpzVMM8KKYEmACIl/g8dZA2tzB3yuau+Q
qWrJyt6Sb2neXgjI3EkC7M+1qgXvGP/RbTMFVnOv+/XpOZ6XEZkqK4ma0ZOVGODQ
TWbBbjVPerPeRn5PnZ7CRcbnG2fPHw/Yfjn5ODaiGmhyVAwy8136wgRsUow2ZLeM
AtdC+r71WSjKEOrqJ14qfMQpuA9MyTbuCUkp1oI8lSIXC7Sfy66gnff+38VTgUgI
7263a4vyRUopCuHHLfpvxaDZ3dhcWpqgWA6kUkOtwvdd9LMBlIkZ3YSwoAEppAWk
/dx8FeyhNdIWluJm5hA5XRMnqT2Y5FPdwmqc87X0k7QBjJ4RW3hOHXkN28lvZvik
Z1Ne5yR98BqRkJrov95XNX0w5slsHBLuC/bLXBpYOC2KMbYISRumGXiN67P8kZkO
71sLx9oQoDC6HatPpYQQjhnumiJPoh/95OqRF1xwq4/s6SfMxwI8F7K4lBPRsz8F
h+KIbUFqn94I6cFgKR9hzRdjw8882QfD5hxlKGBHhOcurJjOLm05xvvna6GJ+pO+
cXtBybhcbO9Y9VmN96D3JRu8ADMj16RQuXIG+3tdalk1PchKciUpRrHfpXPjm+40
nzAI3JgYquIuyrkAicsMgDuGT3mI4dr9XT2OqKlrb21H+3cV1pSHmur8Zed0xGq5
WrmYTyqeJabDoXnxZCyb7uGhmjypzW9rG9lONwBD17fn2xUadQGeaLngv2ekpaEc
ZUdqJl1cu7J8m/HG6z6E05FclCM1ONfhxI1EZVFMeeRZdxpQZR0KHFQgo2F7Q+7C
lW0lUUYxUxRpDVYL9WrOWJL6MZ66Q2/TYVTfRCRnfMCDOvOWoNf4NgzCjgl8gJfO
mWQzrrnZ1aI+7tB2A6T3y1vZjnj4cpDUsD/ywVGTtpo4Dgsa+V4Z8mnM++D/zFNr
5X7PZ7KuKz36m29ONGrClW9++HRSjiHeN6RM7CziFIZEmv3EN+O99sHqOrzRkYtx
uLLjSUjmLWmq9PmpqG65xCusEHmGzgJvw3D/wdMj2pHZY8uMfO35gH7tNXXq/JLo
I58olR+dH658LE92TSeHpSey+ZYfo2em3/XhJrPyWAebNOOgPM4gdL7HIcjIxc/e
aDcavCS6VNqJbBBx+OJ/837oBi9M+1JHWGINExqcFGWaaw5G3R/p6vKKPJwifQOs
sWImrnLktt48aXZBasSqDRj4NsUK9Aha1vvAXA66jWBLc4DwXVAq81vDc8w7RZXQ
5ZJSSYXLAD3EXQY7Xtd75jTbmabY+iYcJ0eTby8GZZSp74CoFaUenzlWRwKnsUGU
ONAssYVVMn71GZzLV7wBT8ezq3j/Vi5vUZpdHnitAWblraOJ4Rp+t8Z+j3Stdfws
qA9nvr+DUKqLY6Wz3XbKI1GCSmOhZKC4APXyq2mtrSUZGHC0P3PBwNAQXYIXodV3
i3ahR6CGa4cSXKITC5QIBOE7uyGmjNXxPs2OJvsVIVFlbOz9k3TU25CQdtV+Ad1f
lK8a7wt6hzfNCF5aFqmFdj9nhemGsdXOWFi4ciybmBHQbTlZ14bVZqFhL0csVhfT
15rBrbb7hX7Hz3Ro1C/vedeuAr+WWUDbOsqCPjV2rjxnFtdcTgG8MuEqoHT1rsGL
T27hlX9xw8pUrZa+xAC5mf4M5oLdd9rBrsEywyCSvXp2tX9jhemfCIPpvSR4ZcL9
aIzj16uWY6fXYW00SfOICYAZl/OQz2H4qdrq9Y/OGECWUKwPE+du2ftJzcy72+G/
9LZQZUV/hwAIHs7zViE+7O8Mt9fNpiqNKa13Mqdj9t5Y5GtcouSDfcCjXmnDKadI
40yUNHC/bFoUJPPJd5EzAqK2YFunu6pwWp6TNnVZzN9CHPPncS7v92jg2a9qo8Iz
2H+7r3QHv1M0CYTVIBgQ7c0tZxj6i675+dVdRd3iWOMJDAbO9QrXqbKiXruK/Zl6
FF4jvVfh2m3K7yjQlTb2XBbB2U+VhqPYfw1yg0ligkm76WvnGsyyqHW7e8spV2wJ
6Ce7L552th5EtNW55v21+FmSlgKuj3HjtAWauuvB7vpyldWy2wq6/dlmzqy3rO5y
NSsdOEtvFs9WM9BgwZAFCeZwuPGKjAue2wvj+vuKrE6Vyl2GxTdOZ5/EDu2iM1K6
WbId5gWV6ke/Z7e7h03zbw5dOi4jJ2/Ce6zdzsVeZwtHGouDMWPtPgL19fDLg2OO
GH1XnuoPywn5nkWqOE/hltYB+ahWfjfMldWAtw2uG8xy/SpmFBgaaNIW4SelxT6e
6pDAuO0x/3cyR/ezzDIUFJIds05F4ZaBfbSEr2IqOOFxXe8QoerSNS8PJrVEvE0s
Ehf738NouooZkYAHv9vvN8aywEd3pUht4WKqUOl8sRu4WpBEmmXZWeNZ6a2j3Vwy
hkyKiSOOUPRoEML7zs8/AdJQDh01xLKTy97xaLNh5pLjLJCD5whG5MR8b/HZm5mQ
nEdG/9QIrpgpCC1EJ9N9cgOmqCybHBVB4YZjOYtGX6E30tCzwXVcz6nVD12tVBbM
x4OozwmJfzBjz2DHRvkB8JipK2u90hOGvT3dtupVigwALZuwgkKAqq6865DmVb8/
zE0PF+mJzrKpHWFl1j0c5rKCq0J3RpGr2su0Uio1vH3ClE3jVJWlQIv28qkt5+mj
ybo8L9gtHoUZLnQYzHiVQcJeOOV3FeSgTAwKlnEYietCnMt7/4GxARn42qTmf1ND
6s/cTZE5ZKT1I9sJ4P219Q8EZZv4I3u4S6RK8t1wFB+P0SzRIpLKG5yFfPLIIL6k
s5YdC78Q1D5yyrTfaHtn9C1KBIWsvZcpr/CifwfFWIvXfcS9KEIGcZ2Z0kUWH7lM
42icoxxcJfELUD98N4wQ+hVYaq6KcR32os4hVBIbx7u2owS8tX++ljoJi1kqNSv9
9IdPd8zhgu1BeDsZZzUGM0sPFoPf+TLmunIxoJQmtSWOOLXCkpjmPhnS01NqWrdX
0HpeT+iRgt2V/tBo9AvHudsAdp+a4RafM1YTkF+klR4qeZrkAlWsZiMNwkzELT9V
ueWRdfoMWrX3qJu9pCxWjCHM/XojXdr26j6YpbdDqO2j1O/GEX/oum+WgkuYp8me
au2dn2EGsp8Cj3hnJKhMftRgoNSsee5X9nQXQyJDdEl4yVUnyYkg4TxjiSELypcy
F26B6QtrAt8iHM/evqLzrFyluxWdHR/A1jTDIgyPwAVOm6Zft7ok33y+GXCLy0O0
p96dhlHpKuOezurspIOTBXnI0h8vPsfR5DvQTYFTgErT4ZChQuPB9ga2RUx5lolu
s6Dgj1IoahPQgAy7oR0qkY7yUusJ2lK7WaxFPYHzgpfW/yfcsJ/qWZzdS9btBWFV
TMJXom07Brba9YLVedMK4Y/EDkT2byHSS+I3qgaZjLhFfUJWNoKagsX55f/r7aG7
VvUwYi9FrEl+dl/9KYKWhoyXm0eDu4DPT6pKZuR28j09i2hGdayVFdi0CdD7oXI/
3p4K0l1F4X8afXO+Rb3WOahcknoA0T58F0qNwbOrI7qJDOkghxiKjEdgmLbnaAdS
8/Mc0JLptn7E2itfvzhnkIFvQ5lquGPvNlLzehwCDmVtVij76NB0eusajB71UPuk
zf5jBNOxcslNNWUV3pZuJ1k1YxZDbAh5IqAmOa9W7CXfYuGPuym+zqnS5Hc1d4V0
lPtam12JtFYDwx9tuyKbMownv6ey1I4uf2zpfz4YBXY8zeDtis6if+h+E4gDvCwC
xOk3shJlNyRtHlalegwb/3qMJo1ITajMTsej/1fCr+pEmMD1gbLa4DqBpEX7Kos6
OedQuQRUy9LYlRu8MPNiEa+I0bj7kJbtiI7vMVJh+FiB6hOLc+totezCMXtyQl90
uTHXWyKrOi3KlbzAcb+pTo6G3BQsbwxKzs6E/Y+BVfD7agdgevKAkKJ7tzX7AgSW
qYIPL4wvII4slJmmwmcHURvbdCDi+yzxM4U738s0bWh7nBWjxFYqAeP+crZOKQh/
sQVjGt9hOf1qb/kZqb7bYCHR0Fh7zj1FBDJqvk2tX4G+tJqRLtUGCG+N1xB+ABMw
v/Vh4Se6eNJtz6z2GOTnDMXGvSTVB3h+R6ufeGaJjxQOLHs3eIg4UVur4Qs1CtNc
UxizwmHZUNMTmyr7DrUn9Fqrso0m7nfK02vucavkL77VB/5aZ6xATlAXEzxCUMHk
S3V0w9yA2Z/dLiYxnRo3GIqmB99pE5nfaksCWPokp1H3883pv6YXFvRN2CXOPXHB
sikCgwQ5IBrbFP+o0LHNkDfOvcdvgjSrwzPq0OqN5aPoVLeckRw22xYPpybYmmoD
uFosTx9XaUXTs3KJYpZdNsCUPf7eQgCLM5kVSvPKqKAWA5Mz9Mj2aEk1q/gCeTC0
bSzwoKZsHwVE2EwfUWMmHxXOMl0SUdMvRargvG5fO8uxj8WhUuYVPIM6EdMQoMwY
fjbYZMa2MRp13tqoq0cyozLOW9CDrv2ihlIYTwpf2zmyLtKzQsAKB+IESs5uDga0
NOaQn1S8/eRVZBoBtTtbWNVdY+QMwMjcXI1hbhqfW8i9ofDbHlD0YyXMo6EQAokj
R5VKzF0hcjK/0LlYMDSoJr45DODVFCl1WOCPbcw7VUzN5FbwVj2PZU65HwVyoIxP
7rGqz4c29j5/bld+2UAqBrchphEFIoZovP7zZ8D0TrcTIAq1artiBouPQ/Bo/pwA
9FAqIr/0ItW7p7j+DzYWG2pRCEhmFtKqcjxELrA5wNhXdJcxMv4nN9dyusF0YdTz
/fz+Bw4gIvx1Opm5pD8rAlGFh2cSWJEROKDMXR05fREvTlbxxwvT7Jsr4CKpNugh
uXOl+sdjK7mAcL34L3OFln4DJqbRJ5whUP4KmIAfVB9G2huEfd1iuDSGt4MZp46D
Rzrq7l5exnMJHu/fViBWT2xlLBM6AuDKTkh8DojQCO8/9TZcIORzfjpeg5pGkuzY
4Lua+E2LGlyLtCkqD/fQnfG6xQBAsANEuzhskhLyJXf6cQDY4mWHKKLu3muh3nzP
8Oj7NnB9FCAUWQyFGsrvC6krwiJioPdnizsrEsfviAuEOVm9ctsE8mQoHk9Yxu9G
gnG25zyPUySpVQR5VpFZWqo950uNJFOK3asD4laDL7MR9mKiHDbzSAKK1E+Fgryp
WT3v/jmfokG1rzCbzDOzTStr/xyqg05xoqxDe+SvG+CIQW+l1vaKQRNzB1czTf1c
8Q9n2jfKGux0tpxOd0fjuq35gL+YdPXN2WDUvx3Ncz69R8JJEPtGURODO9DGjXOD
x/Lu/5M8I9gWQqK2auOuqyh+iadGpEGv9Aaeu66F5Nh5y4mmwwUXDarwJ18zJoA6
XX3QJLLQSQAtXP3HPn6XcGKF6YYCApSS4N+saHzUaDCv+vGp6fzMKH/xBziTv7Ah
hSl+S1mYqNpy1WJjKFgrFagcP4a9c+x99ibyqOJaOfOj15mfjgrFOns3klC/4zMf
ujf9EXycPtg/Npypb1IfhNrLGeLXrJxh7mCG4J9laVPuekdlgmcuROPm9TenpUjb
kytDx+wPRZxELVdP+odrn0XgYKA4SQTJBAStoIH4VMySDDFpMG5XIRIcq0tIaanU
0bjLj51SP49DfVlkhAAs2WYPsH9bOh3o/nyLhjpN3dTqA5hgsqW/RXRTPBSGjoWZ
Phpd8UV4kAs/nuYy/rFKyGAH8+W7UJA916wca2cDnJ4YB0cYMMTQZNiTUyrvidSR
rOl8n1ycO/P/rSDAlehc5bUPLmSWyH70lZ5ks2ejbvCUc4rkQny4c3DWTPNrD8uE
toS75GASOzINH81OpqPShdKjKRAV5N3lC317wSI+R1zSeNMMpj53qXHxFp5AV8pj
ZpmpeCGjgy2zoOmwkmaTRoYf543LRThYRpAnkRvkPWU1ZLDdmjN64UKwtTCzsHs8
xsVauDW1v3HR+r8QbbaKvC1iQ2GIteZZGZYTOCHy3OjRqbUFF74o7RdlapvKSZY9
F7DvROf1XGX71Zw0FhWMCFPx31GwbXxWOFx11+aVeoBqoxH9skkmT9ai4EEPd/nG
P4Kot/nykmZN42rihtK2T/kDmwGzfI7OK0Qi0e8E4XYybQzmIzKXnJ/dQj2GHD7+
ROJjjBRlGFj4T01hT8aPiTwO1H3GSaTzndEmASYmFgC+ok8eBG5oJgUhzgM6zLQ4
c/cEj0vvFeGACELRnyPJnH80YS8y6tXlopNkR6o9BpPiUysSVdlsc8QIb+pUm6Nc
UzKnAeMjGiK2BZmO5YqkNav69ge136tRs45gG7QM239btTUhjNflO8hMv1w7DqAo
vGCuqOy7vhSVmz/xnM2S3yz4USIobHmR1sS2aivM24rn+clAPV0doNK9o5wkHPjV
L3GwiaCJj7kXr+K7PUr5gmHaf0/FBO8B+8DDGNgxu6z18zZhH6IqdqkQkpIatHgG
j1F4Unc3lzCylzkwlb1kE/R6JQZacU7hIMi2YUDrEFc/xuiC4YqMtHGT/EaTCyy1
hqlp/TYvpCHqrLU3zm61QKA73dsXcEQH96nXFfgodjEXlRSgdDWPIVRzp7ap4jtN
an/7UgdnMPxQC6n7HOWStVuv18ucY9hjFhJo7jNi/JQcXrircpMqVBG9RBXfxCZF
aCZvCJvlz9Z39PQfYMcy/sFqE0J7flpO+G3xSOv35ovfArULT4Nty3VULSO7lTXv
eRm5UJtdumX5lx0maudsrZ8GrY9XXzpErEgE2lwXJHRRHXdn+E8Gxpmbn9d41cT8
TDkrfL3thjlGZmFW0IMa7E8qtn0ar3n8t8F6miqWRe0tuprEeJqyCuhngfUuHdLf
CDOlle+hmZ5qMzcNhboYGBUgnG2MSrbchE4ajE03wNneGxO9RBV/+d4Amz75Zfr1
tGKIosqosGQxkrmtEW+x9AcyAZFRy2TIdidOyN+LHgzxk8yqZF1WZnRI65en97Rg
0DhyR9m5CS4XJ3jxZ4xXuCIT3BEvouMWEmnhsSzJ1ILdioYhW48uHBQ1shJU6gGB
nfQgg0uARiZ5AaDfq7P55f9LXbMPYOvXo8YQdl9O+NzF2IJSNsGkdVqHy8xTrYaW
vJB7UgDhCabS9QwaibSuBeFoFcOHLXiQEYf/OlxxkvjPCgslSourAQJJMVMnarj1
CbcrOlJcg25tAnu3ZEwWrUIoQwG8wQ1rB3M1NF1t7SJlAmekBo0jvEIY3dBrtLAX
mafGTGJRBVzaen3zoGgA1Q9Voc4SG4AlT4mehaWnDEgQhztzDg2ku2rhsMiTIjI1
DwFuMwS1KBlDJJalzpiBVA4+k9tWcw5nf/Ibqg+JiOrAMc0ezQxMDq88QdIjnMbK
NHOTrQcgV+IIJob2xfcknPiOEMkf36LZw6UpZzbJng0RFUcKsSD3NwhHElxPue8g
exXmW4XVqeyfIbi48kG82Z8yvStcOYQO5PBsxzHuyt3RN9mnTzETgqcx3dAysHbc
f5rIFNju58hu0an4I7IzoLT1NBjSHNcuXoDDevZENYyvpHfNuJb3RrIOUFFIFBp8
gBIYakAifItO6WgQAbih8xotGW68UfEMyQHdYteJ7CmNYbHgx5w0sA3GqH3HslMu
qvcDBInMIAIgGyqS+CxRKSSVTTEqQZD2mFVF+dnqnqGot9ZqO9fyQ2iON8UXbsqD
KZ/t9vUNnw2/QKA+XqkV2GaY3NBvlYGNdrUvExpNPI1fmgROwWkfDn2nHfGckZIG
WJNC9c91MNEnZtih7SobWCnoaCKJBADwkBgUDbRK+bXeoW9qc2+fGjCu6dZOiepd
Cpp36ACwJ9T66ofeAXNB8SNqgWBFWGB0C/R/pViSNIiOJobcl8ssgY8I4SqDM5t9
q7EjPj7K76ZeGlfD65a8F0xShctPD8iNT1UfIigCSiB4k66pylycCU+5YYtn2v8F
xSU7Xbxc2X6Au1y8p/pLYEsKjvhWPBpYZRKcToNTtFJr8M6tpDWzoH5w5VTPSx00
q0wGCIryh18jKsGqNHI5aer9Gsnuf2BK82w8qtc5KdZ+GZT1RROzfQS21dAaqHw0
5EiczQsV0FLhTtHoVtygjqgz02Z5/tPjVpXsD6UlXMFHlUiCuwNbJWDSseQL6EFa
DQ3LyvbAo7iet5tXfQw6jjryDS7SahBObHWhyHT7/StLuDSxttYsEts8F5xYoDnP
36ReSCvQBYJzQg+JWbPme6wblCw6rxjHmdOd5WRFRUZ7+x23QCMW3igXWpzyH7zW
eRyzUK5MYAKEyMuvuvGk8RiE9CSUHFjLSrlg6MYhwCqD2PlgaY7sqcsp1s5+reY1
gn9UOmZK0RH8sfRqJSzdtGrnZzJYrv4wQ/jXLniiMwAVPTiF1vw8BTGx4HOJwbgt
OzsJ4XH9PdI81vdgxNVs/OHD4krY8XNc5KYiCHNluK+ehFZQkX0lhyrGxND+tonL
N78clkC65DEvYvlgi3ogCNpbePYsNb+C3z6zayHXnLBcv/hEvs5W/c0yJo6olI+6
T28EFkM2VjaI8vakEhaenM6I6rWIsyTYAe4NiKiDeeOoGzjJGVfiCgbFghJPdP02
4+NgCPxWYmeZ5Br1HT3uLGtrqCXAHRHtK3qn6exvaeeMHHbGqRFpZc/GEeHkGH4P
6D88g4AG01ePhqI3fdlc4xRxUOHTF0hGOF2bh39qym0qlsek4XMbj+3if1cZZrBV
V2jpgEbAAdtCshzWSJDxCWcfsLKLN4xA2tqdvfrOvbAX80Uvhj6oS01BNTY5E6wW
yh4P1rCtOVmrgwwEjmHH9cy88kKg903HFY+egimpnYzOZEWSz3PyuAYGodDc+MPE
KiIR2Ulkw5e+96QV6RQdjBZp7Qc5Xp7j3iN32SvBNlBH4M/NohhFDUJpKGfWPK0D
`protect END_PROTECTED
