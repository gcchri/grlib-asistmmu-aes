`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aZO9/JGUDaSCSVIv0hjQgjKxTnYbCVo591ui/LujARcWzbpEy+3VMY8hasmEWnVP
1WxjXXRdpvqR//zbM+PwHNWoxfLiDCaCwWEfx2BF4FoshAaawoERvf10gLA6XWof
BsnYaAS84pCWh5NpzLIiB0uutgACnpxTxvpdoDyITBWhhgsZJGxFPXCcSB7Isave
Yr71U890Lc2dcDpuqnwaNnl4u7WhtMFxDNHg8r1p4xJqrH9JBi7w2YKsUPensdta
3yCyingOaBDYrGqAZ55pezJnXXnPcHzrD0cnhLVOod0=
`protect END_PROTECTED
