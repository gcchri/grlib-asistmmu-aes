`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VLT53s+5rPI8Vq+OOtkDiVDATJ1RztSYWZz+GPiRwxHHLN9e6arXgQJkeLOtMSW4
gCjqEbexSzL9mdCZWvovR3hyXd6YySvQyP61r0Dt+bphNXnPiUTJ79mYkUNUmGw5
AvgkHgMzyoAcZYKBEnmfW3PnFm+/Mmh+SpxpfkiPKAxXeBOaWtTl7wV3g1Sy4p1p
wpvvcbre1hM1uowzasurZGFYa552+RKAcD4w3oXMpjhPgvrweGjF+aXmY7XYEj+/
TZ88EcYxuKA8uKcMyY/fE3pjrzLIZpG+YPqWcspuSpp6Qkg0DNIwp0K7+C46hSpK
7FxYuioEpSW9nnjgurt6vQfZQBhC0dcucx4l838H2/RwZ5BV/ympi1n0j8tAOYwh
qOt1IGQljnnUiQNfi1emRV0hzhF+iHoIPhbD+laOUUPrDQd2o16gZS+SKABABc8X
Q/zZqBMqQLsclTd/4UB3SQ04wP2Vw3mZc+URx3yp+ZBypyKgCSPq6iGa3PbmlBD+
JlvDMAZ4y91TxBUTn0REBFl6ANWaR1nSVMorU5hlMkfsT6I+wLQ/+gVdnZSfl9YD
Tdj+4SKmg+B9XooSiZb01WrfqIqBMgAuIR7mqtKEkO+ECGWoNViLJls37opWfCSl
U0dxjpEwqz8QXSaVIRBOKWomPPUob3kn1+JpHR9ZQSkFSp71YjsSvCkvnAnsmzGb
G9pOHMwdf1llMic6wAg6DWhcg8TnaU6ovIpzhLTiTMe5+K69T+yH2wXYxLixpk/b
CCih9267N6s3H8hfCdLhJw==
`protect END_PROTECTED
