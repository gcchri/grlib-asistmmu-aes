`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NzQjLp9rulweGb2nVKj6ym8UBg06u/yxTgBxYR2eHe8VN3Pb21kQFCFismsZRNDr
eHFysoP5efZVEy2QEKqkpmbPClmCj2WMSuYuN1iT+6fBKjThXPPGeR1m3edg5+nO
AQ8VHOjKMaEItMoUX+c8Mas9QC/0Q8p+eRI43vWrxwaEjuL9791rIAnQb4vwxBb1
fU5/uuFt5vlWAy6No9AR44euP/jHDuQiDAtSNS2JSVhifcwwMb0euUt71g5wVpI3
AIxLQhO33O3hQ8rE31Y6v5VU42ez0q4d7qkYhEnTAKvfPu1tZhLl+huFx762DiHw
ZyjCWJw3etIRmfJckQ0iU4tc91M4S7bo5bT/KSbjb66XoEHYznukHycS0elpE4da
V0bjUpUD0BcUCDRnRhpEp0/ea2LnJ49dlmFvtW87PXuJcMaQaWGegkl+a8SLp2gD
rpWftvhZtsBTkJQMEQJSSY2jH2IqPJwsrNIYCOyXvHA=
`protect END_PROTECTED
