`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iuew8ejGuF3Pp7Zh/iOvYxWVgvTz1Wis02atrnlF8KiJJBmSr/I9/qfxAX5QO0TB
n7oexf6iDMu9CwraWERJCRsorqS8avPOOoOBdrh+5zSC7jqC32oR2kI9aofLTTh0
6EaAyaWdWYBgqX3/guko8d2FgPgjc/kl+WFu7v67cml50tSx/BZru/W8B+gZ08HJ
+SOyVB+zhnUD/urTDSM8ypBHt2TsjXkObnwY5CuPnpSnYQb/kPz7/JYlJFhh/33R
mgzAM/ZXpEP/YDPIbK2HPTKv8aE5qFrt4QIJ7PFcFVUGfeCoUE1uVdrZkxpVH4FR
UD8/P8OzmMSQ5US2Q9N9oqj9C4TWaRpB38w7LB5qOBho2NIhTQ9m9hEeWoV2W3ml
SCpn5xMf3R8vPQJGY6jqWJ73yxV7I/Ah+96sGAPO474=
`protect END_PROTECTED
