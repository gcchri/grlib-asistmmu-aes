`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7x+LL1CTCJRG6Nr1iPrftlbG/Ik/nMBIZt2tiJY03ipYWHEIJPObRs443+ch9wZv
+Fo4/ilKgjKiZuEkKp4bin2aNITG+w7FUjMj2S/PTn1BAnTbfIiS0jaa1uasR6sZ
pG+X0rT7OffUizrPWZ4JJUrn+ePPcDFCWcdQe1sTArMBSJ4mV8GJRY/fMExDkdCt
8PmUmDYuZ2+DfyHDVxtj3vKUG1oax7LiDBaWwhQ5gvi2lu/daVuKDLNW1FFVPqKy
WZCaqpnou26MvbnOFvlKTMi1g15Q7EYxjXSrZp1zd9QUqZrNrfqMPH57rg9ocO4X
339+oLg82z8cwYSX/ug1KQlK4CVuNbMM1P53ysCjJ2ycK5PBkBPchGqH1c2ZJCEf
qzEi9sASaS0oH2fJgeR3fKvuRiPiHIU+aqVHCvkhkf/jXWIiIwV3jN4kUP1BQ2Co
ZNw54EDofmNEweTi3eiDDGioxKzXYRRZXmIbvKTacyEvPzjSmqSWpd/YXdGHYflr
s8wSunP9QM6e5UQhMJFGAUICSNt+K9zaTDZnmvqyut/POqRuU91ITHV7pF7BldDS
d6ik/58cxk2lFx2ueDn50xUMjbRI0CY1th6JwAFWt8g9JvnlFcOs7ebLWYiMOVyw
60ogYiolot5tFsxX2TfL4NXp/LCozG5J2qMdWFB2iWVC5zQS+auaL4oDqp9Tz/hi
QOLiaiKok4lBdforjnxIbdhCPUvmRUNu2GkXNUMKj19AbWdk+DOsU87zdiBJiS3t
VVcv6TGov+kQI/p7lO03rNqKIXNP1SVMYxZRN96qOolTfyAnvOFVdBHthrFTI4l+
PGW94lwrX1bUH/7CeRs66yuRcd2RFroyAQeHg46SwAVtRbd3rJzfL6qJoFU5AF43
CLspgJbO9TLhAIK8Th68k2xxdWu/MBK8JCqah+3J2/+VKuSv4zYlhwQt7e5dmGW1
1obFDj7ftTo+2VkGdeTIrLN4AIptMs4obJW/xvf+DjvRG/81MGyjD7ltPJUxVQen
43QNMjDMOux+vGy4zNfOsqeFShMFLc/Qq28A506awDI90SY1Q4FC0dsWftAgCFtT
ZFu1blCJPIo83qA1Pqt0I1fxQl91r6T7Qvtw6HwywmfvgcZEMxLcqcrEc97uZZhn
xPIdOIRBzlcib1VdRs0ImBcUycsfWimChYn49i/aUYBN5kYLZl1afFAJUr1mR9Uh
mxgR2j8pD9pqhduwJG4vSxLL4kMN7e6CL2uzRxPCY4+Fu0ZYyu7LSk6yTsvFpi+L
2lYfrvurSBAPDcnb3Lf5a97J1t6jHlEV7bljJX7hkji5dxsfUP6sdlZt/MzXbIXv
J2o7mxUh+74opTiobT6038snSJ00cGl9ALHgt4swUeCVQboYn9v6lTH76jcOcyuX
gEBdeGFP9KhidWverxH+MxghhOggFXAgBCegvhZmc0HuyLcV5msHcFA+Rs+vWcfl
986kXpNktfq+mXtzLzyA4QznMeSG8+Jc+1ed7EAoJxaoBuEQSwjo+FACtqb1erxB
c9BXd3na9P6mtrEWSrsRa5iZjcFaIbIWUFEh2hkpIgUqTjhRDdJHRl5yzYbBO6+o
f7wpewZ0qdfNyHQ2v5HIDGkg8kSC4amAKzcvrlt6c2SKX1G69d/Jz1uQ3I2/EHgU
I5/lU4c9N53x/mElxw1sbYrQd5xuQDbqyYX9wEHJkyrWD8eyPzJwyE6EbfsR50Gy
lyxTMjZ/mb8/LneYy9/XvRXv+Xm7YwIA86e/Cu3uglGSpnSshcZPT5fT+cswvwzy
sQJ0h3CHpjMu8s81iOF8QFe3jwatFza5VpjsyhlGdydWLL3dO0kOH/WPd1EszNnh
gS6MERNNARAzKBlZoOINbawFOZx3JP+8I0damahs+x6NuU73FNT8rO4HVi6x7dRw
mZQMesvtUxygH0GiFtFt3G/+IJ7MjpDsjonD6mfGS51rq9hEBWwve46qQ2cF4vUy
MQ3zc3tP2q6p9siHbbg7OxUufyHVJbiEdf/CsEG4AIEiGM/KG9HQXiaALajme8mj
Yu44Wxe/AbIgH0NCQloDBGk0znPW0ao1Q4s2ovKy9Iap42fP599PVZAnLwrA88ct
sobL9zs302T4IlR24mbvbyP589zNBjnWS2N38Ie0k6wtDtcmRj53JUJd97zMjxpS
3kL8io+LSjVqJAgdO/EXn/fIoglth6pZ46u0hoogbnKwJIAT3DHc/gfq24dxVa3k
kbtAXd5YyIdv2TU9kBxjSYsJ2ihtWPOuucSeG15WGq1TFP9EyiDUb4IShHpAfFyk
xiK79UqxIgn0yUHnauqpzV8UCoViMBw3gWmYWQ4TugAiffqvXMZMLM4QKY1d1va4
Y0m0kwOo65R0N7FRJPoKI4psoRDepSc9B3t4aydMFHun/xDx7r5s5kUAMCHiNGM9
U0Hg5CwvZjB/sDCJQU32h6UjgJ4c+x9iMOH9hkcM6coPZr6mFbSTj2niWqupQdOf
zntFcyK4Tb5yWLSkri/DjGdqY/YpzV4rIN0w4eYOMWCAUtTT5C+2ItEs1cV405Yb
w6Tb5fJz1b3JGPNi31AESkHssvgNCe3JHsDkAbLpi0MC9u+OpSZqaWsGKPW2fvXF
5zNEU+BbKI6d0RMFyt4cIROZwqQBWa7A1aLJPr0yz4iubiqMySolhmoDcX2GraJZ
a/KppCf0eH7aH5ClBpWvSdroTWUkmeKiLSr62/NIKnjsSCjtQjbe5KzoK8dghDA4
bwmElOkAG5o//YJSFq6XvGnmlklO9tTnfNU2p1K6rcsQd49vSndaKvTyIATTm3Kh
vNVKUUym1KRAwrpBgjhn7s3vRuJsWyAhw/hAasnAQ6N3o3QsQOjm6L8DoRqWTODB
aUv6krsr4ZGIVui2l6UNQlzXmFe/DJgLxdcTAnhUZswOSeMZS8Cue4OPrzPR0Txb
+kh/UMPITAUe9bE5yXymfGR9a6W0wBUSCmT/1fd6MlrVu1iyti9WnbCPYc0lsPwC
JSRHn7ex86iDElh98MkGXbmxzSSCO/Sha4OmsiQU/yKlVPusChW74KF9QhwtYW7r
Eb7sy6YUBpAih9Q5wR5ymVGNznlyr+qgR+nng7hvuwa33uFoHhD5rZkVubV1ofIa
iIXDIrHhStTxurhtHys0aVyRMwOFoJ2NEQ25xxQZVCg=
`protect END_PROTECTED
