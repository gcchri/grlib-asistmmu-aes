`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QWopCSoXv9uk023nekM2azxhk7k4uRejQgi6uThPPP3hdw3qb1gAeQx3u6m1laHu
W3r2poIzcUfC4bXCOrO+S7q1cRcKvresqbobbR9PI+0mQ+NPME39VRioB+/XYZR/
JmRxDj1c3TWayERMT9pCCvjyiDoDGHvGh1VaGVoFXRjoNLcHNGcbGIXNOOm0tW7O
mYnkPH2CBtvAbdviJZ94CFBWOHd/iTbkMZxgGLi5NKPGIShqhc/NSsdjuOOuZhEy
Jo5WqSr5utHQUjDTJfGFYmtT6RXAAcLUco2cd4EWM3DeNqCGTPgcWRYIFRShhpPZ
TetUWMFzPJw+bf4+UuhsehwHne2A79l2xhVXnswu2de4lJ34EXtBNCVZANNXf1c2
5oQ0/FzU/u9Z0M9mfIB5m6RyhdYoNy3Y4qgNdA+yV/PavkCPrA/KHT3rE8ud6ydO
hbKGLKiXn8tDM/OimEi5Fqhv6ZrRNJpjN4ZaEYYh87XcYgD9KRVxpN1kuqvSInZi
1WLqKtpGLVx9RktAQFxGptdbUW674/PCYmJ4bIib+grhzhQXMA18x4wsjH4wsuMn
h6Mtd+7EqahooCPFsXSxmJEu+i/2BLGBzGjONuXttyqlU6hbKu6yEDCN/309B4vC
/1KeDT8cfgkc2dvD7siLLEwj3YOeGVBecF7F4mg8HDaBua+T266/a0xF0D5j/D+i
zkw5xNhCN6rTnJRp0KmcS8sQALQWKocFrGzsv23DGf9jE4G2tv+ait+TgL3iMpp0
Dz4fDuRll4o87jOmh5RArfBhL62Q8aYyWJPUwpSojQ4132FlkcMwUWwNVE6syaid
L44YTsDa+X5fpEsrtpThE941Ha7uMM6feRMHCzvvnIrERnaERv1LCl9xBuFeks93
/fVPtpUicAy//MYFHmFT6kfGa2pxBAiBXkcUse0ewNZewWtgedScmelohUS9OIyy
xjLGUaap3dgeJ7L40gOcy89Znjt1HfOUoMdqg9g8zgpY8+O7FVfbNFl9pSDFc66k
gGfnMxWRbEC1/PHvev+efKkAUNjSmsUk5T/8bEn3HbHEQdY8u5Qzf1rms0koNcmS
98kI73qTyYkGaofzd891j11zMhqLoaKkKal2/FuI260rs4IoxRuuzLz/cZvM4eHl
3MFoD/P1gBuoX/ldjP5isAAZCBhGr+2nRF5mG9ocwU48/IhgZC5s1nXzgiUGpN8i
Ucj0LTbPkMxSqSF2URFkARNCHDDyowwtxrHBeltjIqcEBjsTKJrRk3NF4vWkM+iG
9hy1VvAOmqpOBi4msy49gftKNnKqldbjfIsufoK2FJ4QVT/0NzTqX2+E3ecEURFX
kEj/+F7nn1EUv4ZnESiMwsy0QisPWVvTH4PZctSY4a97hdv82IkHFOqRnyPj/b+d
UbEF30jSk0Lyxbr1y/8B1mHHw5uBSiiYCAggqlohL2wfPNNGLgjYPlseGVEfN61t
CoX1oNhY7na8mCZ9R7RIJ/qpIhZfpsU1br7udzVUlHz4rB+9kpfE4x3pvhe3oqZD
1+SV1SZN5YBShqgckFa+GNd0I1q7qVkafHzG3teX2OFiOrdiflsXvxVJYRkO+9lS
Pq7rj1liZ02p8DXEz6yu2GVnAmgV8V+xcj9+dYKCktzzvVPlfko8rWEPgVIVSR57
XERilZTnewagq+4HsJNPkp0pwUZFVZplVCJEScljAgXptu0vsA3unodz6k+75AL+
p9w7eTmm9fculbnnIMBYsktKOvtBCRRV980FnW4QDdh0e7xMSvLGKU/HUWeDL3Ur
qeVv8vs5kJg/Xe8IYWOqMzn6IepLgUv4xANrM1Fgklbt9NuXzJycYazGP9eboN9a
59zZHpkukN+zLbr76rxNbn7iUEmQSk0fGGelwf3cQojWHFPulxdHnFykt9q1XYfV
m5EdgPq6Trvwe7wRL82SDkbEssv5rf2+ykoF0pag1PlEA8WmmIYVA9X+r0HXpAOw
D6QnbWHvpUeDukFeBJt+n/NuW8ElJpbGJjGSyTROErCNgZmxEJEm+JZZKFiXlQC7
i7pwo/ThAPFK+eSgsyx7cHhyMEdZEunFBzWWUZGfuH6Ht2YXu25vM98EIBjYFqn4
HLWQn3ss1JJBh8rzH3dwhGls7B8KGa1ldDI8H1U3/O0FnyqJU1mvC4caF6HtJbvJ
wrfuoXKdUHnfFaNW1opLOyAYyDIwMcUdTQsMUVNAPvpEokU44FEo8Bfl5tIbCq+S
T3AkXYfOf1CkygNQWtLWo0yRUebYR+1K12bP/BFNVDD245BJeNkqTjuDWn/B7gzu
J4UM+gS6Guk3pAAtspJqIYJZUI/XbXrMQxxcXyep0m7s6RY/t8FYcyRTGC6qySff
yHUsOcN7tnQEvnxvtflNVutpDB99RScYI672+6PK642dD8nCoINWA7mrz6Oaxoea
3oCL1bUraKHYb8q4aamrUJuMQFM1OzVTKpl9jPbyUreiulyefwwjNoauelUQHRaZ
4y1+LppvdnG8HpBozkwuXsPnyAMlwKQoOSWukPWKendrIZ1vSXm0a2WlevUCbS5x
8MX/FqKK1KaxE2pOaQFEztlSF1z2TKewirfgXrQ49ENBIUeys7v5IU9nS+JJ8bTy
K0ARD+B6T6UE5PHNqPemn2Y7t+Z1+ny9h9AFFfAdFosBJX76odFpiHB5897fSlht
TxhLgzMmbwVuTNR+e8umobf4oPfvz3Vs5NQQcQrd/pDfWj8Mg1PRSYHy/9saSwy7
AiykXhzCYxXSgiewccrh0HfNSsSFKztf5+S0zzOIqW7pJTr+uJevVBRJ9VLwv3p4
SGL23CdFJLittmznicQvG1zZpR+27Qkq8W30rr7V+7RxsrmUFoF35BXkJZELZLFN
h7kOXo8qv82cE6H9I9tJ7JJi95tJnNmh1r0R4D/SmfOLaFTe759iVePIASYGz/gD
j5jHudIdy1s4ZasX4xclmx97wl8naV9SZxoSGOCSl5pgOTcFa3XeuV6DnjGPWLxb
jj+WZh2i/2A/Xr9zv42ZPZUa3yIw9cCwix7+OeT8KCmPsW8m6hTT1Ygm/NqmsCuX
xr6JquMVCytDnxOqkVkwstRPnQV7GFJ0vDKER6/0RHELAAENVcjNTBz9ceAx2+Ck
mz4Ajn6ASoRNmTERMfkoRmBo5pRiiaKkqWMKu+x8SAvdSr6DoKhPVZJb5iD0kYxh
EUYswnCee7RzDXfVX1QmMdKPVx18aeBGg9/KE93t9lxsvP38a3+2NCd4uZcyay/d
bsQBkVEvvcZUsMyMJfVsDWidKEmvo0sCEeBhOXR1JntN62h+y1GeNP1XKIL15E6r
2kurTruKzWETyeNKDXnN/E0Tc5uiJxrcsAMk9oD/MSnolszLr1FNs3uXNomwUjTd
qUytdavLbfX4XfLHN5Xn1UZuAZvdQGLhYNcDHWOIxTp5XeDZ8Cw1ORHEOBBZLuAi
WWslGRNPjGmcxZ0teCecaCDi1Gcb6F6oZlZLo8gv9AVCvamiB5x6orpepfw4XoqV
p6ihj65qOQtqvY9CeAUxWZUUgpNcVwCq8nF1XXf319SDs3AEPv5ikbZzcwNiQ1bI
`protect END_PROTECTED
