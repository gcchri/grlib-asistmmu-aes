`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Xl2DcQMPCkgQuXfI4lwH+aQZAVOgdUTYKx4dwpYv0ivCq4DYaOMwCVwqnilqloM
fHsoZFxTml5xsZ/Imx6GYh44oKQTdK/FW+OCTLtGpl7IVd9Tk3ATZ3IefUNID6+U
IG79lild7VtQl6nCe18XxfyzwlpdelnlVQSChVcSx3QuuxmhMEcOpLtiaSarjPQd
E4VN+3Arc50xYApT2XZdrnYWiyXj7cRem4vYLcAPSnziH9Man1oLclFmWip7wIw7
sRGFiM9h5EIjBInHgYMy506zPN9s3TbWJgMlOY0Aq7wgAPEvmzXJBq6J7QFrky/t
TA6wVSBCt+/9F6jDqjmvnCsScDU25/L5DbieQcHUOnVXo7Mhftlr+GGct72HzzKP
GOps5fUuAUnSvgBIUraS/Vu4yJEhFtf4GX5C/QNNKGYDa2e8IbGHHWlXewJl8Osj
r6Z34dicdM/1Sic8uuHqg1DAnJb1wq2cW2SyY3bMNbR5ch3x62Y04E9QyiHUjvtF
so9FRvcMZmgBDBy7t+yHQMrUrEWme5vnXVHCQ5+70Mr27odRhbyJ9FmBXYpiNRsk
l+NXTKwE94ZfzpFxyibPNhvlbmb7zPmJ2UQubD3XH/mH0qdcQHphB8jDt2xC6GJQ
PWX3tMRqdtKgVnPh/AU2vfxpUtRz5wwdAVJ1e7zOouG3Ooi5UYHs6c0zbmmDI7Fg
9sUAOAPjeyOPLr9+BvWpDhHwMR8KqZc082OeWkzV6ayQs1VYiDFf6xArMmmVzOtQ
Ben6qNWTI3/dXxjMACMuO/UGUHyTdD2ZDbf6HZNHF+WLNtPyyRyHQ22GnNZj50yr
ChrEVtDZ35JwXXOoGtq/GkAhSPR0oR4hTdqvlfGiNu/q7Hzj4TO/LKTAUCUtW6g0
Jzx+zkL0eu0DfYqSBU4UqEnqUkClxV4vIClJv5sZ4jGOdwBuQJAfpdpgcPDbN7mW
IswgyhI6vZ9+LhQzA6it9Cvj2RsYalk6XpibgVrt9BUkaLeY4uJrV2x7tgRu6gG0
ySpJKS8WXETT/UAd3g0Jj3ERPySW7Z/cR+T6D2L7plwiu2XFGDipXTxCGjFMwOjV
e4YdivbvZom2pddw+vtikM0ipxD1i7Unyn2VlujAXTYrHgrq2jz3XU507bg8d67B
g1kRcITs+lrBQZMwI6oYz5CiTvADRVfNP5NlNp6L7u7dsHMUoB1B/uRQE4QDTgFG
rmB26+MlCtzUWQPIpYctK465rfSUPuQO8MFE7sv5/UQtPf3+L/reuFoAS4V/+TtU
xJQFWCmx2cEdyfhz7FrXO3Wc/YvimZJ2xBDjG3elYpqGo/Er4YTdo4cA4SKLtrzU
Ky9ZhDfbHxRj5E8lzJOobe7V38iqXHMDPFA7vgyrcGQI5RsEzJosv+xNIyAMyeCj
ALMb12PCmxEmQVNNQ7K106HiV7ALOuIxBnFefMme0JYyg+ZcEtL+rRIlZvimc7Mz
cy92UiKi54litjNFMa78SuePHKgiSYeopRMq446PD2Y0ms1Twz/sj9M63DPgxx1J
Ie0l2rZFeSbzgndTuGFnTlVM5m38nn5/ydviCW/Mc887QlrQdW03+XsV7smUAL/T
pqIhMCDjfNdZzSeWp4BHRJWecnwXQidjfyFk9Kkk2ijfNJMoYQtW9SIcLAfEja/T
nD5Wk5dh7FKyk6x4H3J6BO4nDWFTfSqUvB75xaqxnMyMJhQqH0+GeWVcZvaVk+ar
d1mhz7mXRKUOc6AGc1hEpHscuZvR9CN/uPvNsQZVamEHIoVD6lSy5t+4lBx+JP33
KKAGSx4RbJsRgQGryooEc0Puqlb2sJ6PMxojb/Tfvj0wsOjps//GPa1mna0NA70x
/NQJWvBwHkSvjLcPPPa3VyGw3D7HrPynchC16QPBDDHpd8m69xpBnngi0r5A+qKX
GY/v5eWPgH/PEDIWLlKohqruealZx50tA22D0Jqdb1lXBLnWDNRtQvHNq4IEm6hi
zPOeJMaIjgWk7+jhJ3HEo37aLisxP+84+95XOSXlmpswC/T6tYaeQMKWQE7twdIb
lkvGTamllIID10twlEHDWDeT9iw3zL+KDeBfdjJXp1l7SlIoe2tlJRJinMbv5ssN
YP7jIhZp0kYNjubUSdZdvUP1zzuOit2wl97IxmDaO2JRN0XY6v813CLQY5n/BAjQ
PdKSP0R0VSU5G0beOBtsIEsCj7Phs0R10BbltDLKwelDmVpTK9cL86ogH4TxO9Ib
NNp6xGC7EsMGJlHdgdgEVzM9swz8GEBIPWRdwSdWBcoCqaB5PrsFu5Kxf9an30KR
8vFrKErc/1k33OajbcqQLY4CvEI9tWG4sin+Xh+0s9gbenZ1Ldwzq41D7WOgSkT5
ypNHzHjnXYisP8/ErApEHEAGdRn7YvUOv+mI0jS5qWLAhmg3jBUE7Wz3KJ/sv9I7
WU2uy+ADTQFsZT30LXvFZ9w3xsp7sQ1WXZ0StMd7hhZvpvId0LQ//PP0rlxkJoe6
Ys8C9PzKzkfAXm6K28ACEala88HzKAH6o9xsFasJ0kroVLgi14shPjVW51DbRbl2
JyZokCdbKip1Gho+jxdxLvrPhvJn3KHzwV9J3SHUsbTRFw3Fbwb80nNxtHCaIlEW
Lax3NIuqYu8zg0QY4ksyUJ1v1zDsk5nPGjH7qif02e69DYlAkOI+sw4vLjc02IvR
s5Q6mAEiUIyb8aPkhihMk1KahcU8dTsktbn1CpRtqt5hxFVbF8yLU5IPjH5tKOT+
sQrV3tidaUlVNu6SV2p+2GQdir0pBp85VGXIE+u9pQJymdUwRcwn933QdKYbGJTc
2p4PrK8ba8+cOCx9nHV8AtwGP2uxZmIM0y9gUi67aYSrMnyVRLjyUUGd+uo+xQly
oH2l73ecQHAxQW49stk237uoT+oBgBo9++oS0I7z8eyFZNHROnWbeUQLBMspmcjh
k/nrAQFxMul4cB01W5Cu6nQ3kV5nfTe9VzYwHHOLyo+z20Y0Dk1MvDuHwebP2L8K
6jVw6TSq1v/iH5EbTz6xX8QTetzAPaVkMy4KMuW0c+NI8YjzajGs8Au/cvkQ3GBd
iU9rOwgnM10wR76nP69GiDoQdhASk5/ppwP7yhtGdXn5cYEPhX3qKmdIcXSz7Yxl
/arHWBUdDVLsHL+Ngw+96t/5EWzYG95VOuYFzJpz2NlOv5z6wohffRcED7w6LkPu
cdbVDhDzZvdGSfdG0iS62R0vkUKjAzk1XX5raYekj10Flm9k5harzZBtuAL144lw
SNUbTLG1XlCuMfMBnlLrjxNCrxpNRElO4cAB6doyqWagLVDTqC+NhwEUOpjYvCA0
keLg8HP6quiUVdeT8YWBNDnv1I/REI/UpFt+1+I8OAYB6m+GQxzVOpO8wWaKk17m
kWttwCNSjcpFomh6fTNfIkLyrZOiCu+fIAM/Wf3Puz5JMc7SW5smYcYQ/X/Cn0S7
zqidsF88grkcxBtmxd5PS4tZthHJvygH1qZWbKUU+m7hJUvOAEr2P787E5fo4r3/
wE2lJdKQWuiJLet9NOPwM07OB4lbntD7W009yBlN2DE9uHiNpJ03LLl9koI8SSrk
hA/pNvCAnyaFEy0cSJmKdJPLrF+mQQUOncclIIi5M2ehMKEkdmfA/3ZPJLmF9KIB
/ytbrdPBkIRv3klpY3j8l/IMDcgAXePvCLv6/Abx5UBQtuW+OF9pwDThBlZz26kY
r1xHh+TTYITLFuCPqKwzfsyrfHErKkzAUra341CulmAOJ7g7BUzBNNG/2zrJ7Gys
9qk7JcC2dJnJGM7WmmGvullS2Z8KgDPAC4zoZRyzlaEhktmeSgbn7XvUTUkoO9+G
JR6LkBlJQwxTsHDgz9rGjinw1qJN8ZhEpgRMlJgILRY3IDOAFknIy361wT5kzC4f
0pMj0VBJTbwdQZLI04q5R9e03bCwGUBwN4EEfyyhM9hxjzdwt5rYcVhtdpkxL/Lj
DSEl736UlW1o2XWFfxkM8cKApAZKDXolh5i25gLqO+GYWfzxI81M3oGMMvHjLZGf
IhBIQI933EIZfSC/NHN0KaH8Os1eNNNRDxEDSb1zZ08PX143phOAIA3nd3zWdKsN
iU8gnKch69Jfcqk27pdA1P+Nbkor1czakA4b3m7/kEMhCoAd0vdfqroJ6IET6qwt
yz0g/nJ+TQ+2vBqGjARvubkILIikBXSPEaJh5xuKjuUtl9qP0GTGegrAspiQtytF
n+BosoAuboWJTm63h8PPmP6aKTVXvGF62kNIo0vF/j/jAXxIo200jxwfqN+1KDS2
1w4wF+Rx4Xic1nrPOKghwVSmpLq7sQoDlXaXwRaixnzsRzpV5FFIEcWJTLuZqtVu
CF/LK9uP8CS4gn2bzAHJtb6RoggWwG/dbeZVHCqWoTbi9mJPXw/c4T6mFYJyo3Ms
r6D6yLUP5RVRD3SzSO9WSanwMPhd2ihQu0prmV+KXXDQWSDkVPCPQpvm4i1Ezqly
ebE4ls5mn1dQE6ZxOQoTiywPnBkWFe2683RX2dEFpMukQQASw2hVWJNp5VFDMbtP
wbIbj8Ubj8c5JmAGY97ZqvjMng/dzEmnqCpksb3FuEdSHy5Vcx/9e8Abj2rtHL/j
OHd0iqoBIUonXu7M2Z2Iw2tBXb9XfgZpZHJmrMRbCPyxBzB+2K4gCf9xuoSCxQ1c
TB9or40WoL6xgJB3PN7JDxzw3JY1EJM7Dg64RhDzJWowvAjBIPmKJnF+FKWODvCn
jiWZbZxdfWL0a3DYJAQALkqft4iGrsb5vZRQKYR2WtOhLfrKiHORQUapgU2+y44P
LwY2czk9j7DBeBO7xg2JEafAXn7Q0Yxdv7ZoAtxseGU/tAKrZ7ANjTvhE7/VbIno
xzC8Dtr68LitxgpZvztABsph624ZABPQwrEC0ekB9zQMDdOC1Oj41F71PRHDeCp8
FKhdZGKUcGTA+NAc08vp8/5DFmnhpU5vyDgtCldN6ZV6Oo187/wHQrTb2EihlFdz
m2WCoQ2a53ba6+zEzn3hDpqOPssdLVTQahe1ufsz95pfsB8BMotnVR9O2Xym5byY
CD/FcjchHRRRNyd785mXpObhQiDnwVNK4SK1GHiuajQ9w029FK/GFS/asOQUsiZ1
Ya9buw4Qr3DlD7zl63MRXkdze6NNogHGMFgqx3eRfZ1QZlt95fv7G6n5Rfjp+PS7
J1V8pJRtdGios0qZmItHpE92jT7LyeQopvSAQBXzEbSxmmSvFN2rgwZgl9EvSbWm
urR37phw7zdxEDzY07K1L6paBlVIakDpkklpF0avUFcuucJqPfUC64nYkZNCumri
MWA/VCq/x4B7kE/+ygCRRCeW6iQ+QzcSZBMjhUO2g//Hoi+FP9yL45dlCEfC2q8c
K0DvPHO+F1qi71utWjz7u4UZh/dQ6A4+p8i5HCFWyNzjIIwNOPW7GRoLwcvGLrWl
1yDpw6fFmx+PD1Bi5fPRFbezwBXtqHguCepeytYZVGGrBuqe+6PxLC32MWiUDK2p
vF8xORpvoeSmJ1ibu93radxmJhQCp/7oWh6f/HGnP+fVA+67Q+Fdjvmwi7KSEau8
F2c88uVLPqhReQzPC7Wd/GxBg6qTtu+HIpjt+z4+BoT2T2212ENr7URvQhttWeGd
4GNNvMtw/pTKFnYwbP3tnUgrUeUpxpJUZVgsv8LIfrZr71dgWFV57zMblDQQNJFy
JPT2Zh9HckieUyBtHArw7qC7SHUdNNGUTQR7HQyZO7/2oudtrVz+gBsS9llxoJ2L
hcAJVACuddJ1XrfieUiyIWSrYBAcSTVZzAiYS9QAhQH/Pm0eK3HfRli6Swxq5nd1
+r7qARqIJzYBra0PD+5pnWCMuotMlPeI88hYyG1ETSemJNXSKtvHFmobgjUuwJFi
6uM9sZs3YgxUrS/3QvSmNGsNWJA5Pp94LAosJ7CNnLxeE0nPt6gg2nzKmI5ITvZo
+prH8xN2sbMyqQP1PXrH+P0MEpQIbfOJaxv7IsHb8PDuWbLtb6qiOWnaNeWFKQul
2nEUCQAB0CyXwrc8hsiZ2H3IAQlH4+/kXa0caDx0sYKch1iO83lIMVucLc5VpFBa
FhK2pI0L6ZdCSxzQ39EEDQ/onUZHiuxE73E0SCfiAPym2/WYu+oPiX1/fMGaET0p
eIsCStQQC4/6gB24hNyH/wRMC0mMB3IYjyEmtRXHbXi+Km5mPm5WYShRa5XXbqNo
hul+79CZYO71ehUrz7yEnAgKVEnyEEkVbOSG67iM5ro07UB1cuEa6mLUpy8lmHrh
pmSmkr6NABg/lLMzb5/4KoZYrfQtxYALqlLwREZ6sGCjdeJC00BpelxnSSMmFW6p
40f4q+6Do3cQ0wZgq7vT2xEXgd2tImoeIHBUEQ/izUyA2+m4Be1qzMctnZh7oRGc
OpLtCDINKcrEb4dvnZ3QLH7G7Q+gDYJRRvgO+1uoIMDRo8M/FtWAAzzrUgd42W+s
rKCHMqDvICLzCvoWIWvU5UYZiAmPZdn/yjlhea7DRzhcTLyVWiYSHs65MXFbSMzH
fh0+rlAO0kUXZT59B9fsokUhrTOYdBu+Fh7ZYtnSFk5q2u8LqHsbrCq3h+3tMrHI
JIthNq+ITQ+6J84i7uaBS3hqTUDRbR1p4DYFC2Teb6P1+ShNYAdwiQmvhYOKOMWB
6p5HhhjsPCcEmOgiItcR5RrkJWATDRIKp0+48aRVlMv1p8KkkqIMLT3TeUhYdvgO
75xMtulYXXiu23X37N/WOXAdE3eMflBZGRm7MGGb8LsTru71DWyBhU3kHPppD4Ai
yxrTGzLmuufSs7oXdVzGjDkwBjPlcVGT5A6sCMA6TCjsUub5smMKC2Q/MzNtfqQp
IU3kY0eUU90UG8LPQxRu1rZzf/UWWMXD23+cjvIlCETdl4MBwQTu8gE1l9+rmoPR
OPagR48fL+7qIu3ky0WiJMuhqUmc+VjqjCnobNTDDIAWzqZl0mGVTtYVoJsUvUvy
B8jI10/VdEels4bAqjeWX0KmnrWNOC58/+UIp9zqE9/OT9GscrcgHTpe9Szdfjpm
bOT4jKGh9/96dXv+U69CSrwejjEH+OBt92tufPhIJc8OUjDUOxKqxcnGvtV9wQNv
zTBR8qX+32JqsM/jCTeMT3PJOzY9QSIgGinzocIR6Msyzfl6O336FdZGV40rCMRx
qkrX6agyORZOyLUna2BgEsQQxfdfeHCvThV2E9KVCHWRAMcrqNJqsMspLvO9eVPG
iymt6H6jJ/U/qZZk1o8ANbYAmq/vdcHP9Wv8h/9T9vt409mkZH6Y3XEoHICJZRJo
dntzCKfKbRo7JgUnPQB7Rml4NT/sQ6tPmdQ3cSe5JWCZvvcNshjyPuBe8Z4dXWDN
HSr2DSTbOKf44HyVhKcDJE5cO3EyMMbnW3H1Z7LpPPjl4O0wBL46NeQJtbSngS4U
hSa3fZEPBTfdGP6OWboHQFwLIA72o+TTOtTCLDgZDCClq736U5P6emcy6d9wWLMc
WWmHViaAFAGpBIgPsrH9ro8Pf8vSYBshgDZNbOyyfpgpX3m7cKM9vlxvqhr+z4z3
tsoCxHT7VrNtMG/OXxBsaP7TL37rr9jd/Iez/Xsh65M8NEk3i6u+m1Fjmc2ptic3
cxAhSQjPCt+63bZaQDPyv4kjBM85ePdT7AwYhPnmvKtXaFnKzsXTgLBMLztQ5fp9
2fpjmeKPsr7cr4i/NXMOq1dwLO9TbCijU+xKBaOIAk70mz9iUu4mOnHPcrr0zeTv
2n3Lh8dv5O166xzcCle/luuPFrjshWGDPWcSHwlQiUt0BsTZFz1hRgvDWKf/nVU0
L7lyozjluKDspFiELkAV5vugMyAPcnqEBG8B25rnWspQPp4NnHYDEyGBm6ba0zLc
bXKWDed1434k2wZ1fcGadbvxbl4yv4kyu6YJo1M4nnBv7qkHEa1Fu5LzT7TXuA/h
LzX1IzD2uvvTLS9SBPlc0LpCVz6CHUr7q3J36y5XNq17bnTVvDv2HQIbYxm5UGl5
5zy8Vg3HaslsTzMG8jJ5TrAGHjb1KoxHB/6F3ifth6jzokYalWN2PcBg6EIaAh2m
JlHgKMDRnyMIUhFhrFI4ACHFX+aSkvZPHm2n+9w28FvF8uCtGkN1Phc0TFSjay8L
ovr2y4gVMASHKi6BlzMNbbu5irT5X50QiWzrJMuQSKq0Yw7y1c0OETMTadRHP+R/
SIvj1XjzoEVch+/U6NGoepPtgWscwqYx0qy9HZmOpigIMOo10baQ3qSqWWujBLAw
D7FTwG3bpU7xuSp7q4FLXxO4b+CbGClF4TZHPk/eUe8Z+R+8dzvXa4hQe+2Zp2xz
1R7w0kaXTQOcEiAdelsIhO9MdiGn1/n7yaAqVm/uB7XjEbAhBJfxvLv8bYH6rjEk
YY12cmVgWlQisPVJK9cADPZgzyhgVl8c6CHxuEwiuKLVCRrVsNiGLs8dXYScde/E
/6QZlGY2RQhRLdJIdNSIAw7W65RU4P69cHh5nWr1axZsX/+GFNLcO4vSrU+Y/V7l
v/HEvUkNbUgMlNJ2OPm5v4JrR56sKUENmJpXHoZvXxyCEXJzNE8n7B2B2AqPhInc
M/QbatqA9qADyvVsOtEkSLrf007vA722JwCN3Bsc9CYuNBhkGYJm8vsUaAtdQ3rD
43+RyfKDbLBBqydQJFFBYyOK8G51T5q9S9uVvwjGsVF2dUedfYPRr/m8E+Jp9k3u
6hnmmO0FgBwdwHkeWY6zA6i+PxndQHGUw1TloVLwdxQI7MNXUDBi/qRQX3gOrCIv
ynOrV7AmXhgTIOHUaGbng9kw24Ft5qUeL/CIjHh3VbyZDL6pDPVA0oLiyoFMTged
ubKVfr/PFk+YyMmHx52iqw58WQE+gzlArqEBytErcCWSciTFUXHKu8GcHuNngPNX
cTBzh6yamF5eJIiHJUqFLx5X49ujhnnDQZ1yFzHXJM465ZGgTBHZ6U+kyIS8OSHm
Q+CtSSHz4hE2BaDQ4U91tB54gbiK0VgwwnEpNtpP33V99en07a1d5chRZZYB1AVv
S0tHsrHbXrfvA3oWLiV/CLmM/8Be0lG423J9PEpW5ARuP0lWgFlQB25pg5/M0Tzg
1xpcvIGkhmyYBVePT8lkK89Qzi0eLYax5J3SVoOpBpD7CNwELXO8Prp8HRxji++e
pjSIqHD5WEIp5w4DYZ5u/r/m5VLHR/N64oCq5T3besDBDUBvk0VYCKzEO1WuY7TK
zRzBAZ9S/Pxwznl6mg3Rlw0o4C5eEUNpL9vJzsrLYTREq+ZoT8PQr7iXFefbqSv2
fI52NT6q8inL+qZIupNnERUBNCNDPqML8FtJM7OnXm0eUrH3rrTUx6To75CC2JJO
gBqGzd/3sYZ2u/8zEwPjio3LuSYAbXkf2Iux8h1dE0cCwKmw8P9moadXbhLGVu2R
b6Lwdjxro5Il0Pa5lFGgYOfc5CjMJYEG1t6Af4AjFuO7iW8VzzYYs0HTEkGw5i//
wrePhiSRHF5JIh7FA6b7LSpbp5nLTXek8yuNJNo2MeVHWiFqIcb8wlLZwFs6XnU8
0R0GJPWHEva4NrdBSQhAaiIFY2Ixf9xvaedBirqJODEu2WQyv3Ro1A0ml5/QP82U
oubd9B8aXgvBNbpXO53i56JSvPu/iQtXBUF3OdA78DTNV8+d5egjWOxnIrcTGdYV
zCDkodD9D0V29Zfcg0M57TwhfmRQ8Q+w+LQhqYrcupF5gR0B3XlkT9+8hhCZW/Rr
ExVueNzdhU4ouW8xTvuRclKpYXdE5F9tshVohzOdJfjL3Emjp6bSnZQ7mu9EAsRZ
BX/PHiye2sjtq+TV6vkT9T9prkIYrjAwalTr8Yx9gP4929NiMLVE6AjFJS2ceGzm
upD4EV8eNNXBfKeU/InCC6EnPg4cZIoU+ZG9MVRqq3B+lhRS/mMbH729KRmwad5B
YTvR0L7rbKJ1lY97Z6Ol3NMczFxgDk9V2UCIjtp9aPhAIWXD9tkIu5x5KvSKrYtP
WkAudPrxBujwKYGv/1fCCD6xDm6QtMHT9tlYoEgAQB+JReI3EPumnPcoilJFXY24
QcRMNhR8qYcJxGR3Aen3coAkCHF0agPcQO4mJAg5/7DVzCUF2iTpvLeKJCvS1d7X
/TUu+VXfuPRYwjkVAD627/xBh2Ol4f7GyXNsVSuhSPVImRSdf9hI37yQssHC4Blg
HFp2Yc+6DmKikLWJaqm9ica9z+M/oyiXQNfwY6YlvYWy9t0Lw4xp0GRlmNup9xpA
3KqM+sDVnJwuAu/OK3UrkFe3nVFCzzRJaZXdOvxJeFSz6veNYUvOBwK5HEFfrihy
XUQ4FTgcO1D1OsX8QuuSxZzxHUQelpttnLL9Phv7Q+jdIo1dTWk86IU6JSFi3RPd
sat7/66xkCPUKlZ5c+9gHxTcpcG95bYZEzXGXgJQwrebM97kxXpyr4sQCFCA3Q34
QAhaYLKE2Wo1wdwTAHkdgW9tGaXi1QmO3sDPWXE93BHs3g5tOVEmtc3L4Dv3Fp0A
JFHOHKp6l9ioxA0x74r0XIqeu9EBQISFwyIidG+uv+OsdLYmGR7rKLhJKfYRqoPM
RtWOwCfmVOoWL8ttRo1QLxdHhhm1t3MsHnSEvFHa4UbqdZ9KFDrNTvGl3zCzaMPV
Fi27IUDkYgxnhBZeb2nVsYPCMG+gKNwtMfIholz36u3vx3JPyKlfOw7IdGrSTNEd
i4mIOkIsYTeUgMumiQqMF3UFdc8cTgazrZMGOHriNX0uFY0IVOme3v1P3BIiN025
RDG3DRHKgj+N42qqZlIOC0DjsE0tBtWsb80OgNLyeXmyqL+n3iAV36wy1UGh+s63
GX6CLXkoQGY0wTZLSwP3bi7SF4XMCudRnRUq0HaOXqjD67oQSdKExr8w2f5GT6Ic
JuCbmN9K+yabIbpwBt0Qs9Pg8J43fBSkAwdrqOFckeBvFqc364KNYrfbjkxyfbek
z25/rZ5x8uWzODxEmuR46sE+JZkdmR0rKGKYf3ZcbOMPArhwbpKAfLqO68Arpg1r
CSt78soRxoucuZ0mJdTwcRZzrwiQ0QtriB8Jh/yscWtBTrW4x43ugDtMagTr8fok
zwDD2HP8WvPZKRRwliKO4nExLuMsfM3w75WGwZlwgbH5aIyidscclW6Ujr5iI6iB
4xne9lh5MgZDd1d6Jv6oXvWAHoTni4r8s3J8Nc2jX2d20QYsPaZdOPyvlHT/1a1H
63G3zPXlSApBa5N+7UZpq2fCxMIuhxwdu9OPKfLygNUwO2exLOAYeAmYePFqiODz
4AmXkVmdoTvX451tBQYH6UNpb6hWIWIIzRhKVwjmfw2k4XPTXQEQ8mmObWxI0MpI
PyEid64YDv69J+jEnv7QBj6KX4yq6Aa/yTgg8+bQcFq/m9XkFSMhWwok7jfEvjaa
gs/FUgcle50RWYiu6PDHf5sb/peA4cAF+4nraD573vJSsrFaTMOVG3pMGm0/5gxi
H+5Pvbb5/AdUDjb6gjFiXl292DNTlS08M4CFWKzV0qdD6BZr60hpNyHhdzjiH4I2
3xT0zOO1TBBq9w+2wp9baPjh+PVeXIiO8JvF0LhIJ0nRsI1e+IOYFxOlK54WJbTO
XJ2e6uYT4sST86nyLvXkcAvLxNAqYCQJocrljTiTzs+jbf0rmvXaG+j5K74AbgeW
BT4WNWELeqtgjRZIsTJgxdmpECgHYSiQB1qeCWzkUqzCAf1Z5p89a5k2yaJKKN+X
MqvgAIvBiAwzUPisw1KnpTNz2vBQmYDyUILtr+7K/FG+GFGw962OzfgeCmYnf0xa
U2AJodAy8SWv1BF4a7N9rVuFW4gnmDmSC+PVJd3LyGC+3VrhxPvRziMOg7cx5dOk
cykCm5I+ka4ui6L95rETLKkJDi9nlUJgWV9CEhNi79sDjF5TcFWgqTPO9ehyHqO+
q5jfC6cKAxpkgpOELdGUfnS5SqiGteWHEPBn0vFrzUlGycRonoSYzysKlFZawkwx
mrJxloxHnxJBIY+T+yiwuXOCL87x/EaXec4ETsMAEvyjTTsV90VAkcWoymBxOQxJ
KL7hz2ONKMK2wePYOR5nO/Uf4OofogyReWEtJHw2SV2aUmOxhBg665Hzx0Vh/Ehb
NEcKK9r+MnDjbJBekt1IeRmGZSNVfUWE6NP/7Gsv9o4J3qPRQUmImqxFguGbI+o/
uPu0G9J2Uv2AYKY1jDrKZaDf9SwR9pMreE3ZyH9xZCcrngeRp8yZhz5JWAHhr4ZT
e3p4OCRvWcTaImFihK/iXuj1kXkg8IGotIz3680xkieVnTh+LHfmy4d/kMP/hkmU
g6QAhZVZ2Rxz3oTnKsgyVbdEm3rVdGiF4cIFvozvZkSkpd7Q1DI7DbU9ZQ35QOB0
RuSDxwEtt6YfYPYpbddoDC2xRqOCsa0df0g0Tgj9zALth1Y+fRFvzCGUmTzB4+0O
NQMR2YWn0XnkQ1YUW+CiRZnQW9dvVu7odnAXEjCXc3hGliDHRugBaLlji7NOMtod
e/uMiVoiTWqZkUiWfJyjyTG9DcXLGJKjNmuTnKC1KNSFyTtYDA/IHeyEoF7Q+/Q/
5Ae1Z21QzVeMGObsD/sEAhJM6RPTUTMGj+aA/NKINPmSj22beOE1+XPcEuyTeI5S
0Jl/u2uAr3ZdfHK6o9UMKA2q67p0ax8VQuRRacPZ8CwToYOEgXVf7u3KgehtAUSS
JtLgjREfBAEsvM4bn9a2BwaQaHkn301KhGN2gAPuy/Dkyvj5iZF0XWrRQFFDvJ7G
BIYj9WnYBSH2gyuTqzUb1HeX7by+K61wlTvP8AQrfkPxjh0yoj/CIO9NgiPvaSZE
59qn7vszJhbLl8limELcl91FW7AqkyC1YKMAvT3yC/Flu6EKIQ95cCZwcIw0gQSx
tEdENoE4mQ/KStI8Oh+uKzwVMkgwEoT9+804fUTM75EhhkBuyQ8kwCC1/6pN7Fnq
w3rF8IMOB8T4J6KCSn+h9H9cMo3Q6hq0fBn4PLams83qdttZYEK9tP0tHnv47GBQ
NkG8veKfYokTydOAqrg7TeYePsCp6mlcUIJwpn0b7qegwFt+uqaDrZ3Be7r/7LEw
Bw9lNsbQZyUNnk4Rf/6KBbIeI9LMslARDpFmZFHybuzgfEaVvcPosnpQzthOdvfZ
zG2OYymW4zovL76pFMVInNnttD0gBKp6wQGh2/zLi3fYzpHJbu6GyenQpY6g4k+A
fpwd6soxtByDTGFyXaU4FJ5KqLvoWqWc77LGvdGmClNc+sEz4X8WJf9brGugVGtf
RVNxm1rFQuzkf6ThhbtbqIoCPjhnAJBiugacpQyavln9ODxmC3bvsK4ks4Q6WwxE
d+AywLHq/Glh9STVxmKE5wcdhHbBudchcE49yDJntbmbiDt/nosc1am0EgpuAMLd
AvdVcg9fCn4NPBZRS5nOiynXIzWuT0cgDZgk95heDgxsg6wI9byGEFtN4SlXKcNZ
hRKJx/gRDIxeqBBYxsutWvl5PUyDNzwelRLLoXSL5sRrY8jMG8Amc0qBkP6WOZ1W
4hZgU6uqlYi5Kp6Z+H5TAVaTd4n0gCH98d7nsXKk7N1P612DNkDDv0P7f0Ef5hUk
Jk88WBAQ58NNM2nRWsgk11EsLpJXHfPzGiaY7eeBsMOIciDN7NMyKSpu92sVlHuL
jpYNTeNlHGnHUqhZQcOTDBfS8N9U8n93ijXSnlcHbg5ObqIRuO1/M4VMJgbvXphd
WY40AMbFS/H+F6GJAaXHH900MkRqY0nf3B4BRnYNiudKQRysdeC6fi1STaDgo6MB
wTIAWCeToboyWz5vW7j4I30jGwUoJdrhY0IBcyoH1sfZiMOFUG26o6afl1rxJ8Iu
YgbskjHk3CGAkvQRuWniM46qyXtphmo9imMJHdB3gXdXhH9SEDSqDa5x15Anwu8D
M1XcOa80nyNjBN3dIy44VFHMvnO5DoKnw8ibugusYghAIkg4vQ0kFzkvxHmE96bO
Hx2QjVDstB4Yp8o6TUO01cKLBYz2t6qF4qXCiQpQtqMxZPMMusEcypkHGkqLt04e
SmVjylJRvsGtVmrRMkgZbeipt+pCELCpD7QL998ychDQorW1GajrLb1gcSV3Wbvb
R7ZmeacxikX50RJUlOTfXI3muKRNeYFU9AADrPfvzmNpU4yTyuhoaXnp57qBkIzT
J+Qo3LGNSbxN5QtjSl8TRA/oGkVqtVZwJk3xef4qDHLO1mzEIB4cmKLCXSk/Nimc
eV9ujbC1HJrRFA8mP4voHvRnEpcoA7QM6jZFcgXGg/tNKnfTS/2ZfmnzaRbsg+R+
gsrB2O55kKernLQBsWhIKxcTGjRa+pFdMnOeeZpie6adZ9ZgntCAFy85U9PI8ZTA
Ye8MWBWMn5Smxkdxgw0ajCaarG1o49/aIBA6qnSGlklMJ70wmrFk1/5Py6cLpOe+
cgLOskPpmk6Q32BnGA8/BbHVDc+OgyjGCKWoTySyXHp3f2eIS8kH1zNkEDi1GlIu
mazhyXdDuXXoQG47ClyEkfO916Wr/sjpi0PcoKmYAWXuaGG2i9m1CK4HExiv2gWR
qx+InWAf6rz3PW3vOgCWWgk9wEan+w7oKTEq5KVPnS5J3u475MqKrRj2ZIhuGWAm
ucRA9POXEl9lBwU0rKZ3Mx6xmOqcafu6Era6lB6UnGZPM3TdHdCJBahHCaayBZOa
zJPDugfce/wjJrq6d9vnPUb2r5G08BE39rPMWTS1ecU47ny7c1y/hs0TrVTXfw8T
wzIBJJfwlodc5ytw1sFywxpeubQJxQjow5+kroC2NwqTbMUPeSxuVEvQ1YDcvQan
rN3Hgo+6AT1Ace5LCMgX7l45ZUc4x1ieVANMi9efM0L3FSNUi2rpoI6g907iHZjh
Eg/HMiID2jKK1CxAngArNAONDJj+Tt5pL4SM97Bwxq0NcM9Ct5gGSyacrIFM1ya+
XVMc2ZjU1zsIOGnfa7hXzhH585zSCIu6TWcFnUbsoPONqmSWuiufgMCdMVBTFylr
mcoSOF8KS7+IrmP1X6Hf5vNOhgt0ibif111hug+adPeQTTe3AjGQoAY3Qp1Yl7zB
OjTODiaJC+nTrcJPfoHG0XUQvI5dPURJsV5JoTb1i85SRhZZusgRx4Lji5c7m4Lm
N0WvHokTpd9s1a5s191qOgAtpULpPUDDlxDxHwHuocQeUCo1tzmSsXuZqHrvYyXg
0FKgEbH3Nj0G1wk6x2CTDA49T0toMcq7N54977rUWDxIHgGDxI4CBTZKjE2Oy2as
QYDjcbC9YdEXPcszE7p8Z25sb4LnnWEm6LGzAufnZghAjZE1NlgXpyUFAD7DyfiT
MXg5t29kXPn3DuYRX2/4/zgr91sSBPxEKHUEhHV9cHDq+b+j1ocWJchm42YKilkC
j6sMIq/hp6XbWrgQsILOzi+YJbFKm3Ad/yp0xC+u/PR5tsLRIZZiXN9TqM71mubo
99KGc/V8b5LecJy74WTHLJQ/uL5rM9Nj8o7VXyWwnVo0l2ucLyhwmr5oBiKIkTQ3
5oxbR1L5ScQgY0z582z65U3YKnss2nyjd8vQCAraqbCkAXDwlH68rrMU2rAxMI0I
JS0F2+9Tn/UAE3Znv4ITl0Bf5R6EDreXFuYfmqTWyYKIUmApylwLFR1QaorRm2ml
Mu4phLkVGSS5SuhqUoE25eL1tfwN4fVsgJZ5gf7J+30lrmI1TRr+14vmlxES2N+K
Gh3hOorK+YX2TF5lD53qHNLU4+XfE7/Mi/cdCwEkfejcdKENCxKmUKaFwtAayEJK
wO55oc90zDsFtknrbqS3ZLaxKbn6f/ad5a3vYWhbrW7F7fjuMiL9QI3sM73kc9/L
4gDRethZLjFdBG4C+PKQUBTBJwKBw8RzbSJFF+aTorQi2TS+yWDPOcIQ7EZgrP0w
wClYioLFYL1m+3UNiA7vkcjT/WgJ+P0F849k026ISkKIfUwBlc1FHdhY4BeIzT5w
PCbfKb30YBV99/4nXZMFWc8vPedLLwd5C1Gu+o4iMirQlnTkvUA2WEaO2TZByh8l
trMykzVi7TMCnZE2Ok7NsbIem+zC86ayOcJB3RZEpCgrg9b9qb1iCVA8ayRlYcqH
eCAGZywUT95iR40rOb7quMt+MSgXXYgqZRDh7GCQ0q49XdTQ+oA2c1LXoxigHJSh
UXzwWK+L1AbyviuuS8wXdVxl4zR0xRdZUJCQXrheWy1nwQ7OqY5WHc5uRbr/xIvV
kaM8DZkQVUGSKMhCt/7zTfk15d0jTA4ogUBtJ8tVIikFQOMBgRkd9YMZ/1FHKE0g
szwohcbu3HkRK4c8jkW9trwGzhYND53FQ9Ku7msES9XvjfGlWet2XDuAq0koBCtm
s6Ju74+yxtAD4DPaN1EuFkWD820Ck9QR2+cUh/+hh/PB4XyFq57Rydhulat7mLgp
E2+y6NNx3grLUmGFhI36WzSr9O7TosOeINhhSDzrvDV17/2sAJB6lQOSgGosnedR
lVlK+vk/B77v6ddUommvqO0Mz8gvno1dXSNoOjvDGtgw7j6JZZdkgclWkj9LqZnS
u0HbcOPT2VpxBVT0jVA35lx5X+jv2ktnfurH7mTp1lu/FFDyujamBHJz34kJKPTk
sXYyPrKoPTREixkpKkHz6ISPVjDaXN/WFeCFpSGwLMsn58w49Yj7tar3Cp0wIh03
UAhl3rJLUq9n256I0/KhM66YvcatMpMN3WLRUBldGUYPJ3P+LfSwyFy0p3g1spK9
pYY0BdBNe9rMJgknWNy14z4tiyQMpxzm021LO9Mn6UtzbtgdF2mUFGOTXC8ThIvv
eNT9cBaznava5Q0clicaiBVXor21LgS7gF6wnKmxinh5xeEJnirwd/P1TDandAw3
VKRss3qEL4HSESLcxiQcQNGmHY8svo4N1XyGSBKVdq5NCpoYAHVl3XASdwPkW/Rd
n6tYLa3WuPdusuDT/wT5PAl723AzurMrAzZLsSKWs33CCMmOV0SoSSfr/cHKpiR+
Sfl1sUKLrHVsiQtYAN3dEXvVhOu/PSakKLLpcqOEOHILRzubYem+51hus3cyTVPA
UpsBWyX2xtpThKVJrpIeov/83ayl+2oSOAZSabV3oT7nOLC4tvKDtwjm0E/eauAP
0KsiiSXDHzKJb7kjDxViPfeda76OyVHaOw1t/toqPyvTBWXVnDQNAzGBWUgwrssb
9Kwn5YVBAaHWSzYbCnEgBsVNPoh8j+P/jOth4GvN5p6qIYduNg3HAftAeletjIMA
YZ46A5Zk/dCqS7thddb76BgDNdWru5etsCyDQyuwCtSlLSotnEsXSZhOuP3khxqK
IHauN71P+Ty8tt6kdxDJBi3aaErmBhbPAKmAkG9tPFglax5ITBsKLMstMWBabnjH
op4gkD2WSSWYJE4AL7BNvWaBybIu5erFpJKZR/3Upq4AdBi1fcaNKi6bOx5wNOZT
cdsVtI3GKsonn+AfZqFcddZRJQbojgRrKNzjM0swiW1T06NZk/LHVQ47Tdrda8V3
ijkdPcPCBXi4GMGSeS82jB+G7p8DfUqGSca/qh8A+YYUDa5qrVVLQqMzen1nk8Tl
vCq7Y79RLTbKrR8zremKYRIJT3rSqLXwJcXM89cbyPpqiQlyLGQZU1lh1BqqxDiX
CE/+L7u3/gQC4ZWxZZQ3l/pe7lwRV1gyFI3oLN3moUWIeK+aDnhNBrt2equdijjL
wQmUQZylJJETabMt+2pE+BFO4YkMClbvAf84NiwcDSk1tLLT0rArUwlUJTg70njy
SX1tOES8KQ9dw7KX6FrgJzC3bpEsegMC00cXrGSC+8eoW2T+OLllMz/v1fKwV3lj
v6xPnl0y9Hhgvwwm1p3xGPNVaSUXgUji/+Ybb/Lh0Azm0QHkAkiVMcctRy0JmdeP
Es1L9IiruM7NwLzLAz4o75IK/N/yb91CtoldWqZJ1/jlfTo+uTxMUeo7QMgEr7+k
KKRpUjV5KwgtUeMxNvni+PqB/klPa2XEHKXUNlAChHWv83CjboL7TVkgIgDM+wh6
TmQy9e8ZGraJlAdMuTkN072Yvg2rwtbWG4bWpOW1lfIowo4ipyBV86bmHVP+Xsn6
1La13At2aUltQ+C8pHfFnGhcs7xNkd+q60gRF5FEQW8ekpfu8z/3cj8LRskCsjM/
P1W9KnIG762SBIKqElmM2ba6ZdnzNgTt2dJf/vGwOYIuQ3mSru/1487AidoN1tMd
8CdYJ16pbdQwehkMGKoRPT9gquwEy3dhPrXbBGVJa0cUoyUoJgk/pU9TzbJPf31x
anK4p+aturLccRwyuaY+rouKNv7+aJtCT27M7bJ5cg5CBlxvYmiSIHUiaEr0F6Du
kxk3h5QrhadtA6dbsHvIUUT5EUBkk82G09EDhdEm+a0dmB3EygQvSokqqwkua7O/
UH6uk5h3plKvgD6R5VPPU/JbVv33h2D8uiP3vfGN3QA+C50qRnsGDXlaD3bzTH3M
uZIHQNBqpLxdDZBvYwuJBlpbwgwXZIr0TI4K5kHxFiDwx/R+QgU4nmmZMBG9P5Je
80q2xq+ytUYQJH6tluJb/gOFG+7/MjfwQLKIHlJzMXlT2mjVOOeJrx+MAffrPqPl
p8ZuXF4MNQZ3cPgyWAIKzPxHGHHESqSvmdAljdgkzsENcfB6z6iQAiO5B3JGrqwi
Rcke9iC3Qh2FUBjI0oBIIX87arxVePimTDQRzCK39GxfT/RO9WIzlGRsWlDvIrOJ
PrLy8L3nWS3gzr6HmFWk3+If50DJE3DWcCLp3+dy74IhCjiP+NEBPWdFvDkHZ7XD
IQkoZCpx3uof+JdJzMXmZEEIxENKk8j//4OUCikING0Liyr+iSCrMfuicMw2HhNZ
hUsfjlu/m3HzrYnwMGIS1TRvLBXztdNRXksP9yBYNuPZevvKIAPznoetr6mP9JSS
0Gqxoq0c6ORjqsdGK0fK+eDc1bAJlDS7aQlfXP2+JGj+MI70UT8n8l/P/WjIXgsD
vFRspIxW152oeQX0Px1TEov1XNFkpWBNRdWpAkyfZrodV0z0pEqDLxc5spjWxfOx
`protect END_PROTECTED
