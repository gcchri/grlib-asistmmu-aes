`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eU5xpx+NO4sJy43tB5y7jRV809JkT9jXH9j0HewczWVq3Q6HSvKvmEKw5p7Q7Wwg
aQiwiXiXqZSiSmINFnhWRjvOHchgfzyclx4OedPFgIf4CAPTbXMAy/8ONDJDvAdn
7WZSLEbcL1VXoLWDJHDVMBfqfy95Ycw3yH/pUcfRrTXmbua2LEuFYMcEAu9lg05Z
PQMsSI3/A5Wh3d4+WToAo2sEOsZ562zmizgDg1swDYFPmPSe0bplTjHOp8+AFxUn
lEPKAUwXhFQC0nkH/Ha046UXW8QFxNfid0fW+iL5+nwZeX/ZmVHwL2AYl1Moko6P
FagFR1Yl80DKZoufy7hzRqt77LbX4GuE3T+U4kYrvrLOgqceZl6lAcOvAzu46B1/
CZ8HJVK7nBAQKi6yxlON+cnlr/Y6I7kE93JRPpB/ZkXKdUm4SZnOTCjedA698GWr
rCwd9k2FNSNFG5eiaQ0ILwdK1JmkvGLQf5WZwVrJzzV/yQo7yidHP3YxytYPkWTl
MWwPbggvzl0ZDJbCUHn4XWr/P11FYBZGzQe4tniDrB4Zs4xfOpqWmkg8aH2wjAkx
r3wC6IL43uUYSlqyV8Ma30N77Tx9lSbblpPFw/blZll43PJrdLjlzLrLi9gpMCtd
p7dJdazI5PzHI/NYckMgNEB/S2jNQU/VfzzJJ1K41OZni38a/j4V6+ChUmqiw8EA
0cWpbUW9beeWUDTZ+GxSIx40mAsmDRUGA9hFqJDOAYu5iotLa3Dk6dVP7pEXGLGY
5RViEhsSeIUVvS4vHnN3W/sEGDOlcdFpgR865FPrn7f9FTpHY0buJ5QVVw2/RixC
NNNb07vial9FBPnxgwvrn2jGWN+Clb0pl89tpk042+DVyR5/s1nUS6eJ9DEy+PG9
HCO2tsZUzwRrYyht8+3TTFg4W2G1NIHfnqA9IxmF4Xd5LHBk+YAG1hTWJ34g8Fyo
LkC5X2GMyEpXrGMRni8cukOIyl+nz2/VlfVQ3PPN5btEUjxZUoOu1+xXTrnKiGzs
YUiIDprzZZvs0T3P7K8vxJE/MftuQcomf73syV+CrSRKq7pOZKFM3WhdTHR+i4yc
w9u8NOgXkYCUpXfjSIrY7tWTXAYloO2QrIh+uJ3w4tPcK7e6xCKsBPHYDTmZUUSZ
yNxnkiM5ji5Eb3Nc3gWL7UL9rqcuUP4W0wLfNR2PFSpPJQVonpRRGI/Sz8hYnYRM
H6FpzJxGkg2uGAfLRwjePGrmjGHAXc1JwTLLc61UbJjBIN8t3Vp+SNBlIr3GPm7G
hxzjtrqqRI3ieVGu9LyO3w6URmmMiMYD/x/uxdXk4idUplFOwmpJA6Bho8WZUp+j
9oXqdXMc7DN8TBfTSg06zn+Qlf9Wxs+lruhGOpX11nY9Bpni7fUd++06HF1Whhd1
iAVNJROhYv5QUPCoihVGyBTbHPI17PitkEO6JeNQNuMCAb4Ook5MNhN86zPZq8Tc
rzor13Sj7JDCzdvJQ1GHeli/gABOITw4KWDTQLQDJq9/GdkeZEWsLSopaVek8YtI
plyOcS24gqfJ5/hsYG1rK0+yGMhyBOibXnqQmc7csD9EZj1AvlVRnZPnKqYujOQO
7fX2sCmnPyf4SsgGohx0riDMuHlAEd+9POgNHmm6rZeRHgSHEqLDfRs8JCNfLX0K
eOn702aR6tMMc8gJ2JCpzMqXswEaYwubenKYCl1JwPf4g5Q3KXBFQJxeXi9v1Glq
swO7mbLdbc7BlVSM54QSHnyHbHI7c6ecGxZinXAI9TdEtb+qP5fYJAlqcL6VldjA
WgJTKrWhRMUNFpc5gW9NaFBEmM7LHr6X9awt2MTKMQPEOINCjm71aVFKEnMJ8NzI
VXY16t7lru6d9HKh9ThkRqldyv97Zs/RBbydoGVO6ZfgyDzCGhiuuPyqegOR4qxr
hKFfOBeSjTuT9XTA5d3eqT9JD8nmZG6gFDGsbIIn12jb+hxrnjPwlYpOGNR5iStR
BwCgtBeC123Q2yGTVfgEbQEoU/aykhI+FybFfIPI2J8C0ZxcRUQUag4kOFiBCy99
jTW0mAIbhilWiid5WmuvHWDXiCe3yPKzKym6zVeYBxI1PBI1nPNN/mYGhHs+prNm
YwOBj0327z1Oei+8a8Vua3EaiG2xal7k50Wfn5Y4lxNpRlV6slVmob1OyLoK/Qa1
WDzqknZGSOYcQDn4ETIJAUDPPPm+2pHGoZZmkvVshdjaRnyMXgrIkHIdsrFvJpv/
PxN6ksL66RR6BdFFirRAHqDgHrDhIzv9MWAVzaVyup4PtWgl4cPca/TcrS1V7hME
TxQbSwBEPbNGmvb6lWkETNG1vJLgzhTt909g9Fjyqc4Uf1FNzOC6AikconutvPFI
oZtQt+KHCOxshN2La+zxCtalFNRkupWRxFS/ZIuI0ftJM2OsuXM2wzKEoAtIp6Mf
J/BJ2qfDDFCrxTehWsKOuaVset3zUBIJZPTjtYg17oh2a10gcyXT1GneneuJYveJ
P5OxsyOrENGcSuyCvz9iMEXpe06/oHcHgew7WBvKLe76TS+m4z2Ah/oadY5Y9qCi
4VERiGTLK3Z6ktIKFSy1lBWh0qERVjluSIzPaK1R4I55yz98iSNQ5jLVRWpWc8H1
0fooFyNTtMJPXzQac+0InqzDIs79Kc+6R9J5IQwG72qGSs3wDepOvkokiKvdnfuD
/pHPQniaXNqjCbbmXmzkQI8dfo5Rtu+dsEJeIoJEgtPr5yqGdjliRtEazFThdKGY
qMndcV+mOFTZcnQqEixiWhOMgLMFEsnSGHAcOoSWcwH6WEKN9R4V+q7D4PROPgLr
H79oryXKNGbif/ARkR4/GyfMFwFTffTgBARjMs4IUjg050+NYgzgh5zi18tRkJjI
q/8kPIKsfi330C13sc+IKupp9LQO8E4KRtNAnLez2UO9WEA3OAOE9F+wl/BqHMQ6
L8XhyGuK/iD9Qvdjpgc0IF81iU64ESMAXUXasEqEIZsw/Iqgz/6tG0Kok7DkIeEK
OZWYChbG6Ps/ix4emO8J9LN29WwnH4TKSyi+oX/MSVf6/oAKNPgE8JDSB1wJzVmE
MPwLAXkLDb3stjAq9tS2RvrPM/6Pu/c9kSEp056TV4e56oDJkl1hQ5DcybB7BUHC
EdoV7GRuscuS8TgYOW0COq8dx5aYVi/oyBOFG23Y1BBWgH8PYR70zTsLG+FEihJN
Zl8xVAkjXShu5tXhRHWcLGBTHPRhsl9mZ2A6GV7v4l0nZIxF4N+NdtiSZG98b+S3
TOfz8qfy5ep+ITDs+QKVeeJtKE5eb4Fj4DxnzouJ7k3bm70FvycKaTneVhxBwnbW
o+Er80J8I+UNOg6C/ETW/g==
`protect END_PROTECTED
