`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IiWjB2Yl863KPZ2qPrdQix5qkfahLqnbSqk5bJzND/AMjeF/W3fXTQ768CiEZo0U
436Q06SEkL4kmg8/zHPXvFQKXqTjqKvoSroUXtl+F8noGqEL0qRbi96qFiKRQMpf
XQRhGqckNnYTEcdVWiYPyxTIYP2ycPgWicHIqb+iGw77LF5gp2x03ETU+yn7ttxC
8t2u5gqG0A7Zhhsg0a023z8NCEwjTBedMj8tRgEEZxzXpBs2F7LDm6xHQ63SFEj3
tGfGk7x4BSlSGdxehD/Ilvr7xr7qeuQoCcnm5x0Cw7PJZktCrBFIlBSiNJbniFqZ
S7cvIuytGxxchOOf06VZUeTGUlptR/+VHG9ju9aTb4KQryc11JK0sdcR1/1kSgkh
SRmmSDzRNrW0702rFaG9dQ3pxdtV3fl9O5G6sr8F2QGri6wF4SmLmjuwBtL2qx3T
fTaGHNRzKuHrRWKXZjjVDnE/rax7mOPrVOKGpATL5PWTPYHbGaWs7XrIrMlcBi7i
p9TjABAkeJNoF7f76S/TEPTpgUERuz58XzYxt+oXXl81rs3JOXH3rez0jjFb3SZL
yHI7SFdgkDoHKjopasNZr5X8fD7Va7BSAzMqQS3u9brmvsna0WvD1x5OdtHCpK0X
9H2BpH6R8r3GDMz2UDn0R8yeAObWpG9eQ89N3puW1383MVJ2syIzASPmrEiJzr+D
Z+G54v+2+p6uyOwv+7IpuLxSmEqsy1fJViGwNWQa+hr680eScpWKv6vOjvVWTETt
`protect END_PROTECTED
