`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1K0eWlNPggb7HMa2C2QeBKUS8v8qe2IFs2ngvkwwtsua3D2RxpldgT+0YDS6+oG7
UB3PMCglpa/+OO/lA5hCBSEcYJMU2dN0rO4xFI/1yZ1R5ZViSHCIo2EqXH0tNg/C
g4M5VlcOIjGS9iof96IXSEoqobJZ1n3d3bhGh4v3ObSi9+ZB76COpTtLFzMr2CSs
wK/aQmAJB3o5Y09pBxvGCCQlLnPOqMUMCttemHpPLxJb6J6PPVpBtDLhWCa3Zc2/
h9YxBD4yPTLziNlDKj8q0SSsPJ7/qqVQJWL2FCjdEdemrS7SwjGs0tu/4RjDdRI3
yckdemlJgdP6gMBsr03EPdh1NXe8VNc3RYVi2cEyJrjkkqlUDiiJY0LZTQ4d7/kZ
KpL++f4ljWLN59pgvIWGIONrpaj5h2ABRrON3Ck0/vBPKSmX4mhR2O+lF+zUcQro
/v/4KXotETFP6e1nkZ5LcdAz26VkeuQe7u4uWSuvYKDNZQtRVGa3U2AMDrGe3r50
SmXVotfRrmmtW+1ox14Tw+0se2aAQpIFGWZOJyjep7wlLuoYblI+94hiwfMXlkY3
JPfpQon/1QgHdWVIhNCqabdDmDr8JCGiAfNh+IfpFPt2qos4stCk+rlxfX1QKCqu
l/wJn0sWhWdz7FnlmG+NlS4uIPrzBAnKD79C73U/LQuIJC7XY68cb35OhdeOi2uq
6mTEHtij119JmFYmqwJmTrl9oykHdUoIzrUy5YygQO37YnGGpblUW44VsBUAlroB
io49EQxn1Wrv0R855Cfydq4b7ZZzTc/BzmK8PUctuZ55JNZxk16DxRFwje3k0hg/
A1sdHKcBlflkLnI8+iLSyXtN4rvt0OMdtFK0hCecAbfXmkrCGozk4Ocfol85vyWd
H4FNGyVD8Eu5ZzDGy34Taz1hA0hYF0XgO+G4fezBRO1doWt4R9m+OfCRQU9hg+V+
90bLoo78WUwDb0AMBlTO1/fSJ5dQpBKo8h4QEi2WoCO+h7SOK3cDS0hEOZCNfjqw
Jahb0gIX+hGPhjFFWopvR4e9OC7YIabMDEd7em5NAoEBaNo893QC7Xj+c7eoH0Cm
4kaDmM28yr00JolF3+oqEkPw8HK2NXcW/3umPonAMipE0nEG12QVMyHOqw8nb6Kz
DDKhpbxuDjYiOE43astJ5xpTihY6f/ep+6t40UU/311egig6nO/PwPhtzkOKBeGy
I8r9H+3Y3FsvLTtGXCHdidG+Mb2A8VqnGKTslfbZrpPJF1CojYLE8y7uwfQHZu0x
jh0maKfY7blXzMrrwPS17j3t+kstPNtF6JNngZcYn2OR37RvCSUWVH7CL2zLJadz
9aTWkT7S2vhqoBUtQn/OM3oUd8ncOBIo7jK8TvtH6eUyNm1+EVvpLK/OFSILO7IM
Z7HR+8oDZwApoz5ZJw+7UNTf+evc6zJtJz+D75reNlGBMsaWE+TB/AsUeqhT/Wz7
XjUc4QvPyDy3SgMkN2tzXSfUi+JbZDEG+Zhbn0lU2SpiKInqxcDSxmJM+jGoT0lK
t8BxrY/p7l7ohAalgxs5MUu869y3le1CHUw1C8yBslDab4WEFSrx52GCh0XkW514
RC4QPiXJhtexAvmg7ScEDDY4h4SFo4J9Ipdb+i6SZiuVlPamihB6dZM8bVR4rxwp
2o0lRwZUnbHdlmheQOPWaED9Ppx8bFFQXN49FuAJC6hdiFUlGHROUtavSJcYxErn
ZKmdv8E3V0nTkSSrfoehJg1jy5+OrfKNG6Y4eFmsTv36l4mvsGcNuZ1k7wIV9KaO
lvxq9l4Ljhm3cj41Ns031Rhs32HPaNa7MY7MiSWdnIsXKqFoAx5aPdAIiRKMc6UD
+ZiBbIzBstMOIXC6jaTHX4d49MX/1saJlZJpG4/N+sZYHTAm/uvTW+AOpr35CUUa
hC+PjLxkR1A9vSTd7rwRENGbSq0eMue6jpdnX2uosmRrJ3tdGUx9uM0NlGbXdWUJ
aGfm1iREOadi6gSZ2kUB0fikes5+x8v19bd+wT60CCQDHHLWJ7bOicKdTFEw+aZN
poN8y0aos6x2rek8Tx4/qT51FZ1OTb5F7l5YhrTjRh6i0ZlHB4tYIH/XgQfOLuiu
dWpju6k/p6O+iTKJ+qP3rfdiBq0wFt0+STEa2uWipLj2QSppiflO7AetJNuWwxWZ
EumXm4L+krDz3HvxanDa4axqAtSBc77vH/Kk49Arfa0LSI+VKyNqkT7MbbqQk9n9
AgUMX3iun1oBGfIHpySwolMloEqzGVMn8V7oUFHkP+rYWNf49tE2wokWe5IYtcFt
A5Oh0zXARhmGNv/kzb4u56UidHm2eB5buE6JIRoWaicTncRot8YgGbpdCXFoEgED
/PkYSXj4jkaOdtbZL8KAdKfy8kKgiBP7amYRvA3wkeY+3OLkodWoBVoHCiKYmb2R
n1r5liBPz9zP6HhLk+tMcarHlhidPu3dqggLxCz65TfKtrazM5nkIcC+Ht+1/H8z
uU7yfbnrO0UOCkG8pOYWelYWP6Xp4OoRfTcmWYy/3mWcMJKJ0TalxTnBkfE10vum
Kq7LDtlxOmsQ0v2uionUXBWiEeJc5CIiejpUpqAhWdVWtxPU/L0gCyOyHOPpa+Ay
CPYIAzNAtCe0zrXEkvRMw8FR/9/kYIEQrESy9TJo7uSvMjNzRyHkY+eC3qoTddeF
nhxoFeGfk6U0iaHr08GhhnMlZaPbq2x5nVmCi+nno2krEI362fk/rHffRrRF/bxY
HrqwE6JXb0MnzNfhQJHOMF5RFSY3rVDbjlQk7EjBMisSxYGLKYfEmuSxOHUWbeeV
MQj9KmovwKN2UeWWOLITEJeaCqfA8B6AwUEjdQUz7We8IkB2yRgoIgnhX0gOoqZN
9kYhYjHfSqNg8Sk1XfzOzBmt4psVJMruGUhgFfHzlyc4nUJQoFIvXlJlIxruSHAt
ofaQ7cGRhVR00B73D7jsd1MsrJiNWvLXbIw/QxXn04b3+TiCG96zN9mt+tX4Rphz
i7wwvLCBXD1O4bhGXQDjC/21D12Ht88Ibweb/Mg5QxwV03Bfy2es4KK8fTGLjt3h
a82jpikCUBB+B4gSbjlLNSk+Z/FAJ1WfecMnpqVpKpyEp+Xit8a9arGOnHI489CQ
5przSh35QRY9r0cuFmBhOaNjp1ZdZ8e0Q22Zfe9CsFKFQ1zFmNTo2dsquNyYiPGR
UMmbfusOvN9gJmd9SF4hWnvtknHFe5K2hjD5Jo7YYMGof5CQZyFabxKjNuEhXKCq
1PyOTg/9teOmOa5iqnLC5QQlMNtYnLtbMrWFDogg33geaxA4S4PNrISr/az9FNlY
epap7klJNHY3N9e4HKp2gM48RAlA1A9rHwZhgJHy857PjpYZQMSNX4/tZ5oAQYxi
BqImCFXP0fq/5Hp0HZwZK6YEvRu6BqlbsVCJ9SSdwWDbG32p5L51nLw06W5L0abt
5VNOqurSAsgRx5gA5sT6vUS2/Vp3AlIjY9ojjwO3XjlP6Osl/lLuF/MWlNrdwe92
7fjI9dXOO/uEOAzzC1OcDkndg861az78l+5XL88Ymq8QXv8sp39CSbz5BkiXKGCV
J5HI1TEVWYVnBq/5z2g8LioV7sWmOslB+iXabmqy0hE4dJU2NtycmJbLzsfpaBnI
2wTJYSlJzLMmdisNAATMQSbx8rvovDygVr+7kSC091w8qbHzvMCkAISXIqTrhbzv
ppQNsECApfxMB/d1SBHQtQke0m2aOdZjy7+EyD8ILcZTvCmd1S/CG7WIxVj1RIJx
5MefTqvwcUPCARmmvd7XdKGZwZUmI89aeIH0tOcFB5pLvDzwAVnte6tOGTBubzed
6zFLczvwyhDF6n8u28v9y53gGmqYKCyzI41Xc5Gn5SOo/ggrj9g3wBNaSWxkx8G5
/hoRkfhdYYHMlHn3jhLc3k8OUAPhOkOvwckAw0kGgT4lPV0/QBICdqI5Ke2wq8oL
m6RHhyhlyYfBA7WkevIYnIcDTHmk6u6+gRSeYVCknD3Qsw9CTrNzNuGKEQbFxNXb
1BBFkVaxWjN+GYTycuv1RakIX/Ec7IrYFsJ+QwSNEm0EzeQ2VR2LBi7elQLYA0Ve
lbVcg+wXJeJ6gMzCWAvHSob07PUmeVTUTxqYrkm23Tq/j3zY4ijKsZSQwvjNkX9W
1JgnjPQAG4wCFvAc4Ik9fiG8Dc2xnBm1jYPSS1HlReKS5ZwLgduK9WiZUF0DZ6vY
wr5HjzIDnZlpLJODJj/JynSE8jJPcouL73QQjw/WOwsMtQDv/flSPtKB2y+JXYKB
AQbtk+ZPO9fT3+zsVTeWn/nOv5tWEp8twmvNJi9dJY2fL3ePxlG1BRe3xqNbeFlZ
WF+3E2+N6GCd9cFCOyLLLQmMaeo03WT4ElmO8Em7KzUYY2+ESjxeUbyjybIWvShH
cinrZmaCHWsK3yoHZC83vXJQpoR/MCHy3Ei/FL9eQ7zr2FuN2BrdhEexbdPp2wEH
XqkHl57hEvHfALEUPKXEfKLBliSnaglwMsBbMGpybmE9TUoRcwLy/cg3xbxfWPAs
OpJAm9ku5Jsu//5iCVZTqmKzgBZGxo/QuwYiXaXO8duZGQsXtLIyreMeoVNPN/uP
2cTA3OxXFmEHH0OoRrn/ub34vxHS/wx2MZGss9poGtZxmfoEkIF9aOmAKFCLIuSy
3f0TAqzJv+jfyPTEyy+zfIFfT0WltQODszyhWEqHycH6hMOHb0oO3lgUDtWCs4iy
TbpMz/gwZbFW9TgqBQSxXQ2dEJVw520Br8TFBQZRxU0HmfjRjcO2qmg/F7+L43CZ
Ap3ioe9/fLNr0NbpCg+iA+uMRemzCoNj+tYcA9r1pJKpi7wMIWj71XWzHlZL9FBK
RL1oWetSuwuxs5+c3AgI3lDlpnEwcKjPOjJgwYePaqKSwmXfO+sJXZByb3xPrt4U
CImQuM0AVnFGvqOcOiqkve/PmA0tXCeM4NqDDtAdHG5Ic4mCRJfO3udJxoIdvXuw
+W4uPftieKL3KFK0TVtCYnGKg6GxoEriMGoSrtTtnesq1KVSXsUgVQjITg/A7ZlB
OoGmy3y3uU+U8fm4sJ7smNAFXy24oUVfnIJXh3Jwc+vnxe89shGV5CbAMWqhNqqk
zOnrADobkMimUkvjzsb/PZRaHMfEN8JNle2eSH5CmenqOqtmYrI3oiGnogUZGdrY
s8kR9P8sUaFHKotXuYWGbzyS/RYeLZirG7rm444WcPgGRKCrfiGOiFqj0+FnjdkZ
Q3hZrM0/0W2lI/VX8UVACuRZDDIDBQfU0R+9f6Q5aGbf//FMD8fDEMHAuAm9gGLk
BJCJGTUMCjP3EOZgHxT0lYr64Vz0yAnx5cvevlm/5n4Zvu7FSCjG9OvPsbD34Wdg
vHLRgruWAXYWGyIue/HlOFsScs4Al/vG6jAZDbCF3XmXIHSVuGth1kkjwzalB1+R
Csa4w3FLu6r39Xe9lF9udlFIc63RdreOQpcFIv7kYkyxVbcokwxNxwSHzUG1D/ac
2T08OdrW7148P33p1Taq7iJc7Z9D9uXRbgt1ESGsuSYLP3wbJpzL5aWW2HUXNFZN
nR2y0eimuNMrzOMFYeg8cWRmy1AAJ8G+6xYa0QU+y9WbO9e4vkahD4a6hMVCVuZ1
92ykMsEjuR8K4mUNhOQwsL0OAMLJGxA4e+9xj8k3pa778V3CboMlmgXFUVxzabWo
o8Rs48QhgJHpZd+0oQysoQE/PAB8Bcl42j59FeGoCptSBgKBvHPjbDUKSJ0KC3h9
`protect END_PROTECTED
