`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XeDqmG5RfYZYausg8cE47IB3VFTOZd7fT+TMkbngKSsjgxQZKbBIslgwfZEphvFz
KozufgQWm042kDfNl/e0RVnV267oMh4SYn5Mdgdsa0Q2IwCJCaHFpxNdIlJrdt8T
OCVBk3IskKNfbocJotUTjb2iAUFX5zHBb8H4whJL0bHH63hw5n2RpRxZ0U0ogMFt
iK+Cbv8BhDv6wwN1b4njHearavP1PJuwYKvRBIDa3E/9tKBhVK1c7aHT0wHgf9FF
1ZBsJEKx5F2Gi3Mjy26w5Q+9/lYxli3tb8WUyjS9xVH5SQPhr6oAPXlCKBDLjW+u
Aoh8GgT23HRA7OkSmumq6gwkdYfZqF86uRoJ/afs95C+y1mBzg9HDIIHnyNNUB1K
PDdkyBiOjyZOYKLARTNblw==
`protect END_PROTECTED
