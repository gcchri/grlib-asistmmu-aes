`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DBg6QFtljK1dFQxCFRhSH7vO8QVPVPyODl9Y83DbfdnernuktglXvP+iv1foSsFR
C7xdO7zERw4U2JHnTycIU4HePcO7k3+bi3I6D7zptEJT/iaw4osGN34M7N1LWe8W
NG7lQfmf5YGViOAocLmip60dskHK9busSCmhlEJvNNqooVeVinPmUyIV2X7VbAh6
n5OHLMzCXLf7bxarX8FTbBNyrCPjtdpTxT8L31vYrXyuMggHA9HDiWxLzxi4lSz/
QAxZkX995SR/42jHEvAhufFGXv2k7MQ8wcs1+KvY8wERRJVYvcXT1DIsrcvXcLHz
o24vHrYt/boccU+xt3edXYSS/zxzZ6kfTwvuQB6jeMRTiptrrX08zxGCylEPnkmG
bOPsubfGd8yRK0W9kXnv4DJMiUcDJ7Bc0XcJuiG11Ts25T5uDox4Svn3fbcSYWNS
7sQLi0FXQUAkQ26PmRaqeeS8/Zhv3e8Z47mGnmQ8WuaT95NcbViJM7lRQKI+18tj
1v6k3YJfQUrpAsweCIqTKpCfGsK3nXj6YVr3rVHo8jC/3SHqM1GUZXJOo5d/ct8P
KWcATCWKDK74QxnxV06owLzgHxUtWfYIQz5ssfdlluoGOCw+UbBsEp0yjRYda+mA
GUNkWMGoYTrWyaowRRnwTu3WJmBrch+MTCgasiy8i3q+LB3DWe2Y+048rR7/VVJh
32EcVCg2QoYm/POWdwGW+Hsuz/hp+ihkQQPk+sHuWw8JZSkawWuO3qaiTkrbMrqi
HySdx1CAAkCXr7QPBzCFPE/N6EpMlmEgXlWrTRwTrzgKomGKCzOT7VJ3y0JMC1zd
k1BbqPnUf6P1zW899RpeM348gPo4bbBIdKFdEZOX59slCZx+b0DdV7PwwtBGegaL
SKO5py1KdljebeMbccCxCMCKbf/yl/c3XH7fhZZC4cZ97m7ROfumqJBYe+GsAxP/
xQ8PkAnosVzrYZ7VlDAjGqcYz2qlaTSLYQ/xJeEbnQGfQ4wNeOkajIfgeW40Mbgp
Yu0wQJVZVQkCLCySajt/lo/hPE07Udi/cXROKvFqfLuJCcVUCCHIMG+RJA3RGS5l
MvzxtDb1Szp37omxbUvtfvnDIDRKrre4PeFI2zukfupD19z1j4b4HHk3uvL1vRAC
CsghZk+4sGWNQ2of/ktLPCVmwupOF88QPCp7h/NxLKRc8KqiWFs0yzNMtDNhHx6C
y1MDJsqkzLtCnsoaxQVwP7oFXKyVHiAqQYScpXo+BP6hLw3c3UFRmCeNTGbF7EC1
dRknY78NHrWxPhJAai56DIRJ0bqB4OpfcO9i/tTvJZVFbZj+7jrctoFGL9bElvcV
3neg5AsaKGR9B7+gI9azQiXFxnB+P9LulOeSPKXUzQv5SiRJZKZiWbxyRBqRWloO
5iP7w4GoYOxhBpd+fveS/bSoQ+Nf+MQu1FkTFq51KABPRHQnSilAE60MJwZPCPfw
FPBahqSTxW3d2NU7Yb3zxZNsQDUPA+AG1os1oe6cByPsaXD7QeT9ymiiHL/ojyr8
a3vicbjFPdIPVfQbbhAlFZ+/sulu4RE+74nde8qVOQefuLkNldNuhmJu/8JOflO/
FVkYRrpqtUFY0YS11PuqxtQUrHyz/+pDdMwfRwqgBlADdHPcAAkbIGnDXnSw/WUM
tzrT6sMWnrAa75nbtS4cDRJF2kr5qP/W5VduHPf2I1ooCB4bTg0AOM0ySsbumQRa
7s6PHdN5+jqXz7ZXqTtyyg==
`protect END_PROTECTED
