`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MpkMGNAxqzpDaqAZv9zv3j3luDllfWVb/zkKk1HAYHi4vK1RxuSKRd7fMCwo5Ine
nMBlJcSnBu8q1s3a73KHgzXSGiLQLFo/M+hdSqhjewjpXmOtfb9Zihsf9fnIGHBI
xwWCdwVJdPHv0BTjF8huvmBeKBKP5p+oSiKxUlntrnDoxQU5BlJKEyME/MauC0oh
8GMnlO0T7LjeLpjGEdG81fPkWe6Z1DwUgz5buc6xPYjQFgBPWievr+Syv9mjR20q
5ieKhy+psnudnSwGNEMZBP+fiZ27gyfRB2CVZmC0ERvux9TE0dJvjTqJNeFeLI/C
rJP96BDYvZG/6OENQ8MJ8VP/WqB1EadXG2NueS2G8hGZystwSLJnkFQpXS/J1EjU
ZjTD/fBoZiTt5VsgTsl64bB3uUxCIieYpPF4rV0QGtU9ENSfBvrQYn8tgbXQbeNQ
ct/IVjOca/m/34EBUCnlYhMm9WVYolr1OcXfAIOumU2yoAJxPrrtl7ib+Dz1HW5e
Q2aVSBBtlNyMrotg8LWf3vuqhDSojen8EK/V9qJeopLyqrtfRVzsfgsTZJTVWdJ7
myrRu9lDNEc48+5KkIZkEA+9xyGjH9MxRVTJBd+Ls1SUOUR0KB4ME/mN0ht20WGk
RbBK/BJ3zhwCnbZJs6jXc2Y+lQb8tCNwkthGZkhPLi1V1J8TTs+h8bjIO+QhxAr0
Q4BsFmYiH0emREI0hHY7lydClSrTaJg3e/dZ25pa+n43jhkc/GmIKoHEHnxvqYH4
BtvEvTrK81ylbkK+OChUJVbJ46YI305VGUz4yjsBwCG1SkwFLDoOgaq7qvAAO9Ug
vbSNMkBLwloCWHo1NGFqLQoBScN1zNxgWSI4vqLv+CiKjRuHlkX+Isfau65Pf5kx
1XoYw0dxV8q9kSa3Ck92599az5+uhFJZixeIZT09+U0TPcE5955QzwU8roVkcAHc
5f0SDfj7drTO339qkNla72z65rbwh3Prn0ldyphW96leVkGoEDc6DC2S8DMBWk1/
x4rZ/YmHxDHBiFz6+WdXkSUvFXRn2vmKjcmjykAVjkcLVeaPyiD0RGSCp1Th6iCo
d90tJcCk00Hv2Zb1nPvMTJtpafogi6Ag1ee5SOWnbi6GipMS1xivw6icvcrnU0qQ
4ih1mbAFKlVreDqwIAyZRzSEUWr3eKA96pFP4d2ukmrEjYVHEIHPntsW/VXSRB5E
JBD9SF58V47MFmLZKkG1nfg2FdkZbZyz2R9f2U/2aRi0Ougw/b5ljoV6rY8/nkxu
q1xSwcWXbrZY4x53opIXM0oEEJQgoQl6m86mx3bSBBJsmeFYpd9B3GFOwTKaBsCX
QwcbLtvDJaynDqwyBAgoMpwxPHdmnDMtoFG2+Jv4+NE5yM/CKaFnt6goQF7QOa+H
pE0IcN7kMe+9hwr24uCGBANCce0o7DkxSkdmeth3ihfhVZj4RcqfK82np3P0tqze
lRsUQQBgJIN7UW5SIq4VKvogEjsl5WNsjei9iscu8fUEDZ284P4iKcZFUVIWSVhC
hlwM1L4vscBWKe8wP0BllQ==
`protect END_PROTECTED
