`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wKh2d1I/lGmKAxWTksMDoqAjOtaRsZKjZeaonV8VoeI6lwdxUjGXHDRowH5VOEev
TN4r3RmrGhy9McrtxQCm0Ksi+NcXUVvXdv4EtCXUwtNt+DHFrIpEgoxV9CNdsgk6
EqCpIVo5EQLVU/5dHpgoRNMv5/fJxn3dwQQ0eWBPpa0JeILw5hqsCSRtBeBU0+uf
g1LhXArspaqCrFbx8+EQ1LGdWH4aepCtRVmyKaZStpL0F/c5cr340WeSiYpcn9ZY
6X4A4pYbu8f2FoHK/AU1sCBymk0JcK4Amt4a8VhZA1/MCEtUzU05Yid+mYItbn52
SGsmoiPqw59q5EeS//CL6chxn06jCGFjrub0TNfkNZv5Xh07NKOF3JTS64pzXWhv
cn8C0/RZLYlu6rNbzmLXK5uUnQ/UtVRgNOVs5UbQ4JLT+GOAlSFc2yoWQNtyniyI
VSRKbA7R0OBbUZbYa8OkuuGiN0TrqAjQnk5kNhIkGS/BiLtEHeUrq0KFnDItfhAw
o0TjJaHC/TmUXqawYTn5MqPj8bUCQ0EkqWT2/YCEpKKiGcifYdNtAKN0yk9iwJ8T
aWMzep0fzBqMDSNwraTwEkl5/FC/PDwu1+puGKd6jaFu8phS8mEBg5z/RVVnqH+I
wVTZwF3JXPwMadTzbqP6QPT6Bx4mv4fRo5MkkIIVlyfFIokedhhpXhD2y0dNuATx
qjesX6SSfsCsgR/DkC0B0I0VmUF3YAZAdtFJF9baoB1rYwGgvjINIO/ag9vVheMk
8OnXxDXHtxcoq3LkCsmxyktGcDTaYzB2xHdL5W4y18gDGS+0t66BAwQSoptYpvUT
OTQ3RGbXrn4178XkQ2KzoPrvz/vX+M54MCIfU2hLePPd1WnbX99tD+sEeCmr8tAS
5V05pw2mZIMMBy3DIgqJUG9ttq/0gTF13u6jJu23wKsn8os3xqzWVU8+CYfWSUZB
wGZ7RtK7L9fscMKnFXbc9DvwdvZveNVnTrP/cQZHyjc+KePT1MyyA5DVwq0BQKH1
kqehcwf7GmfPFczSTPrmduqRLYTerM5A2JglypVyksbhiEjzlflUuUuhIWf7qJ4g
du0UYATwKuk1ygRYjUIZ3mXRiJEFTJcq5+vMVBYfhpPYw92PB/YPXkbUNWZJx/nW
zEYumB0+UswV2aIKA3Vz+pt+dQNj9lX1cArRMeJ7G5AWFFF6Fo9A4PdAwuN68UlK
vuw2xt0obzvXYkcXUWKLvuof58AybeleYiCDSH9inGxoxspLAMUupWJheaAj/FAq
h3XJtcPu/E4tm6sJfjr5JQfKqJJNayl/qs/H5HLNaGjciPcWlbbOrc5OdNXM6uH+
JNKLtINFfnFY42bDJHniZUnU5sniYbP4oOimBCZM8N22cXHxzJukOPOKu7grV158
qUY/yKy+iB2OpqAxptMyAg==
`protect END_PROTECTED
