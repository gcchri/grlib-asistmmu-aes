`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lRmK2tpwBJh+mYezZaatu3/VAHtfPXsoanCTdSWEKGX94o+0ZmykheyVHLfXewUx
hGBONCTNjksBKpNIj90y207DcNl8PrCVTjwlg5bmWbk4xzc2L5YDqDD05Wr5txD+
akwgdiKErunYpfKZTDfxHwGlrvjSbfz0SbzsAIiX9PD0YcdizwD+ZxJsJ5gGaoUo
5yQ/HU65CqjniKNrlREu6IumlHQbRak1dDtPOR1gdb27wFogqrmWF+2ue/QGPzsl
UFi+S6dKUiXrP8JkJGFo25Ts8t43Bwc56jFb5ASYv9I1XUSLYaXr7MdxSgWoGNo+
DWJbk9oIJijLG9sk4TWDIWNih/J3ZAxJDJ+zkgZD1iXicD67kRIq1sDUmZDDP7hg
t5GzZqcQZ+5xgAjoTlpXEkVGQ32A2Y68l722mzbDMGpOq9+fc9FzD2y6xrwP4gi5
17Q11wragniPNHOhwE6bRA==
`protect END_PROTECTED
