`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2YjxZHZPgzOp4pteMNYHnzbwnrpSidyzOHT/SCzJqB46WVZOyk+ooOPgVifZIMJL
WVAFfP0Sk+MJFiHSkGCGHcluLXLBEVB5GZ5quqtqIgHkhSfd68bgBdcgGZzwLGW/
c3Na1ExOk2X6l5Uj2c8WC60XasibTzuqXn6QBelTPxMDcGpMHNTizKpXxUpuaDdb
3kAHzheOa1vPspo9A3YfQ46uG7KtNEuQB4VeYzxnNj+YFkriYphsD87ZtQfeFJ2Y
gtFP54WMULRHVTVktxaLFNfq6BruEodStSxXDSPbmjS61/OJDp6Bwf04QKfEqKwx
y1/Pt4dU7II2I52WDpaIQ64aTSpFcEwgcGMGYr3FVJ4HqarnjNOmvzGCMplV7PLG
h/Twsoa8BVUz8wprxsVE/VfplTgv6hZa4S9qZS13inA/oT/rq5T2i6pcvnpgb8pT
92xzlRUmI/BnFa6UYnvD/SciVq99BUSmsbActtBnxPNrlkrduRtPB64aQt/51lQ9
WJju1NYREhdM5p5vjEVzs6U2Z3E8xY/mfHW12ArPQyyEjZh6k2QfHHi0hrMq+oQz
LwgX5QKRMmGhZHvGmNs3/fiXxUodssIHQCooBSf/4E4TJBHx8+r0npWMmH/iz00Q
NYa6gpKYCLpxvS8pmecBhAj51tIQZoryD7bhA6exjqGcTFH7Bxd3YVJ3xe0DUA/w
2fzZYUm5o7HxkMCP9bmXYE3epkjttBlwe5cjbAP3MbrO7+WWYpC0VZc/aZLA4lFG
P9H0AgQ3DwzoWhWfJlEUJw==
`protect END_PROTECTED
