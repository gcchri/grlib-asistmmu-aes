`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
44k7HSE8oaIZXJAQoE0+y5508+8TVlxwAUFcyIgX9OmvO4iNyAKgyI8ZEdKY7mN7
xGBmOVfunCc2WL74iI8fpKfh9U3UjKlE/Dz5Jq4wFMuagxtgKIN20r65Sh7NRSyf
/bxL1pqMEkGfCNKirEkWU2Ev99hfrva1fj2EDeNoi2roSfYydG7yvtA61gBahSfZ
noRyx/A8msagZEajls2mfvSN6jbXTUdtGd5eia0jIHaSR/HBoIHjvIO6h3g300M2
QKIUefdsi8xf5Zv30ATwVRbGuzoV8ZfEECkkztfuFTK+eErtQWXPd1R+8CyZ2S+B
iftHefQSHJPC8B8dSPZclvZFSGMT6X+cis/66Xb1iYn6zx1G/Z7wLv5xei+ihvgD
/WeWO1g/R8tnIruiIy2NMn6WdXoHusb7AeZZr2oaX3KPEoFqJamb/hOzfVqlK53q
CUSFwM/mSbf/MXSWLmLUZW8Su/E/92Yw3d8Mva8NCt27tDeugeyx8rtnGa45Wc5L
7OZwGglVgdxhLLtWBAsrKVyEK5/n9xUUeV+MECuCKcPsNdxBd4TDoZl07Uyu7A50
snzDtbWK93b5IWUytBnfarjucTErIVp53hDj6W56+sBVHZGh5hhqIJYns1A5TB+e
hYh229eggEBtnr5NxJQ11A==
`protect END_PROTECTED
