`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bt7GI3Co62NofQ8zlA/LV5YCvT0jYMAnuETrjCjV91vcG9iXR6b7vWIR6CypyBwK
ftzvOcQw2Qqf2cucJCrMzl4OYovfmqpHfS6PkqlPqygDx5nBzS/aNhjH8R7/4Csk
BQ8enk7IfSU2uUKoy1jwqbOZIDR6vl71Q4DgHPi+oBBYeilPyvhCEGToGst3g0fe
0yopHeIuHG6IEkV9tyDMJ3vDzcIN+q2Ref1A2xD96tQQlQbM9PA3aj7oeV6oAoYn
GAPVh7HI6/GFLXdfi3xTZzkrwVULnLmMI/ZumF08n4fGeKbGJLNS5JEvAe0AfmoJ
`protect END_PROTECTED
