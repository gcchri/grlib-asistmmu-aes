`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lcUdPFe1vBp7rENxeb9IMVG1z5+3Yc9dvuWd/pgiJi3g4Z6E/rqiXbVT4UMOa3XD
keqlynGYiP+/6nPj6HteDDVVakINxvomNCpV59+Dqn3KOiaQjkBkjFsRKB9bfZsj
EM97n9DdpUPwFV6Qj0gpBjygOAddlwfzTFDhtiQbPNY18SUjokYQI4rFTh7mET0h
p/NOIzs+MMREIFZwiOJoXZ/yCJiJFKorzRNJBhDpXvRfMOoJrcJyjCxUvOjU/AQQ
TOmgrIWo08OPxYiFSL5Tca8CHIJHI0nV+9LZlbF13l/8LYVAFTDjM52WhkdNuBLf
lDCGV9Y9iOrRi23Ldmpk/UQJdD+YV3QpF/4W5PSXGNWQAEg0s1vIq/MJW+Y198g9
Ct5efSOXXCYXB3Kmo/MAxqfuj8gbi/q6VZtVOREmCQa86E46UHZSbe3FCZBfqENA
yej5mFpSK2pmzIQcXpp4uFnuEjKhlByy6ZNGzLc+VAKgB0Poq1YdpRMTCEws5ueD
MhgcetnlNUrgPSGe/MN3pTr/eiH4+AtLfKaolbuCznOKT0X3bQsur/cHRcRd7669
pFMyaQDzv0EwNDcGGkzfb+1lRwkyzOncnKlrR010TGmNc1iP0Ei5DKGvifwmlfJ6
BJv0Sro+hXdSOvu4pPvbkKIN+pC5gQZ+FYN83RE6FjACFee6naFv6DzRPWgEkJp/
qBBIwhN6g+F3D8QptACjagX0Qye1XOYR4wYAE+6DC9V/avjoCDReTakf1nMRNuAy
47IQfmHYbpVbk3+k5+D4bA==
`protect END_PROTECTED
