`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xGVn6f0jTssNve6AFoKxY1QGBDA9KNqs3y1HqIsbRcvX3outBNaUXV0XteH/i/EZ
NYxwCff5BpmAFQ49AsYsAFJ1DJJWYtmHro5+wkqkvrhkwl9C9gKHt7uQrzSbBbPQ
QcNXyuki7xLTkDgZkdlt13fSAJPjQyLutc0CiqHbVsYvgojEM+Ze94FT247/nba7
03TryDuhkCb9WuwdogRXo+TPMmv7aZPrUTxgUlw26RQrlKWk4v2nLyP06hP9H2Nf
xFvTBmKpSATkTMlXpI1jZcBokj3mJIXBaH6NzfvvYHc9KZ7Te1XigLh4E/C7sbcX
sopI0MsRQDVda5uWlmsVNlRJozKqTXyr2Ty5DHP9zu+V5jH5rlAdAOMhxmLhc6H+
N9CohUfMRscQCa10Tto1c6aQa4S4PFpNKCqwq1wcCEdMc80IwflkvVMjI+W1c2D8
X/9e81AYPMNK6rijYx5dDK/mKIv4kSlcXibALNt6ib4=
`protect END_PROTECTED
