`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DMOYiOlTsN0dZLqVuXYHaCsuT8GgYPVru9gJ+DMBuoTSt5XraHtjISDROhmlPUOW
/Uif33rRDtr6/jeifLRMDbnSzUCbODHhpM3iYaDuV6f64eS4b4Xp/go7ugYdiWmJ
htZBKKprRjPk3MVT4t6Fe+Gwn0twGHMfnlWKi02hLK0rBP2bmZUUwI+15OGInsiz
OOdHJvJx0BVBojTo2g6mW5bHJsbwWzLydOLQU6w1Zq5gXmvbOFm1UR2krtBJ5w0Q
TZ6N7BfYN0TdMc59hfTkTj1l98DIw+TGTZeEDYVA+OCC9S1xJROssAAXZpUmXc7N
ifpjZUhdxCTtPdPzYH/YK0+Ymiln6OGIJlAAt939V76ZrHO5vjbZI77t5p1DsDEY
qn9BPvVsbvaN0WGJBgvU1TanQLM3sHzdR0tMihgF3+IkFzjXKrwhuHrYmSSoQ8HX
yos9yq4mP65VvWt9OFOnqnTc8n+hZAbM3F/+1NuiA7HApaMwxvI+yyCG8X1cg5tg
DInkZKD0FOyCGvYdOOEAn8gfkLor4BIbrWWfRUBiSq5HGPxL6d42WC6MHXzT5Igg
rOQlEDpUm+NO9kFDPFSw3XG5WX3Ebkr2bjwQtsHSOud9dHZeoszi7Krko4w3pGNk
UywKJnaiSbJcARG7FG/mTg==
`protect END_PROTECTED
