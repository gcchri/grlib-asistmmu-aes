`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I73Ly+QEhhDDQWocf8/UHgcAtrrDEPh3kT01Qlv9HN1OaVfvrutFTy5S96sSyt1p
NMeINtgSi9OTEqkeshKgWlNSmWGYjSBgOn/7q1AsI5Ir+iSQL5sWeH5axd6oqaVg
Rj2/i1wUGrh8tFGpijTIfSKoTCxEHb+fGFwvXdwCcT0+ISO8YEBZ50r40w/neunI
lstknDPcIcbzPgWhUwfMXi72SgFNVgyw6aevPHFt9elg6Kn3V2YggHnTssV9XPuL
VJq/Wldfd/+MwlWHhKfrQXBR8HfHZA4XdL9XIF/oiV/8OUM3ysLygbZc7uDS6ZQ8
PPNoyCLN2h7rLmmAxQDhOUq9exM1U7953XrFKEuasCMJA3lZ8Tf8CpsLjutqHvQv
ZBK0CAbE2jOjJntiNFdeyTfCiW7PNsR4z4ORdKJcXq9X64sH5cEgwWszrT6bgObd
nopNS7WqHsdvbbO1gSQy9LkHGDXOyUeUo5ylot0GIjGyintGmnH1tzgkervQSDGb
ZOCaVd5HVkvMNLxaeW/9y70H/A+KRml7bXpMX129jRwFOsj7ZOuexXxqf3gYYdub
3hqBGCerQCbCBCCy9FKYd6eaufJxkD4SHcRVavpR/BaOXc6Su6/RqinB2GVOtbkV
KCcRRxiL2DpYIs7nx1Sl2eUKjDc1YrdyPTPP6Zl0KB6NME7azhtkynMb+mf2t+Gc
xoPwsq86Fbl+eXY8pF116b+vIK5GbVSZjo+bO+R6hxRa8gStMZt1VJGD0HbTWigY
f1A05cWDDxENORox2/viZv0ptY1KOBKgUhQf5lJYmgjG9/WJO3TBgO1pgFuHGcBi
t3JNMYZjkhg0wqS/E0iTSBE7pb2l8gNSim+aJ4RVjSqEJg2Uj088g8Q0JOBBerRy
rz8ObG1AmhsuE1Z2miYk5exAo1c+cRuwVz+oANNzX1PCo9hEUF2F8+aKLQ5OqJ8x
56bYgAWPFoQFMqQcFfNPgV8KwiLGMMC2EdKjH710aq3FbtPv4Dq6r6bzDpkGJRN8
F9wTv4rRBnYAvaQtcZRWoWi2dVxIrxpxIuYoP+c5QEJHWW0pwseUhoKyTXULhkC5
E2nMfEHkFjJxjSjTPWC+vBykaSxpg5zck6tPCrX8QSK39gXQARs+jRW+q18wMxyy
0WGBxa4u2v/lEWUjaXz7B/aMkkctLBhMVBmllAnlFCGmiv6dL7Ac5Dk3n5qZokI7
tCx3sbSt2TUEjLlzIa3rtNj4IKNqpSlU6/FpefzbSq6Fn+Pa9eGsaVKokmsefO7G
aYAD1p8PPpk2zF7uEDs8QlsRBjKfwBh8QyoeZU/H/MprtkJqzGv+Mu0I0RDzf90N
kmgPUSPu5qpkfOBMVjKusOUvkAy3bN6lDGbu3YuxvDxzVAEU73wdh/ZpBeR6bGZL
mSuinuq7OeX5JcLGwqWFczVFxKpAeAaQPoFPP5Bz6Jn2ETdoMqow9MlN0bQRKgaa
3KhmMcR6afCfxogwuh3ld1p07M/HBG8ifPeA7mfskpo/aTFfiP1f8GvGYzNnzZ7x
pAnXuykPN8atPNmpdU6xTDgdzG5gBDjG8J0HOnOWxUBrXpGfQieA8InNeNR6LpL2
8GcqEQYA2TKfqhFZbXabjj2HbVz05Ysxu+lkE15XZrNgayqhoo/AMA0MzFVwxqfC
/MtYWRy9nOrMlrmP9Pcyavj0uofQaCan5W5IIERpdHuSGYfQM6qMRQuDujsMdi8v
NemQoiyYdYsJRhreKyg0tHA2ovFl10MDaEMxx9p52DK8GivgNn761WFg1abQVMu/
VOfuUWYvO3wYP0fwlpxnJTZfBvmPmbTeKN316gNO+cKH0dj4W/eEtc/PGZP9s7GC
H/S21YKDUpCsP8KFG9N2c3xdxl+kNC1WaGq5NzsR0CPy+1ignirfQJr9j3Sz+HxU
mWYYJxDXcDHb3mrRPI16SjgBNcPdtyX0XfR5Gcn1T2KaSDhbBTThpZVjrUCNGg2j
uNx+IgItzcOceDTnzgrwrwCbz73EvJ4ElUotrWses2BKrLPzHbya61+mgFyPkqRQ
bs/AImoPulQnji1ff70fhCm+alEkwf3fzRS0O2910nTIwrlgwRp0IJjc89v/MOyu
9Qfed27/kn1rYfqvda9XRHkqiCDPw8G6hywWipSLwkzaYC51pRncId+vfX2LShH2
pO19is3dW8UrUBU0zgVWyFrrNSCPEVFFS7y8SX7sFfZS8r/95+QlwB03BqUGzaq8
36lMzqxrRwj5Ie6cvFT1XhR9nJCgQD4rZHUWw31Ufz9FmpKlLVzPglYoPykdRE+D
M+Iyu1kvP643qToXurvSVPo0E2ExjORjTJdo7EwNNCcUNx208baKSJqn1queMy5P
TEpMXIxRXRm/Sd9DktkZzYc1/xP9x7o+m4jLKkbBPHW2CIAttoyKvELXgxUxzO+C
/XV8hhzdXhSHR43YflBHiB/P30iH00tFdqVVjQu4djdw0IsB2+GkKllakEV5dHg8
gB6Is+M7Rp3Od5oL7jyEEc1FMvhZ5EO+5N/MheoNjb1/U8jzGs2yRCVHdmfM6oeg
03EQ1JonUOGlDcD/wdr3SsfPqCaS4RZk+BR8BS8zHWAGHAAAKrbLAmIcb78S+dN2
m8My+Are2LvB8CYLUN4Opg5/xXVLOjtVDhHrVJyMm0OjsEoaosiNLR7zeR2LadNz
dgo9/g9j+JckPBC+jE2FkKFM5NfRlvx8/EExAG9yBnVRRUzbFxy++D4CsX4Hr6fP
wsZ9mCcrARVk+6GNCAbxgZBWEuysAnkI+6rLDxYsNPDaZI06wpWjDAsPUhuwl7xs
RxJ7aj9ERJLS5C6XxXieY1pORvrVNDXD9MsOvLp+DeKa84MIdG8I62YdTLdNk1to
qrHu0ZM1bAqFYHyHlZBvq214qsX6TR+87BZtIL0b1iEOY5GeOi8/wbc4mGykMveQ
d6gs8g7X36LNbGKv72ATap1g4MwnE+++itjOhZQjJsdKoLZnnjDReuw7WZIJOcA/
lMiN9rMiy9MnXU+TVdn4Ue6YoEBVEEYBnhcDxvzoLcaNFq8l6LnAU359FLDLpKYM
Aq8oB8Og4mZDhpAHnSfWM4ftqt2Fu0wMrMBIk2cTvDCPI0qYpjGCAeubOkRdf3uZ
UdQ2jrm2UPEn9pGoxxVgrDPa2biwZ3rDCVXCQcWQQ3VNeb/vLKfk0CAgAckbZz01
TJSSp5+EIt3MO7w5aMwnMwOLXAT+vTGL3C3of4m6fZvN5dqX1btuzHwMKAGFl5sf
Yo/vpiVxpJf+GTC2Zg+w6/akv7Xkd9xQhkKVjcF4Q7l8Us/Gt6/rcnVwkNEeMsUh
yVjY49UPdDkikfvFCvSvGC/Zdoc8wzRHMQeU8j4uTxPJtAsMtXCej5GJnULt2eOK
kNL898bjieYkywkC4yufgZ9Ob0TISmtA0/qhr93YXb7RmVuSZpRuuiyPGTo/N2NK
zze5EGd6FmTYT24kXTad/7vbgXp0bDoc1F2N7JzgEjKYfFBIA3mQ9ysg4sUNNhUD
r0tCMmasL+iwR4RUiDmpoUk7AodVKw2IIQrMTiCe+EjGHUTP3ZvPfTNQOatRmNoV
FNqdIf+HItiJACvfpffMHS+VePV0g/T+N7KgLcPVZgzC/n/H+5SN83bv/nYlAmX9
+XsuHpH55WGY4EhLfXDjtyi3FiGzX0G67vVtwepIxxC9WNtZIps6roRJDDRkl4jj
Q0hM7+ZFPcEh27W+fquO9liNR3/QavynLWSvAm2nC4Ahok0ubvv25s2/2D5xGDae
`protect END_PROTECTED
