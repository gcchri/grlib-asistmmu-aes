`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qKUGwQzukEicB8enSfqj5LJX2yLAhdecmpvoduIKSk0Unv4KWqV8ZCQh9DT9SvDx
nW1aLHJcs2awfrQK0+GswgNwdS3bBQ/6UPnFY7hhT1yBGkCWUjpwbMxwiAKzgSyV
3M7BWVgAeiB2FXKgJMsIIYy5ok/wonGfa7btILplmzgU9+bctmRjuicN0mGyS+m0
hUOfMUnkiWrpIy35ClUU5c0hm5nZX5caL2pq8hoO3utNXz2qbNVt/BSICLsr4+mN
+a8j6ujloLQ47D22AgqKNXDp6VLK3z9RzJtG6vUzwkfNGZxQU7T6wpVnMipeIohp
6lxjF9ngNkX3x621VP7XCJG1sbTvNZftTf5E2MKvLQ0C/Kj8hjdE/h0cdGqZi+R/
iHEFVgPm2fk829Tzg0nlQn5UDYVNj1H/oHqcjZphgfd5/fVKpI5YBjuJLUWF8vFr
Le+2Ds/aixObkKuYVOCc99JVOafOJ1B5Omrvaj67UrWJ+oj9EjxUGsuCPpE87urs
`protect END_PROTECTED
