`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S6CEGP32KAI7rfJC4Z+Ex/Wi+kfS0JfR7PQvROAAYR6L3nMX0GPcpOi2hui+vSK2
8A9sTZSwF7uXJI98PRaqPD8ENW+kaJLJD5Vqs+pQv5nhFQPbsxMcCZY3iSQlHkBA
RaM7opPbyvKrxk+XpaeDasQCUyUwEnGHEfT/We97TZXEwx/cxcQDNZo1H3XPBJgI
TMlYBRHKnu2oBkoS/omm0Sv8pXVzdW4deXiYIjfo83AZfOrYTDPDVYfeAGnqZeFB
NHQiOWn/7eo/i0+fjygoLD7DcbfKBtSQGNUMYo53GlelIEJstK0uZDCSG+QwLCrj
Zw+ZBWorHo5PMzxpxji9bpLrSfP92BPS/ZdB+8dEtEslwhXLJHG04aY1ciriEexM
+m/Klhm4DoFBCF/V2xabsx/v2/8NWjmdddALHHG5TmUz1BKs86Klj1GclscwFpmX
yiitsYLse79CjRsHVwY8Fsp4hd5bvRz4xB9TsEEYhD4m572MA8quYdIyMMlB7I/g
16XPEdqLyxZbLO27UNoN7TddQJtYj+9f7mJoniQAJtrQcbQjJv40dYRKFED12vHN
ZWGMj29Y4jhJXSJVXBv03dXfBF1b9g94+PSpBXeylTp4EMvKp6VJ4+z7V9viInbL
gur46ViB3s15yPmVDOZKclOgHVdWE1IiounktwRNJ9XauFta5A85u4tOtyRkGLz6
4DhHGGp0gqKA9oGjnsfBDWDyRgY8o4/MvYSg5Nq1rniAv1Zc6vckS7n8ASUKb3TW
zdb7euhCny5e5AkIEWOr1W9dOeQHKuxvWF4WXL08+YoqJjwAWby+Q8a2U5KqXUMv
YyGTVGUavZdGkuQSRKYGiAIzsUS79YStRiIUg9TqIcyfaOwULwAD+TFp3roo3lKL
YBevIM3db7bj7O/cJxu1iVB3CJeZ2/LjMlA7A/aCAU9z0IMS3GrJ+/WuXeKjTrQd
H7ggJsZdnScokW1fkXZq2AwnOZEPA6+7Rs02FquktRg01enSZ635GbfX6IbBKlJm
je5BcfuJqOF16drMvqVdcg==
`protect END_PROTECTED
