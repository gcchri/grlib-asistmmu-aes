`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dy5iAax5Ha101FshHuJZVt7OlKiKR26BjZMH9o1TbpCH0GLw9E75o7tKWq5/cpY0
bmVhQKSxi4NE8XPUnnqO4ncEt8dog+yoWUv9Lb5sGuUL8wdbBsOVF3dg/w2qfQ3B
EeOMWbkWcgV5KWcNWd9K2TOHdoSElv31T2eCQJdMwku43+LmUZPreaXR/yNQBWAb
9SjHCaNhv/1k+kj4l33bBLJCiUv0XmvUFYXC9YsM/y2RPyl0RSUDSZmHaeGGwdqH
6WsSHyCLa9lG7XIGp17HPyAcjfGUF0Pd+zIGQBrimlEQJDyswTwGrZYeJFBLVrfq
LyuIGsNHd12cTpSmJUz4l46VJgeXXgT9V2KNORN4Y6n9wMhkIYY5UbwnkLJ8nafI
jlMWeopd9+7IR28gj6+A/W86fxsbb1s+AmYd+SzYUTrMECzZz6nMKCpSLvagtpX/
sWnU+3ET8wlm4K0qkdJhGijKYUzInqp9jqNbs/fO6zCNBMf5/30WChSYR8t/K3xN
2ZPtM3O/VBaYUfcBXHZIYbvC0xmtQzyNNZa2BQWrci3zxUuSv2oEV4vkBDJLzF40
GxJMQKadyheXgagFPXxXYtogc/LLFAclbNWzXcgRPUwG25IIzhLti4vrtXRkCe6X
0HDoCCCKQsfIiDfvg5Qcu/4xeFAI5542VAqmnZMsgREeqymuvLuy6w9IkCdE67zc
6OcfonztlcLoAppRkrgLZ2s5C2awBephqTDugIuZn/e6X/3E45xwIhfd+fuJAbVn
aQZnn+GxxFYp4e7SwkwejK35MSKE5wEjEMjqLQgN3QfLeAm2q4cyC2u/uV+3MqG+
IoiFkp/k6EDFCrI3X28dlpHM6O2RFZZffwSxlTqYq6vunlQmP5iUppBuTdFl4wDo
/V3smx4nJSdbTSM1vzx+k7ta9K1fE50uIy4q7FHBTZRjjsO2Tj2f9zUqCZPJDbLI
`protect END_PROTECTED
