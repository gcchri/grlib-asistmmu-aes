`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bUWTCVRRFaLjN1e4f/v5YZpsLsIkTCM3Ke/Eg8zXr1pQ4i5sng0CkqfIJS0rJh0/
YVQ1qy5sScnXuY6f3DFviemyiqiomRc2WUrhlPKeyD8V9H+1MTlbKzCjeDHFi388
rd0v6DaRBOuuoMoiTsPqIoPM6vpWMAV2PTnoDsZLjG+yDWGzfXN4eV3MqBSQHqRQ
jKCM3pBSyuTzlzKCChSvIljAyJTAljESHvhTSyQS1m7khwds92epxr789E/1koSc
Hl1ZWh1ODo06fLoFH70c7iKBeVVD5JNHnqSadAe/HjLYYuum5RixJXrAxq/MCDvA
nNpGOz7ts0TodAA6USb4dGeWGGgBLvMqNeBxGw+3R7kr+9H9dMqeJOl2g8B2Dn3Y
RV/VnFcvJDcg085xp4rZccR6IlKbqeZ8E/CDZQhnTiLqv67Oy/f4J/sZ/33Wlo2s
43PWBXw+I952zaAkKi8mPeBv/84Yuhzpr1IQFpspmGeUf3B0p2fhKIQmpBdP8g5k
`protect END_PROTECTED
