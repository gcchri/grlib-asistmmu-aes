`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nNtEDzm7vZrq1QX7j59ATuW2yWSJSM1PZFaMauzsKk4S0m95BX9j1EaIsb3wfLmV
W7k9cuPPvDTXZeefUCiSf/HfwuOHFQxNEmo6N4L0tMHHtWPwj4l0uIQaFKuwnwls
zsl6tJ41F2YHYmBeh0k9PYClYWpDBeuE3Igv951EudqhgeS7JvjuvjmKQKRcdWyl
gUVlH2AZcy/xNW2QZ4MnjQwGBXzwTWTjFo38cU+3eAtJ9gm0c7gjetR8YVhl3yyf
LcRwvn8NOcW8RHh227wugcz842nljWS7fVe2G9vaI8+MeT1HbqAu2tXIPOnfailC
OI5NX4d4bkZAp7nWZO2LYA==
`protect END_PROTECTED
