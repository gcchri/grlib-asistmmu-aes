`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SXAnBv4sjpm5UXN325njvILk7xSSqaxACaiR6+TT2dgVsedWkzN5gYfbYx+eQzeO
1sFP+grE1SinMmimIGMrJndVlNO8aw09Jyko24WFyKDqKcGLsWPFsbIMuUWvAhXG
ZfiaFGFcCkUKr1hgMRMkgT1UcQK0jVOhxM9oD/ejg96ePQrwTR+bAbFpWLi0E0Km
Zy2prHNOUhQ2WS3UO/G7ddxpD+nyxkFu19iUX/rwAddSBX/Z9vQRfPPTPHAWK1au
+Zdcc/4Fxsb+ouPyMsgSKgHNCrx/cF1lvtupv0eEFi9s4v7RlGRfIbaHHDwjwl/y
VqGUDLX0V2HKUQf1SF83wYwgEOwwbs6sOqL+qNrycbF2f9LuX502sljzaXpiXl5h
`protect END_PROTECTED
