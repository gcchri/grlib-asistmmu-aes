`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s1+znAqj+rv0rYpy5n3Um51lMGsY71Pq99KXZCYd4/BpUtHQr4ch/dGWH6Wtg0BX
sQIq4nmbhTJjPg9Z+H6n9oaAMlEH1cSjVGZNLThjq/Y5R81xC/R+EMGdk4rcoHhM
ZL1s6yy/GtnzLrjLnFZTeI4gziGEDAOKWp9gHECKVMxmI8+BGYCqD0DQUzweFNGN
6SYTNuPwxzJ3YPwLrG+rTtdxPk3RZ7rDHGHV94uSPEoobfVk30e4jsIbq/LvnmxE
BcHCz7OeCUZaOfot1bKNyaGxcSpK5oLZkHK6ArR5LHr7nfTwFFHudYKOsg64rlTz
TIhfirZzOXt1DKE6ZgbM3+a8vHvvosO2eZi924UjtM8hsJj6d4qxjDII3CVZ6T2i
8GXxL+gokGWMbiJ46yXQR6y6VUpRuT/wLzuERA+3CbeSJkxonXtwBAliuCvWuuym
xDTaDq15VnVbbZ0h4NLr2hPODsevBOGo1XidmjHpZS5491RXW4YAmMvOkWUNdz9Q
fApB3NTcyW5REZsvHCiJ1v/zb6g/Pw57npvn7pAth7vizIa0EGFkp4IGHO4x2s5E
YA7WPPOj5xddDwtNVups/kr2MYxlOXHDa02K9w7xHjPLuOo7hxblFZQWT+eE7dBb
fxtAmDnLuzWBm1sot9xesdKCZNuWF7wlmsv545Z+Bm8/iRoUsQWLagmaX9xfMcJQ
ib5Z0v+fgmMWHyBcvBLrF8dvTjAmVCLLg6Fn2gnoQ0PZbHU7vYsDQzYMs2gXgIaK
JSnEBY+vmKjGhjHKthKFqpX8nc9kIQLtHDSdCaeGDymCZv1zbY1oYzUAGuH0unfZ
dmnutPT7U6IisA7a8d+Pkk6lX9eoQKTOzJCYPeIdZvZn9/80Ze90Rl5iKxND78l/
AehV3CrChZ6zdiN2RoCNLR3iD8wmJE+k4VMt5rR4/RwuVY5wmK4feyd6N6a3NoHg
AOBSQuYS/WoPydARQBV2cPfG2VWCIkNZVjN3hKhJcEJD/nMU9dpI6WbAqvyTU3ER
aOD+CMS9H6RSr6tncxaBdPQX1dY3YSObU2VamOE8YstpuFBEXvJEQaIvGvWK6HHC
23ve795j2kUi57Zx/fpPhoJhHKmQ4n3Ang49znF8hP1Nz6LF46L221TEjckKvUXE
GiLYgi1raacOyZM34wbOZuICJtKAfZ0grzOvwXd+sAqWLTmz+9vw0tcqe3i24mtN
pB9dxRNysnm3Kje5JRt1o/AZiMXwytjdsEQNPVQl8yqYSW3+c6S8HmGWAebIlhBB
V8uT0WRe0RkGP5BTuIqiGWbNfFl7ZYMt0Kym7qMKRSn2EeKDphKRMFetTlZikJAs
3lK23GHqmqiLED0tQwDS92VZNS9KrQC1cINkCFdl75Pck4CpvNdw2x/BFjBTWU1n
6VPh6IaVZeIFh2VLV4mXYJwLe7zJMQbgJtQZTejX+hiTIdLpNgaiiu0kI0vIGsEx
vklFYU6l3jkZibZghLOModAe24L0Yv8KwpIMnhFLLXFjEuVBTq5xhRvsiYSuE4+F
nZjJfl8m+nXsXFd8BG3Dt61cOnKpkH2j9hvHSjjwj8GjK6fUrAFxGdDKm7Di/7cB
kiRyxyejfdd1+wUSQnIoD9CZCwGkEOPL7yGHsv9iGoMhasXiSWAPE5avy3+ehgyB
T21p14T/BP6ZyZ61yq+PCq1/+BQU94ttFBN+LxS5Md3UsRxC5A/szo6U5NI91Uqd
G7AAjstWvl7xXo2L7mc6A+r3s++UqWI875xs9jfa+iJbOjQ5Fo+SELS+yZv7IMGF
tS9O2H55iJV7yebPi8vTimFZ3xIft69SGZJmEZvkB1CZU1+2PSB9Wgt5+i9zpDAr
CORugDugTw6mqLrb23+Cks0czpLjxEb3nu0RvG/rXvNrK9useZAaRfb5cSPt8jPf
MjgUNopu9Ek2fGuWKPeJT5rDrRXZbxmgZef2SRVA/QfB156JVkcbp+cwvzTOlKFV
fejrt0zc8tkoTbGuhG9xtULcYp2FlzWp2NHOKKdGtDh8vzT9ntGt5QyC1J+FHj2X
R/A8fHvgaM3O2jmUtLifKodDkAEYeuqR4pwRSlDA+YKYRZYPcgxRifDSUYAJOd+v
tV+IyQRVkQQyVpwQupRxVQ==
`protect END_PROTECTED
