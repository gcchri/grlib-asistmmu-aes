`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a1C/R8CzuSj/u1bmtO03Pb+vYkkU8a6f1eumzouvdbCm1oXZgi3HhUdbTrWiM4aO
9wvMTREUHCO+h7kmmhqQhRtAw3C9mhvbomS1LjXlqGzpbSt8Kw6zwATLLLYr1TV6
n4oGXOX00oZlsnFbL3QRPv+dAdA1Kmba6zkUm1SI7gwp2nPkK1/+TTqzdLrFoMln
Ok1GF5qWZyNKd7QC7X61OnbmEOU08pC//BBUFQ02Q3ofm3EM29qAqFb7yRPkmKxa
6KRuxbzKenefYu14ZBjyyQTcBKWb2+WlKzGj6Bynod+lQAN9fQI39xDye1jY5Kb2
Qld+/ljc1k2fQ2keiOb/FiSOsbafrsuexO+e49A1j9JqZe5Raten7h/cbROt9P/h
NrrmEzdR2BPFpvy7+n/Mlswdu4c0osuZazE4soyyxvvsbjXNIS2OmulJoRA9q9wh
2bTgbc4l2Ia5Ln2Akm/exfUiW+kTVTX9/yd4AmhSVk+8YrnLHtPAOV8BoRUgo7Wn
UR81I0nPmaKpmRGm5mA4NGReMZb4RYkg2Lk0KbH5PoWDIK6zHIxOwyDNltx3VKL5
`protect END_PROTECTED
