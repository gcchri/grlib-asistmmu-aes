`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XXnPbL6jvMXMoJ8o1lOvsHPlEOSB1q64gVL0z10QtIiIWZVhf+5Q0KlOoGBqlIJT
QIwmuVMMRPthC0Sffi6jQdnxfJC6WP7m+rBWEShAXTM6/cDf8RMzr2TZD9os318/
/rn/+2BUwOLeiFr1BPywV35PN+hg9T3SF3sIbJ+u5L2SvvhiS/MVl45/KwK6ltNX
LJeKzh2PLeItlW0X/ly81DkjIpp7MvvVkG0DDy55EZvLWn3dwv6OYyUPomNI/RRZ
vXwlFt8kG9IOrZT/8AmREQqD+rqgtbuoPUUfu6M60JHt7AeW6kPnPRk098/k+baL
yytr7zKh99HtGhJuabkNuHyCxp8kFfDlyzlaxddTMJEMDzMGivEZ5ZQwziljK980
mJy5JDcpBxT2IdIIa7HjiToiFZtX2mc1TWwOLKlRkbrLd3Z+k/C9dqkjsCrzSW9F
nDtBRGJhgwzZBk4N5rNbutDeg+idbMzUTyBzS8Kk+3uEwOsciMcz4qga1u7iFKCM
IlSA65GGGP32bjrqPTBky6h+1Iu5dXJf0FrVZM/gWA/Szh/UD8t5mQXXe6CEw8MS
UVjfpoZT72kKeni7uhMiK5h0ssIfJs8coLxDUkJTuKLBMqI4/C9q1GNozvJJVHMG
LhpMLq+A2fzvD/L3elfOZA==
`protect END_PROTECTED
