`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ogvEuFpzBlpA0r02l/Luv7ev/N8H5/1UOrZSrtN0d4NI6dhAm679FNHJCGvG86ga
FgstebgaKq0Yg1idWnMlljsxKwlwPSoYyuuiXsz3nWSGvEnE2wDTHCMN128SDV8T
fzvpuXXSag1oknxG9T2F85E5go19eD7WaajoXhwmJNtW2PFFKQb4mXqh5r54n8jy
D/vu8zn4UG3b/RLyiHSS227jfADIKKY/TJARumGUqdyDIn65pO1JMCBFfS5d3tNl
v5eX7f2dIgxPnhY1z3uiqMsdHDp0eh9fOuYFbzbGRkRSU96I8nfavyPiiGew1UP0
FdKBcr5zJhTeRZWvZ5y/CjexeheigXGDyieFVgUfQXg3asAyQlsuAhWKg/1ZirBD
489CGchNYzAwAJFqfkDw+R7GgX62YNsxUWlZGpwvtTpI/L/tdQsadTnmTVmatCmu
YlFriCaPxqWbTGekfEkHgtEX7TCnmyxjWjsxsJi8dhPNZafuC7gXYqalMG3JIsY0
hf+Kzu7CzwnRGQkHm3YJIGk30YVSejSOivYgUxOvGOAcNrx0ljzzoS3AQ+ZGNphW
b0mIpQ3MzO/bg1Ded6zC7KzPuF1Yfs5hLoVkonN5my601hy6RNYvoyxZ17mjDyYf
jXfuiiy6haPKwXgmJiAAhzOoL0D08a0pwYyVS4jESNuuqAfTz1aXcYVafFYZt3+J
UnA4VwRsnt69nDg0A21BdO77Y2c1KIo/dt09/0xks3kIp+cRVRLbep7S5Kd4Tsqc
+WzlSjStaIQENuqbMVgl6Okkd3hlXp61I1kIXInVyAq8L13DYO7bRlXnhJAV37By
vDlS7McDnVlFTrML27cmPu2mN2i+DtgeaEFzoS/KxqjPdyfnU/x9N+yHocyaHCp1
ep1BLLmyc9n9We9BSUJnmoxcc5//HdX5q5wRJ1UwNZVGvBFJq4wacuY5DR7UMQMV
zjr0oZhkfYawhPU6j/DeTt3PsJL7iV+XOQ1g6DSD4PMH3ZlnjrwZsKc9cim0YzLP
Q7oIyQ0AMSaYPlMfVMOJGuDYY3JSPhjNTn/WanLYx85FOPMn6zrNTgdBtDG22J/V
F8g1ar80OEMBAnfxcQ0ArcXuCeFlMTTNJmMxgYLo/lyPPs3TPQDmiPLkMv2/rKZX
uO0weeL7EEf2PuccucStuI0w4x30/m7p1XpOrGqp4z9RI4MYkQc2nJ4wmxdaDTAd
pJbAqeN8uPzzmx1nfkT2OZ0ddIsTqRHqfnjvQVbhrqFNOjnbMWPX2yFpY6UTbnNc
L+/MRPDhRo7VJcB10eTNZIynuFjOAjU0Q5RGANOFTXzDvwo4+pqgAuqs7axH2yPN
L1DR3z/gthcxVDsR/freDw9uO7pK7DI+Qda5FHqMnysdm72lX+McawPnqpEWDCeK
clfswN2DMOIemepfluVFRXy/6Hm2niw9NMVlb1Y2ZmXI2om8jMondrDtJjsomGQy
x92mK1cnEg7xpx2Q9BQ7dOgPJMFQLrUGj9CMIPH6KXIb/kUH+SHUmMMN6y06qoAk
VpDWhG+ORR6coXkOWJ3XSRsVYUJ+KAQ0EJ6DtF+Kdkvysn4Bm9rcLkaFVQ2yVRSM
oFQymhSLp/QP3MGiIq8HIbdoXo9Hi23+pkC8L6GE5GtzDlU9aiJkgRAd0Zq+/rkN
mL2sDzFrEFIH6sYnBLJOh6tCSQgYlYZa6o6IiGkfZ6tBqYdWiMS4KBsnVmZv+ujT
AANeEFN8+ihnRTrp5yCzCFCgWhS5tOG03wK/9PCYY+PD7P0rYoBrhlN8MMoUM2mT
QBmHoM2/qkTisJMxLTAhR/EK8ynlsLVgExgfu5RBJ+vfjOGQb02sjhsZFmaRhu+F
lm9EHYUdPqjahaJGQrTPNQ==
`protect END_PROTECTED
