`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qq+e3IM9+/3w+/Mivcv2HBuYF4hvzcbV7b2Pq/nXzALEIxEflPV1sEniwuCwkWeN
LqO6nGv18WftobhGwpMbKmBwCXVp1u9Xy6OcYC3jOjx5T7XGgGBwgwLviy8c1ZhL
1eJlNdYIQCuTGoBbdtlaULXkYKEP9Yrjvsq1Nm6nOChhl7xUfhlemLHwoIaCCcdE
2ViFGATLCP9b2J8bymEk0BSLYJNW4raxmcC5pLbuZZOcuHrtLAHkmmPH0itxynAu
s6zyOG74CO74CSyGtM/j5pfHRR60BWzNbziqKo8tDRGmRNwryfFjPmXiI728t6MY
x/GnsFUYq1E5ukKAqnIYNxXKtpr6/p3vaFeJUuVjbKkfHXJFpjGZCf7pdwhBthWA
Jc9FQUW+IMOhTNGBSjVGYO0ecCYqCC26ODlGPQtXJb8=
`protect END_PROTECTED
