`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c0nKw0eD2+ywwtN98WKT6q9OEKhLnn00LMYZxqemXf25rguz+ndZPUUaHKEW0uMR
U0QDq30vHkXZHRcJvFxuKn1nKxDlQrWxk23VDgizmqEHIGnMDHPImbTkE3m4AsXp
Ki23psMRJzBP9EXR5nBAkQ+2OVswjeRZJjnvHrUcCIcRzIx/gUCEy8aBbSfejaQz
D22/zBxaOt6p6uiSerKq+hPsbhDDVHJuLVD6UwGNiMq/Bx35bk7S4YUj9MzwlhFq
Xb68IHcg/lpteEBze5gzy058UFoSkuhD+twftUFMd5eeaqDPdhHygpV+u4riZTHS
O+FzoicChv2d2Jw2Kkk0+v8gnIZxIodypQgWsLTIWVCTm4QvrAxbOI9/eLGstMiU
cBOxrfb+ztboAT/QCplgxxaLR6otEbbUKCLw744ZwM/QRmLqu1IYoOp0kxXaHCa4
v63P5syhSvCVZ44OHBwZXw9dVtnDauC2vVfqgAwF/tumuPH1BA5ge3LlxLulCyFb
dqJAQkrB1EUDaFo32X08v5DYQWmVV9/SIGSbXSgjc9kDHfDDDzCnimK9JWP8p83g
`protect END_PROTECTED
