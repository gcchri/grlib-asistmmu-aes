`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MdZSRZVZYZPkt0TWYOeyBQ11zCytLbH3ZxYWQSGDn64MWi8xp+J0J9iH3HA5jUmE
yH19E7h6iSnjpZm45KMbmCrToTfXRtwOgJO9wJZgX2lpmz/qVv7Y4unKc3GP6WrO
FomvOkujs70K+iLgqLPqqMXN0QFffkbG/7+XpvAaua3wXb37G3WhLn1lxEioHkh6
cxLhHpPCRTjHzdwb0XEYIqhNRu/1V8gdq3yNJlOdrMLSjfuURfLJ3V63xhyVA4rE
mwewHhvOOWAmPI74n1Atwp7lXPCRowHTTrejeCV7+/9ogpnmAzmliKjsvLB4hy8X
9Lwxq+5p5PeoWcagqHSXYiZrwjNuxytRC5V68NsWKt5RR4FftvMNXWGgdSqBCzv7
3PaUnHZ83skIf7w55u60JfGnDC32VNoj+ZIpqR7Ulto=
`protect END_PROTECTED
