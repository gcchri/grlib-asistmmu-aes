`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dzvgcb7yfKm/6RG4k+8PBKQht7H0e2rpzMNFrcoDjCXvhDmbMA8/yIV4DjWU+sL7
xZyRooKHf80lZ/xH8gHmKbrXotCoquqQBYhhiSLMfFbtqp/2rKiqQMemXFrvvr5+
368U+Zyf/9iM72pQCpEbzYxqgNEiVYzEDdorVYTfp5WUNX82KXTx0k/lEygKnc9X
tMmk0JBt+qLZqKTUaL6dubjuH4xEFP3ZMUz2t/UPDN0nkH6cZwi2OLbYZ/NAGQ2w
1MWiMow5dYou2wMKZAk4usAHYGc5FNler1lc4gzNedMrdWlZ7LQVlfGdcSSF75DD
kplUh2wrj561aOGm7YW8sxFPM+4ObhGb60Afz6EDilfT/ZVFpB8wA0T9sZ5DFyHb
2VH3uGsVsqrJ+2ZeAITm4sjrh5pHdPMUDAFpo1HJ5fjuwZ+DiiDwqiCYoBYE7aZQ
CZC2fYGKvEgxcqlb+GDoIHFRaXto/J68oA5rLrGn8Ok897w1Eh/hqffeYC/xwRtA
SB8LNqBUC6IRNw3RgJlBOeLFyeHCXSa7CQTgfCuhwg4=
`protect END_PROTECTED
