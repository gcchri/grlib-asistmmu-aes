`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NrR/1ZNS5iTxk9KmYNUo3Ve7avKHWtPgIuZjl0V3HKmt9wrg9zq4UGiYGgzfMIYm
jbQ3sl2amInlARyldkNy+ZPnjLfI06gs2px/SiQgLozNfzD/yDgOYImZhjS9E6iM
c6P1/2pD4dPSkYY1cdc10LtXzcLwq0t6eapDE16tpA2QU6iuM//t/53YktflL/64
NWJsEdNoOLPvhHk6hoQSQsEUjQYYm4VykycXRuQneqdN2qZj2iF8iqP/yfdEMEYj
Elz8Yne5ktpN1OX7qM+gH3pvjGo3yd0b5d/+lsY8uk+f7vZpM3KeVbncoxcgDkOf
+ruxI7KDbmMQL94Ov7gtTmXpxzjUiOUbpMJ7GgucTsrHI+bEoYqrCvgOaMHgA9zK
dllKavbLI1EyXZBJyQ28iedqzyVi6GYB7h/305ayZICvYTGDf4YQMZEj7j4GCKHb
SpOYUp58iY5pmbK1/37f283zpBhrvhS/tZYCOc3NfGk=
`protect END_PROTECTED
