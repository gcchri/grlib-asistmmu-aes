`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+0jLuZOe73N5lNU1BJoGUPf0t0wy0UJL3j0IMvfL7BYtRte81DtoAzdbD4iT375n
ZyhzBq53bHJXUaW/CSHh8iwS1PAJ0Wt+xecu2LRYLDrDsaDGVjNNcHhkOQ/TvTEX
4FuV7lewAW4ZSOcv8/0p4qwt0/cM5jbHTRqsNlJ9Vvxv6GvQEntbg7+sT/l29UNP
B4tsaQJxyOs+fsaywmUHp+6o7JptRQIFpHTXDFXA6AcRRcmFLPELBP390Mi5EOXt
4eS732rQLn9MgoebPTc9M2mwXpKsmTgPHhSw3VhYBfvp+AGvcisgtNw7EnMS1TPE
`protect END_PROTECTED
