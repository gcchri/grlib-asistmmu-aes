`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8VFZ4bJJ05DNfOGbEOz41p68i4iZE6DeNbaAz2AHRxRDjIJkjUfzqVAxaM9W2N+6
JzZlXlYv8ovMqJAtwuqr2VjgyzCMvTsCCgB0KqDJWjlPU20c+Qhe7Hcu3jK7ucdk
PAt444iUZN7GWDpb8T5rJLBezt37EI7FCSBTX5VpL/POLoPgmT1ufom2wAhtaKIR
4hu+6rltUn7JVyiK6kFx3EJd/gv6dnc4Ngvs6Q85ClIr0H7SJgh3LyF/tDSf5GMb
mT98kduB8Vqe0Qjbo2S6gWYxOxl23yIRjTyQ5GKpqEj4oGguqVUPc7oSOeP8Bez6
K51QCuLHZ6bFl1oVFXmq+h4Jj3JK0QxIdCY2eczKxjB8tMpMDkDGAPnDo0cAsAn7
dwWdDksOt+aJ1EWMdeQHQRbEoS/e2rC+RitBZa9YdOWCmnJpO+jv6fEimH2Xz8pZ
itPUeDYwgIZSJLCpGLw9R2w9sLZ3Bifo7O4np5p/pK78TW75R2R67bW0rFRMMpgm
1dXi14I19XXkMKJ/EcVk090pygQ0FpKu4zuAQbAfYOpbsGJy0YpqEWWoQrOTdwBJ
`protect END_PROTECTED
