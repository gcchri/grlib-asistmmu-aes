`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9vhCWbQ+ZrOd+jNGT9nV79X6k9ilHDnDWvt42XA/9/iPMyzTMD4vYe+4MGts0gIo
Ic6yOFu19FPzD1vnmlqsrOtQvwgjkuIkcxZdmUWz8uNOOO4wb20bzWYE0qaLKoxi
9iEFMAW5fNbWcaH0URIWMZzSmvIR553mpH1c4sn/5wsRjSjMHmyn7NwQr669N5Pp
RzEIj0ELtTNZVs5AhCmlF6/vXqbycQjpxE9pNuI/qxpBQoFu/3F1GO+qGQU1j45n
2SVKX4t/CkLYQc8gxdWPlyjFENzHgIlEffF3ERhnG5kUbL3QjM/33XQiX+elx+rM
bY9inMlWpTbTT8Jn8Z+bRBbJ9XCLPwoEIcNZ6SHrRpOytgf25SVhi+zs9uFQiPoq
OwzQoOGUZyuj7zcXuTKNsvdW9OKoTY7VsJjBLsM2TOn8hKqepX6TcWePTfOH85qc
PDX6qDf0UHUZZdhRCWgHWUgKApz7sfXbdKv1ZzuFSJnKpK73MhqbBQtWL0cSiz/3
UuEF9LlaFS7DzdRJY1kPw5WZ4mmIq5WQ5Nm9ZjQD1bgU2GspWXIslhKk8693rSWb
yeNcZK/KoSa4lTBlufBq5B5Z5wVCcSdooP7WPJsKC46V8m62pGYKFTlpD3Vvy7pJ
i13E6AFZIRRmeRstERULrQ==
`protect END_PROTECTED
