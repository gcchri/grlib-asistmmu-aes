`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZjUw0oG3NEhsWsoRvl5jrLYerPj4scWr4i/g6NYUWbYqmxmCM16PclZGne67N0L+
55GMUFUS2EVy97Ukymo92XPs1hRHbdXOCr1bz5nw6I3Hfd7cpnJeQN4fc0fpLHKs
/JNWvKcYzSmLImQXEuZ71oqznIH50NJpZQQkYj+qm8O6ieqvvIQ42hx1ClaqWHJP
Ro/xCy6J4ML4NW+nEzNsQjwN9KVYqx1CBETZQcBQ0agMFxCVhjqAnc/yG8wCthvN
eAv6Ixg3l91ph+tfIhfR1odLmtNaqD5d4WgZ52ktR7MPQa76HZvRzWCaFg5ByDFI
UeSPPPUt9wihx0XUgFH6czYBNFUry/wLmQUP73Shz1Quqdn1oNvmA8bHAMh/hYM4
mZkE+OZja+wS0M6kBbz43fXkEV/8lC76Ei4IOG7kjd+FcS6WbRJMQkAuKUe+/Tip
tPNJepWn9WpFKd+f7Ogeg0JIHMk7G6dQ7wiJOXGBhR8=
`protect END_PROTECTED
