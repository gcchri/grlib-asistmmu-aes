`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qdycsxTzKMMlWLOXUFLtdt6vrwiA1CLhPti17zNKPtnFXgiyvTj/PaUfeCOH+eOb
kn211mDvgzIfd16q32lQ/Ds0Th+CNY38Cobgp1kzyElEc9YMeLeIGyK154WLVm1w
56k5mLVtFshs0sFe1fPsrY23YS+dFQ69WCy+6fAxCzIEVyx6lj07SNE0ZM2IYIE2
WL1l8azi+o+WnEJu0zj4kYlWNE7oef8hwx3KhLi+Cwchl6kVsm+rkFLtn1H2RrN9
TuBHEQdbPQoZINss3AWHJcYHm6wp+2mG9wy+lI/YD+ebVlLYhGFaJYQo3aGEWhJk
hFPy/M43xJS8xvgGKu7y5surpUTFJrZkeuLJZFN8YMGi3yai7BzpUGX+xQA48nX0
50zpqyOpjQsXez6Rv6EkVy48j1vk03HhaLtkENdPg5TnuDlGSuMQy9c6nh9qKQDf
ff69cJcIqx2EaNjRbVZPlIVf3ub0toXHckgSe5T2uEo=
`protect END_PROTECTED
