`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t3cc/mHGAzsde6Jlmg860CBDFZDsuJ8Tk/j0EZJmLUep6UhZtZKYl8Hi4mKhBSZQ
yTdx1VmN4EW8OK5bK3ZKZg2/wIfOMKfKhrRe9tXOsBtcOJj9DAdORAuwj7bzyCk7
k2j9Hej4oAKeTo8jj2SETg9RHWZo7RRUWMbjS9xN2ssr1waqD8sIPKjoOoZyUorJ
Lg3pkXPrUb9et5YsD9IZZc9JmB1tdAYNtI/FKxxG2+x4Rsa3LglTua4RTCXTTdXT
hxYJ5l605VCbQWRKyCe+7cDflqnLYXzP6imE685YbT8a53W8d4xs/RSJNeeauZj+
IdQJcECgYpgt765DfRNNCvJKSRL6eMxloLTrJIzxoLgpNO4lIOnSeAFUyQKfb9MP
4Ynv5uvcged8L8EVtNmSOV1zJoJNv7tZYnv5cmdlLwa2nWqk+OfrGpBq+6o18Xfe
GcmpgUTW4H4+LUESd8jELxDYqVj/lPOgk+RH5KRPDdEfxt0QyH/Z660Y+DyUWx+U
Ri9FdkCEYOglHLHXrv7TTSYYxXa+hHtqXx7r5HzogT+nxVCZnODYk+TzVUdxwL5r
awrXhGAOIGWPnC5x3T93dcEUKWruFZJyu8m6V3HwX6hXF5E/b12DBnzwyJgGSQ01
oRnkqpkbZWKXCpiceMB+gli2yjY/TaM9rgoGe5sOu6MPVp3nakby59wXH9hZas12
W5vx3uEIDDDV0V7ou2+xvw==
`protect END_PROTECTED
