`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NS6COzKauzkKNLZxtnk4eFvaSgIOpgb5ngDmSPLN0faE4W0cn9MFu5P8jNctqksx
gFsYN1SXY/6XeadwN/Rpd0fSHbU1ZPZPWi397G7SfnmSMqVcfstu9WY+ZdV3Gi3l
Fp+CKe+ea4LAew9oK1djCFrg/vSeNbwHqsa/5LqRdJq2V3xhSlTb/4LQMW0XzmBS
iC6nDZw9mcd5whRa2g3b99JRcJiZbqhbYEHxzKeHg7wEnwD6MGFC2XHsMTUst3cQ
Xpy6YEiFcpCNT3SMFsrxO/aNuTCR6S6fOnOEmQ+SIBhmoT7HiRpiIj3HZjUhVpQv
H+TNVSsDYg++Hn6ruJkByqDda5AkfoE3ivZbzPPA4QywHIHb+7buwXHF61nJVDHK
JbjXK4G/KL5ijwSpR6wakgYbmiV6K879Hcrca/jTgX3RfJeEhzQVryZBYqNRBRDY
aj5Wf+7Pe79S2+Dx/qDm1EvGx9IOVKZSfKIAqRnopMaEkf96eoYfGUuHrDvnyGia
HavToJymeoJuA1yGDPF7us7kp1NHvH9XlgFaJHj2DCgJ75IlsmjLRYupF5hqxr8s
VnYpIu++2NRR6lgew4eWQUMVMCGG5lWE39rRfcrdZwyiLbhP8BdmdmiH7DAj9+QW
2MANNlhGxevlikNDsRNUOtmGwwOV/VUAg7K57qu2LkhmkznR49tVfwDRCMIn1B4F
eVzgFWbMfT/a2/obWZi72Gf7vGtsaCBquiU+SAyG+qOenoxdumgoOOeRdDVXJRdL
JWAuwhykxa1neKv9jN25uPhYQ46LbG5MT3lWwtWqwP0RgAdbhx1h2cI5jtICpffG
ttIrfWQSpcfUerHyu3ITY6S870hnyVnYsnsQfOqBs8t7n6u571fLe1KH6/LhFlmv
5+jhZqb6Mx7n4rvwgzmGfnyrbBUvLxy6h+pV2uUzuYu14SjhnY/2deRwAdvmnApS
knHntt6i7hgOrz7PctGea3EYS7+2rIOuAzZhz1IbEKxFO4AnYemdK/QMrYr5kCP4
xwQu/qYbzEgZWrkOPqfLF+CB5G8YMkdHg/OpfZhO7WEvUXh9SDW5KnWrF8kEqUdE
ssxr//tS3LFCi6clQokLYA3guF8hyHpzuw/2ZSQhK5PBRhq/wX9ypqw04CBJT8qu
D+PLGrZ2ken9D/z83RCS4h2BLmpxk8DA8EjN43nV25tWSXOVa5lEK9dKh8gUh5EH
d26Iv3zuMpvq4V5iFA3Qw0YmXXKiXzTJC8eTXlXd2mlQJcn2N5bEnSvn5RJdWlGf
dpJ0SP98XPUJ5gOz7B5vdmBXpHkGlAeiJqfg7U6PfbD4NT1Q/y8WjQNjhVG9DFNI
Ss3DgWTFX/yltBZJiF0VXuUviNZ0WbLWuHMgrJFaMRJ4gZW/4248Syya/ecIEDMB
tujOyTe6qkdo/V6GX/QTvM+FIO1+mvfeboxQXlmLZW4LT4hOqhsrzNzfGm00WNZG
1Ormy031SYc+DRR3WkQt4mPZMh5ISBlETKKee+dB5zN2ruNxXSiybFTQLKiU+sv1
jL/3tOj0MT8CmuL9ezQUkqSwWk+UVy4BglYrhFYEAmtVIYTJzqeEFNedQRK9yWr6
5/axyyE1k91nWG962fdHfMxCIdasGbpR4MUOLtahP4I64UJXZcomOFMyvoHzU7DH
xxkwX9oQvHjSAjhBs39oLmMHBNaHiIwA1fr0Bc3x96OA0NGtu9sp3zp5ECnJDYm1
V4od2VWbbat6JhIKQ4ICa4ZW8q6/7M8BOHsxadFUiXgnsE+SIqAY9j5VYUYexIIa
OQG8UewNykZ/kO0xAT8u+u01EmO3gsbuFRxfQoU6qvv2JEssrKZseRT2/O3v5hH/
+mjULZRMwftgN9ZDlBHI06z//PQX1dDvaVR4KVrQlyzfw3+Y8fbUkw3KAHK2kT0j
x8YHBYcpwsHoiBxUNhU2w5PV0AA4TcL6+rHTLwoDNQUX9ti3lr2JsIRtW2LfI8OC
kh5d2FZTR1IFmxTd7tfRdt7TchyR3EWrwaMuxR5M4XMLKHM4AedSGcsym0dtNnWo
inoeulgUfH/CBNwB8eunUX6WOxUprtaJlcH7JAnldiqD+iBySQZJopJ4ThMLnXfN
U5QsoXSY3rla7GYiHBN1YmMyKgJJiG1KEHLg/h3Lh2IobdzltDtWz56+bcExVkz/
tvYiaRhgm/g7RUcvNMdcAwDVZBBwIcLDCj6C32yiS/Sw16sHhrcbeKc1BAirpXEF
/vPE2MDOnKVh0n/jP5xZnvi1IoQEQcAZHNZ4rUxrFmuvo78RKLJ9oE7mcywrQBc2
GmQ+APVpOgLQAPKEnf8kH6I8Nn/O2tX/oeOBp3iHZL7tQ9acrLolPHKwS7U1n+Og
4j536qMVyzVdNJEQm9lYKSghGzjFRNVN5OUSSgiUHXauj02CfzQ2GkKMzGF46Fyp
td4JtoE2Br9YpeQnJKMLwqdoDyPuDW0ZYRTS9qwwQMwyAFK0sHQLwEtifDaUQI1e
FH1RGpXIHirmMTKLNuGuyDaU98WPA9dY2UltWfqY0YbNdvNQCs1NuAvklFPV+Sr5
WZGvliY8Pag+EG0muFbQhfjdBC+CQdmE1f7VKmpIgTwThVWZOKWe3tS+ldjfsMY2
RCFIWkUJOvkGAI/MP3kOAHnvzfOUeiuOPxi7XqLFEHFFWLSiHh+2xwshcV+sirqq
tLbA3ChI0e9kXbVcKdR3bkTTuO8wl83MhfANlzC+oanuxbapgznCOzu3Mz6oBCE0
M1cIQbR6v+rvqp8xwsb7fqDKj89MlWjB3ROBEk/VhPmrUh+CahXmb0x2A2kNzNE1
NpeX1MjekisdpV6F6XiLA4uNC3X+6JeELOi90OLRg55/wJLM7GTG8X8Dyd4vJz4d
8N1qMRrMe3S6tjIqwhrLebbkvV5tXmBuhDgzNmiNKpPRNnXfTC0WcUCRQZaOjwWY
XnwJArYO+1PaucIljkagkUp2A7H4F6l3Yd5REHORzRqou9sJYZKz3w6GQthais4i
w2eX0+H6k7IMG9J918TXqd/V0WIdPk20RGIpB7ed5rnCP8989GPUXxHSJ4By3M0z
gytcfF71BnYcvZ5u6xk27lxN1Ja8n2yhs3qrPYg8bBkuoY1oe5o7RCDwyCdPWe29
5p3fgzh9CJfaEa40kdibbimolTLbCU9HrwZ8w2pT66n6YT/XZOVoT2515vCtpWyW
fvHIT0LoZO9+TmpvY31Dg8w/AOsr/s/l8hVsbHdip55bvKzIehWeMc/+pTPN3xFX
DmNg3xuJmQa22YtiQthkPRkH82mj7+hUp1v7h7fM8E/pp39MY9pjeJIdbt4cG17p
u5G6Od7oLQMI2WHkBThEAVw/kFlOsa+GvvKSnnYxDmvl6uUEag7cCczIArw3B1oa
VkK/jBPoK5mVU7gYh/iD38ToPnJJj6+zaLGGuVJmtgmTBO69CEFEzjy7NQbneii2
4FVM7PqTr1rNr8KwtJbyMhrBk+sF7fqXDDhXoAw99sMVcbjzmBPEwUpSEK/KeNi8
vU+gm77IblqWabTGJcZxAKB6T2t5jqxdd3yLbtpn8PM5ZaumstxgYul7BQk9jRFv
PVo5q5NaPVRpL8XgHdaB8scVzmlR9NZpCe9dfrjs1NgQy9CIAa9mSntJ+0XePE+Y
Zmwy7XR2Rn+jrYhg1FQL9/s35j5O9h6HInBiWCcS36SycpGdRnx4w0y88FM8bPYJ
9GMpJJ8uc6z54/EVGiHBAqyyTocCl9KelT3R5MsGanueLfUQ/Levk7uEMry7w1DN
ApBDuMb2xsQETAeWnznOLwNzr/BI72sJA4Sp7Fo5H39EkY8wQ39Bfgbh6gPqt9Nl
+r+IfGEQfvnb6RCVZeHwBVcn9zrI/24tRrzJ3qxIlML+We72XN059HY1j3O24PHu
x75c6ks68YavT9I0p2Jv+NYfaoSOehMgr8LgHCQGcQ3xb6lYlvkq8u0ngmWqptOS
eyWlau9g39yVTJXkpzzrqXaaKhy1waeeZHIEB8GpyvBRxVKQbi4Pvd6Nu4ORJGd8
zubS5aFpBmTxASZCC9vju5e1gUmr3RRW3B+XxBl3Pw+N6Kqb09E+9d35uJqaYSvr
Ufs2NeEJ9bqHn5Bs9sehv8CZMH34I1sX/FqcmAW1hMGFKvU0BIQt9D6jT+wIT3O2
fKazXtqQ0Fj3fLKd1rw4pC3ObY7+RrBkdDpuMyggzyh2YrN+98YeG5V5lYFG9OEC
axFrBue45NxEYIhy7rhvOc6L/PFpCz/bDR44NPawfT//uaSU3gRuVLTTQN04aq8W
t/tTzeILjxbwWBBqp74iarf7u9SsZn9JH5pYt86czUb00IjuT8FLApg/MTUOIkJJ
TkG5oNqoZlQB9o8YnMMKJTjfbklF7CCoe9IiIvj2Lsw4qNhYtS/LAC+ZUZVz4Irc
d/cIgegmRI6/Of1IDpqXi2NjQtFul3Cv8KDi9xsoXUOQzaplohARMzU+3us5dESO
GvpNQFs8EP7RzOVGJB9qoI+CQKG0tqPi/XeecJmW4AXXIEAMJccVA/fNOy6YFLdd
XTMmQG/CErKOrroL5s2EmNnSCttfzeKGEYtK8A+TM/XqWbmZ1wtEcXNC6U2spbiP
KzvO29bbbgtjJiLhS8+ggT4gNIpTPtb8tJjhQzs29w1yV/y9bn4+tursFc8fkUf+
6q1DEKVdnkYNOS4Xgd/eUflTDoSpThIhjvagU634SX4YakLHZ+oGXhbOzDje9zqO
kLDuLQ5wzFJMB18QbXJ2RpE/I5Z6/AAKz8gwqY7HDjU1kgSFMlKDhuk5jGaKNPEj
YmtSoyPuLlYHbI+x4PzQAES/sr4jpeuipC7zmRyD5is5OkhNTb6HvdGOXs0ra/1c
+uhrhIubYKxFy7qM9ejfKgpJnBLr+6T7W8EeEVJE2YXPTMhhFyQMpOwGaoe7wpWF
nXQkX1MqlvBOq9L+KCsty34Eqo+ZLgaUBoVREaRF4eYgmLG7b3JxZY/fzjZ85Khv
1Nl1BuKVzV4jGxrkxGiyBOBdQN94KHKJJdyDtuQ+YO/Zu/HBTJ+caJeIV5AWWY3/
WrJrJ6zkjbgY/1yW60+eXcieZusH/6Q6d79deyLrjZYsPM5716qGcy9u1NeqC5Yj
BqZ6DfEA4i9ElBgx85owIqhv0N+bo0y0yr5F30Ciaj0LLgGUTF+QJKaZmbYKiWFx
kv2hibYlw3cCGAFsbPeh6+NykGnzj/5KZYNDLVyfUc1nx8epBfFnQ+112XiPoHT1
SU0fIAz0GsgCynK8rQFmyTL8Qz/20HwGKPEAhux9XtE9SGgdbucOGdvpUJcbgyqO
lObADnc136UEHceDNfmBeTkpmoKaH1OwCGyat/U/Ugyi6FuzOtHDd4oEvl7A1v1K
Ge/KI0JJgdcqHfGbWbRue3P0y9sG+9O+al0u7OM8FnzRHSlCHydnh2UmG9AK5ciS
Y8wt0BZoXDogRYqZYGPCnhXVbHTxPmyzcy5u+wqnt1fCMbH4/NJeoA6Jvwt+fV0d
jnr2kMNk8j0xYbY4wzWotgZzskSf8JpQTf7Z9j0m/6vJ4kk5LCshVvXaUp9xB/mr
somUiDkHwbHZoUxmaNPPtC4ZFp4oJD9wLzY7LEIm3xCbwBXh/469jpfhLQ9LewPS
gWnWuQ7Z9IloDOc+4vHrnZQxlKM7nUZ76PNyOtyt4vV4MGywBI/WSjCqzufXf2AA
JzOcATyktKqGCuJHHV3PhRFwqRz/zXZxYQwU3k9fncgX4CimhnN4SWAcGBRHOPaO
Iefz7/iNLP0xMXy2B/sfwY3J0F4tM5+SzWf2yB8BRqQ8Va4TaiMghiI6ySN4/fbG
5ggQwK+uYJ/9T4+OP8iVAhi9ivaM1NRVOxfqiyWWkdEPi0ErPSITN1FF4EPZns9o
ZsYhV/0J6aLXaFefIALlL8uR5j6NRXEonbGPt1kY5kgZ5no+aqHZaqOyLpbxk0xi
3j8G5n0FZVi3Ye9b6I0IDh+JZX2mYMW4kABICWaa/CKOsBMVxWzmgWBY+/+9Ca4j
K75iL0FdE4gaYhI72IauMOyOL2kM4FerpARwAuWEI19C8RuBifEUZphPOGcsgYgZ
cPUSUT4apqsOVW7bpmyuGAufs8/EJD/GG0N7XdCkgNxefpqp4rZaEtVr40jybng+
/LG/5pyHkJcYbUDEKHCCJgVRyFTzOWXM3ukSO7in6oHcopSXw4TSGUcL8UB3IGRG
BpkP6bkLNqf6d/76VETLW49O5ygQxGlg3QRoaByq5EbnkbZZ0bHzsZu4mTjk/+hV
R4ZArcyBffyCgi5w5ZxCcAipLyB+TiM+7+UG9TpPxa3/GTuWj/BsUVdZ8GiaU6fX
xQvlDlQOW5iuVqOpfvcYtemlOj7X2PClVXjJOflawEZqpP/NsMOXV+II0sLB/BTk
8B5Z3CASTWhpN9hAme3Fwx17FVVvuxnqzstYo5rExDhrlVZhhu1dkI40zyl6ofHs
3LC6ThkKLlMnZCdn7uHB8ttvSiukPopx+c4DH86OANzexvsLmciQmq3Ckq5v7t56
iswFi9XzNQoBqrPEjJyIKLh2T+iM7Ayq/J9BDR4yuQY+xReR6akwwcxMXnNCPuiO
aX9IREm4a/Mra8ubs3S0endg7jZ+BXzmjpJ/a7HdErZSfUpyTc+jKv4rjiwBa4Ot
b3fxRVkTTj+0MDpioNCVXfpsF0PPkKsycJPE4E1DIIT6YSLIokB9wMaahjXpECsj
+VjszoHg8RIlhOlMYSHXgP4zvv+A5seW43XUp/r3av8dm2kqtpmXI5Wx7JhYXF+V
89GYbnDsZ8r7SMwEPpQpzqEyw3FbJaSmrwGf27oWlqPJhy1bV+Fu7beOWmiVJr9j
4UtWGp4TumAhu22RpeL+F/Oy3ZRTnN03aTRHS9kFcHgepUD4SAughDPs1d6Gj1Ie
3LH/xSRUtiP1R4iOWyPIYJVCSPMfJFpwCE8l5lgpX0IZM9A8zgDBJomIlrWGsUGn
Xmq2zOScbGEQFUntQORK6cbYCHTeDuYBIzGbrthoB8jjgMn1rWpimqPnDWguhYyE
ptSydFS2bl0JMrK5o3WkUHRXuhGRUdrtnsNOKM6fmliRpXrK7M71kSELzOjQ1fo2
dfdSMhVqhK6xFEFjmwk0AWsLiQOqGf4r4tlbcAsptrXw0gs0yOCZ9T8QapCgFvMg
mI3W4u3tXg4hiTKeFVTbO+77/3/kUVOiF2LmQ8GJ56WJfIYL2lgvd+1Sxj9AZ/X/
QGC3KujkCeJ5fZ++/wzv18DuPqnudJH68oT4wFYd7fjtrRtmtUxzy9SEJVac6gwv
qC2z8D+66bjM72DVigfzCczCHLoQP0f6pQwX+iVEZtRLqLDWNUGzZwwNfMKHDtRw
Yd0OOU/hc6t+uUDF/0SwXkyK+Ul/plLhwNF59Gd9hGBvmeo0WqvJPSlZKeVAkzqD
Zy4Z7yd3IFJRYIOd5TXx9XNQ1eOyXic4GDPwDCXJe0c4CE9uRhbyJlxDusHRe/m2
/tIr8mrbIc8RTDZcdZtVcpje7UdfwcTNQdtyglgd1vtyCLJsZS4ZQwnLfpk8STZy
/2sLCVEahJhkfXH5ov2j9dfsGUYXAZVK8Td8ItD1k6bBYFfAaWih0AzKA4q1BbVh
yzJ60Zl0sjCsmDmVOpRLVEkVNS5kAIxuLFF1NQ7pK3sEe7xoVeVMFV8Np/Guj5Ur
B/dWMiKpe6mO0nZxgft1LZNOy6xZAlSqcsU4R2kuhnS7XVj7aW8hBVwGCqXVMo/l
/N0vf2IELjdceiJ3m/0BiZuhDVduWjO91LB1VVbKCjlHOGZ99YjAJma+5Ixlcw6C
l/pKlBXq5sUL59jD6k0LGNMEdfK7wnoDlETGDYOvyUlqNSAiM1P/INTvhW9P/1DF
ydqlMu8JB/OmZdZxbI+IvfklA/D09Vm98UYiZW7OdAL86L+CNiJnYbf1N3n98XAp
T2hLSpI1ws1cP5MaZi1u+nF3aS01N1Ej4DG7/RSSk0utma01+dEE6EpiNmxuX0fL
QTmbIkbDlxvBr/7DSbat3OBdsMUAe2Vy62/C8sIGzNIdd6sryOCGAITG+It//ojp
nIvZZN4e4vnnB7VgMYeJhlJsSeuqjS4iS7XzVv9UdqF45nfh2FiRQnfiDRh9vV42
T12KiMPrLtMILnj7rDx+Juo+5HtInKbiueWZ1yu2JJQc5wdjzCG+wA2W3HfNxHtt
8H3x+XtIPlf5TDxd+u7sS6bbZK4M8PEZXytFJN5eSBTwBZdW7eVgkVUwdI2z/k8c
5Y1IR7T5yMC35c5sCg7xuSSWPBkoTGEJ6N7eahBapkwkLr74Ucbr2NaYfkshk5zm
nyMSXCZn7b2JHDuJd7wGmS1V7QHOf0bL7aJBPPvmzCa9jaCoFMa1oiT1fOcTcSSP
y0+XwGfD/IagTyei6OMAkkUD2aOOV9IOGUbJCSLYgXVN3m9wPP0zC010+S+IvqNu
w/XUprprTt1us6BeKTKtQZwN8yRf9uMXUUaS8Co7rQi2gmVn/3DTeL5OV5gikBKe
x5rJosFYsenCgqfWb7dbsQfbYhVMhXII8S//KaPwIrEnd6tzWQKNAm2DsZv2ZM4c
xQf183Jni9+m7OkLDPpOrjS8wIj+FhTbQYAN0oBy2+AutKvsx2ocNUX2rrlP31At
eglRNmWUvKE/VK1RYNxqHqUNEDMby0zSUNrAcj/yQhSEHtbLt6Qf7qIlvnsdc1zO
OVQM14bCIfOogopNOHkA8moR0CnwFJd7njlmb1RGIJFFcdUgWqvT8YqGZ4HvF7w6
C7oypYiinEe3M+9FWY2XlwxlxzduTAGv5/DX53c8G21tPlNzwW7hYfoQgEhRfuac
N4o38+J1IyYsBqW/Mop81TwW+fs6me5cAMtTINlMprBl80R36sBxO5QjZXsJtKkl
jXEZtduj15TYnFyBFKe9LrDkLc2vlZ19RNy9NaiaNB3XNVQAvBlkO9+lfcwZfy8b
PL2K3fELGPZgpgF8t1xE/yYsKV7uaMoJ5uPT4cdGtWmee2UwCJv5Oydg7xmTINim
S6D+I8+LwrdBbC0RqzAZYhhZkpZiHbm6Dr+w4PYXL3wPMpEgrxIN4I7GOenIJMxo
KB8yGTOVBMw+ZpRAEeT/5bHTqYfqnZdJ5PTaCMCuz0N/MCV7tjZp3WSC0OUQ511j
wXo/pRXiRYU1hanlSDWjN46TfS9jCFgXJo7fWmhfqIr9r/puDqE3RBxsj+jxS7Y5
pyj1u1Ly0FaoLZK4ZvbzWcxD/s3lEzVLL2lqBG8m6Ewj/Hh53K4nZvxNaaRicepA
rdr7521GH5i6P9ZB0CpWvmJ4CxPocl72IxXBD7YNAb+zKE5tYxVTLqZIia8R6snS
ZUyg/XovMa/ZIHmjf7URT8n+LqzgOzdDQFtfb+kNyEwGCPe3GCC/UBtVSVDrBTKD
RHmpjpC3mNmjvFWFkodXwOw9Dm8bvbc781kHZAXTkdhkN9vrBpoegyGwb2q2+fK4
BdYkX1QnXEJPXqXuczywZAP1esZWVz5f6/bqR4hbCx54QtPJ8LMb69fTOHEcrN/+
xICFlqR/IY9/AhlcSXozMQED4q5st+dJZiS9sysIqBtCnJaHHGbqc8WIEY3h45oF
PAZMDDuxq3DigeHdmwWyLR785XN8L89NKS0Y6MeIyphCUuOfBAe5/gQqMU5ZgeVs
/cVXysn14jsetMoRMb0ZleeAxjzCvlXioPdd/kaNL70HPL0t9FktTE8nCpDI+/Ze
/2wOYsQK2XgkWgogLa1M3qAlWUUXnpLSs5AFLhZvWFKQhZ7Xe3yOjxNQDtx6pAKl
HSlNRiSLJeJFZmrzj3UaX1Q0C5SizGwfXx1lCMXEfJWZQDepgdJINh2L7YcSRA0N
nsPCADZQ34KDD4vew6jFsH+NE1d70ycwG4i+7AFDsnWXVdQ3adWgZltxnKrz4U98
Oauemf3AlxYebo2hnb2FQjbt+goDcHzkXCxCKui5ID0SmUVyPcJOyQBRZKw4EZx0
CHK5W1zjtxNi6EtRTAEABs/EVByTSdyaUvEpXeQ1PNjDLTyAxTi6KjYixnUmaRLJ
+9TzKZ1hqbnEal6szm/ppzhGbB4DU2u7qNNSAmCGW6Lc03XRjz6hZqh3T4H4ke3X
YIR+kr/R8CnQW8LTe863x2SCcMZNduxcj1qU9qROBraLAtsLoe+dau1svFRaz9Dk
qAOvPJrIXe8otSZcXjBjMXpvo2agEgkR9oo5oRot1ld+MoDJP40oCXYwsegRJBMB
oLAjTBneMVMvhKOS5KifP9H2d7Gb/6B0lzF2BeIFTrMyPrg2UoIrLfU4bHDOl1eu
iWc1sRYu+j4jR1gpJDrhlNEY7ywIWDKylScXshIPNBfP8yyk9MoUuFv9BczhMZp6
vsfNOB9e0vHIFAUMeORs8iMah1yuUi3VUN7Jv3mcZ7MuzsBSFG6OA3cm38dswp92
7JaeJI1uwtbScEiHPAQIL3l238T6LAgCetNLkoKbSV2RrCmzqlTk52cxmEL0hdWp
xCpgAHJvoBzrvrZEU9FINLtsdPCCi70SG+vToTxCZkUsFovtd/Vt8hweNNqXD5hW
1vAo59NCF8xXeVE1t+UO4jr7ab6rgvlWANEkmxRjGllz+rMy/4xYKuVLWmD+8yhA
S98RQr/Y/ij6pbN+wxdGkRQ8X6AMIulTInL811n9ae6GiIdGuqf5DC91QcZ0FuQE
5jFWAgx0ZDpZl6VsEiSc9ZGrclXpkRlmyRZKLV/PGB+JsS2QMEdvqE3E3iE4iol/
ZxXfydBs2x08m0JN8fPMd0UZZhmeyNAbmYgBrLMUgD1/f4209292RoiwJHb+XxQ+
qHTnhOIyVRpVS4fh+/JgUj5NQCaByvd1n+nQGIyjVvF2/LIV2d5mEG48Pfb+P7Wj
gWsnq6tBgq99VKaVXCmchiKX9xI4orwUzf0MjMKJ/CmcXXO8HSKitVseiE7V++Y+
0mkaibOuvJQTJ7MP8mPox3bjKTXKfpnT0ZtQnpxr73EbTaXgzHd1uRz5MgOUzRoi
DSw+LcMToE4gzs/vWC84os9qDa4dzeGTuXU+iRdisjOmM0G+VH/epzlwPuw9hZ7B
yGgfTgdrAS71iBYHJL2//Kvnji6JH6Rg6PME6+oqzitvDZJTBoT//lfV1mzDCNDo
pNtTYws3AakG6z//lmqn02eeH8ACzVZ67Brguh9RuU9OpQlDJsLHmGXmXkfocIWB
TcuUSyyYt7og1MKnFZqF5MFMGk140jTsH8cJ9jOEKL/hb16NZQDSzaDleR/RG7SJ
AjmGx+pFI7lXWOvE5lBR3JK1Q318SmYr/KlzJkn+o0X3W2qBqKs5FiI19zKpWRhn
Elw4PZQZQpxdIv40iYcCkcqtSawQDoM31BwhFAXXqBzlTOQOsRt0+LCufKaH+npA
uoGLNnxndf4XyEaR1RZ1vUguRg0itkgTHGpRHIRdOc3v7VBEYPQE0kKt5I99/PY/
bQgw6KFRe+xDwoJo9tmMyTK4Zz/KCrA6uERCeFrfHwjBDZ02E9mywGUU65LxOoW/
Kt7WnHz0h8K/bJMWSPBd1c5gVIJcU3iNUpWiGzKClf3e7HH88lNzHdtYbFrA30AQ
8xsa+5rUYEdOkdCkBi3RXYIc2JqxEP48nGDaq8hbsKSqZltWsI35sBDv98B1gXgk
7hYVQJfQVyQSRTBGB3p+d0CRu+HPeD+30iuf7cJTM1moqY6gTiaZORj3q+VWAwIr
OD/j3L13yPDW32D8sV7tsVAn0jupx37qkTbuX8Ekm+2iVZnKzwWuwLVQFvQWhjqx
AyAgHPr/gS4rCSQlvJiLQeiVqa5grPi2dpgBIEU4ietwyWVJ/nVpmiNYtfXkyb2T
mCdr0dj9yvJ76eYHIAKA3jMpFhVM96QawlakZglMcIFWZtg8eqI/CuemThuVrFD8
HpeDLruKLnHzVhMore6EHslC8E29eHEVbmF0wkXggL04QCJwqqt7ZmX6UYSlINVJ
U86HciFNLBxU8SNgx6YcgClaV+FsxDx6a3gFjnnhCpXLVWVhxpFmd/b/8Q++BmRd
wgpaNu2qLhTuSKJt21p5SPCfcGjxpsb3L1EKknxd712Odc/Vp07mQZhiqQw7dJRd
Xb1S4CG0L//A7tvEKn/r1nFHFxOOqmK9ZumZISsnnpqO8hF6+xRvHLLv4z0NafIo
4WaYZDGNt65t7i+LD0UqGF9sQyrCQKU+aPHyCHc9tC6Xtf3a/dzSsSpGaJc1K5+a
PEBi8RybXQRSaw100RpSTmssOQRvJD8kFvvXFDYo9xM0iFT2RV4LbLyVzXX04XYm
vqAgKG63Ll8VkMoh4da5QOortkzao8vuYtbQCWnHLeNlvOnSK7PAxQeDfcEimSRL
Qf2fXO6G53wAifSyUHF95K/syaDjZhm4J0jYj6/42a55LmCoFwULJOXAobvh725N
73rw3uZr/5SjEAeZlaC3UtlfWPobmR+lGHExKGrU6UpUtC+WiTo15hrgtikfxb/M
iuGPJPbbm9WK3hl4Y4gsTaaDui9sTNSw93/VFpHhEwjQuo0OmltDbKmmxs+RS88z
zf1FKyhFr34Q70N7SYHYeDJJfZsEUEhr+GUOZdR0E6wHH/BdtFwxFlviTM+oRJOX
uzeVailkZ13WEUmoEDWALtFXs/gH0GsrfIO01cYWCVcAGkz7VKVGv4COUacLUETB
EZO2nlP7HLGmKLrN3A2OzrjyVaUp2RPtdNu7Q5Dzqd7TOfUpGAvsPFBpCDx+LhEz
WC0WuhtcFzQUKfUSod+OIQNzwnv/hepaEPfqLtsVUu6A4IyjSPLr5kYZbtEnTcIT
cXM2DOzFq39rlovG9qd745h9zhPd8Sau/IGpWbTjG6N6fRVM8waj3JiSpqalmT7I
VxiMxenUbN+66VavRof1L7ECBzFEWYPoqaQMGeEK7g6oBtKIm0yy0GaRUFwpJAm1
gbgh/i5D0PJzzOEI2gwWz6HH3FabrNTX6nNPSbCERd0RcM+k0HJv3B35AnuyhH/K
qyb8BuH9zNPHYJH8Rq/PAhOB5cViZdUoUOK6vjJgpcA4fJVJGOo01rE9XRr5Yyd3
eQIR+BvVUidmm96fJ32oH+3TozDk4knb0Lz2gkpOmLcBgGqvs5+4qg8by6HMnLFE
y3dfvhh/2kjUkwNHiaov7zNadoyHPA03CNYYkrOjbrwYn3GVJRH70lwkRmWg1QRy
CthaOY9aKEtPBWPnrkz+P5kuYnvFHLqipS1piro7y0vs3NJYaJgPxyz/gR5Eqt5r
bo75nxnGF0VLQFjP6Ai3fG7YEiY1sKpfvATpIwYIZ75yC5Ve0Ml6FihsPmTpjFek
tGikcbZGijNWN45hyrjjE3Hp7AYPlbmXgMIJbf+EMsIl9qT3dxcXtO4tHJRlEEj5
X6XT93QceGwLVWIiS7yVhBZm7l91x2LDL/2VPCOCZaG5q8orlIvP+k6lvCn90hX4
nEU+8trhFeRLde7tRiOxugxGGpTde9DpGKqBBvE9Hg3VBAb4js4PbmoiVznu/coO
dhP7M8IAFDW9Q4nTWTXdDOd/KrxmrWrduDY5e2Uvt6woq5sWrAhRh/oGKfQmtDKq
aCn2XWeC8fFiSHozn8gtRvsWecZxbHgMhv3YOaiGVjV1F35ZBE0AyOHHdojwjkn/
rU+nEdis+fkVvemitGbQbg==
`protect END_PROTECTED
