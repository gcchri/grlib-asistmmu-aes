`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zDePZ7vjMpN3ekRHk/7A9JZIa0/qZw/0l/le22+8d6Q40fF7zP7eeFM3bDNNYFPf
1SxjDbLedi+vRxtxMI1KA1OcNzyvhMQJyVy66cxYy/6YCLshkhMsaj+XlUHDwTy/
iNUvZ5I4Ii+InXrS5tvyQdLjWhWImxj8VNOwdIqp7YYd4vlxek+AUeqzvJxxwE4K
rEsg3i2SItIZ8mM2kEpTf5TRbYbGFfDuLjjGBC/Vmnz3UXQDEJ3/CWZR57EJkOam
ABoOMk+SFZ2ktLE9YgGNrbCbAsFlr6UQPB6X7a2GvzMc3Oa8J3LP4QhTZG6YRXqH
2YdhtdlsCi1uQbpObJLhbyIJthtkZWRN+2tAONojFOiYGLB3uBya8zISXaq3x1oe
xHbsZjDeVLBr+gnTFMzFlg==
`protect END_PROTECTED
