`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SYkwhdTpKqU1djl5JpfxRv6QxKBIDLSeBKsYttBgH/klUT03h8J+wxrPHJjGqn8R
nsDxkXQcsMnMifYV1xOT/ykZrFYJ5YHfyfpNUoL2HOJi6YFNE3J4k4XzHpP9vSSE
EsBKvOD2uZIS3u/nAXI1ZnQBnBpX1zyYPUPNQA7qGy5QkNFviJTCWgeR75+Q+UZu
elxFw7WL35IGECZxNXUfL8LCeCi1VDrbrTRPjePHCliuzYa+FTQWFQRtuCwDQ7B3
2b5VfNyO6y/iyBPUGBWutfcOW+5pSx19C0c7VcTLqG98KPEJW96BF+EJHS8C6iih
JxrU4u9KxftTb1xcEwJMOrb1BMNtWvqOnWO5g1Hc7Y+jrZhtaNJJtd0SMtqElNgi
Otr6qH+yz2gIt+TygN+FWt0uGp8hxgs9brMYctbV3mw=
`protect END_PROTECTED
