`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C3mXmFWjPqXw+j7U6nNxhj2BnCk5GP/+ne8FyuO04XuQYXfR7HqFP7S5ozVpUlXa
jCZDCwibBCaPp3LA1DQA9Upll9swoJ6GtiBFxGevIlmPh3P4CDvyiDZA5Y5yCxYo
DAPE9ZEwouF9E12vsnnNWK/bh3RxBYtST+YvWETDki1vipuEbQiStnR3reOfMjXj
YXxD+i993cLJ/gbNgSwdk+zoNz6gNPvBsFLHJ8n/A597zqHynUo5vJmBXT49QdNk
Zb7vcDRmAhZUNd9q5Zp+YSttW9+8nAR9nz06OdlQe9vJcPlFN+y8rmuANrsgdwE6
eQsYcpZZkLZUHi8QajjBrgQ+2wpAPsf66I7Zx2U0+tOn1L31U6qsfTlkq12aia5W
v1vQyMBTku3e8qG+IRkKhrwiePgcsO4NL2ZX2hrDGiZR1BXlLRJNsOHuA3JIaNXo
HhF1Y29yD69OVVlp5tBBOEDgRCyAVke6rIYCgCKFzusuUOSDQZPI1gAGAEEmkjs3
UGBlzoqRgX80KumzUnJiJDegzo5W0eXynLznfR6cN6X12qZDEwtFm772/MmJOj7H
W+FybB51oS37URRgDRx3cBKOlVGBTyLM/2FxnR8hogzI598FSX6W4EFaQ8UBi9q1
x+yET4tr1W8s5fWawN3rzQv5R6Xy9DKGJzMFJZ/2IDH45wDEqWYIKH0ImJFahO6t
a6ds7OkMYkO9TvEwU2UeUsHosTQvuJdB7zL9L0dJWzhM3Rjc9ZqnZvnCKEUvni4X
i6az7C00oomQHeRI1FmiHTuzuD0GY3EhFLW0tZqPVrVcGXt/CnWZAl5HG2CechK3
UD8ezVD+vLdghz04yNWT3u+c72qlZnLUslilsZg458kZMeF2MyE5ca/ZwuN1gaD4
+bSnBKLGiWecaIbvgyX2NNz+6kN2TXYre7lyusMXcXGIlrIOb3Cwbo/y4wURBjMY
`protect END_PROTECTED
