`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6IFKeJggO1OIidr5LYsiiaR/ONTFRtguaB3cn5HNhmm+fsBIQZjIKrQaBOT1bdKr
R4LrG8pmznLsT0YIt19w2DGlEBVRnsE8QyTmeT4T2K+vcT3jLt7jRsJXR2f8lcOW
4+3Cjq3wzKcD/Z8HAt/+GWF6hqZO/QSr638zmGzGLslL/o+FCu6N5OSMjfvKBXKE
jIu8yh/KpV2RkAErgoAbRyPKDGdr3moMtl0c4+u2nj8KNxaAyGw1CWTGHXvPfJIQ
g/O0tlQjSWjGsjkiaxUlpJVnpuEQ2Eh9TIwxTXGkqtDVgBDmaLgFWKXhRhKPau0r
EhRiXTt7g4aR2xwQOPMdgjz8mKxk3VvbU5Z70PSfb1wi0Dq5YjX1FSYZTgLDFsk4
L24MFoYubPNXnjDTgEXHvmJU/jq1EYtpb3D4TAAADk5NAsksCYuIUhTpC0jsaGLm
0PHGkvWgJE2Z0ieWznMwwEResdHJyMMGJgg5Q05bdWrEsd3Wo46g3bJxTEqT3/QC
uuQDG7CyU7zLWnGb20t69HrQeUBihiwARdDOYMTa5oa/hHzA1ijw5Da/vMm/+M0d
43t5zkB5G6vji6YMRcBpUMh7ZxMPjlhayf9cn5V4V7EY6jVguQ8PlXxlMm0jFL/s
GAANjkN9VrVli146MqsKsGg30m1uswcNYBYVSpiycESw/OUWDu2TuETC/tXgoz1q
degm4ayPba4A3x0okTKC5wWZyzbNXtH4615ogw8Ui3BbbRyVnmJUwdCfDeTTmo27
phR5kIWzuQybPJwjOiJT3hVL07DhK3DyFPuTFMgVlDS7Ik+QfefGxrE9fdkqfURi
uUPtwOEzgGueUKCGjALTKDbMzMf2Wm663+sIXxDw39ssnT4jsy60JeiDGmbFNk0c
QCcEulOrpf4I5/GOn3nGtEVNfPzLjeVbG2H8btvepURjnpf3R9zVlCu6/KQsLR7J
++dFAMw82QYHRvAcdjfL/uieOjN+cbHoOBjrx6A8Skvb4IW6v/SEI1Rrwc0deOr8
MyYXz/FQp5qsF6X1ZzkiGqCaDEskjv4gFmxikOEzeljmlTX28IVQRAd9xW/Z2RlJ
nFECfhxKbaVjlQvPQt6VpukreCfqvjOiSzIg2FetN69/godB2t5GZe4lIWbjRg0L
YrnaJZ3RB7LobRGeH+HFRfB8ZzQLnSWNyvmCYTmlfOhWGZ+ffKJAjB0HCjIYpxfl
tAVquz9I+9dyofZzQ78sRoPXgxEwHpAwSjuDAg3kMPj9i7ix+fGNGb/UgjiLIp16
6cAeujgfigQ8jxHMRsRo2Aix7PKt0baLy9nkvWp1O3Wx1oILuBQm5ZtzOk0pX6AO
Gj5Kjt5WKqvL3UbUI1dX3SpFW1flwzJN9Pp0Q8RqFNuz76KySt8XvNmT0X4WejLT
fnHdbvXMgpNtAGUYX0wEGHqGvVBGE3N7x6CuYaW+iExvpLpK0+Fwy1YudzaMgn3h
ociak0T3S4mSU/PeBtN579rOT1avMgRJ/XxJbpUs6H/xxHODMLmYB9HEURXA/1hX
7Ebz1b7rsqXaRbbTTZSgoojYT5ygkQV/tqVzUhk1qL4i0JQ6dTZvpGa/aYcaHBbg
kC+VjJdZ7AYpWRtpEblzAQstu8fz+omSQaWR/FGUZX0PWj25Le7EFMP0D5YNT3hV
MscvQIk4BAJkbvGFyBFUpVz5KXE9SJtFNKZTkiz6019xol7KAQcpiVpop19759FV
8tIZCxOQEBui/l9JLiKPa/ru8Q/D9w+oDdOvoGdvnoHXoNWtpCp9/XIas7F/SlsH
MSg85iUm6+wJJm/nQM97o5wG0mxbsXIZu/tqBwQajVp83QfMLL1rXJIUPRitSjr0
JLPqiVSRUjMKJr47frYpO+LsX5BNUTQ6fXSE8TWVbqqXAJwO7J+pAfOkRkJbb6ci
VyIa937Tchh9ivRAfN22FG6U8XrcrXgGLN/JH0Ax9xrzGzZjpvPQNCIaNHo+ta7X
`protect END_PROTECTED
