`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vjQGh8djCGTGwHvOB5ise2ez7GXa3LwW3YE2J0vxPjANWPNjdNuNm3OY/lalbeSV
59HZqpuJl2nPlLRxZUeDNd2vPJ0UBu4bu6iUXUhyzm7C9bzuv+bpBn33CgSfiaaS
1CKFZT/scMWi4GpSeZicYsgbh5OIs2e+l7c/CnYg6KFTZP1A357iq13OlmQTbpWR
YF1KuJRmGHjcY3ynRXPjf1/i9624i7YARd9OJ8yPU9/nHHWmajYb+5G6zbpmr6YR
Jbs4V3BzFkSXVupQcgxnOs+x/+7Wy6JXu/Pepp7rk8oJ13zrXPdXphGSCi8zr1ao
E7XygvHhXfSJJdxBBjO4PUT9Vy/etJNyYDu4End1d3we1JT0JkXfIYfgUlOS2WZE
op69nSkQo6PqVxTisNjmGNFQtNSduPdnYLNKFpr+KO638VuHeS9ElnsLTrUM1uIp
d+6r0ZM2zvjC8GTlAnUvQ34QNWdDs3J7j86rhE88Q7ti85NFMmHB6lwP7sL9vhnr
`protect END_PROTECTED
