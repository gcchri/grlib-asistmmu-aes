`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9pMV6lihxHEMTF6UGxA+aluPPLXANTqL61UGBmwFNnK+AsQK8cXk90WxvW4mgWV4
DZ5f0NHCQZvEf2+ZYScJvkLV5BfLgRO8saK6fbgJ/Y89JjE5mkUe9Soj1YmVVHyg
yvsxDsZQQmj84Y3fIMp92OQvcRf9Rwv0UziD8qPF3ukRUALior+HIy69B0nFGc+a
OTusEZAkzW2PCK+VdMK9mgyggAbFdXo1KTha/YcHhB6/328k/iU4BJ0tQKHUHkH4
ypzLd4VNsJDilI4m7TTCHGOHErV8i6bSYbpKBvT8HNHQk+/iwAan2agSweZ1XM/W
S8Bv65q9FM5TMTrhY/OrCyezAqaA6R3maBEn+QjX4TShB2u3nBlT3YYT2JESYsVT
Bfp8jVpz9SMq3f/4ZiIyWsWi92j4IOE8HyJTGfAZlrSemjtIEitkwT7uqqq1TFuM
tWh/vWHzNJeipk1G5OW8woU15ZRhH7HUMlhfMmcXifFFDk4ohxYuQdJOsH5G2BGu
8m3et/Jfz4KYePe9uFhIt3FsCYhDtLsaiKSivJy7j/CeUumR7tc70GoGWZ8Ylxe2
DhfVQq6z6HByEC0TMv78y4/UhthqFRJx9UTYEY3e8DO04oyoF0t/V/FkAD5VAp+k
ztOf+QlzLSIzEVpsK1wHv5AZBb4REurfM0Foq19YiDtO9IFLm3YVgsYr7CNDeTew
8lt/7lQcdOQEdE2GLanFHjMZrGXzHquac1zlGo47DX85fvfZ5TqW3KapShgj/y+X
kv6IBSbrb9e1CBUetfnIgA==
`protect END_PROTECTED
