`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BkmPvLAf4RS+v14qMu3FNR2VMoB1NfXAwJVavWgPuknFriHB9cta8qVUqoG/4J9J
dZeD/tkIkmYMmOq+gimRKdt0/pnSY+GBUY69DMr+WlUncV4xNqBOZpUCC69H4pLB
lDHl93n53N7myINdaDgnebS9bZKGfUihAkKvYNfqtXxBGbwA9fXnwP6VhEql8SdM
J5kR1ZjL041FkI1MT8Q1+GZaOdnDcV/MOiO2pEsShEvtuCPCs2GBgwCU+rE8F10E
yuMglM1XIz5WJHRJ11D5tN/Ou/lhKqG8GIcljX5pEXg8q8SssjMBiTNqQcd9ou6w
Qy/NjIu9evSDD+OaoeMPLVgVDD9Wbm6lJCrkxjCL0ZQ0oDQhKl9jiH9W+ry/qMNx
ps300Bv3bUOU5Tjd6LI2E9OQgv6maSVCpQLCNDLFUvc45LcUXIFDDqBPFITKb/5U
`protect END_PROTECTED
