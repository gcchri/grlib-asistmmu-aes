`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RL3BVehu9e/zUSa0r7ikVcXA7ZZZvqki2L52vy754KBwpvWF94gUqWP+qXyFum2C
M1kN7xhhkivGIpnEs5zJ2AZgOIcvTnCKbmDBi5YEDQzMVSfcKcVHwboksN6UgwrA
n1UJ9CZMELfmRpRtFfMgtKWCDKban8XpnjXvsnIkrsOZ6qDvmxqFDmxyvKStn+D7
xbTbGXDi5XM87FKyjczSNRgRmiHSC86lX9rg9dOhHMuZr8P9enLP14quUBLr1Pnw
fWXeJDyKC2mGJ4KOeFN0qK09PBGsvbyHzbCM7I0Eyjl0NfBELPCACceh5DII07Rs
BiVP+a2ohKfBF2RW+C5ibwfV+ix55hHLJBdKnVooxXMHeUI9T0/kONzZotUWrVcw
CfJBnDT19nf8joTJWaUc3fy5F+aJaJASaoPtu2HyxRDuhXvm8bMxP+CtxQywt/SP
c70ZhGl9t/eWWKhW01WcZi6rVqt0zAjW14YT/ltheaXJoa+QtvqD1xddvhQv682r
YZOIU39zJ4JpExLdzBaR+tl1MReWGQ9x/E85PGMwVVTK/xPOcctSwCMQE1zCqKrV
7SEK+cWoVaMYBR1DMIq7Aqd/CwrnBAGPyGmDiSptiXA=
`protect END_PROTECTED
