`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ph//dpHpynJmyQVTwaQ+fbopP6Pq4maMNt1e5u/sGS8xX+DqPhlVCDLvmO7t1ztf
vddwPp157Gg9mFyOcJX+szQ4lDuPHlQaA/S4P92TB+t/ROf8mykDcd8Qek5vYbFL
Um1D5n7uG+FMm4huKRmHxKuJRHtfona3s65fPT38uC4XAcRhB2V/zbekEwIdDENY
tSJZjc8czn3pf65Tit1EpdFEaeVwjAw8dbAP9lDVLj5hYz4K4egLoeDCVItnDjH2
Li8XzvYlnchOBpOMPtVob0tv+FtgsHQ3mtP7b14k7VK8KEYdWL8nfSptMCEZG7N2
jvBI1/M6HUMdIVUtieWJsfJSggFr7H4NK+KY3h1FfJfgmdfLdowpJbGUL8cNGue3
ww1HwvWcfctayGbqAczdth5CfF4nb9AFLnLeN8Lty6xFR8mSrshBk/T8lYXjQai0
QrVRlj0s2HlAM44v3h7wDuZQX0FfxFBSUPegFNUkYpT6i+FPUleIP5FYpcJMJzl+
JentgEmnaHYoRdyho8+192dYVwYwUl4aIp0ZftGGbQ+Xz2X9uzaM+47C0108NCrh
mRSdqsBj5vUufPmG0LQrP2yQ9JV9y7I7bVhvnTrHw/Jt2UbyPnITSpmPeXu3bk1s
36T7NSVrfCGfPY+C3t/ixFJuNoj7mpU8pQ7yCP836Nq+vdg/TfaGh94EcYY14QIV
/2U1WFaP8hWZc07uUj9p01ZZEh28rkxGTFaPF7Wv65I=
`protect END_PROTECTED
