`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gsbKK4BscjxBQAKTp/jZMNXK4ZJ40c1rlqOlfdYNnWNk0F+0/1S5ihpUkMALfCnG
LPolNUccMThwbsQ2xmzLXCLdv1Jlc/UzQ/9z20fcofRDxO62vpsfhJmzRJUv3r0L
Rd19wBAYyyjd3syFpDx1PUcWz3gQGUOIIA9WshsXLdEWFrpJjX+yTta5r2rBX5l5
m2pcwVGUicA6Kd0TPEFZvWcbsGneM2nwvxGhhol0bqllsM51os49up/lZMCQyIlm
+7tgT5859u2VOToZaE8c6lliIIU/R0JYftTCSAQdDfTqZ194BESTtUTmzIqW7fSe
jiEdOhVYliGpM2aGeVc95d/EoxhlpxxG64t4Ymumi9E=
`protect END_PROTECTED
