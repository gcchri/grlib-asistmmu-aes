`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cYnWeoyH54vPrDLoq7aDN/rBG+finTdorQ0g3vnnzMMFJKM3qYelyU1Hht09dQoJ
bAYa2rfVmTs83a+kd5sJEk/BiwLugKFn8yDT1v/gmbBhB+yZQGXDV4I0ONz9JkkY
GV6ynuzOKGxe4ELR0eRoA7nwRFKGtim34vYa1QsI6zHHAjAAuOkB34IgSFH+Z625
b+THmLT5CfjabnRJFaFvXRTj/qxGX6GzrHDZ51n2oiSTPvMAeVMqDmdWnW0xvD75
0uMTvdRIIxPM1a+KlRX5YEtPwMjzHkJ2RTRPhVvDVaLJnuVsnFvUxj0I2R1vVXnE
cE7XMZbN2DgY8IMaj1pL/Cj+GvyHn/iZ9GqwHzVjoBLojNu+8A1vz6lNGk0Bdiwk
ulDrCi5jPfm+GZMMWk5zCFoPzCLOitiiCC6tFoD/bIb+dyFkqBiQbUHI90Lx/8+5
`protect END_PROTECTED
