`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CMh29AVjTqPSreCyu2TDecpP790XEcoBwZLyZaDIfZJsyrYWLXNRmyFrEm1re8kg
RGUOVpay+ByAypvcr3jWID9Hoq3y+7PVWd903tW2KInerr27sV9b93QlRRGsSSit
pEqiiiKLCV6RtVmOi7F1V/24nRgmmI/+NfrFCPbBYPdnVqdrqPISnN0TbmexsYUU
yFT0WOS/rY+Dt44XJNFJv2+lvmkXzd2GBOOe4H/NQ6oX6mn/qdAAT3KPwG3U2uBl
XYakp2QRXvZTT/9A4n/BkRf4c3hbFPjowe4urrJXIvQKXanBRBWPERq1rw1lCwcc
HWigzHS4NNLOscDgVzsU8z5HRqS4akjn016uSzW/oNwpec7NrOifB0+FetEEPcc4
0vQwPuuOeUvsR52IB9kTFUx4z4fz3wC8hko9XjJ8zlKlzp+YUy2K+8/DTGRuJDyH
`protect END_PROTECTED
