`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lVOZLn5BV267PDsNQtwrs8eGLc32Ty/lsavEaUTgSpRUxLiBRHb90ullyzAofKNp
l6YCZ88tFkmClbObRBL4Uvk8qn2ird4rz6DRZCWIIMLEnmVHajSmxaIJufjntUN6
DvnhiiuZ9/KEYDT2mLLEL8OW4TSZ3SOvmr0M3ZH9WTRkeDhIevo6dlOTwtfDNaw3
lSiO8zUbZUzcuHsMox0nHFAiqkQuuf1aqkaoKDRNAXgSl8mQDtF0mjX13PqGxwbX
RdheoFUGvJs3n3TztzYPGdENMY3GE3ebYHrjB+QGmh6+/MkMUUNXpd7k4CXaOaNQ
Oe/jtTfBNFNtCnizsE95YB3gf0RfxG0gDPJ/uxyiQtKe7H1kBwM6JbtvpnEBqPsh
AU7anRD4z5ojb88+g/oivnIwb1iPzK5sOg7ONPJbaF/zcqm4iqMFjOSeZGCO9nAf
`protect END_PROTECTED
