`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PCryn6rAPWZd7zcWTPJYFXB3B3yEva6EBbh+aEdmIfhknONeAfziusUoaPg1NSOM
mEdKYXpVsbMu/juqp4+ixSv6DvW1NGmgGd8vGAbxsMpxjW2r4NqACB+LOYg917Nu
iVezvodOxnymuGP0ng4az0Af734Rn2HDRxOxLpAi40O1ANAZ/yC7BY/U44wFEFEL
SOXJD3hVUdAFPY12ioGZRVQQlVzozHiODboNWEBBG7TDZcRiYFN1aR/rHv9ZqG1R
PuHLUgsgd9pW/APfxdOBgolbQC5jMCf/JcSSiwlhwKXVLrdX+q+dmlKAPMMJ6CJZ
6TXlTS7knD1ghzun/gzrueoTkyJ4ojuSrVP4eMyuKlcVRm3M2sLjMjUTzsBneX29
NU1nN09AA1uBD/3+aaUNw8c+FloyvsLb4nJF/lfNTW6sendOyop/fBpto4ThJ/RR
IGgn+pGL5SeAMgVtRqrzj2COhGvKEFAsZwbomAdtFa5AWAhzRY5tYWZhh0KFon+9
KfKK0EbhoeregW+SYjJr203BYO/1u5V413ITKaM6zL7SmxcgGAisuJPf01Nh1Jwu
a1trqa4B1+YNu8ddhRJzfnlqthPw+F5FCCPTVu4Q9zHFzVHtBjKyoqL4nJtq4euu
Ka4klsVepBYC08yK5Y4uIQzkO9bXLih5Mfy62g3qhpuTiAeKhvy3Uhj0Til2ReU1
t28BqvTsUIt9lJsyW5drEjkk8uzNwoAFl4Po5qBw6HYPdpTu/qZEEaBEsCk+v+CP
2TggByNTSdS2csU+2DVLCc3HZ85O/qWtq/5fcFwcnaqPf6CWmfux7xRyZuxK82G6
zGMqxiCELRM58RUZYs6b8dupXeRvtIMmUM4TQVJZOloNAT0+SCybPLZ4ASxPWddq
Vm9UvcLbwgsFerX5rKB5zpuTydBYjq5xB9h9HIAznV8XwtFcPEAsBKjHnsvQvwv8
YQqNn0KS1yJTOX64psR/HnZcv+ln5+eE/KC/B5MviplwvLiQfUmDQNJeF10n1f5O
UGLmc/9RcTZjkd1RWLDM9ubpektxo5j1pNohP4TSiLmRpSJwRXXmki6kl9//amYI
LMZB0FZlklZVbJXLQID7eo6xkriE8/nmrIOHl0jnGdpitnmECIAODok8CPDjMz/J
ehzoQhl8cu2VkDYg7TiPMAUKXfW3qG+hIsy2z03tQLr+gxwtk9ybYLt+PKk3t8PW
wXbCbJ9hcVQHtaXaJUNBnVBBSJG918ZoX+rYvAR0myzaVYkcdixQXz85xMAWQ4M3
JF0PXp9FLtOf1WPJA56wLCoNHIuNuKCGjU+3dTZVafG5W5jn6368/YjJY6MeT4p4
/XHJ+10NUs+sCxkvVQhw0v/UmMFwddnFnAcuNYCxl3uYvlkTqmLiPOM99xbWUcPe
Ok1UgZOz6KIzkUFXoa2h66cW4UuFXWr1bmpDE2HwzAZ3jBMzBCHGPWI+8zya8pkU
CEwFrJiWvArbQ+2mSOSsm0goF1uXwtb2n+/fzLkL/8XmIRUVsBHfG4118HjuMVfB
Hv7jQ0EcIOpxRXezHIGatw==
`protect END_PROTECTED
