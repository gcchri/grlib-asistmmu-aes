`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SBH2FxbhG0xsYCeiMmuEBXu/Z8OD/247fgL3B3l/SOFzn5QxQueUdDe96sR+eHc0
kdTHC6qyfhMtsQHrQas3GgB8WUfl3ZRqZjR4WhaT2W77ux21gsKbDlZzPqPt6OVw
tWk36ee8TlTcSbtjFzOZ4931u6yfEXiLmqZNTUgwG2M2XCwEcaG7dv7XWE+PZoxs
Dg1TfGyQ/+So/sHehBMg0s2a85/FTkKHSvZXlIYGIG0gNiRiXMeVI+zNyp5A/Tdw
M2k6R1ycN1GTxMIWUcbdhekAZBRFZ3tKKhISMloxe492B9ogbQaE2w2wGIrvLWsC
4XSl4gRZ2yIlKyGLv3NyyMwGwYBgyVgoERhJEmq5PjMZdhCXOFJZ+tUJgD6JE5Dv
`protect END_PROTECTED
