`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wgAb1oH1zmuXcvcHyIRx04o4Z6exDAS+cGCfnS+WTtJcDghoC14y+d43EfrZVwM+
qXOd254KezePq2TDdbnxR5HZNqa7wdpKQqJSaTfW74ewFrdldUmayNgeZw/l9F1v
t3DOsM5CFCLUAS8TzZmRHdpze2PXJcr6KhHhlD4LrsgXq0uGkzXEtUcWwWFI53Sn
AuBZWxwnc3wPVkqVIcCb869Qts+9UmSNLOAHox97dlMfkeOmX+Xmiz8tblBAUee4
SiW00KYXpOr3f+Krz8FYSWSlLieAeab1BliRJclJMx/8YRvHhPyDbUUgyII3bWRv
54AWv/WdoOFeiHDLkdOCSQKTYvJpSoB8ibO8GI+SXAHV3kbzsEvNNxRIOkiTTSYN
fgxuyfCXRYfH/MwBr8fT+uHKhJWSvpsaPnc5z86eE/k77BLZbwDzRcpRlWDjTcKu
8wrLKpPvwtDc13zNd860McuG76fy7hwaVLkqIcw8jSLL+E04ih0S703fZ9OUeX+U
LNijeRE/RyAMowLwSRfEl9Ny9lzoTfs2fFllPoHZncI=
`protect END_PROTECTED
