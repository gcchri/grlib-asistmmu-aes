`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NYxHJlU45eHBsCFnD93a1Cvxqu5l2FXZYeifdNzQAlNh7XzFjPbGsZwvIxzc/Dhu
FZrJFjlVaos4KFXmlUPhncpL/NCU0HZuTpqJtqnoBp5RsDezPgGiRFawb6SDngOT
3qAP4HK8CSB7tw6E5ZDClR87mznVxQxInoeW/v6J0nUjRpFa1KxVQlhxfoW65Bnt
syYpHSJyc+wQZXAuiPFO3utMbLvJsTOhEQXDaZzsTNilCA1mnA9H6/Tve0G2usBA
LbqFgCelUarVQKDrDqK8nChkM7iZK9EiRyoFdq2yTkafgv/G3/8IKS5w0Let110b
ybyTH93hA7COXEQ3oECin9qS85iSC6TpxA8K1bPCNGPs/ozF6Pyadt4muo9jef4v
9ccDwOiddSNhcSwkN6hGVFvklcKTrHfzw3iXDcQ8FLv9jZ1SWkaZdmL2quPMI27W
S8QihL6Lob30Yqc+/8ZQJ0LLcZcyWd78DTYiiNiJGNNT93LKjDBj5Usexq14brtS
1hlh9ZWEn65OVHf8Wh6UyCT+UHdFTs/k94f1XLTcXXC90r8bvbrQLQTva8GKuKtU
nIo6EtX+pdZRl8cSN0OIbIc+Vze70cMlGLEtxbg8Cr1qibVTseVsu0HUO/YDKmUU
dun2B0sZLTuS5U6GXqyRpQszBq57Wx3oeT7ZCq7dbZvMPMoEvUtjA+heHEmhP6VG
3QXU+rDmVTl83uoyvYsgxZHa+4ZucqyUxT/HxZsSwsklFttNAm9+t7QVjo2+zQGe
GzKEbWbbXpY+BIMbawy7vde2eGQzJY05NiYOMBW5Z6O5b79DhXTroF/WIfIfT80v
0d8wYnpKjoASEgeyEt+MySstacWoHJ8PQCWyNhcUmqCmGq9rzp/7+f/r9uw+6WyU
iFnVXCccn26sjA4ecWfM7bk1IkF9URrKK4kWiFzEZ2/4NGLAM6a062u8MTYvZRDs
`protect END_PROTECTED
