`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J8nDULj3Xb7H3Bp+A8fsw7BCtmXmuEIHr1lh03UG55xT1i5v9vc8soBMoDwvtkYd
yHRfXa+A2DPjtgBC6yXXwoMSm2ZyUI1MlUJnapvuYYRzInWEIGXgyibmsYaJYC2W
dpbuWgqDpelgUjAe2YmqpI+sQy1lzNeLxrlA5uadSoyeXAAJlnti5mh+Wtpu1ZK1
C+RBBd+FF36anDBjtgOrLHDRPkq1vopaS/D8m/VNnCAqBofhg2E0iRikeoNZaoIZ
RjBOI1Ugp+h+Yc1C1d5e9evyCL245+FXfq0CCLRZIkcrw36pEzQbwwKFcVc7n4SM
1JhEQEV+X1pZyyKytFWE26RK1FEw9g97ZiJ5L6WF4r6nYz7ygAZvRbKLmpIMRWH+
p3TfpluRxhynNozKwB3xE5Fc+D8BniyBilpTz+g3SotKVSpRuM+ERC4fSNuN4Q3U
HYnnJwIgMAft9xzQHgDcaqWkAdf64owZNtfBhUKrd2+nseh743GDlCL59Lmz38xB
FiCTjqxbcLm9xGjqEGRvyeRqZk2L/DwSyHeIJ+999rnxpbdHPzl4rnPQVYCu8FG1
c8KlNdGtxAH3EtS0Q79N7V8aheRNmtnEHTrQC3AyVDop6lFYwWRKsnY3xUDy2G0B
gQGMahPATMjEAizPoXeybRwj23UYB7EKh3ubfOCmVQzOer2FLmjOCInHynVsHQBB
oBg/x0IXoQ8Gmf3MGo2NHXNB6daXLLoT+6TEuNFbUvW1Xm/T8L3Eyug+mU/1fSAE
N3b4l8lhMOIacJZZi8jRFDBx9pfxRmlY2KmYtJccAAf6DFRAUtYyxXGn6pq4Ozzs
yi4+kdBmpSWAGDT1DhBiG9hZLOBeIVeF83et4nNVmPCEXYZxyiqERIet9nHttJfv
nMTskocKLkIvBULQLSb/v+SRjjVeGCxNoYvuNyejHrBiRUmV0bLoqF6ab/8GheSK
lF0zStWHj1k4IIGglQBpghJ1sC6bFOr1nBOjvfe+VUc2zuCBHujCoyoBCXpc5VoJ
Z06w97z0uGVKrh7foqqR5o6vTiN4aPyGdwFFkjdwr50dORKUNhzrUh+HuJPmg+V2
ud85JJkQ7gKji389z0u9ONNAkt6igs6Q/S5k2rG05pzeXBB4aaPlx7Jm9U7Qf63V
0t4esDbj8+7aT6Zh9zl8IMhe+3W2pDKxtLCsX2MT8IgCH0qW6lPo5AOFeGKN33v3
0rMqHngm+8pRgj8X2i3vf1GpOp44tB6coA/BYW1kG5j9BHslTOXHqoYSQ8+fHNaA
R0RQbZVyUl7VM/4V+lWd4MbzXIMZx9sPoFYlGmizppyqvCiuvexFxz+9xRKMPhy/
ROxJeme8NkdnF5IYin5n9+DBqIebZJYOZcvRJy1yzHzffil6yUsVo6e+3kwza0jy
wNQaWUdxUgJhx2gpwgeKAH4k63bDsSjSTCyAQ+4VL1Tvhkm3dPDy/9y6rD0fMVej
6K8RnCUDdYly++pQnY06HW/fdqiypm3gMFTddNMYLF9Zn0fmJQTSupfE6AyKiv38
si1MZpjzFYx4PO+4CBaAo/zNc5BK1lw1IoWjB9Pb9fMQDGXeWlEqattAFUz49IjS
X1gyWmo03ssVWV20kZph73n2cEg/xiLnzySZuMnycXuo0IGHvkGotgqqEC7MQGVG
hhNpXjCKGZKIDfCZFXmo7tFyk21hRr4D16OiB3E2HQ5ucOHZlSmOb4BD6LyNLrKs
YWzdUoo3aMqZujyp5D0dId0Qyubn9Or9tgQ5N6+qlCgMK8htfLc0//QkADmtmwqt
ntYZgYQYbChZavZknCJMZ6c2HGuar5845SxZqYvpSCcrelcQ9seaZm3v6x1KKNis
d2WoMNiCu/04om4q6Wq2yTlv0QhJc/M/RclVlVwAPubqayS2J+jJ72cfxI4ELxRt
LvEQ09Oz0zcjUegzZIySMUXhEp6lURzrHqXYc6bddtAiYmT4lLGw2Z0bCS2gDW0w
0vvM4+qgK9+dbrb0qx/5hEQNh/6FnSHAhrC42pdjnhfcEaDBPnZQNmFqZY3xeh6i
3jcKeShJnQ8ODnah+Mmpj9nB76GADsT1un2iKDvkKtqHsGqiGDNDyhaEGJTb9zRj
zF0aNIiBHZensq4ROn7GpeIl6G2s+LnGiJDSkiMRSt1JllswRkUcl6Shcrz3avm9
FBzrGr36Nd8LpGzgzajFCu1JChIvIF9X7XqaMAmS57joa78UcOGUeqyHvg8iZaf+
WL88OshlwL6U3sZl7MW3fz2MQee5thtknTQXCT5BQirAFxoAOXFKh/Jd+AVLFJfd
iyWXGsNF/8i5NL5PMA1y5vDb5DAdsE0boYDDMDWQtWOA87Cihi7uhVE7U53GBw5i
LuxQMowE6XD23wJPNkxJjWzUlD2OpBwuPAd4B+xAFSfxOEorTjKygOvSgNLO7+rQ
XjTmqy/QmzPLUoXskNprujFNldayhjDWM+Ks2qt8SailLmcOS3zw/su1Ehb5+ym3
`protect END_PROTECTED
