`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6w0O/oEMv907lWyZGoiTT/wEfh+0vkUE683GbU/YboPiGcDUwAXYbjJUUcAY+c2l
Fw1rBmgA4DRv+el6po1sEZJogT5AVWfZ0OpPd9e9jop8jhifKYN5TkguEQBiKfmT
wRTtc6JVMTboe7hCak5Nw5q6cUrHSeUUfMR6whKOIxheLUHlSEvFmjqT9aLk3927
3SkpiG4Py+G0YW9fSMtII0pp5A5ODVaMaZoivQOUTLPwd3EPmqw/4if4OOgGeVen
eZ9JafaOJLgFzEkqeud1c9m2uaTjT+9WSaivPV761TIN4SD6V+1iMqX00tLTOfcY
Wu9arwGw0yyxJSTewStHsUM8mgyI4OP7ze3KG14TWFkLbif4yJkF/35hFRHAYgNW
TWWkVTDQ9wlM1QW0L9AWqSznv72SeolyZBKYK2mSsQkrnR2G/0W5xyH87MrNprND
uXnSJHJDbD0RYBeulLVKWsgxiWgv1dQCpqvMbjoKhIDn43uLDwYSUcQk9byhXVpq
/sod0heDnVTq8edbEK8ep0iPShrELLvXNIJ4cQPjDKuGYFlJ7DDU5oRPHb/1XA3R
9y47mgG9svzDWJrMoVZ79Ly6pmDhEoMPPhPtQ1zexCRpSE9Eexg9jq+CEFD3MA3+
/kknT2lnhBOnC5HPu4wHkBc9MLZcCOXuGNSu3ns/6HlQq034ivVTQBgeoVwFh6Gs
7HmqIW5sursmJmINi2wPgNdHCbZTu9vsEoNyuhOAKL4dffQ1m/FqcCOnOg4E+DKW
JcA8T++866900kmSWI9ehEsv2FbzgOZ+sx+nU4ZHmxytRbtte//skFNg3VKx/B1s
PqwewXSw7tUBPr7lXNnrPzAMVv8Tav37BJm7FrKm85wwZK8I9L1KfQvVYzBGhY7q
9tHlnympV4MAARVUWdKD2YcjuKiQZLxENcw82+YOf4WDADPCcqDQ4WK2hOM/RPPj
+vhqw3Ly99fKwrDH1ys2XWSkAoebj6s86/KzG4FJ4m0VlA6w017Y4IS1G/nJG3S6
0E2C3+dIDRmNiqzzspmq+qLEoS9zrHMVasc5u2aiElpfGut6qYpIbDdfPZ9O8U61
Hhla5UlgfdQ7+kfmmyoV5Zx8hfjILcL+w416TWRg/bq+7J3Nzkfjh7Kom0DkVT+R
Wliv6NR8KkXRz0fzcwVbYQaPWyTPui7iDtIAWAjvQnI5MCTVpS1e2AeVjO1HYHyy
91f5CgztRaiJikJH/Or56AinpY10qi9uN7/QBHwV6BuNu92eBNyWdY14HoxRRohV
acCzI4xMj8/RJ3QV8j15XQJkN0Xn9nmVUGh8yX67kcrHapc46sx67XasLUQEIbjC
MY6VFICqi3Mwu2r9fNgp6JJnNiW/nBGRQ2XSNagnKM4XI6Gun665wnKTQnqTjykF
4Bsx9bBW2rKJ6WT+YDYGE9m/YEkZWmIublrHqPwFPEG/d/viWZO90bNzZ6Oz68wr
FPaNz3MP/C9d2vnomVIkrvLQibHTYKoa0GVqczCEI9lvr9phbwZlvU3FWunpnCC/
VPdd7g6insbMc8lYDRBVV+CbW+FVvOnmsCRNInR1FODaDjrczDgHe1g+61WFTO/s
2B1aMiC5XCkRljt0F5ZtOl+ucM57vig+57DYAamLvPYj4oZfFcJixWO4Mak5rw30
Bm7WaOKqaIEMFp07BK1RXdm5HLhDlNUrBtLB51ieElpTRKlWHXX6VlDIAWRxn1dQ
Lsvf8HOmajKbHNWN7WFIOQxygeMYTfL0A5JaKYphJ9Jy6+iV0OAnPqHsPpiE8t2A
htRcYXsRDYbjUf9DSqgrC04O+iepe7zuudhNJpoDZkMlPECOe0q3rNPWLBz91ZwS
p2WFMckHQ0tfPTzJfOVVE5WaB/s6eI8FolRcATQ8F2MEYU6laJVppA6ngCznmC5J
fd9UEpOlJVDCaOi1kGqfsYjj2lu5U9MLD2Y269HoNHU+xsaTbJSo03wQ2980KDpK
ohQIjDWlbiBvqJs/FbWn1rVdvSK3fGgV/aVKWR0UNGLqx+PtmNmFhVMOtBvEYvJK
xlixy9uoN55jO8cgSiD5y/Nl3JT8vWgBlNMM8kk2fet7J27UlU6dnEFoepnsMS9Z
JC92ErqAhgy6O0zaQAMHOKcUlqerTsZuRC8cFFG1n/9xbvS2DTXGnVF+LUPpof4z
YB5dULG5lDpC+afw0ySOFrnI1Vnl14EoUry3wCdDQpKUZ41FSNle9LMLAb1MROce
4zoHVFgubgBBeWlhwT0kb9YwnTJmJ7u2EEfB3B864QnNd8kEm7+30rFau7v7nov9
kwkfyHoRwxv+dYG0r4JUY2t1z5soIxFsm3LNhCETxYWKIW28m5qNlhYgPF26UKOr
4buYVKLY/FNZQ9f7ZfNz3FzHI3LDRvDilzmCwdVg3JXtvUQUFOjev4dbdBXZ7iFb
S6c1QkRgkxnHYOjY1+ygRtO0eYEXIvofAJophhdcmy4oRhZZUKYNDwDlgbjdnX7y
R6qIEzTCTeNV6p5J7qbRhTzcC7tEwdFtFhKw4yhLNQPioPJSQpwTE4BMofgXhHLA
6luzNVVQIvWRshujhlal84Xd0vqA7CWnu/4HQMN1bPYrqyR3RXG0Trmkvu2aJnCw
F9/1QVZahb2NsrEzLYfWA7kmZ8NqO4eFXfE/CWpS3KUTUC2p3Jrbo4JrI03C501n
z818fiTuPqCunONS9Yd+bwXEswYvR4RuVQdnWO1SmTp6HxtQKztMUv2zpOT+1tVl
vbiAQBzctk5PuhMjgeLS0YEkg7hSaWZhyN3QsvaHRCYWp8kb+p7mCHVXh/WmtOrS
Q5+Kc3MyC21LN5trI1JfFOYT49RRktYvdVLCluhHsZY7VjaSe2Db9k8NAhPkwYPw
ahJMiUQ44dHSqe3xt0lDCNMDI0LlmQgqCN2LvlRkNF6mOpUUejmmK2sCragusgCJ
9Sc/4GNb42moZP5JWOzTlklu436Nvx7vphwzAURHnkAKLFKdUBJji3HbkDDnRgJB
MRczh8bG154XEYutjuj910tq4NLglRpWMY2fOB8N3jlbfAMcwVHBFWo9cxMvVk/a
BfOwRJTas8XkU/iOjAT4Dq+4tW+Uf/jcfUO7FNrY8Bliy/zinQUEv2d9ewVq3eGe
WTBZt//ndWkgByrmMzNonbZgsy2L9TdSPJtNNX2NH4WxW7bkzqee/pGZC20/J0Qy
KX8AxdRFMPwJsq0hrckkiW9U3pcs2YvzKqT45jkUbWUZEtOtvylCOOxxVhcF6yzh
oyrsxXyH4A2ifPq/vh7f2V83L5l7oMaMkNDKyO01CEWnsC5yXZ7Q0RG1Za0yHdjy
xl+oYhFrMnuaHxkjdMC59ABImSkMg9K77QJLpg176S6KXLVDxH9PMOJTGDCKG6X+
e11NZJM4qBS66E3B5L57sQIS0IUrPXkCW/rRMEkAQEA=
`protect END_PROTECTED
