`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1cVCq1a90RpGjPnjZO3+jfoJE8ftjPCXJhnkyuNEz3msZuIx1JhcNgTAfs9LY3jv
8OpGhpcbIsK3stjbxNZRqDU2aBTOKyX5hMJpgSsOR8PpjnzkKYxbCBw3xOY+7Vqh
fRhJ575H2xKhV7gAYid8ZK1xxfGXMB5uarlhYT6EqZ8Ndp1bSgOtGJrBdH80a8AI
V6EABNNukjYdU1JymA10BLdoCbS1W98oKoI0hHMpsUvBlw4IOakNuV/GNM9carij
zTHlsBYhJcH+HVkzTKUlqJ4lc1+tKepWjRfbPMTZ/PU14Jt2ko2eb8Y9RsTar1+H
7reJrao5RUhT2VMvjqTRpFVuZXXYp4qKKJp+pt5R4OXHzq+mkO9h8YjaWi/TJAMk
`protect END_PROTECTED
