`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3EFxAnNt4DKGvvr/h80EC9DN8kgDiPfLvCtZ8kf5/lE+qKr5QHsXpBJujxtI18ZA
C93byUMCra4lGL9MXdixciq7L5zd+FShr+zozJNa3OgaTQOenIvdnbiofl9tgKAM
5MzgxVKPTYbESegYlNOH5XvwA9J6IM0rVPtEpXPv+4D5VNdVOOPqJyMrpGzv+l+3
yHhRXJ1mM+mpvzrT5Pub2iwyBX1Umpz2uhjE9wzRK0vjHntO66KIi/lpKbYoaaVn
GVQnohT3OvGLYdK2BeYDFa+ZXrd8C/rcBJUh+KNNns9i4GPbPiQGErwoqJ27iXlM
nQg0fwvzBkrIisb1a8f7Sxj65W8cIStlKnSwZnUGP2amOAgXELTAGrl/8HlELKYS
27pQgjzwQWoMbsnDRwfYT5AWBklgFNgIHktzNdvnsbVsGRlFBhQLnnBS6Mnwbw90
Zfcmw0Ixxtm2EE5FmD7JHQ33cEqKea/6MyLJbmDbLFop9NEhA5gQwV/FhwGHbucP
`protect END_PROTECTED
