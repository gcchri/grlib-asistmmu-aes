`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jQh8VMPa10KlNMZYCstY9wuzzvGDfVjlz3483HIjAwLSBBzFIJ/9c7IkYfjFgz8a
0/goB1EREiyUicHP16XhykT3CfsMFWQNltK4foehtXi493gOm9aPkjALw6YqgXJp
FfUDiGTlUPDvjtzSyqG5QzKRkxxfdzuIOZgbk3dlzYgumGLglLhjhJtBCJSCd6hq
YcgrN8wjS5NSdjtmF0l+fGBmqdEzw9be+x5S/s9dYxLQ6ec2wRZ6xZyni/+jBSwq
2I36Zkx/DMv3sJP65qPSPb80x4gTS4RKKXQvrzPCZqBD64lC9ozCeS/L/qV8u3so
`protect END_PROTECTED
