`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QebKvEAx0QERn8zbUXsuGxp8aXSJUy54KLFhav/XmMd1E3JlQ87/lStNhldfayfh
4T1aK6UCYY9Xsb5PDCOX77zXMRoTmVHQxvgjr9U2HDRYg8lan2nKjY8pdirEhMZk
J5nEG4dPMgh9LxrK5VslWqIZvWpQMVUuhMdqWxCnHLRodDA+5guUzJk4KXWrlXNn
jOqvjlDjJsbPeqv+uSL5SyeEHPWb4Q79E5ofx8V89ES6bskgj97nF4rBu8I7xhpu
0ZGsAuyOmgDn5hX3rSM7shpXQTA1oWLR0ET7wKRPSrl+6vhwK6zl+IoA3st6mJhG
kRZMQujEj6Il8q7O1x+AqxE27xVLWyWRQVasTBf5Vr6U6nC7Z/W1IXF+PB/yYMSA
4JlqBqwKVZhLE1353kzgxC9nphv4Wz8To2iVvnvw0cEspLR0AxX4eW8I+kPg8F18
fA+FCFGGuW/6QsYG+PtCI+j3Ey3kA13Bv83SJcWomG8RTnR4q7elT/8mrF9Ubiux
5cPUwtn4uy4qS/DLYb10uO6aBAUYpBmLOyWn8W/8oSH6tRq9S5AKOkHPy9OC/BbS
rBlZmVb0S7yynSy1sbYpy93wBjlXeKZ4xKseTs8T2rFmnx5mNegd0Y5y2hzsDie0
z5qN/i/MP1BRawE71quxlK0Z5MCSeWy4rC0YtVU6MmBqTLgV011ajUR0+hV/Higd
ABxSLB9jJPky/xgfqmH+ZXibYUQVRgcos/g73S7AF9MBVpafzV0+YQq82MNXbwRt
GWlZpNGy4r0Q7BsqxJJyAHTKfIB9YVV1PQfjjRQFZUZG13wP4XZ19fwHip5KYJon
8K5QLJ3Owu1jgzO9f7q27kMuM/H7/B0LVDw5qOfzDAEbq4R/pe9WlCu7TNl4RUWF
7nOxy8uE00EKgDrcMAhVUOdv54yRmiAbGRTonJoBIj+qIMtbc7M2NtNmGLCFfliE
V3v6ujEjHbEfVZetOo2jE3Nk6RqWf82SjycD2IfySv+1vkxjC5Mmiq2fwG+MOgGZ
u+R4u+Dm+8iBjenHCKuVJjRdAQNkcRO91WBhQvEHS2ka9LG/JDudAkK7DYrAXtgx
sOgA1fs1MV02gerl2LylvZa/gTs2Dbfqjx7ukcxwaLluvWqu6vfjAwi7QTCCNvKA
7XwjTUVNiAQyeCxCghYZGq4dvuWuJoo2lk52QbbYCLmV2uzQVha5cDRlGNbGVk0D
8bwwfcnQZZZnQvrJzqBb1x2QCKgNYk0j4qMjKkZbPCLnpP/XfxZG7S4fFvZByOT1
3eCdXbWRlcu6e9IxVWerGaZBOJrE40HuZUt4IETdJL6vT7Dmm/Vj4Pw/FioxEkV+
QyLtStql8uGGUfhVUME3TlC+ESb2Mi0NS0VkIR6/QxvEAv4/2rWniC/vpvpYG3Js
ZSMLIygvO5OSC+XpZkiIaHMmwHrudRqDENJdd33U/Hp9+p8G/WsCI6MqarYRoFtN
9IQCqlpub1U4nUHBu57/qdpiCLLdsfOJWudJzqM0w6/Nqld6WTF4AX8dFVif1dSG
lAQVrQ6su0MYyJIAkOZWxp0ScNb58+n/HoS6cuicDxjmKk8Lm2kdz77BXzhhOaBg
MHom1WAAXJ/X3pqHP199oxL4m9i9zIpZ3AHK8tKxTUKcQDQtLkOMlHpqFnPHRmvt
OEVL8vpfS2O0EpoPHFSMEZL3j/ZIojhUb1W+Lljj7VIY07YtP7WWjFu9MThhxwSq
CTKGpsM3nTQmU+m2iDZUCOvytyUUuZmPZFk/gD6GonzzyyeUixIf0d5mo31uOuPX
1GdLP6Z1bZEhg6DHEGuJs1kb6prpuPcksOHU//jKwe23UyZ5NLDdzQnRgqxLws14
`protect END_PROTECTED
