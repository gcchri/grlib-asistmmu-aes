`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JMqdBiU6hsTBSm0d3Zo4cvEEfd3u84dM4d/Z8qKzX236dznDDb4VGJDC+T32kLwr
Uj6RoVOG3CMlkZh9QdjDiJVJc0lZ3KKCGyiV+bxu+US+SveNF47le7V7Sz7yjcC5
218gXZV4TLRIW0HYNy9q+JjkF7pT0GY1eNi9M7miwzvInEaQ8mj4AVMHju+vcdnB
dF77JvP4kT+6qGQYWXRMlQdLFk3iN1wP64g7cxQAEAGjLqBCOzLLPvAzJkdnEw9a
6sXfiTUQtoke7OrmH5JFF0BWGdHkMFDq/rQA1GkalR4WUSbeC9YURPJkfntnLCHA
7/x8cNSg7FodEVGEtikY5UwPO/n448hVLIi0YralBxCdJQ9U/pZJ604l3HlQ1Djl
bQPpeKJvSBfnO8jghR0OlXy5vueDb2MmhrX4+OLJNp8uoyBBuANaWAaLZpP98PXx
ETbVlRBphHY8rzs5E+uRCMiCW8cbohDDg5YxxaXxQqbu0GmCF52nPojYF25fEDiT
p7JgwQtvy4m6AhwnkFbGa+k9x6+yu2B9Wov/1q4h63D/UUCRy/YRWghNmEH3660u
nQSNH7HbygPyAuReDgXocREPoA6Qb1dh2tqXAIpQMi2WxIlNXM3FmSMzi2TE7ZSY
c4epaRwCSFE9lx7n6wolh9x+W0+lUg4q4qi8bqsMrLU=
`protect END_PROTECTED
