`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tGXIpHJJdvC7oI/rfIOnlMVZSNBN2R3uisFyFOwgfuqWcxdBp2nkXMkjTzm0Ok5O
BdvWAlZQfFRo4gGiuIIU5grelHYeCo2N9dTs5s5TrPff8Yn0hnMxSDFMr028iB0W
JcDYwz/wewXws/lfH7lfwJFUwrC1fKhsTuA1rumrb+glecrSNJw3Z/lqInQkRl6N
CZ3hTJK5tL3I8hPPg1V4C5Kr33NBv4mvwwML6HUnXJQFHlcRal1ivSrRqIDnCS8P
i3zyOxQT+D9w1GVAqyLRm3S7FF8xTaN+LXGfl8moJswCmIIxxGyrw+vqqPEngRJU
qfrRlM6l6P1c5TPVrpGAoP0soNb26H97tkEdD7Ni0Yt2/Ti8Dt1ZYHmKlReq+Ngz
xxjRSHBMNBFEA7Vygbuj+1llkCksiU0RQZX3PblgRt176UfO8aPeXEQFmB/WcSQi
3NrOJ7yW293O7WGVV1l1Xlk1pLhrbazIkzeLEs9FbKo=
`protect END_PROTECTED
