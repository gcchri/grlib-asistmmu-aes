`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0DyUP7XzU8PZ8/afbEhAy1uooRJrParHX2I81d7ck0FwIgA+cDS6q1D4mxSBprVq
z/CkcQ7cUlKA0Hdia1K7JVzkk8MTDFpCDjdhJ0VRfDauMOH6uqIzQWvqBvndFT0C
kI0hTvdVFYZNJ65bZ4IBK/8PrYbPLGaZFN2Gy4owJlucL7RDbTbzZXF6CC67qM9w
08gysvKFTztt+Y7CqTHqz+E+WREZzE36394kjTlONr9xBft+kQR4+Ra3jf3FWOBc
LU0okv5kEtjWM7UtEjoeu4+u4FS76EycTn+2uXovs59heq+JSy/apIgM4zYTVUf+
v4U/jiMKwQW/dNbXWD0IxpdrFELA1g6fouS/o2Il+FiIVcuLttVbGBIZDEbCjNUS
nHnJ+qnrV3niMWeEyOV8hFuw4aXqOfJEqF8SqPGY9jKrtQi9IXoGUWU/B3/XGDYX
4BNFUC7h39CWwoXeSd4dp4Ja0ER1NjaFe9aegtd1oVxJjBw6JnTZ76QyvZ3pWncc
eMjODYl0EuYiU3QWY4q1ZunN9Ix1Rwn93wgVb1YIgaY=
`protect END_PROTECTED
