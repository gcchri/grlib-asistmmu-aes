`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
csaYtTViJRZJSgfxQ37ek1AO32IS3ISgeYw4Z1OTBDTBR+GKlHRmR9A4rULy0Avs
4HDUWK638+jJoRVGSppMiCfZX1CJ2HzmvhP2Fpi/0KIwqBK+AFjH3bd9iR+XDkIQ
YqIHV9oJcICKobAgTw4y/sS19qlukRiJ+u3pWfbkVZZFP2GSCOAHRQuJ2erN50n8
4HLAIHP+9Gi8t7sId4LVjGO3ofdG0KUYBF7T3DeizSrMDMCzSVuwxbsaIboqWkEx
nSHoXcI0ovZmv88hfhh5DhkAqBLxvqKoveyhAJxSTK6d+nZVUQasRfmU7VdUNGJr
rkI0r3BaPiUF/Oq+G72apm4dLcyPBrEVtGjQpGMvHbp+dY37LDNgxOqb46xP5MB+
s99VV9CIwWq/JtGnSJ7FbLHXnHpAQPIqtUjplUMBX6TFAA6ZA29/c2qLs2n366pY
eoq6XB9cdaYaSvwiH6dpthDoch+d8WIeV/H74HFX+6dFMnuiHfV5Be6CvrQJWmFl
+YFlBj5Kmc/CYwwkG529AEl51SQBJiO4BHj8oZ2c5xD3YWw9cDa30rTj8sqDn2SN
`protect END_PROTECTED
