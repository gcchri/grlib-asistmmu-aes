`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oKwZdcWY756IQmnEAXzA1zLkkiKoYe2NkKbPYdtNe6DZ2nymDH9LBrTVgtr+xcu1
Db5Fka2hB6nilvF+I6pebAbG3+93pyUtKOw2DTlibjqh2ESNWGNC/UnTO+s1YFQt
LtIGsqTNRmQkfqQmyrUzoDsuABTCXZ2HM2iyBnU1Cu/pwmpEKC7YNgxyxJku41se
T08iaHzXAIg+/7tr/YwSc81HaM3pqg5loU7YYX0a30c0dyAYqwTa9++ONWUqRfoJ
zq4W85Hk+lUvsIeiP0SMynvrfTsi0+TyJbhtLnL6CE0p+F9A+AoVEbkUAgaG1AEF
BZkUoeiYcpiC+hGZ2zPjoetP33n+XiJurNuOYuG0JtBIx/7vZJQZlPt7LMzPiy69
gz8KRtnHMg04e4836qtCjJRywuU2pSy+0h5NpSVf72PLf1KmN6OK/7o/3+1JTUmP
qvCw4Z/8G8C6QdpulubnUmuyhG69f4RFJ27+dYnkHN4QXC+Uuiv0YanOEl0HGQQd
`protect END_PROTECTED
