`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ibKasqoyGtsP32QtEBKx4tQsyZyNYdpBHUaUSiI39/FRab/qM1eVfKTytpA8ONKy
1Sevrm8I057MECAcjSUdfXG7I53pJMS5ifKohXjliD5xmNpnS1yYXJgkuVj0wxK9
ZT04etHUwNAZefUq9yHDZNO73VIFvLi3d3RWVoBWDipToLkWRlIT6t9txSiZJ4Lz
LawFLoMKRczwbCOWql/F1SeHv9vQ3jjJQTBjtgrv6GqoFRc8OK9avWXgE8W1NbeC
k4DtIF4rFpbpboSRZApD37OhmLCzZ9+kREArnmbBSWS0eBDrE4Uipxal4mmJVDr4
jZh9Ec9J2DA0/HzwVgaEW93PlOqBD8Qom6k6e7yFNFQ83E1D1KwdcCm3tBs5hHIL
fCxHxD3FcxJ6gvNT8RQltdDSfDFx4awIvV0ELwwDhx3jaFwuW/uzB28W8U8gxpeA
VDvmHHOhrcnlD4OlegJLHScn7ud3JHCC/GpkKpaVW4O4Sb03XiGMjyD0/sfYm3GQ
ElDWZentseUQiW5BtpNyWe3qIBP5uFUpfDCGz0MDADjISrhQTRa9mCCWZrTp5XHb
C7gJkI12HLkZ8IISiZt3i74xSzshAxXR/pozeLsmiqlG8wzSrJP+8EKY+KaNSNPi
oy1aGspLPkNLYP1rGnnlEu2aNV6rPxnzPLz7sRF2tuUixJ+1cqVcGB5BGXKc9iTP
CQzuI9cKAdLfpg10Ju6PzsdWzJDON6JfAGHpD+m2WQ6jMse7O5s7Ldxl+CwDol4S
fKS/4Q7f8hOK+AWH8ky54hIwh5gZuRp2B5MTdRYcBw11xGHZ/lDqe5qpw8px95po
Dd2qHnmKu8kcC/y8DRwoCOeX400c5Vdu+nbx8Zlwc/m2vUHSDC3l+QksjbOrz4de
KGohI7x+GUFM/bUUJGnqcauJlWZtyxk3k58rDBryYlPEw/F4XW0GGaTeqb31y6a8
WFF/a11u6xQ+vjnISsoKYwCMhJ5TelL6o/DzMcIBJHdXXWUVyrS2UtpBRfDIrdvl
hk5wOate0dMukTkAgFkiVYeaeCbYuYsj+YMA+ns9fYMlG8AnIOJFtk8WjNFnvECe
RVWuaCoBWLoBU89epKoekglHwABxo/W6ma8QwjBBKB9hH0W5kOvDMWKK7fLXMpQv
5/acbsiCULS/4nnATyJ5c2DSfyS9s9hdBuwotkgtNfjOpON6O0ygJFiDudb1/N/9
LobB0Vzo8b+Ebit81hXrRCNTOoUJXtFiz7kVNN57ephoJ7rRc9vIlDy5i6yCEYCt
XyxGEfr57rY99pmFhmaHdVA5LbdKxrK+TjAJJJ3C02muUbhDHK+4wuX9nqgGqJae
eAp+A70Tnhii/NxLszMtI5vvbsDElwtCHD65wNuna0y+epImpno0bZBs6aw+9owr
wGfAoZqxfSFO6zumZhCNUFobo9krcarPoaOMk4Hc1TZcXlmSQIDGccItH2gDY9WP
urfgH75VMDIgDggELXzDV5894r61e+qSOtRMq6zFY3GjJVvraGv+5QesFyYmzA2D
v+wPt77or0fJQGSoCCJHBXo6GeWFRbyXPIhnXSZd1inSmIR6bZdjeL4frXnADlYY
VxmVn/XgkZE5NEnMGE2RCFINJxUfI/abZNSmZqw1iYFgegxtlPI7KZGFtvmFWiyW
sM2pxs4Kr5M/ZnVdgcl6AJBHoaWQUk9JfgSSCW/3Wq6ngbJ//l5UhSeTp9Ysh0/v
vRjLl84L2yHme0C4iocYWH4rrG3iQT4JP1JVlM7MH/3jcB3rsjX5d4/MP7nPANI0
xSlfzT2WkLDZEC41WXwDQGNX1Llj7VI3GnUoVO5hMPMksh0Vtp/aP7COCLYK6YIt
L+9pBbzYkSpIiEz/gXBcSZ3Tjjh8zuX7IGEaEL3lp5sc+aTA9+RxswzSHbOL4FXa
ewloTBpk7sGQHd1h+X+w0EjPv24dzJ4HcB9sJsO0vEp/6kIaZkKeLIY4NWWqKv3/
LqAhMAltoQXdou7KeOzPFDnI6wajAwxSlwlvOkfEvClDkY8Thpmlmr5FuylGj1pQ
6THnrrFDWpKVTZZSj544nIaJxodJiRAz8F79F2znUKUMSpnSL9Ns4/jpexK7wlkZ
lvrNIedmxS9V792YjSJFjz0QMWLRn1gBccMiCJI4ERROrRXQuJ+5ItUvwOmR/6Ql
9kN6YwIRJA7oqh+mtpOgbf9+juhQ7mHUxH4rJVVfarqRhHkdJPLMAlDhtSlTOVQN
VeErNjEu92gRabW9u0fd5Mh2zVdvErvWktgE1NWK2oL7waSkUEzQayQ3rgKmi9SB
hUpvbQgxmok1jKLyG3xSw15fd6xXXZdcBowjxiZCyoBAKFt/+mP3HS9/qmpxXW4r
ObCJm62/qnalqx+LjN+rFMNH22SU6YjcW6VDFv3jw//jmuUQUKTWfmcZhuQSYpTc
j2vR3FssCVgi2t+74PWZzKmxwcGtpGvwX28UwBSAnJorYAjqFBuxmhft6TmuNe44
Fwns0YLc1l7r2LyFCSyyBzItpWVzOagme3cZKtPeFiCh9h/70qbzUUltnsFNQ3UN
SXQVwFyweEfWZmHTQ3GKNtJSIdXt4wflAcdgjVj2BG6yBv0fS/blIy5QsS8xbjDE
Z3/V8BDahSyiIOyUr7urTDMBXZDoeLyWn4LaaLXiYPC/YcTKCgXC+GYrJNnA1JLU
SnEX4MMfjNToguvtd0wEP1SaUSurHVZhBULXufuxv0l4Va6pFpz+q3SrymJ36XeS
TXZuNDBP7pU3/PGBsGOlYMsrBoD8l268/s1wzkDBBMY+AFxNG3fEBqdj6S05jjIM
s4o8CJvZBuoiqpEg2QJiIWP9AItTno+rAj9DXSTuXdmC8+RBvDe4Pw+9bCcm4+nB
a96j2mGB5rNNhItlyaNZ0lfXUrC4wF7CVKVpPQMEVpSrt5R4OycVDat4MHccEsye
PxAakuuNRwi6/ygTiQDEZVg0g4LNd+9uxj5rGHJiTVFtRjgS95dkAuFdRESGg0sb
o4trV6Y4ho4niccbSe4cU0e4Xh/QrxtlpOmjco855n3FAXn23zOcI92+6mzRLcLP
+BhbP8zqsROaoXGtj03ebCaXJJtzSuwgrTAz/H5rcjFrC8vl5OQBT8myQ4nGtMdw
x4WoMmuJgnFI1CK46TAyI7XCX99nMcU28D0fcyEwTzMYfToCOL1qroDyIaM84gjp
bY5wHuVl1maz3XD7n9759dxJ/1lDwEWdb+MVEBvGMfnhEvsxB49JyGVm7cIrj/gg
Cv9jVUifOPlFuZnlyEa20iGn14Me5UXMk1cMkjMEkmmiNXiLm1Py1KkTlo+ECI2O
MGf2datDI6OfSMy8uomGNsgXzn+SuOSCxKpf6oZltEyEztgeI158DhQXVLKjDuAt
mZHQpzp2R4HDJjOtDnnvSBHNSGRfvDCDaPRgShWNU4vctpk2C37uWFGnKfJL/1lb
zk2GzHwnHF6Nens8hI7YxOkkRPu/TugTwxonUDihEgPXSXMnJqUnsMxPduRRhpoW
WTDaJOi3CgS/AT4u4FfuRTadk4SXfnJIq7Ul+yBABS+G6qbvKx4jnbENyYTGFcoU
di2aEvpD5EAJo4WWjIl2wdT5TyD4++22fjghoxQks9xsya7gSFzV5M1cQfUSKitN
guJmx77kqbsB+EOZXkAK62U7NpW2LHnJ8WK/ipuGJxe/ot+TzcrvI7ld3xU7yVV9
XKTcus7LBbI/x5kiNVeNEeWFc6C4/mvoyz296hCu/fC2SiPzOkWYnMmuRkqn0ujv
xgdflJ2drlhOCXWGggHsI9jx1tVQqakTMv+gxKnveUe74J4S4n7seHS2hYOd2Nls
q9uJ1fExS+hXazI9/rz2rtGDkjW02MhhT980B/2FQwvQN5VdXoky+uhb2FYzzTsK
lrp4wesbMicgPyII3uHHbwUklkFQlh7S/Y55Qgc9DylE9k0cy8vRUXS4ACb8k5BD
g7K5NRseLohBc22qlsqXtb98IHKow48YUzP/wbcVblKWT/CnQrl6d4xQsrs9ghWP
ugFQWq6p3lk+cZdY0a9Qj815dMN6OGz4rxUyOhl7KTGiYr2SbVirFpc9P2HuzXEp
AED1dTDRSxibs8A+nxdWRU6kFyjdbOey7qZ4N/VIiaQhawHG01X6RdrkypecnaLN
mVH/PgUan3Ry8qvEJgqLOEXiWABYqTsRBcFl+t5eMvWyL7QdV1srzZGNkXuvnQCc
QBreckfqNMTiMhSAFiyyzglDaHsIv8l4EDUYdZsVwCT+KbGeBTtTNbSlmtOixMc3
YFH8vkEFtVaqtFbAugUK7ht7fQHhBNQR72W3GbLnrjFu2ky7/69dMFfItwUvGdVY
F3FLsjQrFl0UVstBsVFW+qqHlesgubX3nZ/DzKXhOww5Mu5SC0grOeNVJj/hSSzQ
eolpoqoqxSO83pCliLCU0FN1vSCl1eWdGtjCf1cxLNz5XBNeF9lnG8fBYqGSkqoj
fSMJ062Ui3Em7HYmZbLmQNCbaSnJt1kiIuyfar6gD62glgCfxls9PM+S1qeNFZcD
yPUYeMBfZ0VFTsIvfdfZnAos+c93e/+cNL29rLdNRS1nDMxoJHrP31C1Ys4ytusU
Jpp9rf7dq8T4BtTke+88foArAIhBpXTOn1jIikWfxE+W9U7fKy5FI0fhOiu5VRzv
FzgGkmT3boEwsZo2s1P3IUN8g5kk0SUAunoAYP9Wv8YERbKRwp1vXbbJKPf+kacN
IunmVCTpb7cR+KrIA//zoL4npbm1uA9iMgAIcc5H8CGwlyoLsbbX30igsbpjwR2J
4tLITfRdHY3bdBcILtgiPqd5EJf9VGxisS2vNnuPgP46A7bp8H3D/plpNz5baRbc
Od5NEA2l9oDctB2jyrjSKu0cRuI155UKqixVXNGz9iCy1yD1FIPL0vCoXbyIaC+8
BlhnLaB4qqfgx88gPysVGqnFmaXrbtVFg6A/YwYuLOgw81zAH9DJsQmMZa5w/e3n
2WFgvwxJnqWLzOlitFVH+K2Gul9vPQJTDDN0jn95ysFAlnhZLrhfUAesFcRSAwvn
LeGGAhkTniA/PBGRmCnMPY2uuxruGjr6zTrktbDzPRTUwoM3HeTLb9xdOazPkyMq
lx1bGwc0xMAv67LEYyAwocbs24dKrLl8l5gJ2AxPm1TlYtqQkObuWwLBh1do9Jkf
xI3lnUdQI8puea3n7az09hd5MfHASg37Hq688BjclMN0kuVlTacZSBgvrOyls3NB
SIgoraNsW2LKFNvQ8SiJq+pikpQjlavc3Qoy5zVrrG+jW6+z9h8X/TL5jQOY3LhS
VC5J/E6AMAS2kAHsze/0U6y5Oem9ZSBgCZ18aSf28xINYr+944Ut/McW7zDSLF0y
RIanMeyZaX+AtSn0vXemI8bpI6/O4a+3mcCPsvwdqdINYay8q8v7uORvkfpmPxLg
uSjinRt/SqCuBqjwSk+xU5R2DjV8uanB2B47ctVe/uH4umwAmZ8wPwwHpm8vHAfA
C5OOB3P2qQSrZgKdvBwk35hFfrT8sGMWNEaJ4jzJVmZ/msq0XtPWN+KsijTz28dg
GPWzgvW//zc0u3xMq1iGAXroa+sAqSSryK8/LX5Br7OTp+Jky8mIm4jSOu1XGI6h
xRESwpMX9yeAbFBsBGlXcKLnlhrJ5tYtphfdJ+iKfQTGUTooPA45u7urp1fvFjS1
nJzklhwhiT8pdd7+nbEfQ8xm1bfNKfrH7tmFtenHgoPrfp9bpZ8zgKkMCuWqDSCV
Dc1oSb37h2wZHOaNUETdQLy6Q3aLyebgL1+8K6ZWL0RqJXIjEFXExZ4woAHNK5At
WcASgeG9aYq7heZdh9aupL0OXIahOBxQiOGfW4wGu4xxz+94HHtQZYKvZ5pyIDfd
QarA6u+c+t5cJpywMzWowYGG7r5XqkTMZsCZWAmyOYKgLs65eT0sVLvYDAcWccMi
kPGym2eGRyU3UsuwyAI38MEUt2R4+oVUu9zsb0SVWhwvBP2DK0a+zFeWnt6g7ZTn
+Bi/OHbaMDiHeTASwOEutbDVYgWKdpiD6OAJvBwDFuS0lO5V/0xMsKHZzN3ppQE0
nlADqbOVnAdKZ8cE9fceifdiY8LLqLXISpJEo7u6Z2dPs2nPwGzcgvD/kSREMSpB
4dC81EmqUMQNjp04XTLiy7qqDH2HqiDtfWxuG1rXp51bxzAEjtIRGPXrdv1iAO2+
BVTlZErKhkbqyA3C0lMNJATIyHhinqdwc7rGoIGeMYjhjb7Q+6hJZfc5gQXmG9kk
1Q3Gvjm3ErC1u/WSuZjUt5yVG7dyLE3bqUmMHac1Lo6Bp0IPXQl2x3K1yz/fGBqh
2G9kCwR8EH+nfIu4+4wJbg/5Oq5TJb7PhZtJ6WOCoWlxBr2cSzZClU9mgWyGZ3sX
g7tQOt49VaK02DJygpj8PPGZAvdfUpPPK0IHta9AFNTZR1pZpdfAH6/1yh1ahKkw
yiY+iQ4ZiK1ZHe2Qase0/WIB/kPPUDBx5qVDHcO2vxtI2M+MNCMqrFJohyrvTg5j
VuY3lSj8W1glfCbeQex1rAklRX3fHi5QUZ79iNyg263S6MtpohmFyFJGKYEgGvL/
VPpyFC4h5Ppz03vI4lQSWa7+feldhfm0KpyftocrzFt6tkfVmtv+Y/fag1A82ySj
l0Mrkoi/A91qI2MZ/OBrdPjUa7ompstQchOeXWHfW+VPMXNoNfdCJWc9cihlk+Q7
EVdGa24OghGCwdOscSJWgg03d6Vex+mft6ghugBPC/mWnSjaAIoevF7BOfMrKbx0
I1Q2xgpgjAIp0//x85pYy7N+T6FAGiVlTI0tkgW3+RWdrY7AgwWlBPFVkDap/udQ
BxWL9Z6YBYkMM3Ay/v9HrFWSCQOB2zDn/Bu6Kn4pM21TgostfLYY6R9MhCwC7Y0J
KCbFtbU03ohM7RhF5hK1nCtgqwMl84kqJXnMz82aTZtp6lrNggC0FevsqCZNI8ay
TMM16wfO6k9ajJDnRyijlNqPN5bieYub4gKdw9+8q3AZvYqzwp06Ghok9mcBQDmr
oW6OndPlxUZvPxJxF5YQf5ZROIlRyNp1bftb3XM5oMiEmDTJAZ344Rd/cLXhe6Uc
ycctBK3XmBcZQl/7elbH3STL/aabrE5G/K/6GODhQKjjhUp95kwsxs/qOrMl6GPB
`protect END_PROTECTED
