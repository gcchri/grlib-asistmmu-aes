`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zHNPuS6S1/0H+JSnv+iKk83+sC/X8ta3hZbafoRN+YfML1Fvu5rsEoW27B6xFxkB
7A+9gOIPhq5XAwknSyqlR/ZB3n+G5DZXEBTGkTx5dYz/MweiHa/2FUY5NSCxg4PZ
C3D4RLkLyi3fGE36HKVKNUmMMaCn+UjUs4RsVb0AIzl3SnMnYQDSCZoMx9IyW9PA
GFhit7OOj9OScj8W5B2Mr+KuqDUbaLWRu/7uJhTJ0YBKJitwnL2eQXWffKBMjNaE
Othdnji0d3ZM2SL0Rfnh+/QLtvll5tMBTlzfpqPz+6xH0c+C4JMT4xHNlyLfzy6v
iud1vJVakRNh89l776k5MVQ96i/VnWkYtALA3FBzAD+85mCtC5idIHiLCRotBJEF
/KIf3Ydp1mhZIwPvMVdzjPTM07efpV8EhphYHE/KdTLMmrE/lZNM1mVauzUNN0TQ
PjgzSaJUDngUZPXLtMBxdUCnNUTVRdU/BMe0lYOejurJizqtONMCV5gnAusmsnkG
YR9a3Ud8+wVDslrfBU0/oJatc+tW/ufmfr8+y2eeuY918uB9f6Ik0wMfX7bsV1Xd
jr3WRx7T5TfQLekVxzqmgvQTA32cLb4EinGfIgt05X4AeGnfa+DCpaGQL9cuVdpI
kZyONz3lie8pYTINrkpSjRvMlFv/ccAHbpYEp8eMo234ihx6OvcS7XqGygW3NgCr
LGk+RwhLGCOXbor5rU7e9vQJGL0BwNQgVHu9r4HjX1Jv1GUa2WMLrIMAGEtpJCTV
zkiKnFz5OrA+gQL0+aNtzrq7eSGJupfTofeCzkz/60EGtIVVQM42p0ImiJ2Ui7BZ
LChaLgk1vrzF8wnJhblxHSxu54AsjGfU4axxJA4ccMbWOg7C/WWitZnoSV3/G27A
96VvjZ1IVd8GjH00lFoqX0XkwqzVRU8AzY1u5sLirSZHllvf7ytYWe8JF2Nxb3uP
dJaaYwMjIaUAxPn7vXqj5Xidjalv2c3YuSz6XhzKxmH6XembbVi5GtMJaSpfze3R
RW3Ve1vnumvFh7Bzn/4+hVge9AghOpPsI/79cWEmq2PotNbZtQrxMr3JfuxqnoYc
xG9im09l4v5yS5rblTFfIGMa+FmHwRNCEDmWlOD7IGlZUhQIXTeNRYkQhKtLovPJ
JJldJrsH8R9s77IkGIAzSuihxH6Jdm7ggFYhXfCjHmSODpSDCPg3XH1YIfo8HY7q
abS4D1SraRfqtvBCslukmMR3wuMTvI0MAkuRBLvEcJWtU8i5RrlvEBU9Pe29HKm5
ZFQ56wcmWSQc1l/B7O7QLf0ep1XrslXNvJfbMqjfnTPrrOvlMItzmGgTm2JtTWcP
L9i0RjpGXPTV1prmO+6dczBHXqQKl0kk8Cy087y6N232CGy/QfUASp8wIr3nVmyf
hyeweV04NVyIz4Wnx3S4g5tZFqfJx4YOxV9/jch5R5M5LNPTr28ZsPDTFkZHjjUJ
u6zFDq3+7hD7eZ0ryPuWiD3rBn+752KAZVSBV0w7uH4Kg8gbBnUtApUxaYEbVnXa
`protect END_PROTECTED
