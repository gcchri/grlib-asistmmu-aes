`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T93kaefn+paqk36K/0TtbmYSJwULZYcnpN7l5RWI/Egq5l4W806kHUxB20iZLxTJ
Z89o9ifZYk+Ugc4MxgZMq4J0+ELcP5spZHAKx7mgHh4BIuQO2p1GssblUF9cuIKw
hlZ8wSYXHk6fzz1qta++52dRDsVIhuVOtQanqxAuzsebDgFxraGsaVs/ir4e9l9T
UV2hUJvL1rZStcI150syELvepyO2q1YOwPnxgIAoQJoCD2EK/AcetNdMPJw5i8cE
5l4/8ZsCIvOpaJA5iMTF3jtAsTbQeeK/NC2tKQ+6J/jbkyLbHg2cGWCXZPNJ+JbR
tCqO2I7c0epUW27vIpj6U5PPfcaIba9gxhFXlzquppekBFcBcb6oOMfajMxNxZXy
rRNVFYodxyCPZQ/lkJydIgqAQSf6mv3mFWBDlxoig2OBXzKeglD//Qt8Kr9Szmcz
WbdxREaVE5iGT34VgKQDte8+68sypC7Yo1yqDAAGfCwlpryNjrh9Dx9o0ruCgd/B
ccwefB3Esqgi6E+IoPkhdrDNLd71IeG6h7rYmKoDwTn7uoQhFu6I8So1vp70bnA7
eUsWTb7WaIQK+jf15Otuo833gjytNQL9B+0APGDP0BZEssYy8+L5E92gHNSC1jNl
eMkbUPf2n7mcgrkroeZe/PRMYb84CgeoC28gyO87HQ6BaKDp4LLcdTmvr85W40Z2
V/sbrROYKW8V7NcCd8KCTjLJjWiYVtEgIOz0WANZTf0K2zq+TF1T3QK9Kf+yMEJA
lns0IKgwEN4hiNGnyh0ovBgo/iVohieYsnAGOZC5ACS/dm2HSBwDCWnrDB6h48X4
eH9u4PQnKgibzrAmqS2fZm1VdrTUSyn12rRi9fLTuIYQpwVKNhgv5+ypI3/LXqRx
PfyIwfqFRFX15PvJ3QnhFFXqyuofV6yK1OOcZO9dvO2n+v9AhMuyuoBx129GyJfC
4ZycW+QXMh+GEZYc3JVshavVkAj0N686hYkN52BnesxmJ+aENPfL7ZC632ltUaMV
X4EPWwnZdezrIx7FItCrf46vkfVwqT9V0wDKfYfo72uYpdGft1gZ/lVnA+NKGdjR
punCVyXOhRzm/btCyQJdjbwvYneI8fjJMFHrRmZp+WtwAJYyh+EJccmS7yZrLdJ8
XGpTOL6TnwWxkTDmiPu8c4Zy6vXuqZ8b7t7AGPWitn7uLQvbDnU93lY+llwIcZl5
633Vm9j5wHLowJIlUCOCRehCf3q08p9AE8ktOL3jfEqbyWTj1eRWqUxnjKamQ8xS
38T2A/EBeJKV9b45gDLuH+5zkW6ikIn6XdoMby6Uz0OnGG+0qamiM+Zw3QfcXM3Q
2tG2buNNVuh2kpUJR6k8jBqo/2pIWNq6jlxsvrUGUywo7cjjHbPQKhoPMCHcW+Pm
lEDJa48EsAfLtbTTazPcbQ9xEEC6BxT8L/JARhZaKyGp+Wg6E8aPjmFNU/ntJIrz
U19hUC2K2XWludSEJDKWITufWAMmiuW9q73Pbaw5Knkyc4WXLtHRTDjYiC7RYdFS
Vd9Hp5sk5aPPCMB/Fyd4gxe4m65+an1yIK50+csYwUf6HoLAktaNin4Qt4a88ALn
USH011ou6zCqCz9HD+rfdACHZ5FW84cav3vYsYGYUd4hE1xvp4lTZB5/FWK5IO4W
UN2EzyDQ71c/cMed2ZGBKMrEfiNB9h/skL+NITXloN4TKiAoTuKOLsz+gdB0j8aJ
TOmHyPb0tD7z7cOfVi/ps9rCwWuSoJVsffAi3ooco8j/a42XviAURfOGyphBqF2c
vLoULpLDvKND0iG0x74IfxW3oCbpSb4dwhb+ubcnxiIpQQJ3kd5hDEJK2foDbZ2Z
BoBW/sxROehY9fPV7J3bSPPkHVsJ5XBxltxKSyTql6X6bIYslP+zdNfStq153jLb
2At3OXv3LoN8Qi9CP6EfA7x6KdIwrxQbPkP8LL6AojrAwjlCfeTXFruWFouifJSc
6sG6HZ3m6U0m1dV/KP3/BI8tdv6rjd1BGC2mhCzprRoCIWqwBu6PzaG3pO9K5q6M
L7Qjl7SttXdWUSmnKjoCVDpEQFlWfCK2XDEc43UnlCQEAYBDXmDsjFxHgx0YjQOT
6bm9CEECubelS1Zu0ISwd6iPFwjC1QGJ1dgybYOWeRXdgDRqtgSGaa1dcpaWqyHF
2oR+mGjPb5ElmmJJgfU+1+mH0A41BdLXx5lc1ONI1/hDGcHXMHOIPzr0YVSpoe9j
TCxUAisud6KHndjEtIwVJMIJ0dCag0tMFjaQ4WSLZwpZiYJt+RDMWGcgIuxG1c7N
3Jo5USTi1oI4yrE0gzqRumuroXch9Sqj70aGAr7ht6nt94ECfbKMMZ+3Xo6wBReE
oXTs6QhWiT7XTXOBjg5k2MQNoyVN3LJsVJVZ5wSKQ6kCcDoNJ5dHk7FL3ELH5vw9
Haf6deLSanX3pMf4WFeOjRLbYx6mA2qhGpNiVA9QmTeZvCCCVTb4jZjtScrDmGVf
szfLiqUOVn7yuhDuhV/7pfGxMqf7xRnQDz7L1TWER/dN/4qGk6fYd8P2u0A+BDuY
Ve5h6zPJ5AULMXrScOUl7hCJwccHcXckbkiEk8Xq3pRX3lw674T/5qq2nzasZoxH
XR3PuhSEeJuUPC0PDY9e3XBB6T/pw8mHbuF0CdFRjXktVrOBqmgCgfEqO6nH2oxN
YFWbdQTvRkcfL6TgDh9uWQ1/b+iFJrfzOa/3iUVzB3Dsk3X3H6xXNQu1qxrJaIct
K+Zf4jcpdalowwuA0lFkOIk/ntft4b1BV34osES4LBFXQbaVAZ9amejpDtlxtwqY
GehIJ6xYqoYwB660c4mrml9uJpgmH+LuqfhZt/bDuXBMC4hZPj88aa+Fg0Sn2dO4
WdMiB3IzbUfLZhNzsDQThuMqVIGW604XMXKROBBS12vQiVgyuoiPBC4WCoKE24Yo
CWDeyaZEkACL0pT+91bThvzDQIXrFDwBMbZ7JthmEGfz0AOQAzZ6CLBK3iiME4Mp
JMPDlSL5XPZ4QnLP9Su5gOFI/bsiNN1tH2ghPx9VosF5lmVXyL+iRGCUqIgrJVOM
DS7v6JvMvtYVDe8WaUAzbNi8uUe2nPwD7B+gIbj46zZwMzSlvrnjXhbGI7Of47ZE
LtySgiOftR3B+Gw42iVi8mEkhPl4fXrdq0SukhcPwfu5Obzn9oLtT+0s7uW2LenI
IfJPqORTBo081U1AAFdJrdbCCnJMbR7A5BuyQ/5CVIztKjUEqJPjdgFK6sycigLH
94UdsleyZQtgeesiRqRUVTz5YznVEfQN8UeaS09pUrnzW/Ob34O1LifyPB5FHx/i
ymWAyH+AeaewQI2BIzmP9DGkWiB7aVOz51z1+lILjzyW3O48PfuEZgZYc3F27WOC
ajId8F9Ex4PBdtHRUh1G4JNwgAAOI8bdgRGXWQjOhV8WsdRjSM9FMPgg2sGeuCeK
Y02XNB/UHdomL2C51YJQctviYqK7OaGbJqV/aKqG7wKbvgr20ONc/PDrEfP23GpL
wAX38sqR8qRqcG4fmDMHBI2x2GuRFCMYaQeVkAHyXl/48trUeFXv3XYgEAGGtwQo
wPLtEU/UysBmgesKjsKIEJIqpAqUBQ88ih1dm91H3nqYLmLrbEFBUm+EikTiYhLs
bTO6kK5nipFlFD79p4NJY2fbgsN7sEdHU4oz3oDfw8J82WGmhgXGAENWXbbvJlhl
qZVllXs+lGxStTLEYqE8of0zaeG+dLYFVottsLHIjHQGlj9tr/1HUhZfonkKMtiA
d1xgDQm5vy2pp9TGIxQ2XlENh1Opu39wxtdx76gYEzKJ9MDsh4DqcvDI93JiOtEA
Itrli+Kubl00TK6XDkauURQBk0DPPV2dWMh7ThgyZTX39kbMuRjPlFV5IN7nsC0t
LNY2Kfd9qwcBQFJeaQoJndx9hbyfJo05M5Yphfwzm8jwZraqQuvyXZzttTj6z/JW
VUeVvoYT4hLPoYcMfzsU13In8ZMAaPzhHEBJMDJZoqZkc+sP7Es1Kl8oJac8Y5r+
vglZRKYvVgcRi/5I+93H5DIlCazJapzdx8iVxytwvjE5TkwUL3v2SdcHtCgtNnBG
HoBPYeetSVLXZXbD9wwg9ZydiFtZJp4JoaBHGjzSA9i3/n4VmFGc3MequVbWtjWj
1XHGqN0lF2XWA95+jlF5oE7opqZMF6VgwqIJK59tJY0bhQ6elpBS5/PQIjLPyJzG
Gy8x7lPZFvA+ncojusI8qIPlMj8g5MjONKtQ+Ery4+VB5Redmpm9k1u/MRMC/mY0
EGB1J5dYaXbo3dWWgkjhEGxazJNbDcohkHgTJ5zUan08RhLTBtvWrtjYAMb/Xy3a
lpyTsapaQeXhh3oeWj299azUOpQkcmpImMIySwpSdJe3DHuSOu9Q3HsFH0e+NPfe
whvIive5bHL7Vdiyx4Xft1/fjix+qG4mwgttW/DzHVtd8G9RoTzvRYqnQLcc3MKl
VO6URjcm7rkriQ8QhJF30wfOISBRaufGB1VXz6h8l8y5DnqqPnz3XWHllarzbrLs
fOAi+hzk3EIQN/up7gq7cEVNa38OixGkia1LsN1ATmWZ/zxlzRHVhCqFgyekzB0v
Qd8ETDmZItD3BmG1TACa3nvBlB5Vnp7+WgNKAcEzQcQF3/mY/xYREkYvuQLtVW3c
Q7OvTtkFDfgnxaySLT7ZgeDanHSa1VgjwllxUIvy4jCrO106pVXTDp9dYJNHRbpL
89FlRm0h5W7/VoxVTXb+PzyeDRWWl2JJR2kigY0jOnuuuXqnwkAS0qZi6qLzORyK
tpD60EafVDcb0HC7uXze+egG4qzaL0cG7yPFODFedTfcZEzgneJNCrzIWDAA8gss
EwR9j/fiVUYd0/ArsJRLRAxI+7A9jxjXUIRbw0Hr8NLQJUBTc7UtPPRr+3V2ptnf
ZYXRjvOgSGanCWHTAwNRI3l29y170uXySvGplDxzGOC+7l7EP6pONg8ewoWFVw0Q
L7MLeLZejmU8NtCmseS1qDj8hpUAQNlc/vrdvej5adeQoQe6cUxcIrCo8GRybIQ4
34NZMfjz+BNPk8y8xkdSA8YETdPF+CgNx6NTAMLHy0EJYT7azqxe8A1+MI6aY30G
NDFUDqReM44/6l2dP2aU6mCH1Gr2RUb/yObbiPIbQynzTCXjIqn9sv0YVRfEkqxN
OmLk3sMMyUEB/Qp/jpI81k9FRCwAMGsagxLnEMOYeQMT4wHlje/2yf94DlCwOgZ6
fa2WfONeNF7SKecbCgJSTg6HvvDmefr3PSqq2J4kvV5jKnKbod1LjIrw2RBSai/v
5FI+Z+YVwRPWrsloktGY7i5wqsAix4Q3+grOVmpc7zDk8YRvDbDuVTeKnku37sVo
PYmB90joMShnCCCAIPQo2dd7CaCIR+tn0+GXcALeGoYdhs8tdjNJmNglgAyGnWnv
AZuDuP3OaHCJLN7/PF7aPIBOqqFEcOWDbp+9LCr+IthLOPpuAZ9k1/Vy9pnLWfZV
r5e4uNTfRRHahE7ZaJGY9CenmPTn9vg7jA4WfiEmijlsKpF0mlj/v61D3aguZCpx
kr4Nmf42o4bW4nkhexfCnzR0Q+vhvVoiMGI/hETFPTSFAYQ//vFIPNysqVMVeRAt
cn/efVdwwCfk/xYg9o3ssixi/6FK8qB9eY0aMYJRe9iv1Kxi5Px2yGVQn6ccAgMa
9LBGwYu69LEvXQCGshhAsrIwOopcjWwYzgtzxPllCuAruTX9coUzpMjkI/uJazeP
jnmieTyAI9UEac2VSF8pKTsa0rtM4MsaE3QG5mVo1RODCX8007BpWLQ5yOHaA+DT
pRBNOaM7uPwTvRnSSupJL1E8K3nw+3U0QBGVM0RwEaxinAmVAYAvtgd46UwWUx7J
mlLumAdYrJpbMtovsR/q7IsH5IwobH9PVh9U5ZOWR8WU5vEjJR3Uhnxm7X1eVW/F
VbpwqZ+Dlz+NIagWPuoxu3dMMLx6h0A7MBbXkMGoS9ETcOFTK0HlusIrJc4eQQb9
nsezPVlbDIYm8bHroXG+IeCVPnzktC9P9HkgeTZTjExBFtmP4I1H2tTbL9ntPJry
cYk94MUhg3yi53MUH8jXBegLEXc/9KDgdzUNaIBWRG3pFKv1bfHrL5pkJDHkdrlN
`protect END_PROTECTED
