`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z9ECojjQk6Dvar/aEkzU1wOPd3D9EQYms3oCu7PuAVTo9QBooXAjZ6RQ0yYmYZSX
lJ2iT9WZLHOpuD1TDtcwRzA6ul5tOuHDpebSnzvm8jP5UvlgEBDfIIMCxzIaI09H
SfsxvEh71CZ1gbAjKaL5o+iT8rLJ7e17DsGJ/S+EaV7TK1idDP2F1YjKYt1HpSqa
9TbFHm9oaKZuk4d6apr/N+6+wU800+U7idEQsHYLjpEVbgcVwcPdxbwZLV/U5pcH
GvihLwIL4BVj2D6WO1IdGZxbw4HcresUpsa5D7iQCbJQrwPrkahK/wCkYMdLTrHU
`protect END_PROTECTED
