`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J2CnU1KMRQYdIOw4Z2vU1b9qL2r5C0pFKYx2E/C0X4WvMhxFTK8xqYzqWwvPJccm
CBmBLJqzTqlT1/rMZSbg5jN0Kc1QwSzjgvk9HhwzNYHtYkqJXf8cXHulI6x3MAr8
80oSwO9bHH0nsRShtmc4EfWNJwzfUvjyxoSuSmbQSrT75yvXFpVPdMCJZ+RMQSNN
71u1/aezl1cuxoSlVperYubpQ3hYnQalQmz4+8l5skjxj5RQxaw1LqvuerBwySag
b7yqqyh3DV8qFffAJuLclNkMJRLyxYFwJ/DYjr+sizTMklXasgOYJg7i+TTzl3li
6BOM9A1vsSIo9VhoNdQ9bYyLSV2CPIYSm0fBsSdg3iKoMQbgN62NJs3/MJOcM9eh
YM4KuNjJ+qDSltxatlv+4eqkVT6o+U7FIALZ7OmdtCwMi0Vtg6QVuSfxi6SLhGoM
bYu5hr+ybb0+hN6XR01vrdrlcla54sDqFQBg8WMOK5Rwnxo044xIensVuHHzV4Vx
syVvObTbamP/SQvoYS+Rtsl/1+Xardvf1Q3h4Qj4la1D9u3VTBuN+JRIIddaVsFM
`protect END_PROTECTED
