`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/GUP/mHu7IjfoQqKxh/jUd4+hcFpeb/J25ijDLDrm/qzDeuOTZ1VpuXMQIM0HJAR
C97zi1EeevVjSqA7SAQmJ0CgEsoZ66Z/MK2NCiX9TRPvSbdNA3lJBWwb6lppDCZ0
arK84CyoWfVTWmv8ZHrLV/tzHztft6qWDjs5lhxJW7QLXktqbyaCjbAgX2/zoVeX
FVRr3BhbUQ+Iqkf0UhUl9O77FGpZBWZd3g/awa6Qz0oAyPwYHfGsrpEDlHhpp6FG
FQ4xlOH037mKSR72ok5pnQk8KUT4aeTTnwm6FMMCXZCXoczGwzF2AoZgn7pcYqma
asLmUxo+9kxK9FOsu9YlgVLCNgoqDSu7Ci+JeURkHfL4DpDBPK4HcIDjaQ1yFmpN
WgFJysr6yJfiZZahsivix7QuOnRK/LjYQg4eQAIKWRs6m4kuaPWEJTT3Qsh7ibeL
5Zrxl2dyzUnmuRt75JLqSH5r6B+HM0VPUWEQ+h/gwle8hGpohEgrWjG4KVHWgNS0
M85fVfGeGPGEEqdnk/z0ToOXgi8saqh2PYtCYNAT/4k0z5OTtIGvtI+PhLHQJugq
Oy8IogPRGW1NvaJ3QgYBxHDNCBBZzwg6WM3V4E7VlElpScqDx+WanKNlmIYm2ujp
zbuDagSDDOBUKeKC3g+VNrEed5VW3tQn752ZjHTAYkMbcLGhsY+GTbti/6/nGH/W
4f9rYAAlIAEZBQCthZKp/f7whbLIVvyKVJZhI0/p8RX1Z5kwcGt+PfAy0LbGKNtX
4JCN+5Yyz+dz3aysIe3pxPyzDSHXg9GHbCx5sjSUJxk4PrNs1Ljxqh6Mm1sGjwD1
g7GPQKtsdp7Pu3UTswyYwhqXNtml5aI1Ksh9w4XIKXPaNdgdnO//9W95ynUsDkqf
g+Qf2s0KzX7hKKfVRDYyszpZsXAnVsvgLRIihV46TtDx/fRqLdsMnWgkf/3d9vFK
5rQn+87I8nW3MBH8FUhaLP/KRw/ZBfQrM6oY51lnGZ/a38zFMlxi7GON8wDDOOmT
vLoSmBeiZ0rKFMjqJQ0PEilfLoSHYHE2QuEuWj96461ljlca+NifeafDYU1IixV8
Ms8unsNcN3azSUiV0LX4yw==
`protect END_PROTECTED
