`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uK3yrbBEfs+Bebe+H6x2AXrL7CSo9CnDtRYr1R34a0svPgoJ6xdJvwC2gMSMdN78
fNZa6s3e77+aT0jntDPIOP6U0cjmHX04AyCL3QHgxyM1lSndn5YcLVbp13Egyz3p
cRZe4nBEBvIBs1oo2iRCyIlcV+noaM7e9mKFERCCrkG3KL6MFcw4INcKjEoa88GO
tK9bePC5YyiKoj6mpri5wTr0fpAW6rvK6xVeI7qr1gpZZCx/3flm/IoxI2Di0Oki
m6YShurdfBdZYq19FQt9VC3+nFaODXu6LnWcL4KXYniOXl0AC3QHn5eZrsx2dL74
9taGmCKapgFhpQx1snzPOdCBGfZQCoFtmNQpDdDBeURRB8ZaAYcYXEObI2ZkuoiO
eHvKtUaHh91/zFuXg0tJ4fqDOTKI5FPZmOnL6lyOZ3sfuCjwAeplbo92kAo/1awg
sQAsj1Kx15YI0EziM85HzMmmxt7g3xNl7XeoL1wzhG+HIcU3ZXkNgvXBdq6L2Y2w
`protect END_PROTECTED
