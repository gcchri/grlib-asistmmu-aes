`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oBI/yvgsi39Tm0qe+oolSp1wmwbVGospt1u05H1CA1+OinmnkBDO81wM4UZDaxkz
pZHS9fzra5o1YmgiFxrcreJWHMeyCR0XwanuMMXEgGZ0LreLaHWQC/fHsZJc6FhM
OJr0iwYbTUgPya6Jrh9kuhA2u4HJxUsZET6RV0mikxl218OEoP8u1tev84T9zZJT
kLw/PVnzkqbRvcUdOdCF7j8X4h/jgMvNntt6739SHox5VuFU4PCL/C9tTMfnZnyN
qezZMGFk7Bl91agnFcmych+1PWNy6kAPzNMHQ/v9Ux+GwshLq3IRF9+lBBbTUbBD
Zj0yf45JNUtZtnqIZt8gCdQssIXLR7MjD+g5O4wLUY01vJcO0lKf4LdIkUBH2hRR
6W0c8PfXAAWLCnHrYEmNkgRP67U1xl+0K/HVlLxbuuGfCTVzYaxlHWpJDBRxe8sA
p0tP6LZSzU/flEdN7/MJvsZX0WaaeexNDrBj6U/k6O8gvNSLmw30/bYh7zHdN9+J
vfVTI2FZVh1ZYgu/7hwaSv+if1ijZQq0oJu16zA9QIOmUGdJoWOuYkWqR9GQaNkh
yJKBh6gTJwWRcS7j8HjQ4/h0XaQU/OrBIX5nCCZFA2urntpRx4diDKxkLBbtbSCv
5bPJ9KXHD+mBvqHzbP0izoRn57yx7JtG6CoXJg+YVqJx2ZA9YWjp/R2Dvrs7Nkzh
svlhhy1jEiuSqVzc0INDJs9BeZiViBqOpNNzRaZcR8xiebTQouhAe+bpC4elKfer
cJJJ+HP2uFj91qdATkCbh396W0WSTNVTP2GJpkxKeUhhmhBScIZrRY96f5ROoC9k
3B2/axe7RUZqdpKYka2eSZOg/vJxdl5kU0e6/mEsJ8EoKMPNA//1bsQIxO1jWKUy
4iuustbvyCC6hfnCHJ9U+SODCa5UJvgONnlH8u83wSjrwbkDr6RUSDiRL/NE6gM+
jd99yMnErCkLdKWlv/A4dqhJ1DpRY2jAhww2RlSQRb6MIB81qfBmR/+pYmv/j95U
lsxXYsdXWcjrV/PulXUTpiiZH21+LjiF/HHs5YaGcr+wCxOOVVzPyWYFglcpVIEy
lATyQgdEvDDIgdIvGg8GIq3U25mLvnj6cgho3ie83R6qlP6IHgeprhnKDNITRwFy
1qvxEdOXVqLcmCHF6mcelyivdXPlxy+Ilv2O2ot4xmCDljrIxoiu6nt0JKwRpvDt
V+inu81To82SVad3U5HgVnRaGASM5lahuVk2VYaxAB5u5S1PO+4pmy2X67vZoOye
lIgFjb9w5uTJfHZ5Zs9adfwGq5gd0y8u7xj7emNYHCulr2Cap+1tGy+qMriNci83
MmZXGw8NnYbEJesbdRba2A==
`protect END_PROTECTED
