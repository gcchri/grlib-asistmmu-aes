`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/DsfV+AijYOGRU9CG549zRs0LnPLrRYSJ+9Jty0LZqfIo3cJwCsm3XI2n8crhXKr
SC+nVk6AH4I5SLWey2CeUWWA90MAmikBZ9bZYzgAeR49QCe8h+J3Zn9AQtYNVJ+g
d6pmrPiWk7HRYUnzGB1V8PFV+lhvVp9HdPipbY0GgNodcPEdoGKhZAlyruc1HCVu
Hd//lZ5NmIAftYnjq7FZTbhPuc7n6FDeC8Xaszp4udCzb3Qjd9F8uEldmoEaz2oA
l1JNwrqyg57rw6MJ0lo3i/F/dhruX4CI11N/QpeZa8v0i7HZ0yi+uy9aMK/pElr7
vwJ4OvLuv+oChJDUM/aoVw==
`protect END_PROTECTED
