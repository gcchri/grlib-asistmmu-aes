`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WVTL2Crg7q7yUAOlsvFcLg6st5w0uFjfBpUuFj5cwLbbZWDZFGp60GTLufGJusH1
8r/h+H0wuvCVu+4sgeusshrfzQvbtL9ecqDgV2g7SCvDpcElRhO3YPI5ITwe5D5t
kvp9y9i72/uqfj2Xth6bYIZvdgDOKVkjfj5cfLSYUAyfEKH2Sw3iCUIP/5vG7mAX
aQId3QTTWh6Xavb9tZSXyuEPcS9qZ3/4/j2iA/p2EDFgRngO14HyS6D7QgmyoXBI
NqM1GKbLdIUJyqPsZfuptg==
`protect END_PROTECTED
