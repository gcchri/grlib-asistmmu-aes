`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aXzqXzjNo+VVDKTEIHtBQLG+hZ3xsKC0ls1SoXbchhF4PoD8i4IdfssRPDnE8aJ4
xWz+UPDCInXE531flrwR3eEWrGcwgebYymMfOXYWRQuiWaxx0bjbaivqbczVHwNi
k7UI75Tu0MUr4P2CVu0p4Qk9pd0tg6QAbKk4ZpkLWih8Fn5/ENsbwHLcEeatxa8a
iuY01gRR5gjPBYL7LWmGAGb+qqxDhrnsqjGCsjaynAVYktn0CAl/h6BpT1BrqP//
QePFu2nMsH64rOTnILx1moixEvBB8+qgsk/AHLcvXtfYNEeeKLE8TBDhYVmb9/n0
FAHbxyjP+B+7jcpq6EHVJzYadeOa2/tOh5g0ZJMKZDbH6/AF5cgLeiX9uQDXylrE
v1DbgTuawKiQVkMePmpUYQ==
`protect END_PROTECTED
