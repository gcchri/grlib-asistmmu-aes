`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tM54ImnQ3GyaJzhFaQvLvLWERr7NiH2gtcxpa4BAsU1E/aJS//T+1McxY5M6vldo
ckTcus/v2xLmF8aDWC/L5DNT3J13M/8KONzQOsnfC8CAfTucl0vzgaREBu6rh2Mb
8TkWowGZjPyTfCIP55xojZxjrVzV5qnoU3Fx0VML9HMhJM/ijQm5v7Bm07QVkb/h
Bk7wqNberH+hOLvWTo7lB7D/eGqnrUysQQEpcKhVoD0kv2E//gEAhq8lNMxA5uO6
AOmnCOI68w7iBAUJp6Z1e91rgSB8cyWFKgeQkD4RtmHn44neO1FFaYsQ1HvRJz/V
1Gfezin0XW1Wq1CL9bfFxZ9wOYW7TN305tXfh1NcVvT5E5rP4uOiz/M1s6qwJdRe
CGdAsRMo0FS594uK3aAU7XzimU8jP6ovLZlOVv+ffRk=
`protect END_PROTECTED
