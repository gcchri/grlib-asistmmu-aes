`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8KdKpeggTaWGA/lOvOXa6pKj+6GpNWQCeSvVpVdFcfyEFDlK8FbuiejgVRj0k9o3
UWCXl21RS2RweCyc/KBT/ZXQKYuSjLrsv1mJJfJUqClNDRZ3HIq78XAw7a60WkS9
VHa+2GdNyPsNHNkjerFPGfwHu+Z+BNNcSN0+pFpT9ZwYlYSWQ50ZLpSA2DrR6r+U
S0F7GiWHG0yN3x2tNe2opZ0XhSiuAIO26hA+If5vVPQbdbg6EMbefE/he/xvAk9S
bNCI4Zq6FKtyoaH+7PdWUmVgD6xRlfun2a434UB9I0kyRzUj7/MQ987FDxUsH+KT
0LTbpGuBd659MWm8GezaqNMGqT4IHTDktH245LyXKyZbRtDiaDSLP5wC0VRVWiAi
xgMwDQIUYPzdHBZG+PMsgQ==
`protect END_PROTECTED
