`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
60QqGMzFbyf11UBFg+CJ4H4Aah9SMCYjUJZPPQ0yd5GuxM8oiE6vNPRd+9kFn4MX
/XtgFzu6qIXdDaC4+SznZAhhBWBn/CAiCt/WysOEQ/HVeKdQ6D08G+fSKs0VBdBe
2WDP3IZO32VOWIqFB+engGhVdLjBOhIJM9uUGbl5qCejjfTg7Xq1fMuyfTYa91gt
Oi4SVEMB5hw6B0KcMjxLcyw2zMJy7HP+9npDLuuBv4/fGDLF3xb9jN4WOfekfRUg
NHT8bsVA3GhD4LBAzmNr9Q==
`protect END_PROTECTED
