`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xU7FSy84YyhJDqVcOcfBxR7/YmGoS752edB7b502jfYJSvRbElf5T0oNwn0nwpqh
iZw1s/PrnQX35P3el/xU7AkOWp+sh5DZyoCyQSfuK+rEu1J+TR2RrQqDMU82XjeE
5x1aYDA8RsnzEKO0GTRqRTAItgfnNKEGrVjXtAOVxzDY3leFMPwGxpNSezsKLhDd
a8CNbM+GjZdWClQXxcRusbDG3TCPJ52DgnO8MX3CGSw3mmzNq85Q7Yw0+k96kpVp
gxSlazUOhvkBlp/E5g7oNW/F1Tw+WVMeVQz8CuWhZ+bAReKM5PEvMGZmL2E32QyA
DtNU8me72HTWMG1T4ifoWbX4FDLYhDJ7bcm9z97OJlhkbSVSK+PSgC7CD5RwBu5e
uye4qwEiUXLonh0V7H5n/xGrt3lHD26Ymz2KMrtkLIP941/Ky4K6Wy8Mqgtqf6AL
`protect END_PROTECTED
