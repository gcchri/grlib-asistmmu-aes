`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fg/da83ao0o0GSVuPWqvygD90HtvRkIk93mrIjgZpXfE46kKSAoKzeRLJ7KsL6Hd
QV7YVWqxy2pqXSN0LpYDnTwHzIK5YfsmVlml30Ht85Sr4YpRaP3xKno+VEd0gTAH
dERtlLZkdNBxUpEi5aEGXoz0EG7hhKXkD9jf5C4NT9l5BNfKadG43SygBdzG4Q1q
/v+J91bDbYjHX/QLP1PV833ZjHFMoguJQxWb/bkIeHnZHSwhsTX8RdSfMq/UG6eG
20FXv3mXLWQV1FnfunTQJXZnox57Km9w50kAVRtZH0ZYP0ET3/d+PL2FmS2zoWoU
7+y3cexiG7kRCqq/GAu8mqNxgUZfupuo+nRlQnaSpCsee8ORmFQj9Zg1UFSpSMU4
Z5zMU7JQm7BgLCTe0ZfUB9HRvhRueCDANYDxb0kqDFgWbnL+nba8dnZ03cHvPSQl
YouZE2WkgWqXK8+FiVEHhsHYJsfkWCMcS6jVsn4+9gm7S/2bDd8wTn07mTLfHQ6N
Bm4cdpxuKjT1LRP9akQ/2ju7E25G+x+C4s3u1jp04Hsza47nBQp/Ohdllkva4E65
249dMqytMnIzoe3CHOdfqrkQjGedAuT64DEXcSBV58/RC5aKkoyS4sxuTCHjkupn
hy9S064ieHyKNrV4jFON8sO4S3u/6O2STxfXzuA7t/7xXEYFf4s01cUuEgZv/Idb
zZm0+bdaKa/8jJyQwBf+jkgfpx7WU5oQkYMNp2NRuBE+WccUWiQ0oZd++rcyeklN
kNleN8Zen1MRZgJ/6hy8JBGf8gRRTprNPLvCzsRrOQBw6L5KTER2cNM+ovgWiqBO
gzg0BWwDh8qdMQY+KxdgFL9v0+Zn1DkvktWTnzUfgVpZ80u+H5uJHNtHtsyBe2vQ
231ODGkzE6hAStm42OyZrg3/5fPA51C49juc9wXxS1b0m1AvoXoVa4X67ITHcxVH
BkpkjVIiCJw7VKkemAHsIG4MF9fDzyum60cPYB2CDZkIRVJhor7ChLZgEzrtAzph
`protect END_PROTECTED
