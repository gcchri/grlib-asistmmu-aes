`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
08UTtPHvbDGsfhRoTy6G2gB/StUUwhbm6debd8uP+7U7HznNSH2PLkEouBvqfbd1
Rr4812i+9aPHb2brwdGFgcWd+gTBdx3Q6OrnHLXllytqaWkqMxdi6EJhCuMpr3Xh
tk5OoG/eY+uSgzX9DT028lcWaXmpQ14Vsho02057Og1RmdjOikiEPAKjoylIlZCP
QAfbFoV0lXqGTZCcE0JGc7/G8lZnXe7y2VApw0kgQ3+XF4kPS4dZ5su7U9vxtC1T
X2WLp9TwXohE7x9L3y0jVs29Baya8KBMUmC2cdsMjGYoH9m7nB/mEK4nOqmWcjVu
097K+1t2F5l/iA69r9Q1ZGQXRdjWNtk2wrUaQaoYcwFPRM9EAwBnF7lEvfmzTMAx
P9ZeD/2hQBhI96UuStM24xAzNehKqMACPzS9M4CfK/6KXqmZxGBrfCP15qbe18J/
wqELIKjwxW97UuIAUqngIRlaiNDf9mB0DFMbsHsAphEqXSCSNyuAqbtqvemSJiBM
N2ecx1JaqwN64b3ulVnAe0bif4lxqkQXfg0Vpw6oRXNu2vEiCzIU+LOtuw0ykS97
f5L2CNIJVhPzfyKV/7YbCHZTHe7o8vQlu7cRBrXUeR/0hHr5x0sdpeNfBFRluJ8I
QmBCP4MkGh3qQEtTe5o97iJqii/mdQjX+NeBSVVNjXfHlXf2gKi/TirjBoGi9jSY
5rhqsSzeDUEcyXDPtst5G8uDwu8WRR9IqEsd+YyDGIZ53oFFNvuM2tQdLc3jkAUd
SOKOw5/PEe/yHFqIA80PomqhHHO4IgayeNROd1PT6I9nbl9MqHiwnSO4WRXYTLaV
fZdPKORdsIScaSj8paL5ht8WyRO+fcYi1DaWB4ndGh4aLs6bs90v/Ruv/fh/+XMA
yvUFIIXmrB6c42KOw0T4WEBRk+NrTnjqt43gTpPuQjneqYEflqVfa7G1L4jlAT6L
jUUvIDVJfoaxy2nmisBKEM9gS3w1lGQFSrZPkU0qi+OF8AG6RQTrKZKAW8/eLluX
SzuuBRC1APG+e7DWVyzKBFwpTJ2vLaqd2CZsZQO6GZlPtsakM7zYkpuu2X5JKq9d
jb1p8ICaLyBxzG+pG23dOBgj96Fk1OUlWTOyXIgeSGHHlgx8AkMmADlfFvlDtMyO
pzjoDoBaKJynQIN+XcENcy4HqYncMQqUChmq3GqngvNEZqRqPPmQ9YnttXFx8aSY
2JspBVcRAUGJBKuZbuHu08OHTB8p6uNfotWJc7j+8U8sVSN7DnSMwWVrARF1d/gl
SBFUUv6rvOkn9iHrSoUZYIiG51kpcWcOvEhQgkoOn9v4rMFiBI6U8swhWJT2eFRq
Bvi/PRTOw4Ad6ulhMAdXQGRhTLDTw6ltRr03xNDzIFP0cklkEwtaXPIu0OMT9qVC
eblGMDmDXD7B23H6z9pWrtqxwBGgiwdBNYK6ywsXaS3le4J812G0lJ7z3/qlIXpA
LCc48KEoxW0NNzDmeMvL5Q==
`protect END_PROTECTED
