`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IkpQw8W0oyaFltJQOe45347O0VquIwkjV/rTO4XX6SU09/WikBg3OUPzKCATpbEN
0DKiGgpjp1i3zIRK8c9nd85Yr3xkC2uwhp7yrNg2VpRYwwYFZY5oUAjOtmvV+lG6
mjt8u9rBt68p3SPZDDfagYz/Gpe1HH+koL/yJFajOPHOsYGJGDTIY5XwK+gdjzNe
u2eTzQF7koKLveV3zcV8tSm7ous/Px7RIxgRbFcmnSTCHX61pmaPZA5IvJBZ3Yxj
PmJMjkuAOTlQYl0WO4qu1LYsXvFOliTf6JYC2Y6qEz9TkNOyBkUoqQCc1nLQRqfA
tfX81+H0OEVf6MsrIAbOZTuqeUUrpR8nD3lzK8MsN03Cxiug+jC0ZCyL8bqrn+2p
Lrtmy/l+LMQY2Bcg7XhxpF4zAnYnR/x9yMASjC+uliHchsa0AK0mgWV/ngfocVw4
`protect END_PROTECTED
