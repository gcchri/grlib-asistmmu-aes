`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rGSfbX5eOxrFx3jbPj2QwbYvouuvlVndcWWm5hwKNknCmHksGbJEUuSk12TnHj/t
FJczbPpT6cnf5askqSJdrkDEV+EIUwByMKh6E9xvAgdqL1KtJdr/0PKWsM9Ja+o9
pLRsR7MZyKpCjkUf33JgMlq7i3eEPIycWW0Bo0zYz/pkYGvR+Ty2unZUulcTk1xb
3wkIGtYiavkpRl1z93zj6sqKgx0DbbsxTAJ81ZafoagfGsNPMO3vcgnpZijgHZiS
pUfQiPYW1oGhre8JXIFks0M3hpm/wX7lCllJlj3Nt97a6qgg/7bL+23gxWZ9IIiE
4sz/QM/7c2C3WQ7PND6TdBbxGsQf8307qgS4ccl8J6P05xB+xmqvxELRtgUCeoaK
kSQkqNSqwo+gElx13cz1eRq8w1G2vw7AtyvePIwnzgk=
`protect END_PROTECTED
