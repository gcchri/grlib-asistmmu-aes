`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yQWt6ryMFWMclEXtFDRNjclGTcfCVPsAXsPXt3/mPWfYhVpQ4VdUCe8r/LTWd34v
o/lfmpzZcE0RGw4WmYOBpFfsMMHKLwBpVxJJROuh5ic7ikPMtKQ76hhdzFFn/hzr
w0l9DICkxo70w2abAp7GzVdSLwZU8fyd2jW4cH5UUcKbxhXUvrBMQQqCW6irN/9i
J2hIX7JcJmEiR0fWih/kT6CZg6oR6s93omRDa+RaDWIcCg/nOUtzBPWOXOVg1Jya
5r1EdHxEOukJFLcLxlls327RtfRheKYaM2jQpnHTsbK8wuC0+wo2M1l23AllEuVk
W8EQiQSSEXSW8ytpbs2Cp/Dfk1ee0K9DegfS2xg1WlifOarhX6HuXUvBn9GFgLAQ
i3VDIbENYOEtwlDBkoyLnjX3AbR+XnBOrenGAQVEXaItY8ezjwY/bUu9LjYZtK0s
dT+PB5KE0HNQ2QdG+W5G9nv330d7n3BRgw462Mu+8Gc8+6act0hAxulgDcixyQZ6
hJoid+w/QA8p9/FYJyzT6tdWwPTx427kZJv2Rpicx/HgILdyttP4O11jrI5w5PJk
pn23nw2BLspbhAp+RQ3gxpxGzqw2tX1PSvOV1qWao7zcpBOtTTDg/RlMNn7WCMmr
yCuehiSvOpt9eRt5ci8nDYopdz29zSyZzzxhgnz3Tc10hhEGgZQEH72K0obzWgN5
fRi9HkFOGNbXazUvKe7ifiqrnrRExGds2aVDagYAS7w6RR42UghIBXjhJQN3xcwF
1EW4esuoJVIZLGiE3vaKNlaF5gYsxDIs8arTjX2gOD9PGNsmpMfLlhi1yV1saVf2
00najJd8S/SeEfpxyWKI3+Oeeugb4JeejWVZNytY8rf08CL8bm67RXUkpCUdb+EF
BGZq/zFezfM0J33TBQkjbXoYPZ2KNtD18M5heVAkIJdw/prKk8VIiTvhE5t4Sxq7
tPp5qJruRReoj97EebtepS9GqU5xkk13s7+jUwLYBVh/RaWEXHDNrNIcSsq5joNw
KgSys6n+wWF1gbAv8vUvHX1wh0Anf9ng7WyAWrFR+6twQXr2DX+DHW3ISeKx07uf
WaSW7wa4sk0hXT0oxdrLyLCnIj9ZfBWxarr2P+rqg8brIwdStH+25RK8bM5oj+q6
dNyVrjCrKRVDCsMDXY+tje/8K9nxKLLrEmsjFl+2GVGqmbugZVQ7rGSZFVmVtDaj
TnHqkfGqHhpWqQa3+d0JPlQ5zHszJ3WcFdYNhlSNHL18NCMlhTQwCD4LTgHsadSI
7i05KQ4IWmSTnEqrCpCwTCBXB7MVsIzU/eWjj0CYYR4s58fkMfnzT1PiYxbMyqUj
OlfG6GI00kLbJIuqgcEdbcAEEImw5z7pW8yeowS9/D2VWfGC4EXnY0RUy6jgzx2y
Vr7V5kg7KJGUGW3RtacAYQnDGzGhfgnuoFwxRmKcyV1kqTJeaO8Q3lBpVPPwOYNW
bUSEGyG77Z4HlNmey2gprXHUzUQCF/AsgPsNiNpihVP10WgzUIZnjvgzCFS4SfpQ
`protect END_PROTECTED
