`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qcyZoMgAxHVevxAZE9kBljevEeLAvgZkGR83v2V+tY5aC+UWnwsBDuLDBnjn4dSy
zSZiyjLFuq1djUWkAnO0hZP9QbgfysNYCAEIvy2W2d+Jx+lGvCDQfhgm357bNUMM
cDU4ct7+0JtHWe0QVE7HKYIDVcGqEkQjx/MTvaenKLs2S749HL/2RFv9mHErmqC2
maR6tiByUm4l+ymRWYv2lLNdnyMhZ3XOP+5kjSwii91nSY6RM+TgxOgqEPcefMWZ
sRqi8/c3Av9Y+YB+7u1MgJGGg+7Bu3KfZjx/pwTm525zfITq0qBt3RNKAHDc/UY+
5ITvZWIzd1w2OUvEP6E/ek8ynLm/+9bJ43WO63mgMtggtMJ+zvnnIvK7ymtycrLP
eA2DBZhrXzjUL+OrDqaltuUFZ4jzbc2Daoq8TQqQg/7ms5SOfpBRHtolIwLa+QJi
H1UASU5wLav8BxGd6n/ifCdHLj5ec2H3MyvwwkcBH42yyOz4ZSm6UwGrYSogyH6k
+BkBtEOiberh5hZP4Ty7vR2UhBlcaqyWL8o+EzzKeIN+01hInh9nf4LGSWX7ExHn
YhhvngSTJiOOPro2m8DGBe9H8TaVywbqU6Jpagp2MNJhxd2XaYl/NpQUzIh9CQrK
YB/aIOWNqdcQfSy3L28CtUEHZls96dsF15cj9S8dpNsGADcyD7cD0ZpjTqyKk7uZ
nJRPZt+ccQW5bd6xcPRQI3b8wUxOm9hyZuM81kwuqKapZI/TGU6kDeb2mJoswxYX
mn0Ki98L8x0xjqqIFBTKSW30LMmTwt4jywr9Pnnqxtif8FBLI/poK0DHAGKREvis
2D8uuWjgDRiNcZx5ujgC3XGZ3yyYyCf+DnqUdfLopjkjFBgLO/8YL8emdWN2i9QG
r6BCB/x9+YFeLkJMvwivIHjA8qygfmhPWfJ1iTr6H80j6QUW5UUD9CNOlsGRFVDn
HbmK8WhdllhTw4jyaGhe3NPsBSWCZqQPO3+fLMek3id+twGwFYtHiJHzdU11YPSp
NK7Cf7pzbVLdq1lKXhN1Xl9ZM1YfwW5/zLt6LwO/HNUShz4wyCCx6ZH1nLJKB+Pb
VQMK8cap92NV/YDqo6SNLg==
`protect END_PROTECTED
