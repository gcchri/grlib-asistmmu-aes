`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FNfxGJ4ZtZ/pVaCu5zxu9dYsMrgjV2YXx2x9gWdOcvh6Gxz2y9vhOJY7xQEFjFlG
Cq+dePwlt00CFQ1Vf3KdmJyfHm5wTLSH1VdU8wScNTXKvkW74wVvLkGcT/7Sl9vk
hsibC90z4WL6EHCNvEM7/WIWPOTUUYLcJ+FOF3lcRhz4MI4izHZVDT5c0VEppWCK
l1+UysFH+ewzHhR0cAgDvHXtsjxWMuJA5vFv63xh53YqUvmjWJ0vEZNMt5BVa6oj
eyBzuhBWBS+3Or9XKfhPeNmLL9KMwnvYDC/XLdwFq5yu13MbgrH8aL1EHGXCWBYj
5AOJpkqSwsfqSuRJQ82JH7zipDOV1ENdKmtUxRaEZ082HgN7x1bniFFSqCsQ2Xtd
+U3lvoUtb/gk0Wfkdm8DEPMU63GRj+jFkv2I5PeTa75eV+0O8aDh4uRkUeXw9W1A
nj2Sg/T10hMVfNt+O7K9t0fITVe0AVnmYLWMwIzox3mvf5oLtYIC8WmhefIMyT+m
doblNYPBMSmFwspYal0V85vzwW4HV6b60gs+5WzyDrAdkQLpF1g6zi6tVCfONKMA
yOQQGJXeZ1+3SbIMbKZ82XfOAb3bQ4DeGlINP+Vwuy8JLwJ1RkCBT0bKh+BnmJ9S
PYPSJSMqULeDlPzLYgq1FwUP0VGb7cKYzFH/9uqQZYar7Tid3t7ECBXE4ROlQVNc
2ngP1jIPRBMjFqBgCJ9CJdEPMt3c4zYxv9ZvVlW1hwe5K0EfSV5zMTUXg8wsiH1F
0WRNDm/1Lf7Ak+dZZtr9cRtoHVUCqeJ+9qufpoR6I6J6t90UwmjvGIZWXXcCZiI8
ea0g8GXNlCU2fS4ouaSw5SXC9k8Rdr1XLbHF0fVFvlm55nbGjgnWwELGL1SN6uPU
PN84l7cBnvlaitT8m6IIfNt42n1Rh9uBo8vKH0SOpzk=
`protect END_PROTECTED
