`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xpdoloPpSy9lnGDq9AyFbNzfK+JZWJ8Ba1E/Nv9bJ3nW++cgYScOvrpJXJb7MbwX
u49KCqbLSBLD19SkNMqSfXOE0twkBw7TTeg/wDZlNAej/9Md+iY8gftmfj07Q6YD
kNtD2uxw5CbvqzwLQkHWLsJF6VqngPWAQOkeS3WSweXSi9u8QbMQlYbvYaMaqzid
ENgMtKaRnYQ49o2shOLVG9qravaba/SsQJ7Ax+9TgWMTTdKoeYPnR3IxllHrY11l
lvU1PPAAaKleLMDGElRWf3zMYdqZCHqrrPwmtEO7oPlhkzWUa5WSZomNImHXA1rH
5cOP3xIMuulBXiXoR4g0mhHW/EY9npa09tm2BA5sD+HN7wHM8aMC+TS4qj+xxInL
6mbXdbS6qzfx893cWiTnk1RHDmtraW8qryHrK+S8D20=
`protect END_PROTECTED
