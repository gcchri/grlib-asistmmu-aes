`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r4rlCuzUyoapJkSGzyHcM/oB5feUhbUQRPjxDz3N2cBh0K8GKgYm7NMcuL9mIa17
XhbjT0Ns7VCVxfpKdZlOsZf6Lm8AF7hzllhXdTMfFj43lDYZU9sxcUpzeH+i7ZWg
Pysm+hwEg467fQwxvRHQ/ojHo7WXVcCKUTvAjxr+WKrZo5FlSOD87WbkuzURFwZd
3gvc0R+Jdbn7Z2/FJKAUpm+qiNJ7LZOZ1n9ucteDe3TW5d+21Aa1kXKL47exOYhF
O1etOFXG6pdQJ0oczg/czPjlROvmAy1sDXAASgkWczVCgsdslLZIw2fYIyR0+S66
sFuL4+4SMJ84FH3yNxpA9RZv8Bjv7YgMmj5HtpjEj6311I7MpvwKiHElFK4k3UTE
jVRVaEKkvLNZmgCacUB1SQ==
`protect END_PROTECTED
