`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QCXQ6T84qaiXz+TFc5wGSsL1KTMjlj5xkhBZ6SwinfF2bLMTHwBHFNW9yz1yOqlf
tRO9u9/rovFLGZJ4sFYsbbyYK7AXbDcUzBSJwqifKya52XVbDG0w9ikmqqWiTz6q
gvZgIfpoZ89FXUh45MvK0ZJ0RuLBhTZhsTguZHEFhQqx7VTtuL5JA65zmjdkX1nj
iQoxyqXAvmoJ/wciJryKslXwhQGim1w2AoU/PZ1MwnI65eHGnSk7Bi0eHsySD1i1
fN9+rJG47AsN0BvexY5/ko5b3UXCNi2ZVWBsqawx2vWrVhVQhm2IKIEgO2pX4jMw
pgKO3jcB5hTXSb9L/0j7GvXGSBWHD30LHvNqN5X7JaqvRYiPdf/zIm7OQq11k0da
H1cj8OrHPEP0H0bPlZeVxIYwM6zoT6D7YxdNUJiAo58aYGNNKgXs405zv0m/gfUA
g7n4y3uPiYJ5m6hp8AFVu2KTtXCI8VkQcFMozxwheqRIA//efNR+aAUa3mOYfejP
erd+662O1n19KpcYB73E2PQMmOi51TBhTmaprDF9MegMuXs7Oi3AHgZ6s6Dpu/nP
dfPCnNEMWWaINy+NNeHwQOTHVsXNJuaznC0plZrldXpmPfvDFOjDAs2HbczvzzMx
FugUCofms0gxxHkZeYXe02XvyCKXtC3LYS1uY8kjpC5zhLHPWhNmh2nqpqAzccPW
KhOSM3VHugYWk5B6gTNc93Ahx9oC2SyLHXw0RK1F6Wmz1n3RjeuUN3a61aNU5G4K
kS2m6vBbY+m/2JHnmEBB0e6V0OaSTja57tLIHUGFrFaCmIwtV2A0PD5zEp+HdDXJ
dts4Fkgo+m0n0vjKDEZoiYsBOK5Ul9jfxC0oMiNAPZAPiKy5D+3e1U9S5EAFbLQC
VfP4I3nIExrUnXs0tVjfI9vLHjCZyjElYYgLJYYwqIEv5UH0b4D+j301IzBu3s0r
eXUDgw9xkaRIeVWHa1PI8oLJ88tXoG4/CkvguNowuidnqGxYLCL9iASbYeFRjqPq
cWmaUutXLGZq2diVJE3mjXX/JugC6CjPuyAdCIpwEezlrggRMX3z/8shigLG67jP
Tafe8aDRP2u4KvNsYCzbPcqsbt+ovUnoxLYSQwkhVj1vkBBHWsMFzA0/BymLdzeg
cGowp1888NCNBGczvDvHBm18XHtV8HaO6gu1GEHsgB/1fCdoITliBKeu5/BnSJFK
lyLQBEBlTwo3QVDCGR0gaVQjXacPoeUAHtUfSS5ImQE1iXykd81uU3Bz55FnPllh
vvvDSwr/OAzHXKgmve2unFToTum1j+FQCDetxeL8qrVaMSM9GilGHOJmVL4/eFVQ
0hI9R7q2IWQhxqlIBv+qTMoO30Sm8w4bhETFBk7ilAu/TDsMC+iCB8+I2OL9KxXH
08ia2twtyHwOMUuAQB4ng7c+uSCmYKrvyIObFKlyxtOjtKZgeRcSbUz5s/4p5w7x
N57IfJW4sCBOorY3QKmXoz5MH2dWLohwF4uevWwz67L46Nat4/jBWzKcv4EgxDMa
N3Wm4gspPcAFELrxq0kAL0+/TBYcxHxudBZf+BTb5W0Qr6fBtbBdpcaQIDaAFNOj
sEPPCmoG9DSJXOHKeNl7VgpiZvrlESZvk/FWDQtbXPpiZgSaWjEK/jWuUytrvEGW
zz/7y+6IP4o+WPhL9cW0Dlhi0cN/i774kMw5tF0jQ7FPxK01Z8U5DK2VuWW30tso
Kq82B3y3ExVcb08C/g/3o3MVc5UiH7FZJeKiCrVASu0JraYeIL/KQyIDEf8K3eqS
V4agDxkJyzIQPk9kKMi8epUXqF2SfVqz2EkAw+f2WyEfKlSyuvBedz3k3n52+ZzW
cYIfpS5OUWTYaA6KioY6DsbvBqriaOlw0X3irK5YyBAkw4TAQpJEo4ajFpAGc7yS
sVZc013NP1RRjwmL/uGyGPO4ZqNPEyTruG+wwakn3WIBkCBj0E19NP/o0L6JaiGM
AAi/yURnd/sZpDUCSgDjiQ==
`protect END_PROTECTED
