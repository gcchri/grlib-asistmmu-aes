`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/tFBQlKAzNH2O0DPcmO6c+Q4eR9gLMEcwqNERo51LdJvwdJEy+U8logzIcK01dpq
dEkXQE+7W9tUu/46t65/5vJtIQ/F0plECiQW8RXmaUzGBxt0FgmMuwsqIn08oj/L
b0eNOArygaeFMDsikBNAa6pnid4SDKkz+iEd45C+2OUfKA2YNnIsIyWEgQEW2OhB
V4HQejuaDMtuZmVCuuDan4yJv9xaN3G9Gn4nzDetWcE9EZmbhjGbGFr27Ragxlv4
5+5+VDPTMzmmttPrkl1EoNBqoeEjwvx7XfervyVPn/aupgNIYPZLhQF8O636sn4w
n2bZhddbkFNzXWmCQwcSITdgUwxsrmsU3l9MUtfrUOLAO5lbooiVdCPTQE2Ebu1Y
RdX3H8ATSHLvlCoc3ZSoqGwPmDMehxZJm7t1P4R4NQ472I3AOxuaM0x6cvUg3s5d
MlyorEOHucjQgc3IUzokb1YT1MTF33wM666zRgPO8s9Wrvaam2FgSgZgGl7TAZuY
6UExDs4pPMDCmwzlVPwMY9Dtka4OaiS8Y7JeyKm1VfDfQXWa/gZWOLf15l34Trx5
M8HgKTRe5ok6cor4PHvPFI1s41lzH3S50hnRhL99pCar2iKC4gZzaeJWcAIRVPIK
rCs5S9KOn8b3SFmgZiUCR0jZW4UnWAW9OeoTQDmB3/pu2Db0ZpWWcZg4gsv79Xjy
ro3PlLJl+wiqRiQhzsAr1nWuSa1wvqKZmYF6sNXyTxo=
`protect END_PROTECTED
