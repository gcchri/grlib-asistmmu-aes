`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZfwsgUSY0SlO84cttSFX/PPrPELBmcxCAuXzkHlS5Pe/lL4Rn4osmmlmC9WXu49
M1oZLrogezpi2FKcGrn3DI+cyh7EiElRmgPfsJu0xnNIJ9BC8iH9den56dQAyCoM
lqFxGrK5q7dNMA48Xs+W9JeduRB1Aegk/xaFk9XuY5NEFCJSCZLZG+HJKvRGq/Iq
+GIRIfoIhWl4l6agGqByUs+GSX9nAQ9THKH6fg3TsFq+Y0W+PTQIfmDV/nXvcynu
vdei1zp3yMOaQ3P2UXgz2ZqNSauqAXY0GEHSosvUTpCUE80NvyyJgkvZzQlZmbbw
GmB+F9ID0C0urzJloLJeJ/F5Df+BVANTj6CWdPXft8Cxz1OxAG88pv2GS+ODfP3p
qKYf9CDB2Wu+IZpqj59wIJVJDolRQGD3BZFKjE+vL9dcZEft7my/HOWydhAG65Yg
`protect END_PROTECTED
