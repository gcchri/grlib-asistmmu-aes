`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nmgm+6eek/WrvfUBQa5A4nPPTssNX3eyBB2yPefi0hhLSC4T8tAh5oe+loElJ/gt
adQ+KI9tEZ/pBHpoznO4tCehZV+Bkkb9skNLK1pz+9hEDABhtwpbLTCTeV97tU/G
gE4jdPkID0oDuOTbLuuYmkoapqZh+8lqeKMDfLvbQ4ccFzHBMQE9ccL/sLR4hCOK
ALhBRXx+7RI6mKnNtK8wLRh0ggO0zl0YvxH9V6ZLR34bVtIsuOjTku3lLmbED4tu
EZrtWapHJwlEaz5k0Jmm3136qEWflQkIgnDOx9DbmBN8e6RgAdkMuruTEcOraYsL
B5IYZ5Ig9pDeXHcEev5h5POZL99eDDvplsEARJrGpFmIfw0L2dr2oxsp4GE0GMvC
1RVaDHPCNSYqjsN6f47LYuoc90sdS5rXo0gut65GDTM4QxkJ2bqF7wnwsectfItE
EjHLlU9cmcJq9zt3SGgEfhNFJHHmLDDO0jj0Fywu3N4T/+ozpSxkqjcNrA+k6iVK
D2QRRL3MrnOoHVon5vzrOEkQWjoY+ZYILMpmvVRXgoeC6gBjDo+HvN6kS9JC0+il
Szjb+YVqsA4irYPRqo+62DZ7bsBxSbY9H4RQluk98NWmBx5ZIpj5ybBohbVteAGO
HYkPgpCnb5ILgMRtx4Quew==
`protect END_PROTECTED
