`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JetW3VTCvmTqqluN8cUCz3N/i7VrxOH9uPlYcOPyYKONNfzjkCrFlzRF9tvNqGte
1F1Faa9ET6wkIGb1C+8F2snWj1lQKDRGovSYecn/WsMfyO+4q3XGUqCFsfu3PXUC
HFeOQQg+xdhx5feXWmLErQx2MsL8bSfEEYoJJ5fhG/7SDR/hddlRayd5j1pYvBdv
wTIAM2kY1RYcfHfzIQcC4rh4eaHfaa4tkK6YUD4eOp605pEm7JuaKZ/LQPJjZiEo
zpFlAL+NMmRvLsuV7nLSlyX4LR1A7gU/m25MUn9aQgywuLAjW4WxgoXEsfJUfBqC
3Sl11xIJu7owvL5Fi/nI7Ib34AB7Za1lWjrfq1xXtBQWcKq3xVauKe5lHPviRRUD
pBLIxchInwcbY61hNGP9spCSOs94rh19EQQ5wmiEOezqhZJki4e+tOn3KuFoZNtw
BNPMd3E5e2D31ImDl4L/SGp5uTv4IiuYKxjfyMaOJiU0hEuIsPSHKco99PQDVQRk
noWsqB1u3oNxjlNewYAgwgz3GRHCasYIVHxH9OXK1ROS0iSm6o6GOf3ZMJ5DX5MO
J120Kym0Q1IxXyqV6+MppG+90sZaq0hGaTJpa6EenAG6mqPce7CWOuKcKN82AA8O
6+ew3FsxAMDROG5cE4v+GlT66Rc1wmbCSh1HvucuvU0zk9XNs+zltSqSErAGaSPs
/hfXsDwpJhE/nDtoTTnc8D+lNrCZfLvjL3iD+DOCavk=
`protect END_PROTECTED
