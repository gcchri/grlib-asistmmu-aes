`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WTfy5ZHwaHNaeBoOha7vCJsCiL/czo9m1bHJ3j7qf7JT6ahua07wO3d9TjeRPTQr
XFl07gOyN3vj9kYo3X/kO7r2l6PwGm+TngL6eQjTRmWxHg8lJeAr14u8SFYDGMHt
BKLuBYf8/jCqTRMjmKEh+L9uvxwGjJn2Obj2wu21bDl2yKFrY0nfrmjyvTGcOl06
5N7/xEEdkdak59ZZewRKZzOsCCdAFg8eNbHH5OLzlRXZC42CSy7y0VpN2I0rD2Id
qdYKeKCt0X1KxT9HvK6yxNdZCh0Nl6m8j9W8c4VOgnwqo61qBbwh6SX+V1gPm2cO
z9+YDd9YbbwS+D0Ybq76uMWyN824rLg4Z9YmFeHZCqk6px7QZCFUn9lBTBN9BsUR
6J8Q1vbMt7LH2yZM47n0LP/3kfrf/flLEnFemfyCoYVAmD2No6Y1nDC8rIk+g1HK
oYgYnhdLtYrNkjh2ZtYgwxaU5md32bmr6Qbk9snd0f1RBvE9wucgM/ZqMVL1EBzy
ElehQhUVlyL5ENNzci86jSy4vc3HLV55u3pOySKLwcKDrIe7L9IdO6W40szO7thd
cGl+4TeNl604DmVs8bP1iCZONCDWtHfh/GoANdiTjIf6cR4j7WCuMiyStVEfo5x/
q4NDip/g0RMH/NHp2jK656+qdgLaa0FJVRThIZ/WoS+eR5E1t4cIH/by6QLTJJ01
RLrirduFtu1hqljkN3RsqZHZRJaajPSjdihzz5orLNZb+RreqKltB60nVBYwOCpr
vsZeWOZZGIS39X9vjiV+wg==
`protect END_PROTECTED
