`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iY+mD2gKzOoGxUXV5tnM4pEbY3jLC8Ofinkgp4P9dqGpFWdWwKFqyY7E61jDapnH
nwb4S590PBKekwskb8M+V0PBgjz7NE6Bqw5pgRuXM6hMDnJMkUQwhodKmKDpRPep
d/FRGQPmHAfHrKUe2MoNxelHPvNu2FJ3zRhkwcUzA1zBsYoD3tLgC4rOHqxaU5fi
YxQcLhJ1hF9tQtm0FikoSTi3Of7tXy6MazNwza8qJAy9WJ7gJTBxlsAH1WCdXE7M
CCZyQEUltS/Ar9rJgwdDDCoktqIqesSi544M5Eikq7WW51vflKPfvPI6EL+4Br/j
oETj0qbrLqfICXKr2R5pLYut1Q76MeMpRut7HQIlIPYSrjrZxlv/eMJ7nmPVG19f
752P7h/z00rS5vMM7CYfqqLcu3ADpzMA2MJc0zVn6W8SUzExTXjMSBO0kNmRoB+i
HOlc/A4ayFZ1zGoYuokrOv8vk/OrIfIuTv6w00502UZoGpVNvb2DNIpFLxVTCQu5
tG0X0ezoNjjJBbDpc+Twu7Na7Gvd0sE6Lt/hLAPGO5F3QTmN5hHAJiFqMytCC220
bz7pBGhI3F/TpbQbz0lGJWoMIw/jrq9nn1RYuhOJOV/KFDkPBZNjpKVFyrtXs4tG
wUvJQM1Bus+5hJyS7x03B6lBpl24GjnQ/P4ROs4lMv7mJVNZcu/x5HH8NtBLyLqH
KXsDO2uiPn1CWqws3d65jmD7sHob69OPWi5WppVQjsZtH5qetyNVwfrzx55fajyV
YFZfD6ijO8/DrI3ZCjl7vOMZRAg98wY/MLwubBiSr37N5T/GilhDz/dvh8atOf2u
gEu4FOjgY6sRfyymPoctvzA7djG/fgYj0iSQ5+Lkhj+5lFn+SRQWiqNPdj4dw6Ze
a21ynhiTFb9LLkStnM3vDcFkSWXA+VBcqeV/sU2NMilxi+9zGeBkvmN5yTLSgB80
ctaqu70tH5J2IEeKfeg5Hz/pSOBci9hlGhGcEJ8ErwnFcZMi0IzitQPzhnAmoNsy
vWxA8fJhjJiWgXk+s/KmUsfgCMldlIVA+Sw00OzimdF+v0xrOtllzJ2eLZci8n54
qClpDYzSmW3RKDS6QIC2HyDY27SmOr/WK2f225mjluiwF/6djMkFDVMLKrJj31q1
+ZDcGAgrC0sxk2KhTTIkmKY4GtNQqW9LjfJmXf9PJq0Ri9EsQV8PcLtfiSCwnvIx
q2kVHAMIiLYyGi+v84X0Qm/Syoib5EJGl16hNNRecMp3/MD+kyKietUt4GyTbv2W
UzSoV40Ie2TY34Jy8Ca6fR2BZwadCRdbFjS2DBGz8apPi3g2t1YbTQQ8l9/7E385
H171iUlUCk/E7b8WENDJa2DczKwbEfOA/1M/aNBokYB31ULfa9esCxw9JOSLK2hl
yVUWB78pb4D0oLjzI/ZWTDT9voimIit7TFKsPITv9+8R5ADXynCjo9oZWowykWKz
/7+tU4B2TUqVqGGgOCURy3k/TtO4gLN4qkqloJvsZq+JeFgrUlWMYIKHH7rfchts
v1y/yYjgYpVg85deHYzXG7Z4mKPv78g/wMKwuDjn9T7L74bdcZQJk4JOxZHRgJ0L
qYSm6KVOco7o2Jm7ZOOVeoS8lajz194uNcoiSuvZxA2hl4RqTxC0AptFnlP9S6TU
dndHK7MZ1/rmbI9WH+SF4mTJcg82cCySiH1f817WOXbPc3PJxfFZ1dkbZSsUHMBP
c7btj3MpnHYxCiSNp8bL8jsnKeVGOoY/WcVLbxZxKZu8UWHVBbD7B7pBOAGNOGyT
piN9jv6l9vtHWUMwJJit+oc1jAcTQDc3LlS23aCEDf3cmIMgn+S8W4McTMD6TJBu
3u0oi9O0DKwGoBaNmKpi/kX4bJ/LQc1zkBs3cXgAQ63nj92I/XL1GyATWQ0x2wHn
po0K7agon1hBKk+z5nv986RqtxYIjA/nf+KDK6GrHdMy2rmuM4HaeMRvMq0/yES2
c4iq5h6PLqSpPWmRrIMrxpS2I+nW88Ce+/WEb+Jxe2dfLODvE1UM3B5rkrcsCmAq
GotbAOiUGlRWebvFBn031yn1o73iYBWreRu9JRFLPOoePhLVHqocqgBzjW9z86fs
HRacgA+7+FREE2R6xTvCF/3YHcMVU0eczZGg/93zOwggXqgutqFelVzhAfwJjMza
7rX5H64S5z5BLdLCljVtyYJiCkl+/wdO5aNYrlefAJGUa16PdnkUyUZcZMBgWX7a
woXiQpTQStkNuJFtC8vF9hZCykjW8A88B0mg1I3dp364HIvlkwnemQwOYrLZnP43
uDa/fefgoj4AYxMx/pn4BWWIFWVqK4aPf42hAf11ZqY1CVFzDi/nbm45Smz6FCDy
cMGrY8LaOMlf/dzCu2o64avU0Pqei8igQveEHxdreZnuEzSp4CtlxKpVCCc2dEou
DGuREJCqQjsVecrdpk2X/s7PDLFen1pC6SPk1RgIWRm38ADooURrtMyDM4kgAiX/
ItsztcTbsBk2JWNn1B+I+X9SPkoyFwx8mm2GLQiu53+s61+Zh/LJqvKj+Q62hk0h
RgyYPVK909RuwNdoRdjI8WDzIsclt/dD48WlW7H+NiuYs86FUc8SzIeURYVqe1fW
y2mxXCK1X+KyRN1yDOx9yoikupmsMg5S6/foqjyZMuBAiSWiXr86vU/8GA1cDTIX
qvbCRBo5uclel3yYxVR++K8bO3RE9b0R1T3OVBq3vnhbP5wnbNyHZK0LRAJZxcve
/7jBNk1Jrc23FPE5eeX8gctVCbpS9QPQYNZCkj0Eo5ILC3MuaAL2dgpI4Mo2VhLL
ALCjfbAPeLqMxLKfm33hyfGkJ9KO7Q5QGR5MRbHmlEYe+rg3HLFOHXGvWP/S5ZDK
4e2NtKgQ0tfwxQx7NVf16ujJvUtVYolXkBjFLJvK+Cu0h6YQ6G1a22MBVrTwhlZd
+dZAeeMZlfo4f3otScbtt3O9kATod4pXL1UUYYQ0Zd6H9Qdqa9kxRPMSseTwSc5U
7iIH3FUP8k0QYdp8V8AAcuaBypyhOkrwYkiWm/WpUuqvdxExmc25OG5cIIXzQLkS
kWPTIVQsQkvSa572cn30T4hd/lnfIqem5icw2IsOGcgoOfKHHyR35+zMgwWyL/kD
sTAUluswfqCprsIAUoVSlyXn29iSOmN6MkekGtiAD67T/f0gDeZD73svQC2YiRye
txwnMdil6sxlwg2t+eE6QHIkVE60gpsYyhtwOB2E8Iz/QmCOE5ewAmK/BB14oedZ
3OKRKt6hxXoSmE9nLrL4A3Z5dx+f9QygpTcX1CsL1NspePwcwU6STLJfNQAKJ0P8
B1hVCBa5U8ju/KspdI7mI/NPi8FTcB+a/TsrqVRgPmQBhAHGmq5pWn11lvg/pNvv
K6q2+SpIW7YJ1F4kJFIwosRogoCESaR2qN0t5oASn9rd8jjV3xKEqVM5ZFj83QoK
L1h118FIYovDAKXdYvGW/XPTzHc4HuH73jx0U74nOZlZsHw2yzSn1eAa+Shr7639
1/iLOlAHqYXXnrsNr8JTcBqOwR8OGwbuV0TCWwIzUCS8Ki3UKxOd2HYrf8RImGXT
tPGsABJyyifCSHaRZCns6zp4saej/S95DAYwmvgN1pI+4Zmxe0qtloBh7Up4aTNc
xxyENAzK/QpAV/6J8npaGh+3t/6o1IbVZYsHapDvyLTkVf3JhXfmHAmHXRyCOjgJ
5F/N4ifjOFH4zs4G0cjwcWMO1ld5RBoy2mmZN/eoiwOitYCXcQLltRSeYkt/fS7m
nuKvcEF8u49QS6BYrt4dzLGuWZN3+xmHs8dYI6vmZZX+bNhvxwfEOq/VkgYDkmrS
B/FnqBpMvePBbIWKy5QKKU7AAN+yaMbAui9X/j5S7nkVxt4Bp2uUdu3nSGQpyuKY
qpEQNvDfQMAkALcyC/BIYk2/0m06JQ3acwQq2qspBjVHM3Jx1TNz41KVtgLdaxMD
0xQCxaeRELE9rV4im+3Ll8PrQ8K2EzR2vzLcktUYn58ea86GroEfl9gQbVyU8zst
X5lexQAzxfte4nqSFPBnxcUTx68tOBKpBvv+nYhvzqpFmDMU2oYjP67gnBCS98Jk
DUpptS+Gj9ThewWR2p8xGno1KqdktkMFqyyM9p7i+at9KxE/JBJrm/HwxwGFgdW3
yY+sK7eLXJva24G1NZ+Ui+ZEZh9DIflPuYrH+JSgBHh8FBnuSrAbqeWAIg41fiOD
jzpcbaOiAJIqqfVV3wnnx+pk8hlF574hprOtvpDS5eLNbljyVODHIg0k5jNoiDhk
zOH43o94PdCS7D6LckuwEbxTXEwrYk/EeKsVU/Nh8tTvHwO95u5AiHq7my6MzZr4
yDgRjWeGE+vfg4/1utXQ7Vg3lr8dpCB1B8X3Iv7M5Ss3Q01MGBRgWdqwlMiPRzvT
WttoePzyeZbjSrqU3PG5du7/lMGivm+kWXA9gQ0PFdGWoijzgYocweYRp5wdCePT
ysNBTzNBNK5rLAewD8yr36MuF0/N0trKSBo2D163JeWvhuiCGfTtrpUnOYE10Gv4
deyt/kEtgl1Yi8KKtkMrV0XJFpFMPrftMrEH5aGiC1Nh0yOgH8djybLrWzMS34am
/gPOkUdetqHOiS3hymYzAQ05F9FX3W70BNCyqPcbRNayz9LUrCLs06JmebRJWBwB
b0zhtRN/vqJXP+61938qdGGkBEn7g8EUdzmTPm20N/2MiDWbV36YjeX44UwvPvYS
wQ0u9CIf08ekxPfxpETTiZDM9XrTMAk/YtMCZlA3ziOKTE2Ms0kim5TE07v4U4Ky
EfKgwCDOwRcUw8S1vVCwDUTOUIfUWPIMBDPImRSJd6Ifb0Hi6aByd03PHQ7rI+uh
FEbkdGJwNho9y5m1pT8iFeQMUGRlFapIXxvF9vlgRCqw3OmGgnL3idnrsnEy0Bto
uO4SR8jV2uR7JempJBBcuTWy/H4fYdn5jwcDCkclUG75r6dev5GtuXqHVFP+hl+K
01ATb042lCQfszfsA3MB/iLebz0otB/mmJoLJtLU2oz+9F3m5RMI7Hdv7wioKhxD
Ojft2qQFFrqhT0BcaRyHqAOmkYiHEk3k8zs+LDNldgFdbNRp/eYNNm+Xbjw/7Kxp
gyeVsKdbkswqKEc27fSm1gpt7+lnPvx/GQgefbSC/paIiEFwTrAqEk7gTMzeY8bf
EHPuwtSbeXZNbkBmoHOYMbQQCrOvKRxebkpTPQxCtKag6ONym0D/3OMmkLCUVukh
eSoSoI52UbnHjGpde88wT+KuwyiiK8v996031k1myq/lMFiui5lfozY8h/RwvvDQ
kjTZCvmRCAl50Y1a3EX0zWs6QHO487wwckOvgPtqa9E/5ehXxgdqXMC8AQZxWBgv
47YVlpVNR5M2sN1GNvT3tVs2flDsoSPXvO1d+xCJhsjpiap3MI8OiEReG+db9JKT
aXSp4w/ze4XXIBslzuiaxxi0RGWDMw+hKLhDrXVgsGpIxK5L1hoL56L0zlmziO/Q
aQWRTy0IG/HhmY3uHg2+t29czplPrET9qtllkNW6lWvWk5/HOi62ldCZncP0r6Gf
4LtHfHrhXRGx+ZaUwYvrgHNDwcWUMCyXDpufkSDPYWKyAJ3HNkQ0QHa6MkMPlzTB
TZN2V/XtdowUZT0JHd3kYe7HYEcdP1Nyn+KnLroEZq1c0TrVVVm3xgGpqXIFu8kB
dCR6/Au+gvwSKu8/FJ1QDqwKwysRCc6N2sv2Q3Ua6LC9xwVU/akwYPZXtuD5UVGK
tA5j3kKSmA9OASXbJyttXixVVLi6W3dIFqvDQ+AOdt1bDQIhF7TRMW0GhCtAoa7G
uSGozy0/b4lY33lyU7lh1VQv3h8dP/wMpgYnLCqXNRazkXEqKGQnKIzbMeeFBKkm
jhpATmuurnqzk49uIf2M/RVEdvhj3C7IUiaBd7wW0dtNlBpjoHSf1dRg3zxkjZcm
KF1IoFyoPj0vsOIvIbfhuvqMrDA4Kg1jDRCS5BD+3upYXIxFCKa91woS2L84XvaA
EdTRvNuuwqlEr7Uh66eSv2iCsav0Zs7lzjPemPwSXbGlPRNfCzw4sKvS6gZp+3of
E7qjgzpYAgXFpldJc5i12KJ4sJF36wX/+xWvQC6+h0hrp/RiCmqCvoNO/JH2UDjd
gFQvHpmUxYnmE/PIJPEUQpLcfdK7nPCvjpRHh34lUTOHKW5VnO+eAAzU8Db854sN
pFcZZ8ayxjESiSLDuG4pRjz7KuyKx0nEMzM5lg/owcTgEOnzV0YptXSMFJ1nlg+4
3SjvIKoZ4RoVGXazOm6g24TxFPK44C6dq5FHXUBN5uv4eppYEeAMB7q4JV/HVpV3
5EXaZcsrK9/GwE878imcsG5diSe87F+hqbimKhoTOQUbhSYWWIOj+J1ABrVtNY5J
6NJIlrjoFMnW6/RZL6mzfeVhP5/Fk3v5rYbCJ41j8lpyoOTidSkbMvQbW6hx178O
ChdK8i8F0LGlN5FL/g3ODaU42itcFSRwf3H/iD/PBm35F5sFODHzIc7/vDmro9Ss
1cQAjceQua+4DSTUvM5EYC6BfTFx36FrKI2wNVVEKa0rtSETy+63rsFGjaV45nlC
ArE//6NYClBfkZ1yIG/K2nLeU0eUmFpzoizPprJCwe2nqtRERfV8s4VGMFnybCER
jJn8CveznahVpLje61JZeziaRHRPDDmQsf/liK+DS5URr6g6IhNUEswI8+6cjg0R
ASm1oxu6dagOWVGwtHt82TMeecZFm8of0DUO+hkL4nG0G1lXesFDVrQohtEibQpO
eh1EKZjF7tSkoJbRm8//wNJKbZBsl6FfwOlgq9ZHEVXxDlhQkrU9Akr8K/vTAtMa
vUPlTBrcQJBILs8T039ko6rr9EByMa++5lBB1a4x2Kq2JqMU/zyQunKFyGG4qeMm
7vcqjCmECZwgkBveW8Hw5spZfMkh4WHDfvQhrBYd7dgiovZ0P85P4wvEFl8nag1Y
scafbuDpBAcE80oLwKoBy1BdChb6eIJ6ejkD0NiwhN1FmYc1/aMvi4hya4oj7AnA
TLCp7vU4geswdh+13pjogEmkKFrUv71UotjFAi8pAdWEo29+AOyapIapCO6aZl9k
/h2zSi43OqQ2HGUWsLETT3r0OYIzZ6ZUq9RqQpv6tBeL90WKg8GeyrWAOgIXzXgf
Xxir1zP6/b7zftRjzzS9kyTfOQ6uRd7ETvkoXSvCSqq7i0RTvlOqTi/4wy4WbtIo
Zay7m1VPJm8ceArmRdt40QRpcYXDsfkzSLF0pnCJGvdDayDlXhd7k+s5zZlBTMXT
Urw5Z708UNtGK8z0Kw/M2xouEmdcVDo3xzNQA/YvD4Phw5uuz3n88HOM23AdBGRv
Tb3UL1E/W5Gz0u+J6dwLkJnrYmQ62mJNTNQo0xD1360Jwd4GzonHDqo2BUYr7yKN
QWIyAr2wE+ObyCu63toguT8rBD4vpv/Y0EX452amTb8GswzQu9yBbNWny1Xrhx47
5Dm7DhqvKqnTkqkqFsjbFvG7Kl1VAow1MPf+cN79CfgyMjTIl0UXniBUKA0XgFA/
akiSuEgQCT88tcGrZaHyU7NrERqRAbOwOYvjluBAE1AQki0Ms1+6n+/ypA69tCbc
zc/ZiR7/m+u1TtE78AEHEkB1G68ZhJ5KDe+moJF0ETgBnRgtv6qE7hvYBedcLdt8
vRgkamAAQGuYGm6Au9LUSkdK4Mn+z4DiyB+RV4GFhwmpvMuPJ8FLZ9L2prSIEt9X
ktsaYNQ/MTtzyvXO2sSJlHSeP1yZS55Cz9naxvCTsRDha7NX6OZcgnsWfMyG4lkH
toRp6FH1rGZNx/dgLihVhN67AKVGJsfiQqkIY99JGhofgYd5qkjSg6BF1B3M2cTy
djIJmY/vrF7kwSdT6+0euVt4ryYBRkDWDFqL+yUaedNuiYtpI15iyBbAybx6m62Z
UtSlZluYUff+N3uDnTY9D0Afjo06sT/UqMHPkUpADA0vh6UPZ97Cpxk0xU3/dmHq
2XqOPqj6iBxlr9dyldT68fg+qizlN3XkXxIbIia6nZneWWUyKkYmOUDHNmExSAnO
GBYAIudQ+qb3bsfgu84eHgnq2HwqEnCOsgCzuyv0AXi3DP5jPfjDBpkTZSbYfASI
hzeL5HK5RMmpLZPGlo3/LAdUeFG+MnnWxj5MGavwHdajRk9HEB3zRKQT9U9Io4Xi
cxHCr8qJOIkKGFBNq8h1YRdB2ozmN2NQe4Kl/vC7PF7JxDsxv9QhvuaXmMwvSHpx
aJm4DSgwpUXVaW8toobsDJ+c4sMX8Sb6T7nVKpBJ91e06bG+/aCqXdyYZGZS2JrK
j5nyIhuu9NVzQKzgJuZYJkpDFuV+POWmln+5l7bgp+rWzHPKhHgo9V4YXzQON3n/
WotHuLXR1B789KHe+kGVcYjGhwb6yf5jM3ZV2wlQRT/DCkzTyo5gRiNmA+M1KKVF
O5fivguSIv8JUuHHGF6IE8sieqvtFi8jG+Yriwwq0dXJgQFMwLBeF25OZax7j9el
Q6bTpgVx2y7X9tfgFiXTmLLhg6C4n/t6yAMFqZ8Zsv2H4MoNuP2bWG4TtxyYkmsd
uCYk8xw9ONf6gXPeM1O/tcHvyGKS+3C9aZDmAyd5Fqqz3xXmo/Go17tkzfARFz5B
ME6J/59H9/Vkb6gCv7UJrnK330f/aA/SciWhVL33lcHblNaIUKN/xs0CjsLcHUCB
9tRnOvVCaHI/O6mYIRP/yLxsEYtTFAkeXQ6BRwW977HcQ1fgdLO+wOYu7fexOEdY
4iXrOaNsCHeFgAfYlZcAzVeTHNzm+P4qb1jaGi2lngY6MTuiYxUACyGoxj6QEvDt
hnReMVXdYA+/CstSVFd6VvsfrYG6h2qLv8nS8IGpkDyEfR4QYete4GXIWSVku/WG
1zblzth7yafmDCye8/Ko8RylVhh7OSaJrBWohM0U7gI3VuPqTffwC0xyHPdqH/Dt
WHKmYZ0z9rZ8hb2Z8QxhykuXFAYA0FukBpuhf6KWk7g/PRXWXYuDnPiKuJs8+sXP
y6cIs3EACIndsjwgdzCi909VDr5bvpWnHTWwL+/m0lePmHWltIXP/EnkeDwBPBaA
fnI30hVYyUoZTxrhpAIg/uG/Rj8X3sJQS9Jg6zzRn7dGFtpA1UCKVy7PCuiRyfKf
k3321A2TRnWG0GqsrBE3JWYOPfVXHkg4KI4oGokoiE0hsmHyLqr3FQH+2begZSJa
yL1qZxzCvVJ4FBHZU8f2PNwqBvDaTO4+WveIj7K/IIchlc4u9xt0XOMKz13xC+VY
gt77DfRv39Aa+iFv2W6xRpmXBoYOkYriNyAG/9zTM7a6mkuKLnYDjG+i9Aqy/mm2
6M8JpDTj5F52vqcOsseMB2ibgnxCRKZYR/xiR9g+XVJxDIPXp0u6GUcXG8hDdu37
OplbfdLaEOFGDlOiEAA3KbU/kLGfiVRJwZU5YHpdCZ2/qKzjdygeWrJvTU14LTfh
86Z0Z0pqJNwPNyQGr8sC0kWxxCjD+fHVlWOq1YGW3+QzcK/kWfMSpSmQ188lGLSO
aPUfeVH+c7lXR22ewYsHyV6jd8SwgyftB5Otf39QLTgni6B/Y89QPJd9vvIpzpZM
2sMHB4kg6cQRRf+VIafBlKKvlVSVX1tXhkcW6IEXRnd87+rd7jLp/FYQQn467ugo
8VO1ON5ysp6NT4tOz5eyoiNpv84QigoiaC8ri3PHxxhwUDZHnMvydzoYXjCCG8Lr
vLloGXeYL7x9nr1Y5sZM8MDoxDqxxCUBIu5qfvSrJllfiBoT7Y42qrtWzMroBnje
o6xsyzNdHFCfC4BudO8sbNqhqUVQZmxOrZpnNgdTyuNjcq/Iz8Pl8oG54tpsNeqb
LgYWd2GeuulIgUpxJixERj708nLd+0qmwvYlnCb44j8LpTOSiynEwkZEhiinVXR/
PLaE7OiJpK/iKJNbm9q15gNwh7KpsCfXvUhxepu4y6QgRWIVt+b1Eyfiu8Ebc3TS
GuHeifVDJA9Ues/bsr++opxw0l9DFLFliwQT6kK1l9ktLue4kh6Z3q2WZcOBYoJr
xlO5M3Dn9iccnvr2myg8VOl/XRxWRvwyBF/aIAxllnWnqdHSH+qhPNNvpgZrom8r
3P1lZ9SZyR8R8NxFPgLS6UKgFGGKeTKvQkjuVHJljM6aBwRNe1aqgTGRSXA5/BmC
d7xQQ2jZgYZFMrA9x5XcAqIrBffXXr0PQwGYUaQQTf7kj6mPU+Cf/RWC28VzFqst
ptjBC6jJ0bFuM4P/fiZ3fp+L36OwV84Tg6PDrOXB1CGN52rstcDSgQc4Jhrr7Bq5
zfvDU4E3vmeiYJAzeRYwweMQs9g4o/3b8hKIZiHxkxRfI0y5Rx56vm3i5p2f+pfk
3H69QSE56fooV3KYpaBeIOwycljgzpiqGXLU/+r2GalFyg+308pQO04aomj2kthw
J5fB+7yVGAlWis8YEqTRSGgl34f995bulPY7Mqz+zLwtkLNPpM7veVdoUXbf8ibr
cgxZSVGZsMO/Hx29T32Wkb82rr50Jn3d/4F84AZOceRzCkDU2bWEDv46C3g5POEk
KuTckdQPoU89qYPQn3J1lx0wGMVJVekHzo2DMFCnTBFccx7WrWYLG/HUDFQ8Dc5E
bl/EY1PX5F1FKJI/nZKJaX1KJAn/C0lE0NG1KXJk1vBixE0BI1ioPyr3MdPdZ6/z
T7IdPSmRi9G6cqOzNtA7d/1YJeTns3a7vpibkcoz9fwvdApncnHrUTodvtA22tNu
IvjufGMSNxagZRAYYxd0nXWoy7sQL6DgrDZeUnxL1v21d8sFYqMuUjgc1nTorGH+
gA7CHYnKpatQIHfeUjhlSmjtYR/nJOhp7lyX66ygKaHkloKHUBhOGLIaUClKdlny
Szo47EgqKJAY4l84GTg9fVov6DORnv1/GGjgBlgz+M0uyzsasPdFpU9AVrTI85ui
wxO+XCMjS5YCVD6irobGaM0oxxWotwQt+qh4YCCjF2T0dfAbUlR5chz1pVhfgHUF
e6aKCSKIghkQuOd0KghUI7nlD1wgodk8yG/2JRrwWGb2ftjlvVvO4kfuYLvfUvG7
q1Q0f+O4Uqf/+eXXHUjo6N+Ycd5Rk/XVPNX4bR4px8dpLi4jrscVSILMq1HpJy2e
IN5EbpBonOju5BPbuqq2JcFu4TVY5V4N1wCK57eLHMImlyX3ZpRzMZqusSANndv3
2nFc3TRUoccHztRlY6Ap8AhWIQSv+Zbh2w4dWdLMp6JWLLIN0A4f0q03G3/s9iWC
zBoiPzWzCNS8VhOqcugtFm5dvjhqgW9HA8FhinrwkDc1FU1RP00ZfR2Hcc4h6ctE
9B34DC+3DRelOAtArL3YPNZ3tXpJDMjGJygyMQVzoSz1N3Npt2UuCI47kGG+8Dyw
3iCnNvrqn/rr0ex/KpJNa9Av9ddSSQiI3S3zSF/McxP61FCrLwDxJF/ErSdb/JNH
vQG3O4otIMgOSiexowciNuJjTqwbDISJMD7fHIkgest1xkF+6l79iWCr+JWPV1xR
w/nPiMick7uTJrDiHojiClc2+qBmD/ScxriY4499kGBpEtUs3PZJNwtvsgyARhcN
5Kuo9mTlv9dSVl89c2unPwERFWdDA5RJueSbrfMPFJl6AHfScEZIHTlDZWNklaxP
qh/qRAIqkhF1GIId1p2xZG/YG8m79zqHBaTlvb6hiNifX3Fkw4wCYtYY8t8UiNfV
5us9AMTntzWDVQugqOabmv/3bzCaJTNuph9Ap4eiZdXWRyB8S7BK4qHGKmbqMrmL
P/Q0qgJ5tuNyKOZL/ossgWzI8gotidx/vNtGijz7mSgR5uux4qJllhTRVPZCVdu7
utMOn1qbfvegF+P2Fm0bERThucq/zhop180o+RN2pDbpKxSpEDoN8lT2REHn7vRu
KvBSb4VC/ahWfK9Sfjn1xPRDDv3o3Mw/ozKzClBe11tDJ5/0e2eikLOKphdTNMPB
12aB+kVmGXR9xpdC+onsrBX6ngqVyhQsHyS1TJAVcsfkBxOudH8DLTQyDS12shyS
SOUMeKqw/y8qJd/sSXjzxmeN+bf32k8lTu5b1Ec2ZYSB9YC1SNtZk49BZm0EeS+k
KVNZgAg45fUXznEnGBk39voqS7RurqJVs5WGfH0tMpfcOVpO/wUJ1c1/DQY+3LNG
JfYhuE+ED9vI+tceRLw3XxSzEeqoJG70o65HgiC1fYfcYrI3U7UTnhpWELL81YfT
FRzb2APQBr/Gyn17dtLhbPCO9+2wQXCB7208bjO2zia+TI1H4RumEhIcF8czPqfv
CGWmWRKIyliiS4Nj/KknmRgPIuMXO42Q+G6fufb2RrE/1NMG9PQ9uckPb1L12dH9
lBhmofLF+8SN2XdeAmZSx+yyoOY+GHHEyJLtm630UtC0Rd6KYE2im/EvMYBg76Pq
+JlEko/5MSDVgm8H66GQq9RH3k3Yj8eUPCB1GxvPZG/plHAS5HZ+zmiXsckfRI43
ZFMc3tkaSEwCLQALAssj749QSMX5HwUFoqk6HrMjJ+S3vev1YhyBlv7kEGKyQK+g
c5h2difFFLDHVpgz98BJ8vxKF67B0tOgc//W68MfcdNOkvEqzF97879vIVkDFSla
D4Bu+HzWFhMsBMtU38LsCIW61SzFSF6c4JRtLMCKg6/Ojk8/yDxQ4MjbOVdfy0RM
4988+VtMw3JAHcQkI1lWCTL5Pyff4U/C2HYfQal/3xtQokjlBY6e7wZK0BOfmzNG
3mh+FLq8J88scXII2QerTS+/4ishF4g8ERayZIQsRzBV6QNxhD9xijYLpQHpOFnX
UqQT8mTWIeax0Arj36s8YXkvBbnOsUjMVZZ9/YuFQfaMSsNOULr6EElFA8Fbidon
Nc41ZP2FJzRF4WbqTGEoqmVU3haYdOwJiSCI8smwlCbctigwCiWXQpv06fCye3fa
iiKqJDgOYwlUZ90QKKURYlGck2a2LCqUr44T7LOs8HUyL3oCcQPDRTzficHFKAdq
0Bu9B7n7u6dKLvdqOR/3IYxyk7xCTifTCNWjftQ5BeWi5sZ/cAt0ec9MsfhgjQkv
PdEYVVMpVASlbuws6HqsWqyUYYyzduJaXiX0rwo0sf0+uyruSGM1gjyQto5J//R5
Dn83gtEdK32pclgyDhMoOmWE36OSTI6pWg1g9oQRtwpRQYK4yFMf1Hva+mNarcQi
5E+AReddtzpNFpTUOEijhid5QSA9m4CIBESP89bUAwYoKUpz5N4EMaBcWsYyJkz3
3lVo5sQTkHTeVWjXNHMlyedpi4p5kNjiUOqkcQ1GMthnb+6nYL3yRvXwtkOwDzg2
sIaPGAZO29U1PD4OjzvezaOp4WtDoGB5nx49qCbWPZG1EaVfv1peLjXjFQfS3MJg
cFf5yA1wqv3cFGaTwtxghnk3ttim3BTk2zogzKhMNf3BUnZvOmycPXwaysbWoE/5
2OV5Kgn03CaYUr7+QGuN424g9Q3N9QyUo8vVzN1ig1Z5yvP/VXtpFrL1eXrFl9R0
O88ciiodcc0qteGybbJG5KFtQtULaIp7ZOm7n6llCZD8swmoZdgca9SIMYUZcq+V
0cuEL17uT7gFCTtGBAqTHFk+aVTPgpcLLJsu3rIgOgga84Atp1Aacji5U83LS9dY
ewv0wNNrcgQ0BvRL4GMn37V2yA5NsebdUskoM5TkGT5fQyJfu0LLuZPbeAzRF4Ng
63kihLKAbtHJ6AFdw8cPqYrChfYbGr0y8BnadS7U3E0mOFIuwJ14wVCOHx9G+HwU
qz9VR94alwa3P5X2GcytflylhlD0OxQ2DUkiK1ncAdiQKxSKXLIKYr6S2zqYMONt
vJ601/ekTs5G1u0KSIG6JBhDsMW2/BWza+OVWqSYFOIteKCdUshTSt2Z1VCxnF+7
V8Jb/Na8s+0J1awJXKp/IfF3tQLy+OhorHDD4UDKU8P/z6I8IQbDJpTH5PzOsYeL
mIgOssOYgQdqN4ggLQAc/bF9qlZOF0v0mftW2Xqz8QKHEgYWrE3cUWpiupsOwQNR
045nnj5NyaMIk4rrEfJmFdSrEd98Fx1Z2ZM5gIpB526KjgmokvRbJ/9/vMy3gTPB
VYO9sgRIwxZScHRBePs5EmQAhxIKsySYH7/rGcnZe5r8Yjh7+e//61U/eB0yXMgt
+zjs/cKLeexv+KnGDiQZqs/WXSvUl1ruFbDTFRpG+3Uv1sVpuO4BzfsreB2ZlniW
Ld0c/ow/YzfMA51A7RdZkQ6Yac3sU/tfQsMfZaylpgNWOp4j9NZ090MSMf68FASE
7pwFgcD9RpUzl2M0M748AG9AnIxe1yegZSz++ZRTwW2vCKWg4yb849P4its2IckG
xlGYZDHBCN1Dv2v2l0nXB1zTN63ZtKbTX+ta5FI4eQU02UCdmWJ0UF7dhprb24ed
rgAIc9qAgbeaHbv3ODQBSL6KfOAddvo6N6nhEsu4Trm1WCfkNX0PRN9yNVYS5MM5
u7XwWRMeOHYcFjrV1Sw6d/kQmIMF9QUR7Q0LLhpqsLfCzaZaQ1zVsFI1ewTktPjq
cKWNGP5oB1Q/KslILUxlGbu6eIXw8Xf9IhS5rKT/k5pP9lYLUNwwr5ryPwJ8J6hO
bxfPqi85FKkU4mXyRkwTcmJ8cKGWU2dNb81BDGQTAslaT+1D7cBp8SErclvsKVy3
73nZQhRUfnwvxbwxCdE/YF/jk+I+o01IwdmZxXLilHiMDcpk58sclvoIPao7Deoh
yDKla2JcQjU/SEu6KObxY0ZU5cmTg6U4ZCVDJs2082WnTs55KKAW1oB7TBwHtsdb
zBun9NgPAfTGbFBw7mwQv03F2d3EadIUVVo6L1XWo31j0Kn/39SP+edTu9XJFitK
dvEHPo5YDnxzdsNCfYcO9Tvwv/HkcH7n+nUleZWc41lK3bu74JD3PuE063+KjZia
BxtUkyeWAd2jdu6+UAg5vzHgTox4cJ/Ivrivj5yvnW8C0EELcsYbrRK707NQjGEI
pfXJ6RBjNtmg/CeEQquz97tIiAGYdqEHo83lXyX/BqxYofkXPCSn6kTinrzbuB4d
77ElNeG8WhDlOkpy5z20mLIw/l7opFbyuhSDko3P1g0SDvXEFll+M7ZaeONgE84H
sM/MRtOZ9WhsETtenU2tl8fG8FWRiav5ba25ys0vvkdZWS3lpL1ncKynAGEN9EBJ
3LvH5f49Sgs8SJHJtcyO9O8uHKBlsYWejlxKSXcCUN0Bw5gpI4rPtXesc2yhHgCl
MgBfzxRC4y3yLrzXzdMh0pPZAFMfAITmdWUKBJr6p+i+DrSuDY/Kn9vNbnhOSzDZ
VXKg4ldXnjlxYwzVJKHg4YxuePVywhtGU9gBfFMxUJ7EqJSqb9dVSweBPYx5MlvP
JADZLYUIsjnCQ1UxD/IFusOHGMWw2hdmIiS3wTL7ptEKCI0DMgahVwuFUDf5bqH8
VpM0vu9y1kyMJAWjizQda9Rhx83/5wPdEIMGr9N92tk/sGoAJYZi9m5iPrGfSMts
Y8FseO3ZoUAA9SEaiM9wOJLbbKHULKCVbBCG+XTqrzmMFfsKNRqUpw88fiL7LH4T
0i8I9r2i7siHGCnFzfrPOhuk7I5fuWkt6AHTq1nI1K4iY8IbS5yWhociCszt3x6H
qWCSqxoAxHzHIk9XQBPKw76s9rQtyYPJV4jfDuW/Yg2bQyxZjFik2yxXr6l26EPB
mAx2eRwv1wsCTjIgmSUbv7XuEGZ7LQKxJ4oEqMvE26myAYJVT/+6mX//cZwTxiVd
No7lnDbp06vIODSGL0XpdEvULbvPMNIR3T3lAUwQFc/qoSZm2TqJIYpgdeipi/1Q
7RqmkY3yk4NjuwfKkXBSPe6YuJvrpTZKAU1/M7iwC73RV34D6U3aOSc/UKbyMLgh
KoIvPh/AYMRhhgqOyNlhHuEXb+gddRE1Nwbhvw3iGSQz+2IN+4+yaPCdwM1P1CrH
L4D4jSics9R9huXDlcm/C1cx9oxpdWCfV99khk2Gw6Iz4nGtqb9Yu+XdrZb5Y1EK
W3jZRHbZnF7EPHCmaIQ2xMH+KrjnmglzV55I1waTmX/RgT9Nj/kaqsEafqOIUP0X
eUpKLqOzmtDihPaucxiupRPfj+v/fqWFWrBDX8/GjT6SR77H8HNJdXAybwrn8wlx
L5VsoGa//wDqLHuw3ew0roUKlghlLvQ2abortBG5OwW0nUcgGwC1QLoEV+UHkTRy
BDMOTcNLfXXUih3zPIIZTgS2KfCnWR1qMtKr/GEBUgA8lzjggGCj/XT0zmijnSRu
0WazAuy7RSGWqw8tU1zBIsvpywN3ghpclxAQFoznclGIJ3KaJK1p+N23ParYJ8S8
3mS5AaP7+jfv4iavng4e4en67Br2MSgE48UZTxvCzF7yfyIy/Fm5uHIMRHEnazWb
+CuUGS1LfR895oxQ+sl2OhtzuuXvwAslM0zuxOrjAMTG7JU137QSxfg4lXrOPXI1
JHlJeUSbDAPMRfnTeFEYQTGgybMFS0nSCDjy4CjY+VLLaTUL6R97PZagzDEBwcq7
MDGWVg4UNYxur37Qi/A25JfEE5BdFP5bGnm6/B4+VEiKemRuwxXKDZEgddm7uOgr
oJRUG7byRDmKuylY7Fm/F4KJqru9cF0bzi0swXg4Ke7i392k87FmJPAOBMlpMojG
Xib/DSi8Ixocwn4jytR3DWsh2Lm3XtmWVslZ0ZBshdDUDSlb6GaK5D4s3B7g+net
pHF/6YzEpdwm+uJGo5tNuN1akiJgphpeyOc7TfDDoBkCiyFAl/63YY4X19bP3jj7
dKl6A59GevdtunweakOyOOAiRm7wlilYgy63Co/opsVV0zxwTlFYKJfui48y7NCG
tATbhwiEKtpJWk4XIof/wdpi5DPXznheXhUerjyuPrx5Ts6BuHW/ne6jiuebwqPu
Yg1AgH8p514J6mstBXXdvhSTpOuHvpig5MJ3O/EJklHQxPV0P5I3DWtX58DuI4pi
jZQ0zlBK8ai7W0OHQFX9QzpypAik17esxMHagI6c1XMBYcBoVZ82nVsuRg2J8gzV
GBVxSymriC60zgL2/j/tPToEii51WSpfJTcKHEKvU1NV8PrwoWOFzZvekQIH+BW/
qPAvHHIctsaUExpXvv+ihM/ZOXs0n78OTNEIBYNPJSVFRVW8PkL7CubkVCPb1BbN
HhlvSryXqBFsCd3pc4upt00zM5T+DYEKMvBUnQnQQXdLjThAy7P9Hhwc8IzN4pSw
1IJiJA1PqGuLSR08Mu5FhUtIopzHM5VOv+eWAO9iBPphwyr62KLfp/h5Si9+ke1g
tyc9iFp0isYEXLlaLk6Z5rxG4ifVAUHXWsqCSgfKT5rPnTy5WfnaKDIWKYfNCxck
Ugq5Wk5iO550zmfQBadx3hNCXbVPUspAK+tFwOiUw/jQvI2oUStRvaci5MlSoxK4
RFSLE3snOtVbtE/lfMr/4GXuCVR+nFD2iYTJ7FlzhJfV0syLDbF60OUcwnYT+GNo
6oJKVsp6rnKp2+ehATCXRyOV9CWQbHvBksQMQ4pSeMMCKMkS4Y8TsZv02Qk6TJre
KJ1OaiyS0hBpV/+Jt7K2Fvgdqho8hZ6UmfcXUc88+z/vuNUsAk5gWVj2n+yBI4TQ
2jXCcVnIXeWVlTTtZm2tm0uqd91GRHLvnfAJj5Yy0v5lUbqLu1rlDn5meDs743oj
YWMfMXmoxzlxQt21GacA0xEkJ1johMh6wXDTpju8dYiwu9Na/5t6BnsqMiapG6pN
4SehxUs/1l2GqI4wJvHz3HyO1t+MYx7PgvQNAV7G9/SYhVPteLsLqR0RZr+kSNKj
zNbmblveu7VhExHeIYk23edBSkb3U88DdnRedbWxjSw07TefT7SKf/O97FSmwRnW
p+F+elAOet0dKDztPRTrjrgwKmtCHwp7Ic/1Wsp9uCqkfbzO52Xb476LZA/UuHfX
zNa4foO9KDzNVkCRweAmjIYTjt62LoYje2oVBt1HKtUuVzdBGAO6kC+j4UPcTfN6
89Ekbl72o9531hikwqhqNvVnAv7sU/Se+xC5H5bfcbVYWzJ9a0JVHLJxUFtA8JQT
7w3wNpoUuSaXgfI8qmamKaMcjdIMaUoWr0U2WUwksCwnSVP3mKT6vbE8n25zSIjQ
AkhH4fuHPk3N81eJk2tld+eK9XCPcrfWYDWzYGcqaHshMA1E6nq+54v/Woi+8lt1
jysNCHT8iG8MgqauuvJv07jIETmNtqjBz6/C/q47UEupBKWCgZ6cm/1JfU9pdy1e
uCTljo4wCXniAmIcQ1p3wofysYto3t10E2Y7U/+51g3leNGo1CPmC4DLqp3WpB0+
PZADxodVC3yJhnV3QiGOg9jwyTmt5hROcsEvA/7w4ee9Luocau5ifYZtfC2Dveq0
IrvfQZXFvh19tqDprWC80ZrqzhRBXP6iOvo8bNbBNBUeVb/8H7PKatTXgmtp5w3d
tpJX3KlCX3D9Gfwdgxrp5wVzgIn2sIuZB+YQWbvZnxiqcgv3EjLHoXEg5QogwP4l
nMYl+0iD44Ei+Cpy/cKeJtL8zmzqYq0LcUYzrPWW56HNASqwgI+SPuBal3rQpYwM
dxfKD3Yl78m3N610gHBgb3MPYlNj/8larm/wZR/L5A3RJ/v4yDfTq36uAWZ9G1OH
c3GOIqlhG3p8s4tzELFDlSOZAVSlFkGrB4e5ejWXqdUnLpBk9BCMzxxocZv8BrK0
5jBzNCNSDb5WB9lujbzNeoJeF+eH5/x2nNupUQgHUN/EOXrWswtu4SoL5qbQr5WX
DSjC31UC8ilPSu5RtbRvxPMnqEt5cl+9jAXzQoqfxBjvnen8rSQRNw6BuF/qu/QL
CMWARQy6RKG0IEQXi1+BAcAXUDpt6xPWRVf0zOLywdezTbNqmvywKCYx2HnUMI0D
oz6ZKky6c/Drmvco+E/mOTLBL6Neyikc9UFpIf3hn2DdvJvqKw9grGzXu1hFGM9E
q6U3Qm2qYqosf0e0OrnX8U5/wQdOHfbwIwl+5JuRN+oviPzcuGnOtgv9JhhmKRFn
JRBvUkBx8Ll7T1cgDfzD1T1W+xQo0C+MrPzy3jW2P7P9CydvQCR5revlStWyZe7z
3LQXfRE0PKZk7EWw/6vClRmQoTP4siFz6U1rDjpLmwHb3Jlp9/1FhqiAz7x0njnr
rGSVOHVCtEhIbZ8kYJG6Lgj7S9fmr/Kfpz+CXfuVfVV/NDKwGyANiIfEYmc0p81s
42b8tMQNcilP7Y/lDx15aUMaonMkkY+udk1lFSJw1VYqh5Tsddp5ecaV1LmTgohj
oGUAp+hEyNsa/S8jMJiMKbvurRqAYST/gFuGPcdrwgosMPsbcIC3gu6+saoIfOXn
fgqyEidp4Eps9fwN13Z70/H9LMMK82v/9LQuRSZ82j0PdN1jZKG0j/V4B5S/PeSg
ubdRnHTZR7aQT++63dKbWj8CPfX5Xksy4aPtO2QxtYGuwj3L0r768lM7Noqy6XAZ
a8HdkJc+6u1U9M57cd6uq4wdCzBNeMfuTxSP9zJKYv27E95PlHClDZVBRfnl6aQx
HKK1cmYZ1KOLDvUxRgaUZaoY5s0nZ3iyzeTgppSowXNHKLfizxDjMrxsDtduYXAS
FsXGPE7nHsoMMTxRYlrGyrBbv5SOfTY9X1QyRQAgXDsMgYGFLMIkBtqioQK8A5jP
Rl5se0+ur77yUmW1tzh7C6HLfcsRk0UNba6rfbQ9T3fZwo687MO6mXOySBRVNn2H
xxEHupAlOILkkQvs0eNLydbNfGEgWFR/2d+OX3smgE/aFgiicn/QQnYyupglDbaL
E2ARVofYDkI6O6ixsNwZ7kJOyrkYH5TItMAu1qBCTa+DTotzXJGHq3gcTjdv/EId
6UPKTAi5I8ixYwVo6CUFQjcnJ9Zp384GgO7Ji7rYFnnzOPToXe2uzlqbE/acLaLP
QUCUiK8exDjZL7AGgB7CzlDRMQ21454iwnKH1VMpU4R1+sy+V7N67NPb9dyW26Yj
vXP1yyyvqSC+zXfzr56Zl6nvq3mtt2m3ctZRDea7vd1SWUOg59shMZYtD8sa7S1D
hRmcqrQVOdH/ZziOI3pMBnjZXoD+OSjqJyxHtNaKqlDMjSRiHMj79PKkTIRlpFbH
gwDyfAkbqeQj4A2c8omEkll956nsNAT+JubIs3BcELHLgP1VQYoNQoHNPqDOQhVY
KXe6Ji17/VdcUXE/Gl6jPMaD7wfHQSGojR31JZrL1cA+cme3Ym2v31Ir+33tNcYO
sj+P+nHuCn4S5HgrXn4D/IuH7VOkazT2ejcfIGjVPJBTy5WglTsnk1hHw5Lc27U1
lNRr+OGzFCw0SQHLuh4qAGtCexHOo0Ypg7FLL9x1kgaFOp6nldbRRpD/BImOP9mb
kTXWUlrrcpP8vIIyLAaFzGvAIdeRAtSr/Bb0kYBOZEiVDvTPquD7OtIpLK03SW4Y
nlLxw7GoISfbEcsN/+cZXBukzHZ6Ubkqsy8njdxYJU02/Cq8PwGpr9O73WH6tSDp
NVinAekBvwiUb03qD+yWo1DpCX+QznG76KyKlcfrqOSqDPsX0TzTLOylpSeKRGG0
raD7aLAclRr70PFaTtbA+ZTIVUjNkl9hGMs/otsPG1wT+bO8n3YbhY0S/D0410a5
fYNIdjkIqb6RfL70WhkcpPthwTtPACd9MUloDrfCnT72QXRgu9l1mo8SAcvScP9H
VXhKoOyn3A3AKGGZ7tZ1penNLPXPkF39PFJ4F5nJkvK5udWNXnfPHzj7JAI7OgQW
7cZomrJ/6JigoARHb4cvTzPy5+o9l+EksxVaU7DBveZej7OVGMKdds4RiUko3VKw
04NGHcxPvHeShEL4N7+viK/ehvxzcj9BXWkArCjHZvzX83fhrtRPhh2d8AdFAEqo
Ym88I6oGqpydWueTs9KvcmRVlMOLVFBUd7jAGc29OrGXlGkZ2bRpK3655NwkKTiK
oxxT971iK+P3ExcnTyiiAbv93mHcTDY3VBNZo/Fy/FGHwhH1jf20NUgUNrG+cx9f
mVPr7JH8YsHk/JQCTaoqLoBedqGxJ7upBBTyj0LRAl/JqQIayrhrlIJCL+Fgt2kc
/VVcQu/F3THRe9oXlxR6haIr0USNeiKqsmQoP3U3Y7AUhmYDX9WfVEa5oTLC71t/
A1rYscrnEbXEjNhdDVz1BjF0vbVCaqtLSLvsb0SUfUl0J98O59i9ecHAF7ACAB7l
U+uc7kGKZPmabwToahnElQB7pOAw9WWQTc0y5gwnnMd61fXsvMssNo5DM2GscY7N
xrjiIXB0K7pSXiCrtqBH3D0BljUOvWk/PKtawhdBgKs2X4cs4r/CgGxWUUCIscZm
BLH3oD7gaqy4TQxjESSlUY0HFlZaLrPt0+Pufm9tRQJKRka8cmScGdcANZD1YjSi
nFJZ/6a8/yQes9BucpIjVGSPO9U6wBGYNdLGIvA7BL5jcLFbv5WUyxKQ1q5yKfsC
oRGoHuXWl8gCJJd+Y06/t2joHgcbtX6GFN+wigJiPQe7kVS04EJxd3i7jUWKnv1Z
Y0IiaVYOEMv8pY7Fm/pnBxGxwAMu7jXBuFYsEEuWISSwx8+hRpn3aACdhwpq62sv
zJl+zXpOgBacLhrPL3gjqkDA681s0Ie6qE+XOs83pmGAWdYb6+j1K7YB11/DT2MV
vmSf/TuJ4xz1CqCF1PN6U9gKYnz7mkPDGO85lXdogKe1NDgH0ABxGkdvpYopYVxP
TzGJj/AZ12T4lhlsOZa1Ku64e2yDUptC4JyLBAtkeKAYPp+yUx1O7Kk1POI6LIDW
Ya/fS30dD0bsp9atgCETUsXq1FjL5Lwd/V/uaUtFdDmc0gNeTCsIH+a5U36CYn5+
InNsMVq244DBPVm/Xtel7C0LcIq0mZhpME19sFaY6k+jb1/PX5H0xN+ZItjg/QPd
Afhyv4S6zY/jrO1AxsR8UZXX1KeFmcfbaaw39cYO2N5+lF1M+4df97zhKzOnR/Z5
LDGGWghvzNd4H1ZhkieF+26MRJZnJeE9N3wRT+1gWhMSgRB/dxQbEY2HQn0FOZIi
WBVPKRTTnj0JlIanfUmbIiOHWqeJX/ICWZODJikK0uSSAZ8zj55bgDYiVd6Trv/V
r2wbO/MsZ1pBtGh0se7xr+vMbyA/o/L5n5khtPEgxinstFeP1EPsw9vnRij5bOtU
YV18SNhrhmwOae2UCxWJUITmFyxb+ZnQobWCFbF5ZyjO1H8S1cwGqnZEIcCJivne
haRbNTqB5+P+GyfaC1Q9BEHmRGyCumyJfJJgg/voxTwTaOysYDXGAsNcPw3JRyyj
GEyq+lJXnRPBpfIfYaDM40qzgOoCcSivj6Ba87XyKTtFe1o9ASxHw6msEePOZFFH
Re8imTJyOOOn/G7HK1cbMSEvudnj1DaasXknIHeeHdHfcaWyvLnmcAN1StE/v0FC
46DhUlVHLiWyaMHprwQOiw2qwUc5rVH9bS9/jlLMck+GRc3vAF000bHxEyMvZyHH
BzmY0T8OnCK9KQLP9HnhSZhm+Cum7gApCHgkt64QxpX0HbT9I7F9swBRLZyVJvu7
c7IX6jg2uW+pQCxv3WUbqUhCxH9kZNbk9MBgFRYKukq7z+1a645+wnZ3kv2chk3f
awiOUPYes1cGMs/XrGGWSeN5I0y8gLYsv+pbf3/Ceta0AElsCwqeioG7nBqqE0Rz
N0Htnhyj/2SZaeiz+dSy8gv3Q6YYBAAh1ofam/wCISRKhvIFOrL9sg4V/JgCyHvl
7r7DaxbvnzoA6ItYzEBiP1YjV6qvkm0cEm1U1VyT0xTXDfq8AD0xkDzT9wU8pqFv
mwruM0nUCatT/jlEQ2KZ9DdKejYf43utCQ6wsPsKTEVuPrKyfqHXQB/OaAzZItod
0bPy23jeQXF3pZrUsCp0z9b1eeFZRHUbQ6VWspkiLQ3fwr3+YRfm64DgOXrboqiD
wVsLG2vFtBzkhjemo35fKI+F+eeRUgJjTrI5Hx/3WDIlK6NKYo9J4D3RyetRCCT9
IZKlaW8F4TPvZ44Xs7/3g8vd9YTrPgjFRYTeDsqU7C5CgjXvTr1NOVVBiwGXUh8e
HCmyIxTt+ljckvCJwfvh0Azocy31ZztjXJ9TK8CGsukjIsqDQQE2Kq8SgSR5xiVa
qJOWKrImbOhLXjTYc4UQ3t5urirCYmE3BCSqrHjoZN8I7CC0RoIsmbF9/24DJaux
z1Sc2KcLmBKxcTkhH7l1DAlq96KQTWFUcR/4fFB8/D/P62eo28ngl21dBwagDGVb
oTowuWRn2pGbYZrXrktuzII2Smbj7Edr2KyrXhVgFZ0brfgQ0ItgFev7rQWMTi/k
wcSabNJTS9pmryrUBnup7VmpYY1+jmkY6sVHlM9AvqOj7K36S4tQiYKOVbIUW3ej
g93cUNPy/sv3PTO/nmZtp49n+CvAbcmfVnRxwjLnQySrIZnwsSEoWKFDMP5S/MRP
dVyPeucJ2szgJppfWCey52l7FHi1I0wn2uq4XhY93MpTawz7yP1+pTY3ZGuX6X9t
vZrMVvDEODtg1qVOGdyHBH8g2VJgOaJlPJL/PkvBvycdhTcH/bo0rB3aPL5cvKMm
Fq7LtqkqY0ISPV4oAkswkAOX9mPJkLz2FD2ecgtdGHmuX2sL4Kt5svBOkBuB10e0
P6RmpB76FEnTAX9P8k63BdHbRQsZyPYmChKsWc1veymJgkIq0YCaSkhNmnnTdHXC
WNxSIz8k0t6/pClaHKVsL8XaRMfnvi0S9ncZpQbvaI/aBUYN+8AvJ3RAJ03cF5Sg
qzj2DpCETiB+q7Kt5FyWCWxJJxxwXmGyetPP5Y0RZXG2yt6J8SAtKG3pgLfq6JGG
IWCpr1SYT9jJiceUbuEb0XBoF2EeIG+2iQm+XN98sSoxZY5GqM9hSoWzyZKyioyF
/9CcIx7ClXPU7ja4+TSfRdwYE9SBFWiwrlvqv3qeraepsDD/u5moxQ9MLXXlvOEu
tXqac7rxl+xDIe1ai9WJ2DbJOA1YXYnBgkBinfnYvOidfL0ZV6dKuo4QaNRiN+kn
zYC6AsG84nWfWjRALwC05uUh7KHKmrbFxq+F0qXl4UtYrsrIW7mXL3jQ0Odmt4C1
MGTSOalmNmMjqdWR/c8N2fhjaRhN6PUiRMXl7DfkZDckPapUKO2GR7dKIroFel02
3zkZhV/R1X+lD6fRm8tiScxdXPGxLRFxgI81eqa7+zx22lAnSHKi9Z+ZvNmD1Bxs
omWZw38HVEEJBjVqk7lw2QNcfsNqXsJ4qb5EsXOlWDGOCaBeGk4qUeIXX46jlR22
fe1zth8ho1SmfW5rJSeB4u1HJak+rermPLNsb5Xef7LhiWqXl6P008dDrP5OgjNS
Cs3sFb+GnrF6h+BWdU4CwxkxInybBeSnrUuDwdW2bPooyAIV++wLJASLYsrW1vr8
mULCyQc3W3dnHn1nNe29Vbqom1o3gC75cxygKBg4GJWV/l3lEx2Q4kQQlH/57n7j
j7TtFw2rdRlm5pOlCxhArgUCFwfkwkRfWpy4wWZXAt5r0Ayvd7ePB/Kfn5uMHtMu
zlIo1KG5SBPoqjqyCt/d2V5CGsSgdiTc/OdyTsDFbPEc1RAbKX0dB2qFbBBWPrl+
qtzoiGceM4zGtVGCWXAPpUdVuVZoLIUeQXep0K3v4AJM/Yu09t9H5cuHiH+YFU1l
zV9smgpf9F1MR2Q28fT9ippkTz+zhoXBhvks4B1YL+Mn7hvOkfUT3iK7nBwqpS7l
k8xzgzik6dPNLxOCLJtQz6b+fPF3eThWF2hCwLGUtkCx11+rfCQvalKaDVyJaZi7
C1LCPJIvsMEFWeHxYOCpQ9MAzp0WxQERXH/+X6ZcSHXzzvlnCYmFqrSxWK/1b6Ul
V8D9WqHPPFuOMHhSOecnxg30K+Dj1FZ0//h4PCed+rcRTKn/FQgLvI2XgYbT8vxE
UPW3TdTkRDFdVoStSCl5mdgakpdZDlKWhDzARJZEgVwhKCEcgpMbCWE1Esk2JcqI
JOnzTtJG8DuQZDyg7G1HMuoiTS7+g1KVziXdGLHLcm4FpJiIm+gU88rVBSXkcgxw
Guu41wQLqBVB5CfatYXKp12h0g4ZKs/aHIsLFan8W1mSaCI4JlaIbcqMULyVByv9
zsPZBvPWhLZ8m/ZN3erUcGd4S1L/FB5gtG1qEWtyAcwdZGlxRuOzP0PVo6OsJvjJ
NQ99VioGd5oVA4zbCY1ogSdxfHUrvl0Mx04MqcgdYV7GhF/v2zWCO9OfKj1kOKt3
04aAswdmKhWdWWkT+qMb7ocIDfiFELKtt8B82d4hrVTWKfsnpHvvehCQqj44pC2g
uRolLBEmGQm3TEv0OU1Jycmed5Zo5xV/k2bUq3PbH5waJy31z9UdYHgDRDlQpIXA
jj5awkGkfc2Y8jUpmu0NJpLAroJjX7Fo4PK1OQ/3JF1ZoKN6bCwsblkiYLFwpm7V
M0WY3UTSLeFHY251Z/wzektJy45xuA3lmlt/lXiPx/UCz6mLPMPAmR7krLsdh/qU
hv1tJ5SbmLBRo2ssn/IxUh2K1yUBCSE6vimVZJqFiYcjrX8IhcWGB0i9CLaj4WdE
YtyUf6dbRVf7HDKYZKW6YlCxcOeofFcKx98G1cd18l0ZXH5CIB3ZaHhf9dvgtF+R
UUkQ0RqgbXa/YcNelcFbN1SjiQb8V8cnx4hIQCUZWZwwfURelrY6qS/zORvm7Vaj
/WrBJGdZzO94DRrM5z6x4XDUCWo5yEPkfMve1oV7gg2OgjGwRp3nSvzSZohEH2ae
M1Fepzhd0c1w9VE+NtUMTG+8W1cqiM5n/8so+p0mYD2VYOzAdUKfX6Om0piNT3iT
+igsjh7EXAoC7SfEHB3C5d2tBDBE28qmZVvHb+oBTNnm5pG6bCiD5/sVfvdpNtvP
7n/IntZ6/byB2CurKrPJhgRgO3LdxsueAFFMDlq9g3si5ViE9pkLdz7c07VHPYgg
S5eW32i7udROXqEF+raDRGqYMfLJVgCDU8QHlLuStJTRHfbf3nIBRPFHo7w9XwFR
ItfIBYW1dPfgVx4b803enUYq80jcxMiOeIpyuI9Tv7WMJ3ns4AkS659y0Pl0DHk8
g4ex6qfAVCVE7D2tincHX+YyysXBoquy9xAnft6o30jl7jMuV0V9f+RmiIG2iRfJ
j2Zw7GKHHwD+0JBZeSPyXygeEc+VL4tWmgR+nuXR5UxOFa9b/3EJgJHfpxoxzf9Z
i5kcV8UTugwLRaqjyrx9il6Qyu0/zdjlKGbbSYXkP+VBK+ZyWBivFbKwPRwf+d/m
4LlXsPIWDqQhIG8VPU1B8os2jCpkp3kcUG6D+IQ4CN/j5PAhSWoAaILmz2sDR2Gc
Ps7dIVuWJJUb+C8WVR2WNTh1QQIN5YiNTjVdxpXDb7CLYAqbJR4P/9FYkERwic2+
Yic+LjqL6b+jBlXk0WcvZnmSMSS0RNU9MMBbCNica2IEbb3cow9MB23XZ2vE9Lck
5elhXtMN3sKmLwO2PcM/3IGgkduDU7b3YtMqkZV/9hLuu3PYr40jdOS6m+Tzw1AP
mOA2KcYOQcGRul6kbc8aPnE+r5+5foppBofnf9toEK8L1d0oMluap8vd4aDxyt77
RpV74x8FHbGsb4FVjYY4XEp/HyQoozNcowFZZs22RlQafSnJXs+mJBs9EAHGMnP1
97fLFlpwEYUIMIocn0IFaDJxh9HRIjQmAzPFBtokDk+qOGiHhITyNnmLqqoiG38X
hCoJjGAaHRAtZqlWwRwf29VLL1MlVI/sttpWZ0dk9/LQFDblKehlp0XKDg9Uh3Va
fmLyPGXpwo4QRfEvndkq1MQ18CNqYIfS6zWYvtps8knXWNGGOBLIGkeqmPlK8YEj
9BXPYMhMbgFP35OxrqfoDDiJZxHdAFBiZ7YdML7TF/2uxFxy5jPiYN5zsku9in7S
gHOSEV9JdfoLgL2KEpiPCaVyrXQXbWRV6azfDbWDzXaZE9wyLq7Si5Bxe3jVX5E2
7QPXSps3GSy613UTMNu9PoatSBW6RU0Ck5GQvwUB+Zb87uJXQIevv0ntYpvRj1QC
5RMTTW645zYKgGLa3sAG4MOtQfkiGhyBXKLQGXfpBYwn+UB+OpuOzhQYI22OoKsT
rDuGTzYhJHucDBEiTOxN7l8XBm5/0cUA2SJSdRporOoljvyocPl3pmYYEjShldjq
UsZPmNSJ/AXftZ3WFnouhPdTLGDytmJtIYyV72d4SraP9iqfRmXn0QGGaq5DS0ff
y7a76f9DBZzkf2XE92mCLT7TnCMYcWDS/hBQq/CrkFoK53Erc2aLNehHvhHy2pvA
dFjMwtplJLc6BRMvwf0ISx1stYNpe7lAdAvwVu1s8L/yjdNrpXVxNOhTInhev66C
GUx5r+m3pNPo9NLi028Yyjf0Dr45lzPwhFvMUfGJ3TddmRUwhr3mUMRzTIb77ZJM
UWIAFm1mURnVCcLnE3kF084y7dWY4FD3WqP/VOGy/Rn+T6XIyl8k6Ev+viVxxy9x
yAhKzGunXTnlGYYEG+y3v/bF4kQjyczCHZmmC7EDswOCp75QV5pn5vaLtn5lJBod
veuO7c+3mN36Vpg9SW9nTnqnwEJPaxZGhJYStqroCG2Y2wee+ysGvUMN/Zc16XhW
VCQRBDDiEL4LmrSe5aoyo5nRmCQCV2nsYnODl0ilLFTEpVgPs34v+rKEWqwz6A1J
QbBODRzJSQV5uA1tnDa2cm7foaW47fzf50c3UNF8aWPn/IxWzuMdCfGsPvqRHJCh
B4fiy3rPvlOKI4BVF0IAxfN/akkwZOtVujB4Y+W8lZdxa+AyvCJyWEvG4zrCXtiP
dOFBDyl7hm45IX1HTIHjFWUohA7lzcMdXpQEw7H5xgK/l73WZKtdFagYGvoapqHE
mvU/d/cpwKWNVY9UILjXoi1/j8Y60CsWiB4tyTY8jWQzKnyXut/AcvJtfKxyByCt
szBazbNtT7cpbp1xID6XtMHA/174igrP6LC9ykqjvBhFiX7PQOnDbC5cOE3nU1VB
ZdyyRjbHSZXnCMqC3J9c0cO73X04P6jejZ4+jVlY3YmaQlNk8BvAcP6GF0jJJV9Z
hor2f1bzlZz6oP/x6EFRZ0xiaiEPhyXmz6z0uZzy20e55yeU29J//CmB3N7s2wj/
nSmwfdYHG+481iJufzPIPnoYMfWecKn0mXhma9vn089JDdlNb0KTBv+J0awWbzdk
QflgDyOnxVS+8o5RlFItOZUX7wDsD7zqgUA4yVOjrvsAL4WB5rvERyffT8tGopTu
oV1NfFtlAZzEPmorIpQ2FykXcgzw7bkvpN1O56z2ilWfFg7dBnrbsLKh3yEYeg4w
HBfE+T3YIP32VavTTSPXCpghpEDcgLRPal8BpnOlyw9BCy48bOlPR0exKfW6IDNh
GXJUrLxfn+RvHQ29ozVrORh4QLFeAeF0w3fmVYmXRvQIuvTgXKGPGIdunBivW8Hz
seLMDhPN0tcOZYyrEPpSbgNhqvOiuoP/XoC8pjpjnDTLo50OoI/Eq++81XYrt6wj
d+V2cS8ppjNLOy13EYdM1fYdd7aO6u6GuiGhfpCatpY+KSENfnDZ7P6aTJYW+lOs
Egzc8RuxYkNpk9I0s3t4pp0OUGlVD6H7ISr3Tjb8hBSo70FYVWSSpLrNdR8LrSDQ
BGlPjMQiT4LNFz/qPkJXtQHwndrNVbb1lTyOqjS0WJJDAv6S7bHdDpHYNg5iektK
8rwTLdojIki771EjpR8S7sxAuE8BPX6kHk9qrmILQC+pdpKsumNSz8sHuwPcsv9j
MOEI6129pW8em+NLhsx8jhtygu3TBa/wj3roeT6wvHOwd0edl21y5sG3qyjeY8cB
nJCSjNl1kpUEikDjH9SLIQaD8V2F7YmZv5dqYuIGZhBUWwkE8PFq1alt46vtQwGB
79x+YtNc2qenPn199+0zY1FIswo4/109HMsZj2WNGoiGHapPOqxOilcRSjSh1rlU
kRAavtpWSdT4RPe8SuyxjidnOL/7Gic0EjiBmwdHZZ09QXdMytYqVBMtyYuxNM0/
oug0SIwaQO8o0NwilOlAQulO93+pRHC9yNXPbWU97RFIf7Eivs9M3MVE2YBXjBGc
kswHMXRaqFJ7Ix3FnFb5CBr3unFrJkqQPFhvC7gTyD+RSQnDhzoonqf6aIH0KFYa
o5GySVmlhRp8vH/WKrXDO6kQbvsA2pX31299tvV2ft/2ysWZaJW3Dlx2AgQIuA3o
1v5ZDxQ1vePCOum4AHDRbBHmeRP3sa2dRPOnXotlv1Br7HEbHx4dAVI1YuzDBrip
FQG4AR810hgMLPDq7RdWiiA8RwCuLuZxzjNAAc2MuINvAPB/crxqtBJJutoH2hYC
D6T4eAUsiZS7czDkHWPmoi/nvaRNKdPY6Qx7EHIU/UO6CSJexpQKiQC871cBmSk7
yHGt2BhrdlgG1GITJ3KA9vZePKwTUEfVnTyWfx1hARQNkE832WlC+kEzkOVcXSb6
tFPy+sVcYseQNMYLzAC0Ni0LcvgGsedfRl2v37koW8pSD1vL1oez3dg/vAYzTSLv
n+0PO/QtsPXFBgK8kGbvdqqgdrEK2D3VYIX42zzxm1Lvc42OBdGMZoHEAVq5zH52
06CDC5yMi4TVi9aL2VT3OqRDFyjNGuYjlKQjT/MmEqEvgbzD1JKlifsl3xHeGc/i
3SFfLZK8lWjGXX1gdhHJhoo6Sxy0e3BwYMgQ2IB/DhfDY/3YsBRaU5ksqjJp4dja
d4hIHgipMX2VHf95dTAzq+QH1Ub3wexVR0U7ltxyOs8fGWcyhoLIpPPbBc8v89xB
umpQ/8xgQ9bak8WlqlIxnUdlIKZY53gPPYNW+OXBy0ghGqZBnHL+vmHne9bBf5l5
ojRki2TmQkpdECxzrX73Ci8UP8yHkaJ/OsY/z3WuhpKN+uBP0mATLdFL+CMzNrTE
vQgBhthH5Vo0zTq+QrnvbIdQGPE03x3+WKhOXIhpvFbnomBdixzLazUTO7MAGjw9
19dIAvhdr8EVtfGyp++uJJ8R2bQ3l5J1HQWldrksox2D3o58+Ul6/OUJ4zeQspwF
8ZurPtJQeI4oONTabv//750qKJjsdZeLux5WGDbttbDynm/ZiRshWfhMVBvCRzAj
SprfyKabuwizIX9W4iadK3Isshnn6hJgDbCGrPsrtuIhw0BaOPCAYGxU5YeIB4JE
T+UgLMZJSyHNV5xX48wrTtsNja8iev255r1fYEmcB3RvmAIedh5LeuDRUBxRdpjE
tODD8UbsH9/7FZH4u9xJOQiDXzic+6FV+bdPY47DiUIJV6KH1hRr7zB0wWXnVTaE
viBEghvzQsh5OFU3ur0x/hsZE94k9gw1tNnS8xy+7QHjYQf9t+7gjmYiDKsA5+Ae
SKCVbfaG4evbwC/wCBx3RLSXcwLyXAPiorRscazt/AQtRQQvHTk12o4qi+VM1Bjz
0iWoe7YR/8bx0mKGwBSOWyA/IdhTxo9od7bW+jAwrB59BVVbxlZVSnwx0RuWbIKn
EB+apJF7SCPRK6tJ3o9HCM56yVnnrTsNU8VJ7FJ02HkKTwkQAJKpgxpor7Aaisg1
JhT2QTWflM7ALfLe3bOpFlp7ibMpGu5xNAkMcNcVXlaTTFGKNk6oMnVp1POJxs5z
kwm9mWzaRVdkqtrsLaxvzJj/fPZrIZwh8/DWMe6CpQ6gHPQqF0ApDDUwKJDSkEO5
abFfa4jtE0/bB3JYicQ69p03F0npcKrtqRT09wJZKZcz3jxmlDhxmtyQR2X1YYGp
UqyPJIe2uo+x7MFdOBe5lpXlkgZeFPYJVp+Za2NOFqlAhelA4GdVrGdV+lEh4y3S
9LtCw5TCFedOIyJVBEmGtmfJz9d0b2xm8+o+KYQNgJteox8KTMMYQhcaesIPYTEP
0F+YRGBjIRv4H4TmzeuEbsEGuBLeqjTwbRMiYSbn3XtYtmt1KAurgBkWT4uZnwTE
RqiaFcOHPEwULLk9i9wKZNMz8r3wsk4nLxy1P0FtZp0b401JKgD3tDwEEH7+9xV3
hWbn44tu5bxaq8jkAg/5HMsnFyTFwcWzNLORBQ2yQB0ELFu+WlXRvvCs531ja0Y/
zs9rjf5lMYAiqlqnygeYRdzNIzAd3ti4x1ExXwI/GUOkHsznJ7CGcz2X6R2Ds7y2
xMabo9OejkR+m+ZGAQQQS++z+8UieEsENJxTCyFCaKDHL11JKJqzIOwohK6kLcaF
LMQ4ZWkb3aGIQSMxDplOAtJkQjVL+jGgMS+YZQ+b4T0isbg8Q7ZiVikPACFBupR8
Uuq8Xii0LuqioV5tUbVHW3uOolhN0ZASmzTDzQaizuh8f8+gBbejlH0+CAoo1hCp
v002lanhiSvAeV7l/eLkZ9QalSextUv3mxK4TdvvkrHUbubT9MdQqHvSy0WGxsYF
aNnq2YBxKWUlYVg7250Yso8nGzOdkNPWFfcBL/Z4/wpa4I8tYwLCuHikphFmZj6D
GtX23zPmnWiTIl+Su+/Q8lxaSdHCIjYFLe8xxxgvWn4QGMb4RUhtK7UTbnK70Bmm
DsATfG52M6EjU6SXewNL/YU8plg0rRSGSBrgZvPFi+rdHI3OB3egXGUvwWZS3C/0
45R2fuSWSE4acBTM6FahHt9roySaTiekzun4APBPnCIeUKEwpIr+t34ipHWneEHB
4MCiBi3Qxlq6MAT2raDQ/iZEdoS/hNrd0NT+Z/a+RqKs3bYIWXM5qhb/jVv/LvnY
oHbdJebQw5gzdo8+cxeQ04zLyVAmcM6sRxbm2ABan4DGX1sVTeKT86VOQJ8anwKV
nUC12Kx+yONv4TvJ1bTeby1PoGlv8vIdni2NvOFmlOEbiYTy1Lz2J3Srw/c3f5DM
SGe5yXkoS9OSj6Be0nTncEhmEnK+q/MZskmzRZAt9GUq0JzCxVZ3bq9raFrQgNYx
EGSBn9LNFawnKYtRvaAwqeTM0kL+8sKLAhg90X8rg8inu+gEG2GJQynXsVKkrUyO
AtfN/mdtoDcNG+8h+dmO97mdQxG6mQO18GC6jGmyZkc6aWvyr+aiqQ5TjSFb6xvX
XNgdgaEmSRuCDQ/FBWPYWCGAZKUbuTopxwECdpOleRJsBPK2WahSdgd1F0esBuSC
w81m8Z5XD5ZxsnlaWKFqsG0va34gJO00G6scnvq0J4woHTbfd+muryd/Z7y9MVun
AFeZA6kzy3D4vgscaCBH6QipREF7l4uaoNgkDsPbraRnoMTF600PNLdQ5BpUR6NZ
ILu54vvS+5XCE/B/fwjXOZcY/KL/ehZBYVBrAvFx6UCNjykLSRyEVxcS2cZ54BlV
zIHHOh8WlJL0Fon7SildcjPpmWwCMm56IZ/ajfYcMfKhMyNZkM1kh1YyPt5XVOuo
iJ1rBXEusV0HjwXfkD2QCd0fViNFnjgRpGwYf2vue7lke8SKFBzh9zVs/FvV7ct1
fKO/AbMubgfuSZrrjO+PcVu1JOJUhO/iLWhFxFNQwRoZH5ktm1PK/oFeCs1H3g0Q
E+W/H+c2+n4FxtSqlyCYq+lVKScAy3g5Qx0kHFoyyTDuD9mXnzxNWj5cmRXdaDy5
Oktu7gTHaM7j99h3HqDckh0qT6rH3LYMDQa8gmGuO+FaUReZ4LWz3MJRUb6TFAEN
tzEv9wV4pDnz7BkBlQ2wOqyG6MLMuVEi+XrwbzRY+U4dJ82lVyrjc/nLwS0OGamy
T2kiY/uFRdKOsWk835vMgSXDDDRsJIJB809LqA1yTzJM2bCjDxuTBb8Gvpp7OVbi
Q/0q3BSwhK7zWtBZRw5rPxgyJajC80mSUHpDR2nRoxZbCqT2v7Sm96iBYj4C7T0F
PKiokxz11YRXPgJCbO8E1bBHBnZmpfd0SC9C2O7SII8=
`protect END_PROTECTED
