`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/nJxd4UuuOUBsZzLm3Em9m9GmNl0RouOw3PoVpUqmZ6+wbPtf18tkxZCv8k7S4rT
/s/mVhpJs+s+VtUlAW1DIQmKNR3gOXDnG3xdfGKoN3l64kEUGXi+TzlJoEzLRMDR
bMgLxpKqd5B3IZFqGYk+5IdKozw+P5oBOpqLQqg0gP9C2j4M27BRiGJGWMNvqWBI
/2Ogi6pQldkWrj0WRmoOfZfqy12vh3M4hMhGhEwUOJABV2ovK7c83iKlz2rBf4Rd
pUL7gernEr4vWWSrLqu9enkTZ/VE2UL6xsSHtDqMVIyOjxdRCamNI09i84JVgdMU
HCuM8h1Mw9ye8yHEPu5VkhuEtbEBGgIdIfOwuK6LuVg2UVklQhJytPT0ePczqwDV
3eyLbAlNWzf6Sy3UWoc7XyB8l506zZyNIy7l/jIgQ4oqy6j4H28OLpZhJuDwDWUt
+6qcfXXAA0UIVRTYWkvhXinzcDS38pfpBRwKYUjjhQk=
`protect END_PROTECTED
