`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K8AZqjtR62e/Qk2IvmyV7y4FLdyLRaOd5J9P6nOoKo9KMiUjQvLfgAIm/Qba1Gov
GelxVSQF9ZDmiYlvn/U1pU72lNND833AO7QvpN6wL8gaI790NIIMgmrpe/cKfJHu
dPxU2zEha/9dquKvSUty6n/bOrE61Lcd0D3QEbCcTHm6L0YhMth4wTSxduSb881A
maPoNTwo8OVF4TWVPAvLsVfcN740as8SemK8fJtqrAp8vj7cxJ8kACvFFlFnQs7C
0r1CufukrXfVRGsJPW4f6K/3kcmzO/LXltq/kAqaMSA7qlgitwe7Zn8QjorBt2Fn
jiSey+Q0A24Qnd3aNZIDK5ozLm3171gkJjTbxwCeTqey9TmW+/h0gV5QyASid5QQ
ana5wGgNH/Qr4+dhuvJShio/Fboko4QXl1Cv6DovixMleNGJIcQz5VFItDthGJ82
g1ybiEdWnNUU/9iGb7sB1tX2uXcI5/62lLWCkHhYz/gY4eTzvaEzIKQjYncRhx4Q
KA1L6KEQgFdEucrG3WcGJ3RrXPLHsAt0Zwzzm2p8UCqW9ZfscnVyHnuM4FE4WHEh
JNzeV9pvLdQHxhyzFOdFoh7D9Aw7eRMuwI4m3VrPxyaMfOrNjMbcJaBrycviBXnv
g03pKn/rEmRAHrftWO0F+w==
`protect END_PROTECTED
