`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lAYl8Q6IEX1X7F/ni7QwozIjhSduXwVH5zMnW6gkfmPjULOpii5TBc/MuCLhv8qO
OHQQmqcqVLIERo9kVz4tKxebtB38PofpLnNqjk07Pc7HGTDemuMHfBKp5MsiFDDF
0GH3iuvnPS3Dr9hv5P67R1vSKzgNHn5hgqbTapzIY71t14Cn5O+icokzpT8ENfA+
9abGif8Y0twov2oJh4v1rESdK8BMV8xbMym09ZQvJ6d2RFdkN0nDqHQee3ZHLTi0
YNztGNexmhZ90hj/EGvmD9igOWVV0oHjqx169H0ugW6Ck2jcNHllSzfJ/FuPzFbH
N7jHUQHg59FUWRFYrW3i1buga5OLQKCeCC9sikJ7CIBTNV0kHdScqtBaRr24g6av
dmnL2+q/qOxbe8zCQApCANd7pM+PuBlTzWyY/dwn+oh9B7tcmJcKZxTbuaYO7f/i
DHEIFbhI+VG6A0q8kaaZG5k2RyyX9R9fJe4hDJVAapRWTn54O+lMztbr816qxjs/
DMIlwNNbE+64ztMxXxSFn5WZtRzGjgF+TxgzMDeovNk=
`protect END_PROTECTED
