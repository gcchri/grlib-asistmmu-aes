`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5tzDwE4Mop+9+GXIgIXCUYj5jWUgTAQCg2OOUD0OwT6xANiGWGDRFMNfvXlIBhwN
Okl8M7+fGZf+qkl+AuPzWRgLlld1YbbrkVfiL35h/1U7eRF2f4UDio2ojIeo67N4
J6xatQRkITmIeaaIuiqRN480F/KKMIwHK4wtj9TT2UFjxcGBLXVzdLNX1Wcc0ly+
iyyKa9dS01NP7TsAKBl5jDpQbhp3NeVNO67Nf+6T9sjHZZ7OPPJDkXotGaDVMcVy
iOd3c3lKANLvpu9pXYkNYKtzFzwbUj+m/elmqQhW13aw14bDljuJ/sXpHffMIVQZ
my/TlauMr3gF+fTqzDjVc1Gz7rwFgDEeC0oCMMohmxQLibiQf3ZHunF+8JStYlYR
j+OxFjB8ejQxMYbQyrFn/2zWgCrdJFAYOMahhWofspCT478gAoaPr1iu8jXYXDir
`protect END_PROTECTED
