`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2cNz7YWbpcKfXhzEPM2gp7+iGkn7DCicFkfKCZMDHD4DD4CQL/VyFU3r2LVNJ6a6
ua/b9lJJZQYMOHEJEbRFs8YFC9P0Cazqz3VjKzZQp81Ix8YXcx4ZcYra6EMSudm2
NvVaf+rY4pfS43X+6h1DvdFHbPY6FNKZUKNNubVb7Nfi80y/laTrfdwABY6GgT5l
k670lAYKXO/CKV4y3xnW2EEV3gTt3qFCO6lqfVJPc8kwEBtDhj0nAE/drZ5pExZf
UFB/oa5UQV9kbIM4ZYcQ2p7HI671OYOZFe+frn4vru5F0kZbATmhBdnVuYGRQiwi
qhB62wOTyehnlE1hxYbi5aHELqiFdKSZnYL2MDQ6tgg=
`protect END_PROTECTED
