`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dJqfGYIey9UeV5Xyf8rvwhD//EdQyNoAI3ZvdK5Ca8hJvy5lUWRc49EIuw0r1A6Q
V7YgD9n57lq906QyL/5P4d5bKBx8MACBCARpIWkdslL1RDEXGybRx5jVJbqwCE8K
Xq6FfOMkmRwvuUflNqScU0fyY3HbUazaygBb5GWzn3Lm0y7v43qDwb8JyKkRd5UO
7+nF9uPZ1pCq/T88Rdgf8n7/Ry0XqC8XFvhYIo1mCgf2nbd+aAHKZIjZ7ZnuXwXt
0McX6uCUlNY2rc2Etg74LOV2Z2fc7+bq7bszi/rt26P+a1Rrb/7sWglGAyXFN2dv
9PjR9/ddY+Ty2ISwq16qRXcLrNapTjMu3Gwq5ackTt9T4w+rp70K7BtpFP0vRQ4A
Y+5DyzCmJ/J7JludV4+L3Kk/QDqykih5rjVjoUIjzutbYvoSlrDeMBc3oENMALEJ
4jw5ZwHOTZ6RBbEqE83VWeaJ/iaZtD9ng5QtcO0GAgpj6JCV9ZTE/5vRVmYlFFjs
s7xWBLP7+RL19vVpOwgImTiLlW2Y+ejD4NtDuFbY8NC+zT5B1KEwqRRtb04uyGhN
+vJNaxJ0o4OpxUgc4SNc//SP0iIz5iST+BmW2+C6rtv6sp6klCzVO5wj9FVYfTo3
tbL+y+SXH7DkdRC5Pzgb5kCY5E3l6K4aaLMV6B5bxI2+jhsbwJG2IMOVuRo/MhlW
qD+58SUZBhMrK3e/urQwtVpkjMjLsYQ2n/pcLsfCw4DiQJ2HXGawp34xs1boAA8j
D/nufYKM5DIG0kbix5sc5mbHc10wZp/WS5eIxGic/yiXjHH34IBhQQk5ONBJN16w
VzLtLGb+t9ByKJ7NESUMtu2YX1Rmbo1xQpiTLkZld7XKDSAh5PxduFcEhHKREtxA
oXkQh6DQlpT5EpQy9MbeviOMyJf7vnWcjA28OyvkZhlICDPMUtJHYorgL1JgsWil
Fkukq/KMXvpNd3rI55+52URJP7I6UrN1pF/WI7Lpi9w8Y5ZGnzFFXVEw6j3KfMJZ
FOtaC+6Z5NQuz8zcpt8BraGpRho8BYInH8SVAZU+n+8wga11hRtP0BkKHRsXQvut
f73u34x9wXp8ZGq+378Yp4zeNxs+gIg27wBmL7pkZjUFUPle6E0ktDDzocbhpSkA
UeJdEtdkcUXLQZWsUPrewxCGlgT2Y47JX/vgtSESJyDWmkMr0exOOubaH/78Wsxx
xfzzBN+ejKMOPUNarYVKoHawfVEfMIwnF6og3wsKbsCiYQPe82bhWRBYxrhPsKiO
0E0wLLQpRLTXDcD+uXz/Tk0xiM6lX9hk7KSNoc0vWRNc8E/4hpVb2K8nmas+JOHF
Zlb59tTwiTKVa+hJ59YHyZiMSMTqcn5zVoQyMEgwibuY+nYtNXiGl/uj922CyDVX
`protect END_PROTECTED
