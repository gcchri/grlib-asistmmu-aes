`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rm9YAmL1LS0pcxrCU5aux4ldOvOt258q9+emBcx/RtzXzoOPFKqcIQKI4zCjBTIB
T08ajQeC1084VG0Ktf8/7qYC5R/EkHZSw9dqTBDGxwcyKvaRxfyXZAM1z7iHUpdC
HmSjleDh6eSgm/pmAYgwA9sADB77PrxQJvLhz1UXt4l3ZmFyTFR3TztKq/R6OxvQ
R7D8zz82nb8lLUY6vYcDeBWe5r6Kq7ImVxgczpVBvdPHw4oK9uaz0lqZA1XGkrpF
6Niw2j7XtT1GIs75omWoIWCkL/+WV8vFBWESJfWE660445qRoEaRQvLsaEU3PS5P
DGmc7advaFP23HeJnU/lUzp4TJX3FueHXGEnmLMmM3iCxqI31q7bDQhSP04gXHCi
HTgYu+60gDiCQE6WDExwqNRGXzGcvuBDOcZITANBY/9QxDqXKcP006BIZVQmjBLV
8+6S5czSb04Ol+dFsOLcPxxfkE9pDPeAvfFWbIBdzH5W1Ez/fdCdxQdpE106I6Fl
V4tJBTvuY6x3tYe7EALaeRM1/RDBpPNUBHGI/CT5o+CcGDOA/+aG2jWdSr04111W
1I+0a5HUjJ7XbV42SmTD/07Mn62YXNTmH8CDbW70x2VbN21N7WustSRJl7BQOsTC
6udn75mEZjvo9OOwvBSRWeEPwwFToHtj6fZW0Ig/nYGfYAkhdPQWPw4Rin77K4/u
QRCQsnB2FY6Y5hgMucbUHmlgwzKLx9MkshTpvXJeG6uFeUxn8WZML9iGNI/Hef85
jIKNkI4AR/42ZROKwzK/nvAZp3JL8LPzvSRh/hQAu4Ywn4a5tEsDSUHXWh/5h3Fz
aq9Mq2oOezt6UKCg01kvN271bhMI2aLMgbjUahU+Jl29rRfWFB4d6kCYH5tzgFfM
Dyr6aU0E4yjX+/0kWbiZPWyhBEU+r9SwmVkGbF8X4HAqkRqibwFqSWThCXspQ+c9
IuxaWk/cpNm6M7CXhxsswK18QMcH8npwkwn9ZbRT6XoPgRxirgbumIKolpADHA4Z
AsA0/AEBmLQBB5kj7I9mUnZJbvFCR2poIJmSbW0G/qgLXvpn7eu2gvEfOkINQNgU
gMzBFr1oUly09+D2CwB1yG7oGq+wjThFoIJR8/xaN+k=
`protect END_PROTECTED
