`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0/TbxNDfpvhxrwJElVv3QVETnzbI8PJma5TiCl6H44+SXi8b7gXpLOKqMaDtDeI2
aU+bhKzef/3NOu5WopAHUd8YQodo27Oyw0fRKvODXv41BiUw75ks9TCNz0THHYcn
PmLoETxSOUGGJJFpJdipd34g43/LfHfOFI1L3prVw0HYo10w6zLEBh44f5SSXsdU
wRzewyn2w+Jk4feEAOu+8PpaQ6eZ4AwGcF6rNJ8VeI+FbGo92tSq8umWFO5in8nW
k/czvjFDTGBvp7IVEEze9uYZBQ1uAsiPmIIuaq5KTr/v7DbcoshT0kyVKRFUTtyq
wqlaPi5DXH0NtfeOYJnCfzljUEv2XiVzU6ZFNr4Exo1nwq3juHsRBIqboPYHFTiz
n2uA+0J7BNBWLunlLL66Wz+ZY5S013TDGLoFEV9zpS9x7/3Cj3y3OSb/uPBdFN1h
N509IZUtFMEP1UYfd2RePeKwmtWt4hKW5a8TPGIRiwgd7mgBqGMFzZlfVvWd5Ohc
`protect END_PROTECTED
