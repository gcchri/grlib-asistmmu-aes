`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xwR0BUrtoJHF3H27fRxAYPlgvG8OimbRQPEIyjbhd6vfVzPJZdawKh3YUbrmsiRW
OcZZFqKcXdAx9CK0I/HoHYCu4Zvk8eoAJu23wRWNLm0pyg5sVY9TMLXUsGiYr8CU
r2LOSM5MogGTpgooLZmtHcS3zOQHmxeaIRz+u1lrzDVzEKzBl+vTvL02LL2a2Ye3
ckF9pvjMyXGzMUyadGKiisPgkZqZiQmIKWBJ1ycNIYk89LUFElLrV7Lm6g9mnTkI
pVHbJ0YnqS2/LXaA1NQ75Q==
`protect END_PROTECTED
