`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w58tr0eZE6PYBULbmez5LH3oKtBy1oNXhj5BL7ykAT9NFZrsg2bNXnnWxkuFTxId
zmvwE8k8OXRVvbOyw8huNmb6zMyivZhAHIMLc5vevm6orP1FE35kwraljWPodAs6
PsTobx5+6aNiwMCOIAWVIHU8cxf64uO6ocm4nocZxDNS92j4P47pnt1ktYGWdtui
0bLI3aE8Ls5VbenSerLI+RwtYs9CH3LQ1bPGXvKKi4d24lKFyKRDj5qRlFl3m8QW
SA2Skcr0ulXCqOrqcJv3ks6bcjagimPGU5gVF++udtab03JtR8JG9F+1/Oy50SnU
ANfreoEOH2bNGPFt/5BfUfzaJQuv9VuEeWAcHw2aYtrwQn8hboyLmPYdBXxBEVog
LsuwU/fxa8TDq34Ez/AUcE0hr9he/Y0tK8QQ7Y+ynWBnQV8/d/yukv/IRzU0nw5i
6AaQkzi6Efv1KAt9Y/k3TyEnkN34WRch0Wfy0FU9oZXg5V74XjNrszj9JZTNX1UE
0b6XwGW3CUleFvzMpaChiuZedDl3BzPkJOd8F3mtC9JreyREXSg3ZgtL8DzUP/8n
qnfm4fyOEKRHLOGOnK/InZnuDNu5AxNBmWCctCqJ1PEPPWuF6uqy5WZOZ/du6SCG
sRCC+SHEYvIMji3/itoSjGa48jRtWyZPErChqu44hp4dWQPDfIYrLc40zOZY6W3z
/L2vHHdN+vehpvzJS1lNq5UAXYddo+tiBmM2a9gozIJK+HXntrQMU3xiyr6vJufi
cCD/rKaqR0errtF9BQCTlmxVETYsVLKRaHOCtk2qfBxZO18JIsccMGRb5qmXOYez
n4eyQrMmxeOGDjiTpHLEN0H4gGlYhJ5aYgQyT9sFLgQbucKdUh26Z+4b0l2SuH4E
C/Al80Go48X2ZMojV8eU6Q+XufHH0rN2VmVB7MLFZ2WtX1Y03W77bGON8PReqc3V
tDJlIzxvtzMTbtdXra49kYN3YCo0wZeButoEmzm/ptucsI7oW/ySbngcohyz53i4
SKB4wg/xtVof6B/n5uWBnDEoFU/bnZeEmpdyIFGLDNXBBcBSKrotrMqSOrzSNgkN
1PZxqT2QGiCFPlvjnSj+9Ff71yaU5bJJxWbpX6umodaLxy/r446euhxT5g7+1UG2
SsnY2Stc0zqtg4Mf4l//UFgsplv+SO9Y+Ly/0EiVCwNL+kRYYEoap4SYjHXtJ4Z+
APq61Qn7Iu4g6U6WAiAY7fNlXYu+e6LmvfBnSxPTpO/eJPm4O3l3+VX+qkfBFAsw
57BmOtjkQ6M7bJmeVTlFzwQCgYKtFpPbqUXgTSmzfNM=
`protect END_PROTECTED
