`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aR36vEsGBLU4SHLs3fpKm+BCi9ryphsz13VbL+G0GhgnHZT6WjKKroQfPCLMSqdd
GlwAgyvPNcI1cKqTsIqkkPT4YMMQnEnoucSq8USEf22Ig4mQaXrsEWY/6H7nhs4p
lKldbqHPG0x+W3My2qgUwjrGJnqbyg5p6AQ+KPnwo/uU/kF5fZpU0HRVFOg2yNER
dFSZz+sVQRDp02RNvBwgnwGK1cuE4h+nTqtWgXDqZANBQlTxUqv/SrCqdZRf702U
Y62ZQistx5XWFysQ3dGWFxhdXlC9u/rausmjkUn+xXFU5F9PlcSWp3TnvN2wQEOp
8r1Su5RXned4Z4VpGmK2cplwcG5ll8Sf/BiMxxmYNk7FqKxTK/+IuL33Y6ly/jMM
lCCfw+oAoVUN4TCpchZoAbHv2Eyvk5Gge7L1sjhXLKohid9+BG/4OKMXruFLxPSB
ix1Tjd3NCuMDBkwHU951z0YVT16Qpr2r/MHE94ktFNP9yOABu4WgdsAzycWLFl7K
qd1Eg6+C5mRyjOOyV2koYB4w66IrCfAX8PBJR4wjsIPOrga5sC2ilaGdZ/SRagcC
3C8OlyUTawpiA9g70GKVOkjHxmn+UbkLMS+NPH+x51+W9r7XRNAo4ubQKREyGutG
xY47dJXNodMObkmh30cr2yCG+b2AC8Uv6E3LrlXrYLLoXsKbTNPMli2lDpQ5kmoJ
tiAUDD1w/aJhZ/G71ntHBplB2zakiajaP9D0fk0NQty3aJJFbpLfJvcph7Sngf2u
3cotnzT532qvyRfUsSSZcHW1M37orCuPmrAB/jImAe36yz/ds59ezIAVweidPoKq
giLk2y87zTUbAWZN2mV8BmT86c61vVvZJ7J6oNZN9fIxC2jKHWgQCl3IM4+JDIRl
9amgfiF2pWnP+YJAaPoM7tgdYDzuz+CGXm5xLVj81eVjsz44tGvlqyQ5Bolw/ze5
URGhqFP++A5tGm8tUoenZegUfkBLkxpxoIllndbPQBF8C8g8GNLbBA1nF4JxRzbr
HLmCCTs5ZTkIucwWaUDPw1fPneAIQkZpBgJcTLrsaWqVm6lMCgH1GxD5tXIpkaIg
vzpBq8qqcRTlqe1IjjjhDtMZSq8GI80nr4xk9X3ya33cIxklqdELRrZJXBPzwJE2
Wkej8T86Bzs3fBriOzxrxxSlz8mYq95VBcCeYirnxWJJXK1z/yU9e+lhVticzOVk
+Aig/hM+26cjA3Lfwqmrmb/RyXots6Qq6AdIUwLpORh8Vj1q65Vr/UGzZzdy/KRm
FfySki+ZIjASaLptN7sjoVVeaqYbilOLzZ8vAwKjakOh/3WK7Hmw6TQcb0gNdyL/
bg+BdeOtpbkufxlaSj7iaX3FzmuIbYWbk4ZLEr1DIM7K2PU65dh7CYVt4PbfwGZE
0ybg2sB075voHRuXisngexS5vAPNjBr+Ji6/n7f9hr/sD8h3Sy3MoDWtecEOicE+
ecc34SRDSJKKZwXAETXnt6nme5h5xHP0zoNPox5lVm33j0yBmL4jsRhSJcgQz02Z
oqTzJL4/DSbRns0uQNo6AVqlhw0Wafbm9f4gZq3g2YhXZfAKZZf3ytTS/UJ7smbI
l2ZWaop+hRTKQnriF9I2qU4d+AJkO9jJGqximl9HkgyHmkbeIZHjfzJiTOCv2Adk
4wXDGXxNknAS0z9NsuBY84dqV/UYjblfr4o1s7iJ+YwKb4OCQrLV6dha8jmQVATP
+qM8wZR2cE+0/m6wvboOWg==
`protect END_PROTECTED
