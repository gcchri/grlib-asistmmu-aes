`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
twaTjO4X2IEbUl7ALFvLKbMI8LhSIFNMU5QqRGFjI5gdKJLL16NgKK5vyhz5Ia3u
264CZrX09QshQXO6BP/k/1TXgFRC19HTmFh237DLzxNKlLNsamJ3EibgUdJk7EEe
FkwfC6sYoYRoWK4uFIZ1qWf9GhJtIVQQq+ribelzpasafRqcBJDuJwTyfirR4rKN
C1Wp1PN9ooccN3U8+BVKlGIKOUn5UQKyc4o6xRHAHnV9NxiL2Q2QsNSgeLfvOfbA
6R4Ngn503oJbxjXv7g4O0JcYqZFrfBvWY5iV5ZTyHLixcIn23HsVK+v1/N5zZxwU
cbRudAR4HbjI2WnuCYKdFKHbd41fNh7kWPn1nWIedo6k5b2/d8PXS/jrAZd3vwGQ
D7umYnxxF6HEZP8lXyAQyFSdswiXu23qp5697llCPK2YVh8TjaJMQUtX+GNbHf7u
tInibXgNzX2zX6ROcKEjvzxtkBLTD9+Ki7ugDqSJ8CvIVMnwfFDYegi0F/SsrqRz
IvB2d9oiurbXFnA3ephp14g8CtznCJrmqCtKYRajYiufydGEMLxT6OeiBQk50NGj
Iry/zo3FSnCugI+jk84idUxKbZvBsHAOSV7BiKCfs5wF1IBc4dztVMaHGzt52MCD
kPBaKKwgKkiwiRJRDr+zag==
`protect END_PROTECTED
