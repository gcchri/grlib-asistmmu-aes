`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
33P6MFC1T3CuLajrjCXomTwqWx9urM1qS/LdTSLyzWVdHDUlbCP4zEx9g27LBClA
aeX+RTqtVYBpAVWFt4u50MUvewXokGm5yZT64+4g8rQAts8vYr/IRN673IeFBq6Q
8mjngzHj7S12U3Zx3TQyCg9hkjy9C8hHn2vtpySbFtx+bLqX2Apqgq4FiY9iRYMS
SeN7aVLmCRK7PkNg+ch7N31+NbCuMewUdmGpe3vd6+1NquRzpZJUbb2/2RQ0OgAv
E0dYpU4e9T8J0H3OPCJOoUEgSUVyOnUhSBRKymeDZxo181MI/TU3ttj1GZ4RctnD
LIJbGCAUQarkt2X4hHf0sVW4OMejr26VVyQ/KuFRX5zZX9UM0Hc+ASVSjICN5g/Y
X8X2aIGt7VxFxet1nByZvoWoUAv/pQnUQXH540fMEu8cVXbEnZPbMlMy9SQhL7SO
GQFFe1e+RhJEYS3j9GO8ynMsT7Q8OrwLRAGNJluXMyujgntAoC0jL8tL55E9i/m/
X6SnPj6NvVgK1RqjyAEu0SdCf51UorHuempcpTo2Iwug3PjTs6NSYYmNbs4WNY2P
hKNCJcPCnT29/65PJAXGoQi+f7PPf98+QNTotcw0h4xpXcPWMVIDWP5ZVBQXEoUl
XbLHDuX5GXJ6rYwlXuXLR0d/K1HsF7i9XfbCM9VgvsJ8uRYWtetdNI2DB+jvCyNp
JDCbYsVcKqku95Ei5MXoR15YWnzC1S5IyJUy3c/OK84BE7+3tWCK5uue8OkOD+86
kqmCdImv4BL3uL6wx7Yqte6CHI8doi7DATCdL0J+6lHNzMjpwXEugfNKB9VKGFTy
NL3nOAhbFSu7G7DWimWBG2K3AUFsf6tzdJ2fvd9+tyRU5EJPT5JYnn8jON4vAd9a
ZWHNzcWcAn9SDooB+3dwZF7gOGVj8tyog/LaPbavRjTRtNO8HyuHouii0yWVER2S
XMCT3M8EyCUftb9vQ4IZm98pAS1PKkquS+T16MS7CrGZ9qlwAFCn5QkKwSQyLGtS
jm1eYcz5Z/S/5/U3omt7eNRrEOm4q6qG+byNBBzdy8XsWgUtRysiKFxJH5k+LX7l
yCbVuE1MFnjCWf7mU/lMSa8ciWDS7DvHMi5jqvXYhbxIvdvDqA1xaRWuHNcfNIrX
9JPPIgIe55ksokJ2HyUz6KGcp4FuVR5KJ++NT9kSsssap53qN5wJcuLdrajmTDsw
xdEMtgcS+2UmEJITzyZMQxd1K/ZtPrsektPb4EegABkvI+IVVPwidfCkHxieEFZP
/3TuMPmfnx/qtLQRv1CwxO90Yuw0CrJhanpJcMyqwzvicmKdM5pZQcd69B98E+IB
mzgiFJiOgUZprXmFjqsG4xCfwFjOoHh1OQ4azQaK8VKjUL5MQLd3kc17VEwuhW/h
1cVZkBNdacRjAQf75FSiQdlQwgrSqkXElySd732VcizXz2+e303KL3hS7J5WzB4A
g05UIhcNrexQFx6f6XnKPKsek5Trz5ArRSp44A0UpNXQSqgXvINyW9MpEYbF/vQS
phWdwGqcdt9R5uLU3+gW+dlffewkGhjbrNnR+glBNs+YaLFJ8A1iNRyN/UQdI/bb
tEpsJ3t96XniZ6X2EBtltaP+NImrSG7z5q0CVyLCoYhxU3xqAELoWX3KTKPKT82B
qtUE0lzA+b9uL8/JW/7LRPv2kO6TCrE/Uy42mm0qjY8raNQBArDoD9wBTmW55P3E
wqc2chaEkfwBUi6nzyXlnAoPn9ipwRRpi3Gm0+xx+e00Ko/1E59byXRjGS2QBm0X
j5ACDXPdV26bdDd26t8NIz6mvU0hBXHva04gYhUgNsTYNWMYPUN68JWsgOIWFaTZ
a8ShWogJVbaWy8NdHieYu51PFWB/Mj4sOSrmHPx8KdMsidR4GX/eqHDIhPXUTPd0
iiSxUl0XZ8W1biMcQ8XcATPgM4yfqItbhjj5NpmzNudlhmC9042NMkV/QmQfjBiL
96LuP887pgSbKLnRsZRVb2DLWpTV6ieuVgXvrDLX19Wk8NLhqWoaEIQr1CRN7Wwy
H0m7EyN3uyN4fO7L43dqqesw6uqZBoBZvxYauA5FQAdS20m20WP2gX/3YW7ZEOX6
IbqaW/uxjPI9j17Ts7Xc6ZvGxFrx3RBtE38Dwjja3EuytFQ6pBRcHrZuajQhXDsd
g9bkSbf0YuhdNVNUnkcDn59grVpLhzXrg7a9/gLVheW17WwbROap3+OPbpt58h+m
MWcfJIRNANFYaerqdYbm5eDknEpKoBLa0bC/6dWFdIA9hth6jK9T6OlnFErrGeSM
l6G8eKzdLCNjrUUDzA07casrx5RQja+VTSUiTUDAXcT+AAPFJMjoyhFnZ4LHNkmZ
uEfv8KwRg43iI7nJ4Ma1++kFFIPsbd9ZeONF9xn1XgkN7vARFpiMTD4iExQXdEbT
jwKXsFfijWi83zrOkxLKRlxj4fusA4IHfWhJpQknPijos1jPuZbROViQByEkV2A+
fGHDKq5si+KPfV+dCMwfc7JZ+aS/sazoWnSqVwxoSRv0fBfugld4fu6PbMBdBtxA
FvHuxQMyYjGaQQPZaUsFM3O71+nhJc7kVZSZ/A2KJEzab6UPvyfjn2NBWE4VAjfg
VprFXJHw5hzum8e/vHnNuEgc6vZwe2yBSkhcZNkxeuBOdYNLt8xy/GyveGtzHfFV
kaiJf3ZaOBxuqPe3etrR0hICeOzscsXDlkpc1lttEkK1DNFgR9EbQiABz5zt13ro
g4TloCl5J8BBsdqgrrGhp7SFbw/mAkOnutVzHkMafl2mGhndK9qnemkYSq5jUFRI
qsb4qSmuu8PSw1m8xFWOywC35d7wP3puxzeQTsAbZl4q16u8BJ+yBKIgZzH70N9v
JAdSBLg3Sa7BsIbxQKA4fPicgIYuZ3oMM7xwFdHbm6H6zBuW1GZ+Xr5NM/8mh+hN
pOkgd/Q/zykUpFgXd+IO/U2uGvR3w3u2ppRiGQR7KPztddRb+oMytr3zNkV6j4oq
MqfMuZ6w3jYwTTqfj4zAyEE4esScFNZPkFa5o8RYCBh4Amx2WWtb5ZUBgRc2N3G5
fXgyT6pfbo+LDtdNUNm9N5K6I/unRi94FcD8hBderj9LE5NAdOSdvKIVb+a1Z6qH
BLGyQclQ8g5KaRY7RiF1ZTIqXGgUTVqeBRdboK6BtFEFmVMqJhD/dU2tNadWz+8q
vZG28xqrMXNZLCJJ/86hTjj7C9inIApmwozLc3E2RE/9priZ1ncWrNgAqeb8XsfI
cLr1oGQRStGpl26nTjAd3bmg9d6ZLvyJ4e0s0+pucf1PgvItbVPePyq1yEZ6T2BL
CulJ8zRAOiVtBYxSlNbv5WV2hArmtIHByA0QKW3TYFZTS98iQ+3yyBCUSf7DEzp9
sFbq7RcWQCM4SnXzPIOi76+BMUZtNseHmh1FcKp7k5K+vHpBY+XGGg/sXVdrbrs7
6JhlUYjTdVOFK7naEZlERB2Xvq9EOS2hFqxtNzrio4PykvI/y+hU4+zxUFTdC5qV
gvyiHQ/e6J9w/gHI/SfB+LtM8/u/z9IJk3XjJkTu9JyfjCrf2ZiP6dMoHKcIbdOl
osPtKEPauir4F+V9lTxLn2TVaar92U6CRoJBK/yJT+mlHU6/3vSVXDMd7G+dNr+T
XBA1W5QJtjWWpLiZ2rJFHadHyyNeGNq7FkRThPu9GMhhvqYAEYZoR0zMQG+RslrL
ZvrPE32wN/Vke1EIfqrGuWXGMntK/BB4kLgIGvjin3fbkR31XXL7Gy4x/hcXIUd+
wAM3TkIHl2HqWCMoRNOMh1JDJCk90ehwo7v9uTgeLAOtC6JpBn1tppgsOPbtNf8O
oVjv4bEtTJ29paeVlQmGmzcUPAsFkyRUauzjqSnJZhHlT4F/BDzluuK+AfMd0DnO
VBo9V2LWVURxjn5eaosOBx1vNZCdGty42rFpNjAMpRcfr6YBlgK9rrEjZv2VPOU7
SM7ccgZhWEEaq24sAJgwdrvNt94At2CwMjZBW6xyEYsm5CMN/2+BLRREVbZ5M8EP
DRA/iVRxlPF2CK81F3X4M7lsUvHd1Kzpr/Ku9+7Uhyf6fUYghMVFHA2yx6n8j6mQ
AvNDZe28Vh1FlXnzMzmuHYPw/h3L0SmvkJhKpsgSfqzdCmQ6PZnV9Bw6TTr+cHWw
UwWab8ECA0hUInoHEy/mu0cO2MPKfgl3CTwxlTCoo4hrWquf47uRDBMeJoypGGjn
7I2q7tAXa+B6/oyLzKYGbY6saHsdo5J9Z3XpSjVy77D7g9ClBJ3y/8zI7NQZjO0s
u/dzZMGDWUJp8yhkk30brViHkQrralScIEOtShAdpO+wxaudwEwuDznoB1MRwVZC
nIL08AxeozqOT4s4LN5ZbmbNi1aOVdrFUOZdbH4hbxqGIU7UGugoH4e0HbYHClmc
EDnKSb7BrvXbvE5CDpcwhISrQusaaxsKyA/bgeI8gexHbk3BX+4Ul3OJOXAbJ/X3
4K1WfoHpS7OeejCDNzbu81bBEt37kfWzdOAlbvpd3P33AgfM59ft31KjUwC1WVR8
I8LY6yZWhOnB4pxIcnK6eGV6d7GUfQFsKGIR79Iu3nxpnzyTRmHRJhVQSaN6gEL7
3hPx81YFIaNlt7+JltHWAgcvbdNLtakCgAhD92bCT453HtP1dTj393oFpVjkM/Fl
qYBGYR+bUouI1QuVyN5MKRgoqy1KISRC2Amr5n1fXEyRhm7JFsKERf2aKk29/zO4
miAm9tecplUZerB5dVwn/KcRrOUUNhVTDHUKYu+G9xWN6kl8nuvHyM+P3aJ6/Z7k
FPw6soVsVGJ3Qzr0mMoNDWwJOQI0m0caEBjAuwfwiLOWasKW+8fdJacJgsQ6VrPw
oboTb5vXaIsEd0KD8FceD2zqQqnhetFLqYD3F4OO4sS5gqbHVMPLLO18N9+Oapjb
lkmeBcJQ+adkHhonqDQYQH48lIl44VNIfU5z8MEgqfNEQsHcPxQkwi57jlMtFdVv
ozimPXLT4zEM7nhXt4Fosm1uXVUg5s6aQ5TUMVVENAlNXF/p0PuBuS0zA4FTwUCi
fp2uSFNLfM0T02NUGRSgiyTGe1jBRBaozFlxKIH2Z+T/JgC/XLz/Qp0lKFOoAwH5
hGf49QYRa2tD+q34KtBkCHlPYhXP8CxZwFwBUBIBnFzIn6SYHrWr8QUOrV5jXsZz
M1HAsyYLiYZbYxrZGZF3fOii8WY/ZSEC8rg6PU5dMtRn3g0RsDrZ8kE755O/tx5d
b5Vi/uf83OOW9ZSMGqyTZYifNFkr04XutxiEsmRCQwW+Zavrm5UhXenSyB6msyFQ
q2eL8O0a8oYsbujTWuvkQhn5iMzEAxr6Icuo0Vtb+jvSn3riqzz5wSUOvfGb+hUa
1Ixdo62lm0WmsQ+qntv0d3FZoCgXK70P20qIp0/0SBd8cJDJ6gAVA9LzOuDZgGcX
3e/KQIJYorNNc5kXFgrx4NV5H5UCltp0oXZnPqCHteKo5d/2ePu8hIY+SSLu5G06
YB0JLvNMx5RlSdZpLre/n7WTqqGE317olu8VQrO+ypCE4Afe5wtLpgDf20YLbm5a
Po5eJTERLd9UCz0WSNzBnrAUB8P0vVgLEwJPAN+tkM0Hsq2Hh5LSu/7A33WFeC4H
9nMctRHi2OV6W/gKSKPpmJ6UgFc7M4zsaPu/hJOMyZHoCo6kh4ulAFCNJtsQAM2x
FqC4eK4tExSXfyM9VHfUbYOPknvathG4KlEw+tdJqjaFhqX0pZCCcm+9Zn2jPrTh
R6ZVybAHIlK1RoKFbBUohIHQjyYQujwa5hOQA7ID56Eg33yP56qdi8KKgRtbsb9I
7HT7qrjDvvnkAVnmkkOXFtPi8U5vlS0z1Bq831a/iCKM03jNOuD80WHZ8u30z1LY
2J43rsf+l3JNgKU2oP4kcyS82XzVjO8TIU6EPA6ewqpfBjNo4Cy5Ax28cONDYTyJ
6lu/6KC3FrgJIMV9UJEKt1Tb7GsjsJ8q4rRykLzo14Zb7zmJs70WGDwn68gTljAX
`protect END_PROTECTED
