`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dYN3Yjf+Bj+C8kzm+q8o5p6EPSdKI5urZ0gGUPc5r9244eBLrsFl2G/UApvEY5Yi
L1unnOKg5hsY1y1v5yDT2OVp7a5xlNRUBwCMjLYsYJajZfAdeRAWVpSmGAFokaVt
49QdYOBwKgAx5qDTKZS84dO8BAbuNP98zqksyIGqWasXbEJUlSWKIng8IrXKv8OY
56ObGqh3C2Ub7jdXdARYqmdgTmKalYHeeDfMExEJcmDlYNPld4l67ngADyNHIrzv
I8LXTjo3A/QQmvF8XWKVRZzUBS4mZLgrOL0JX0hkkVmq+rebemv2Vz7bCADN9t4C
NrQtc5J2SJGVu6+K3pU44Q==
`protect END_PROTECTED
