`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
icBr6b/5grx9BjoDweSCCgQ43SBgkJupdHglgFDVdiI/8Oxoqw/pT2Ci89+WGcOx
Aq2BTpAWBKc0A/6AP26vJronvsV54EDRYk7AZNFEC0ZV1VxhyVgUCyhRPL6NVymG
wA5X3sammB4mWkjHnr943T4pCcIUsGJvmKDps03Mc5ptd1HEnUtRm1FoNdeG+AiX
NP4PCppw7xh/ugGvOEadfQTyG5kqBSlZngkiYkx7IlvwCrq8+kvD7QBAb9eoNeeQ
QS3+lpNS609jvbfaF4Xlvu8xTDD4D7qF7eLIk8cMUyxiWQaahhouplRxX6DfGYcx
kxqe9usoakhaISmoJdtcrAAfwBh5/iJlvRjS7bD4jUbeyFG6oSR5OADu/QjJihj5
8+m5lVashx0Gzugymy9b8IqGHeekjbtsrZCEewHicGfkoja/trBQcJVnBgdgwBLA
TAHViYlVHx+RSe1/vtJGJIibpZxfAI9J5fZ+C0VVHs5ukr6+q8ZpjTqvh1UJXtBZ
zp8McNYrYSgUiTT+Z3F98g==
`protect END_PROTECTED
