`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5y+T6lmi20DQiK9pxhD57D7m1lkpULAJQJcxizHwaoCeLwi79BKvB1vnA8T5B9Vm
O5J7U5Dt2nfoN1i69WQNpWpoDBgsYADPzugaL0QruxTXK580ofj+peuXwoyQrBdD
iXUXEM4ZV6i1fYM0DQHmxjBrHq3V3c/CsN6VURzdS/xHSU/uW3zV/gXI6P1mAA7M
8RtJ4YwTQKULMoD2y9h7Wj0G6+SRRm43tuDU5hLO0no/vky6DQbRNsR/pMXqFQ7q
b3+Ngok7gKu6Se/fE6tmwfo8Dm9CIRlwaYP8T/a+4hj6zzqz0CSqrjPJkLg36k7a
62tHEiGiKL4gGaBVLmU+4AXj5pysb0dUduk+UZY5HWVcVFrTajftdyCfmI87jUBQ
5NKVJp6VDg0d3wqFy8jMreCCqI1VlU3u0mBekzxwGB1RJsrkLz2NN+O72L2DQn7z
xXAIv7cdo5rMzq/F36VKLuOt7GKx/XscVgVUtNMhWaHEZc8rA6zCfQTRfgfatOyE
0+iR+nToYhKSWX75zkPJfJlrOecZqC4ofaXSr70zU+blBj/SKacPDVk+8Yi0SOHk
BTv4ssGL8u8wS9x6LGPBni0PfXI/y4SQIJXfOAp21lmpyx67rNLeldjbuoodd6Pw
C7LJVTg61KgJihMbjgw8Bb1z5i9CWeIb9cy2s07LFXkLBkTa7EUiqxyo8kQufklA
GiBFy4sgZBQkX7xr0LG5h17+nWp7uTMA4Zfb7RQDi+k/uKTONF7wXc3SqzcMm3sw
R2XQ/UN4C3gG659oKUTiU/cFwv8JHOvgI7LvADFpVWU6OnapWZ8MyCDTi1vBoQbj
qeCduamcOqLO1gHpVPUYlh8FSPXuYxjMxcrWUCM8iZ4hL1oF2oOrHiP2cTuFOTaQ
3d5BvOpHyygjcpVq7fdZNRmmGUA9CRdVOH6kCLQtw5wVC9zQ8AOtJ4Tz5KGjSbRE
4NJPK5SWuNVLcvvoQ3mVtg==
`protect END_PROTECTED
