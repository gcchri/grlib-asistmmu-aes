`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sHYJFI9cVRKIIyyjmTNf3naBW44RZzRZFQ1o8yOludHyKmbEhhVSWvXT8DUHKrYp
Rhz16qpdALyam9HD5D4AqdUsb5xP/WRqercNtBnsnfnCI7M+hqSjVe7OLg4vAdHW
tyZN+faexZlpAl7hERnJlYgtkzzvcZuA0u0nQSuZ/tmTOG8hM5L8oy/BNbnXOfzx
Ag6ePWV8M5bFwl7RuGRuffWzjDhfGEErxjaoBYSVDTTRyYm69EfLAP0Bk3u4wxN1
91oNuH4y2eqBIeWjzHoXWMky/huzO4ehLWatNDpm41Jr1yexVHUeNSEm+izh9uW0
7YQxCcZf5I7sB/sf9AiSREK6Y+ctb8Ml0/piHKxvpAwXwStzgErtBCfie45J0Fq2
HOSBAiqGrKFXwF0KMWQgNU9JrpvahsVH4lqmXOqF5MA=
`protect END_PROTECTED
