`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JAVy32vgGvIX+8oplHTSYoLALR7vHf25RUzFnWuaIT9y8SUxwIFmw34kc/57Bmk0
Hc/YyFxkpfuBaP21m9iA27encxqGkbtWAbq0GMHWLZw1+0tjhCLAMsEDTUwk50C+
7iZW7mQN5cmCYJxqAj9iB7uFQ6OsbXlKLxWuozOuJcTEiSVGxBVFRaK3kcWS00uh
PcszbsfjHgD9WfA1ywM1uxsDAtI5PfnT1fcyULnRstABlQxYY0e+GaJV8ORF1xnA
i8mEt6x9KzvahKclbJGQQ+t/F7Ld0g87Sayo2Cx2aEiY0j+BY/nACGe2grfNyZh2
JAAarj6eYcc+Avb32rR/bg==
`protect END_PROTECTED
