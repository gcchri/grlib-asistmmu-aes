`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
67CKyKGt2bZkN1S85DbyjmZIh4x8FZlOFwQ/8Th98x3HWuKn5af3FBeRWKFgqUax
poVnG6A53bGGuVjrlnSyfLpy1zWvxGMCG4IemsfykuUWyYMlDBV8isvFEGoqsVsb
J3LlrGQpPqqjgbL+ItaG7IGa9hIV3fDJjjAlLwCnfHDJmGvFZAKrriDRInBlWYKe
Pz+tjdB6/5o8H9JOvOgz4XABCYUZxBhArGzDC7mqo/Cib95ah3o2TITDMuIl81iN
SDEIeXDgeuiZ280sO4t8q0Tzsrkj0ivO1R+MT24V0Viv2OZZu8qSR/hvd1V3rgkN
gMySp+W8/sKiSEkYS4kBQoKH7afqaMiojIUn/8dbNVhafmqSEOX2bfX797dM7O9S
gd+eOP9ThCfaAcXe1XM4X+md3WGawkktz6UV7n5NINI0fNdvM1OSPXibMmjXnjqn
3fM8B+VSIg5l9uNLbqnY8kHPnoggWothnBMrRuIyDUSVx6aVV8z0Jws/fCSubD5a
`protect END_PROTECTED
