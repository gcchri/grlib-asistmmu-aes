`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cU680RdCMhx+I2kV37+Wv7oPoZ8eLy4ACAI9CEh1UYtmGCOz4Y2OLnbEfjCq3e7g
CpKzyunBFR2d12tYDKnnCLXZkNNlNYxk39XvCETaRoGbfpbAvlHiSSA04wAG6zqr
G8NffpM6tBBjcd0ytCn8PwFS7LJiKQ3Pw33Kv6kzsqilUutF8X96gLccb3ij+Tpp
0eyGBqM6xwucxiBiHXCq10d7Y9/dE8fdOaiKh0f6eLxZnZ/ktVuon32o2CnN+fvu
b+4vey146ix7JJdrbrhEO+v5QI9BVFEGXQ3QdvxCfW+Qn3JctzRyjurISEirV10x
t4AgPZGZ0Bclka6b34FGA9Ir6P/Yt6uu1DlsNhMZIf1upD/ya+3eBONg3HiJrvof
3pHZdSpN9/OpZQLRZzs3rFdanVVgjepMFxlijSrK9F6ptKpTLOwNEpoHoc3NP+Hk
lg4Xjsqq4B8aKG7ugzU0tWJdKItaHUpBW72yL1c4mR871CrZjiRyBXINmHT8HUj+
Icq+aiPB20DsTxhsQm8c5sOW80okgUphkjk8MqX9oIRIhIsXCZk8YyU8MAuc54nZ
rS9erBlIsuXRIXS3SoTn11pUrp0/OJgbVARBQUnYW8xOX4b2GvYjU+CKUMuExVu/
Xa6rVfBOHSRf9FeMgYV8GGcrLG2zJe0z9AtjgGGqxze/RA6vlorZYfZSd3IT2zw4
Qv5ZwekGSgkqPmlyerSAyxGLgvDt4voWjWapIwGQulWFTeknIf9UAfURCw6UJWKr
MI5X53E6lYvX1HD+l3H/0XWOSVon0KRDEzNW9MB3dM4dPIo1DUxUt8LnDx7PFmhD
0RGAueuEjYuXbzXnJv6WZHX693/44q65/nOCqnLqlc9PLCpyunDzeHV2CKXfZk4D
WXBKDtT4Q+YG6/EulabbpK0ijM7B8UrK5ywHSv8GruDHTZErQ/lxNTjrkLHGOgUF
9vtSUMH7rnoNmuFyGWxn10olRd/NnYNP67l7Pk/JEo5dJlTgyegeV+GxY9+AJfoC
9RWB65Nn/0xz3jVJdTs8XuNAgtUxhKyWVd77HhFQKcsSmp/w0u8e1zdyk+jYzUhq
DYIkKRalFVwki4pbMYq3tY6rQtAuO9dDcM9XqruUCShfpoaf8lPK5Uenzk9NQC2I
UyF8DzI8aDajbEiJ8FVCQlAu8qyJJKMFYqPXBhALdw2aWuovudGi+Sb3J0xMS19i
wWIKe1mYirha+x+V7fNBjmkitHC2PZlR4upqEjjYX4lPSTljQznC4VbRRyv0R495
jeHXkAwS4egbBRCicDYNvCnksOz/x+GjroL75AZ8KoMa1g77fuhS3kLbdH9WWOAK
aGweUeRs4a01Rqlol2UxqdKN67FVVkUFqAg8RRkixiDPhMPiiNc/UVBsCJD/mRDp
ZBOX2Vefp5ElC+9o/q0JKcp4nlyR7de8scaRKixsJlILxWlLM1AEigGAeAHl18rV
f6wIzwuXQk05GyPQE491PVkMhH5tPYGWO2kP1w4oLLcAP1Rmc/yxm03eRmHhkinx
c3oC1AOsdbsLTVvgDjUZoINzEhQ0QXxGKi4M+1cZNMrSVThUa7jPBl8JPyqZKNCB
eh3cVCfECC99BplZYA07JvpMtNgscwr4a74LPYoJqHO4Wvk0CdXBBaYm65b9LlzG
uvgOU0NGVy8EBq6aDsQrCHcoj1zqQGhCU0t6ZPU72r+tx5+nowZVhkm5XmZE5fvq
LAk6GjXwqu/JpyKYjgetDA==
`protect END_PROTECTED
