`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6fkQBPwpkhxRaaDFpxi+SeocimqZSEUfo4HXmH+gEDVsdsYDJg4fGWt1okqarGcP
LI1Ubxca+kLKdVX2zNTXcSAAgc1aINGE2Q0FhpcT8kTdyNzFiKgKHv3EWh8XFpso
fHrB/r6kxR/IolUzJVKCK/7hEVuNPtBIzJi0hYjprqZEp6/7kvmrNK/SclqwSb/D
HGi96JTcfpfbLvcY+RhT7OLi79rrQwxP8gwfn7CSVKKtypsGcAvfFRg38uguHfr2
bNycUFBQXM4Ki4ems6AfGupforEGpAdIwLiWjPgcMy6DZ7W1jQTatpt2r61DWqbF
2TIWcDNbLCPP3rsacgSZS972NJ6siD8L+Su0Wt9Xn5Iphxe+XZ413C430i/azjP+
EDAOtVdH+V0k5TNFT+TtHpHHPqtaDPdjH6cf9tXYuXS+i/qWInNZ6ZAGNwi6MHs1
iZ2/WlSifk+O1Ea+8klW3xhcWJeLHIh7oTZ17xNjquiFi7ktzod5haVFdKoHgn6T
ugh0aBstKoDFHlxUhkS1jjH1D07N96+LlOsiotJsuBy0ydX9VxDSD2LrbbqekBFi
1QzsHIEdyde9xEyvTXLI6h6j6+nOFAGwxiMGCULtd6rAG0EsuRPcZ+KXOPcXDpDI
`protect END_PROTECTED
