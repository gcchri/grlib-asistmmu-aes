`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HA1h2+ibgJyZ0M9uv3ptBq+C3ty5+S53mpe7dL7+7WYFWTI35Nla3m2qht3kDwkZ
LlnqcubKqAkMjyILAb2WyyOl9Idny5JoVwCtkTOcjZrZmEWSkvyR0iwBI7Uf8Fqx
EI3Ohog7N9MOUs1qtvm8cQwBkgyDrRONjfXDcHwbaCbWxpDD7DZEc8KfZuYKVhBS
EXsdoB5Vup1Fg3dG/sloQM7pMUrS2EOpQ9ClhSrkRGseNPNtyodVCFNaxEtG9Gza
4y0mFnES9k3czljwaBHNepp122DNg6yhu76o/4UYCi1ohtn+tHKzFrHDND5igTd3
VWB8i3hGsqK2QBAStXNnXKK4iWn9OCoi37d8ECzduHuOsJbML+3A9yih5QmMrxN3
XbghwM9diy78bChXxzsgWLKOw391uE7QiPNlgB4nk6f/C0AMuE8bv4m4zTSr0HMZ
OEBJLosx2P6omA37SLJ8jjEf0GN2+BujAOAiv/5Cceqk+I7w1eFV8GgrhZho0Fyd
w9f6DjZbItyBhqVaGl1I5A0dPVXP2LUiD2TfRGhIV6/dO0Dp0rTzb+zjIoOWpndj
rNf0ElHHqyCziRp60OfyXRugoRflH7Epy9lLQrvBIl1+bj3gxXjrUgL6mSvq0h5r
Y604fgOJE8V0UFwqRJ/+zo0c+N1QQ4Cf9ugIZAjq11gxPm46DHWtNmdIlujiKQVi
zYd4EchIYtKhRKU3UXGL/RTDM0lrJsKZ6AFoU+XSQuXHQCHduGfC9CtGsBob1bOR
ufKSkPxHweYMeO3bQnsdwYRVOuzwRzIFgLoRmUlRM3UYxg5LIGlWcFY/bkFhzynu
DnliwRww0JWFA2UyTLgeVXPUoXGF9ib3bTY70szuS4nsXj6fwwKGC+EulBO8UfgG
MDXa38ACcb1kicjCuF7Cuc368DvkvbnpxVrRhq7ALx+w0BJesql3eN6h2krB1uwe
pk1BJ6bZbjRg5SLA6z0aB0eyxtezSsGryD9PB3KQ1J9xF+lle3e1QC79YuNH0zQQ
v2nR+Av6GaXh2sFrN2N2Eg==
`protect END_PROTECTED
