`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gh5AbbwC98K6d1u4jUwWSjJMmJnKDI+ZZ2gh/BgyZ+8CJQFnS1isvcDFeUrlW3jM
bzi/1FTpD6q5qHBSVDoj2EEi6qgkmcUhIRSbUatL8by+KNYl0SCS+4qKq8Tp/FCz
04znPxCLPgzSquTzpFCRx31P51dFm0fHjCpX3iiiwBUkwf+iI0OAEMQ1XBt4YM3i
1meu6erbIBWWKiTSFQxYc6n5p1wr3WJYbQGnq7doVWpoiXqcrs8B4PfKUhAthlHO
CIRuKcYou0LF8lTxOZDMwEhf17JTauIzzYNcqt1pvn9edCOhYz5dbYypMiSuwHEL
c091KxAtQ7R7NURsHtqggmSeYVq9UdjGcqqn87z+v2L4frI4xKdQBhmaW3+Pf3TN
7W3svVhhWH3wzclMr9uD7Bc/F1zPsdCnV1qAzQRCQmAw7qyjuvsVF1C+kxNKJytB
jai96c+lXgLbbT02xGbWOGE7xK/FrcdmirJRDi3JaaBiEmXAiayng03E1Welezj3
UXNgJzKdTymoYiDt/Bkbb7TFBF6PCyxteg1xvG1Y53eaI2MawgIjEtvjL2m0Yg7I
CGMJPU1LoObqJof54gFowBDeVhG+k1iMQLvZqyyQrQlYIzFE6gmfWphQk+ZAnsBn
eH6zlz67rTuTx5G3A89WeWmhu6Ku4qwTQ6JtZnMAObtcAJ7f8dIyySXociZ+Yxlk
XwkCuyui4xECpYK1lHaPWUJlxxvNA6cRQLEWRV5CyGEo6l7SjqFvIzMe3H0xtl4F
qxYBWcGQheoFbcf1kj6Y1ygub2NxqC/M/IwcF1LBLGWqsOfYbkME98twlspC9S6e
X/Iy4UdEKZWKoPnIKZ+gFWn/zJRnh1QXg1Ur6VBsB9b8ikZnjNlPFHR6iw5yw/sL
0zGpNf0T1Yy50jSzPQ0dXTmqCXzNEwXumov52U3SGYM0KyZTuOMwK1GKixIDWZrj
AgK9KPfkD9Ex7RSQcl9paQ==
`protect END_PROTECTED
