`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jhJldrgSyCVRZbaGZCms71ZyqGhre7PNLNJ0wScduXVhHAnB6ZKOfeKNUxISgFob
YmTrdAtR507gOXPXEUHwFJMu2COk2pTvSKQ2+I4V9GnzEUvvG9Ea/Uib16Vh2m5f
6rS5z8RMeNjLkuhrLR1460OJ/pryZ6DVb0qiKZlX/w9L179IUZA7n32JmdLnd13b
wltTHQz9Hd2LWa/5oZHRYHBCHCWx0yRpe6N5/vhYmER0KwKlQJ4Lkobv4O3DcjFF
UMFOTNzyOZzgvHiTIZbOyspUdrQ2DCvcLvAV6uij7Je5snfN2VdRODwclm5uWNcW
gwh1685N4kGDFl0UQuMtQYohXhkqUSJGV5H/q5mni90Kn4RY/XTHCLSCbbAVIBJS
RWNTnXGbhtbs6IgopjSWK3Jq1lRlBr6rnmvb5jhSI8cYaEJLinwJsdBo4hO8l35w
BWWAx5IjGyHFMkOorV1moTdBqBML+kt2lzeBc9DadWwuAV7aNPZUloii/kYjCrZK
g4EyOUZyMRwNbeDKEQBe4A+zmf01B//sgY/9B/fbV181x9AmRsKNaZHPSCPJ8Yst
2XXBaFDPnlbhRqOlXI9HeYpBq0ovEviF1lF7cIBS3gxdsPZZi044YenN2Aoes7K0
dZcr7Ybya8F5I+xEtxFVcA==
`protect END_PROTECTED
