`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r3rxG0J8mwTtI/8t0IblmqSPEwMMNR3Ij6Wb7FKdTQy61Z9PUUHp7K6yaazLIc50
FodGaWKh2+zR3KxtgyE66rKfMY590FeuvNq6kYfGw7IVoOlhlGfPQD8iHGcK0APs
/05Xs9I1LtnXqY2TCE9y+RMrdDaMyadi++j9izq+48nkNwNfp/XVSMos8HlpjCAv
jL07fL64zM70Iu5wtAsRGltZYWq9BOxCt/SS5hBHX5hC5C5w+XAvXv8op4w1Q3Jw
uNi2sx6FlhQwCydJSh8s3QZeLBKQqX1NR5VuoMb8eghQClo5nO8w3lDzd0jkEPQc
7dJcqKIGl2HERtShtJry0xTQ2/yNjIWxF0DcnPOIbP3AiZLZaMxZnRqSMtLC/HeC
uVBrwIw/nw/ceeT/t5o+XxnH/26lyJOw7Yuh5TEe4wUTWMrmqT1AGVSCWJOVjAcr
BQfPoTQh+ASF46bhw1/s/s7aKHiGZJpZHPWrs58zh9YgCfeX2390EGx3kBG5/BsL
pcSyfqeseCQei9NZH2kCsCFIPNfvsaR3XDpSFcrIbkYNHYAySIM7XOi7KFxezjlp
8J116+lLfYGgi9jazTZqAFkMQfplYD8jtwn5LZWzBSLFChPNqPlABsc3idqU70fN
pJAITP4PggOmnjXqXoNRF1dIFeRYAHCnr23KRffNWUds2LQxD764eMmqz2tRlhDb
ACPcHo+6p/Lp35NpffM2NiFDlmF1bnJGxygv4hBFB2jUC5H6fuN7PO3kGWh0/Xf5
FWPH6n3k81SM+LhIziKh3nApeJFoUYUWA+F7iucKgm9NqGfWCNfcJw8Y7q26A3dt
liZKQ3qDEkHjJSqLLFgvIV9Kx8wv8DtVc643GTuDVDymCDbUnRAyBeb3fGevYMHY
nGo0esX8HlHw7wsjLqwqvdlVXtsEaEPBa73MQ3VxkDSt8Hzuw1U5vTyq1BA4BAao
fCuhuQlvfVNiUQ1NqsigZ7DtBNY+PEYktoV80coLDLr8BZbsN8VLnhPJxN7VxiA/
`protect END_PROTECTED
