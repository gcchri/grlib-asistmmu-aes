`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d/JFHCDj0c3Y8cSSd3BMIWjv84rLPhfdXaUtU/UVKF/Zg5cVSddG4IIpdZsBfa1u
pu+y6Eld5yuwWkE0XFjQwVi21nFcecfLXaLZO5yZY5p0WeG2IhwHczVHXIfKJ4AJ
U7OorjF4C1eMNwjHkCFtTAei+zDVP/S6g795QVlCDA8rYTi7JQDOrfD8YD8gPUkY
KhIBuaIZQOQArg6GE1OxMBAtrCGH6cZDmSBFSptjfapS1wCAnEgmXisxw5M5t8UP
cEDGCf0fjENiYxwrQ7Zic8Pk8E6DPmO8+ItruR4w1IhqdJQ73a5gSQtAJVShm4uK
9bS2gy+XKwe0nxl/SyP/rvoo87ycAk7e9M+laxNls2XFcWHpc5HrMNAe/db7WC+d
LWz7D5vgtaiNCYPF0sdEUS2dwAMmxbPOgOKKyIZJKesTodvFQ6D7C9K5HcLlBExV
nGeMuKTDSTR3/omC1cVqHOrop6yjHdUHcrnRZZaniczd9oA6F3xVbvJK6DTmBsj8
SRdnHGOwSyrjIUyDh6acpW/TpCWQPdFKKt4Kb5i6lsUejQmg7co31yd2optox4Sa
BRPc21RxwpEGJc9rn7Y7s3wny5f022C7DGSo5SYojZruufty3ggRamx6mRlnxQ0F
0caVba5PzaUQMqPtolhpaywLnBqdcInjkGLA4Y60LaA=
`protect END_PROTECTED
