`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Shn4NHTvd/dMCYclof5uRCsfpOSx8LYVaHWBcRRmQBpaMWIczeDcYwZWp09DU6a
Fyc8vKeZcA+Cp1Z2Q6znzIIBEn/e6mlN7TYOxa5BZnqWdgyvJ0caZmIwN78D/NDn
DcsW+74X0Kn9imIQwG8a7VKizcKdQHIYxfvD7zHqBrfv52o2Uf4hptjrupKzbn6m
dFOC2dtWHc97p4TTuIbKV74DWpkDuTpFTPQ//Dac4aYBe1E/I1p1c2WZC5TSHx4Y
vOfpNOcYtY4NbkMF3LWe2NTC76Esm/1nna57192WtJ2GVS2+PoyAgD9v4a3z/JLb
a+mSJW209gxc5U4+Cm+lhcEQ+5PP7DIfR5WXufO7Mj/bJeHUhBzEAysvyv+cwSaq
64niDtstOmZui0OBHZruqdwUcya5IYsNY9NBgzLWVQZJ08K7ocvbyHrBOXnoRHTF
yYJ8XO4eq2uq99dJsNtXhGQ9s1CyeG76T8BlZzqBHgYZVjoRAOnZbM5cLCuHd9Ke
u9LHWucP04mxcDn+yFBs8Nh3Dp8ZNJq+X6bHmYn/hSOUk/P21Yl8QcJULt8inR+B
X9TcVjzT2oIUrlCveWPdmT1TUB42ELjFhjm4mjAztvebtEAEffxUW0uzELI2Lqmd
cBQWIOX2YvH4B656dlx5bQ==
`protect END_PROTECTED
