`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aMAwZw/HilS1XBkUmkj5tLtR7A8DeAs92TmjYsJ2Jj8ZF4ipcP5xDEhYqTad0ZRd
ZPlExUSxpqC2rPeF2Pi8Op410IhrGbHHZsOl3WHnwimC+/IGA78PaKlXw2SK6JcG
ciLq9F9llNhtkvvBwmgP/1NN0Vn48EHh/m88PToBKZFoxiMnpFfsN3e/gjjZ131n
S+Jrjwsvjn0XiLPlhAq2nqd1XtMn/qP/OPPsWtTaLjEv+dEK8TOBdhFp7YQDQhWo
pKHwFjBtA4VlccbJocWXYh3Wb26I8uh5WiOgiFa+zA0Ey2wYq0PqvA1kikVZp9Zb
XFQG0g8hzGpyEQbKBURwe7jy93uAxuCANGIQTPRaNINr60UCC09qFizGmb5s3QqK
BeQKfne4q43zkcbDUi9Kw05ls65YKC0wMD3Q0US+yT7VKnei0BDoY5kuzsCkyC+v
fGcpW823fYEtAI5+KBo0ToKOOio/lTYSJHMYW/0bIEZ48adCSJ3gJ+AWNPsuMqGZ
t6SgYdf7YOsmRfNnc5j4gIlG6LPD5uZg9e8XhRl2GhmFfodI8PF6ktrSesn8bw38
pLiRaU8lrvhEFtLX4XPS35BXIFXEeZMS6MPA5fpIP0ttjwi+qzky/ppEgR2FLSwx
4PCkZpjR7W1wZuWlzkWThFyvCr3VXz57NhDlp7wHt5Nl3MxyrMZ+LRWvsFX/iQUu
+UP5puHIFYeDMdJQaoaxzfckoKaAtPsKTuHXOtBw08hdFvDwNRVcrbSy42INw6QW
vo3g36a4Q/adsWOF7A6N0q9eSwZM9uo5wnRqMJXwu4PBhMOgQrT9ouoY3SlKJVx3
Nfwp6InZJbWqkjkSNRyGJw==
`protect END_PROTECTED
