`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GRrTC/zJbO61CrALStKUjLQorTDi++hLvuxDngg/rW0p0eW4VUivkJn1wLd8rwVL
j8gtZpIU4/vsrpgSKg6FuyrSI2UsKqxpxLSd514fqYpjqhCh2KPp+eKno6g6PHNr
72ivV31JumKhO9oLbNgrqNSrh9DEm+doOtDtsurhP4UuZ493uucKfLc0BQDCtgzJ
khRRX6RQRYbiDub0ti/AoZ46cyJwRf/bLhgXNHYYEWm6kxTK1F0T/HaHpK+Q5s5m
d4nBQEXfR7xbVm/wq1DmZa0lCAqa2GaHPJq5Dg4emykcVGTTBH1H1oTLqI58ABQS
J9vLeU/9mhZdifg2Pj3KHkF4Au6GlhOPy/0kP9XnHZj7U0JHmoY82dZ3rzrZrC0R
KiCkkvQbTH8y3SWhzsFMUMxSm77jQMCMgrc0V+9oC+3PtOqJgqcJXZhvxbdWATgx
JB40bcmgSkKpNSq2UZOg/eSxGQdSccIOnw7wR+01t3+eEnmVVHKqM8QkfQpvwqoK
8MHDKaG3qkbv+lIvX+J1BemP1Wf72maGRHqwSUh+4M9mYjRZs+/XE3809ZsWhiuF
guw9bveTqkfVa8N1rdZoXEUV/lwHmg1K0zIRvFkCrWvVTdzFFvUJcoLzBemO5A95
`protect END_PROTECTED
