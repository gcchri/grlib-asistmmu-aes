`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S0mUUBTQS63l52cAlf4qFwa6Xwk8hz5wmBHgNGTLmW64HwBfN6h7KR5sIuYW6MI8
r38yKIqeHr5fN52E3zbmaRJxrKhJsOO9I/ZKS+DxrUwkqXy2jDqlns2SMeZt2lbC
CmSqZAVPPzPcPgfbfsQxkreJT+H+lPqMWtWw69im6HRhCeHqS+ZuQW7if0aFbVqR
hEb7gNu2rEh/YYTU2uQxDGN0eF66JJF/qjNKzGqFQYKONmB2gf5H8FJptYOe9SiP
cpdEhqwkGxF6pwdoM1sxycu0O5Ft092k/VkQlJ+olF1kEdsBDf7q3dIQA4V1SVse
CBm5gqLwtB9VjyKdpUcRxxXVdw3siPp+4OXekb66bZPPlVZ8WF53Z+GwNIq9nt31
HvDmfm6l33ys50S6NzPdNGdbv5cWyyA1c03stdNkZH4=
`protect END_PROTECTED
