`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gtzvMWNIjRNELF0JRzPIHU9vrtrzbJqsteg9zoAoIxXZg/r3u82UZa6gC5xPOIaJ
J2Bb19zjf4uPDtZ95/8uIx2Ia5MeIXFe6e03LDjh23sijUA5BXMdEX0dqNM5Dj/Q
HnxdIdvJP6e1AFUtrs4x21aDNnJ2Vir0ZWvwfsET65gAOf2LL6wx5jw4fOBvgeIp
d6nnEYh60HfSinTqDtGBWUbv/uY3kI0fnkOKclsWFtCdWP4Q5jarNDl0o93lnYYy
TMPRpoCaXs+mG2gJcAHiufoipwrE6o8PUWor7W+hxsUBkcaBBqWagm1uU8wYAURS
`protect END_PROTECTED
