`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WPToJFDjuN5VtB5fLiEtV+L4OcRUT23EbF5f2rJ4obzDGAya5Pal/dAm19AeBjXd
VbvLCE24VGZjlRW5pc6yR6mY5wpbBHhBxNSOQVwmMl7Pd9gOB4X1/0h8f97o0QHa
oMv9FYM9/Bjs9O8O+yJyI7++ksyor3e1J4/+d2IdaXq85rTR/gj76G/D0ZTKpmzA
8wxatp6dzpJZCfvZqka1qPyFljQn6F4x3lMNGMGEIofkB0lToKNLY60WgvrDc1oc
7zJK2lZNn1oyN0rKpOMiYtUDs3urBCq05iZVnMCTXSwDXBqPxxf3UtiASvCX4WwC
mLYCrpOasdgA+hoMhF4yKVVg+dfrtJyWMB1N4raekgM0qgl8VduGhgxMLajW4ia7
JBL/2qaUblsi8QQ6RpUpdSXlOYYSoban0DDTgagM8ZOiHmv0TvfT/W79NqxMiw9x
10oOub6NmxnCfgbsAuv/g3PjOjKgIJt+9eQVR1vOsrzhqpSgaZMKnZNdParrtuSb
`protect END_PROTECTED
