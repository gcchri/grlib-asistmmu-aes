`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rwyTc2cAIBARrrHB5OeRWLfcQoEzAiG+COmiiYKH79mUTaF59s1u8qGogGdaRL2c
ZAv/BgjpP3IWrqx0yJaaWO+ZGpX+8GUj9JvJLiaJsrHMo76azSeXZ7J5aIDIXicd
kMi3oA+wdSJRlQEcDPOyBJbCE9LBDg3M1fUpESyFG0B+bQE1ztfdqX8QFYAmo2Fe
xt2+z4CPNh5CcPEXLwnKNX2Za1ZoWXqAK0IG/g3hQirNn3C3S9h0uOqB5ueNtN4O
QSAYLKeFVUly7FUcd43ilLJxWsnKC7xajdIma/ogBpu9lXyYuHCr9+kcjRpACZ3q
qtOYd2HG1xMUb8mLMmsK6DcL4g+lHAA8+T1g5De5pA6Ugd5uEFudyNeXZcd4GG67
3G/dAdS6V9amSSjDAgnZoK3nR0CjSjBDQROUG3hz2PluraN/Dwpu+iqH/PHFbhjb
4y+KkJyFTMgpc3gZrfcHzrmxwY7neDXYzPT2vecID8z2Z+hjEsYTNCsnYbjPRE8f
ctjHEPCFSHzYDAQ5w9bk0sobV8jnIIlJ6fRKNeOJFaf8vnaeQpqq4nZlLqbyO+Iz
ED7PTJI5VTE/LhYd/BNvBqdDcvKkrUPIJPUGkqvjUIk=
`protect END_PROTECTED
