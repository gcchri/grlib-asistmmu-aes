`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ezu7Q5y3l7UQkPCothxa1Y/mxKor3AiZm3HePF+fSXk67K7SrGuMt+EugQErsNFq
zeRJMB0Nqg3WoiZZhbYtCyLqvdL/njh2yfyGWrX92JCTg3EHzfcljQp4np8pQY4G
iCDmny/PyeM1BzxtvZQzxyfss0CTqIh3aK5LTKeEaaxwF6+Nd77Qi8qTvDPPka0B
iLAJFBkmRBTwEusXVG2cTq8Ql8Xz48nsFOxm42ntB3PKDcy9auJrAcAd3cty9Puk
aAtFUo2LBjnVpwTw5D/dl5d/j+yeVqsQA6MEcB9bCRxukfU4vLP99MpN/WLIJl5j
2QKH6B7YEFJX5XOPQQbyXMuIo0rGE2Y7Na7Za8tAA2JhNDUO6dTU0TaOWa7G8aHz
Hk9yWrRq9wm0b6awwaRgGdcCmfR/Z886kyPAL5e+Sqr2QHxtKLYZzOf1XGZl7DCX
/qA0BcNxXHHKX7uIP9Agvt63UcLecm+27GvfkE7AmFe85g0FFqEJ83Ytn8kCVhG7
y2tSTZ7+y7pxH+kQ7W6XhsPzsS5mkJvudbFrNBYpPraDYbpqeoQrI4qxfBuwiKwN
7EWJS+NZZJBRdoDL5Q6rPFVYxekgA2F9m0S+F+ljfNJPpRmKwJzbYGt7OKnxZWlw
`protect END_PROTECTED
