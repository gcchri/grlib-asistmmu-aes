`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XpxH7C4fkMzPbi0rtzieKHVpSSJdD73/d4SrGB5LB1qpfo+dRXSzJUxJHvlrdWHx
Eh45OELh+cyuBQalPEiHPUGV9AXf8klvHrtJE4If6uwB4Rtir00naXdAAUYoi4n5
ADYSjoaRrZLnwYmE8iJmmTFWw8h7F2PKPsDi1qrkmK8EmAG8NVoBalheO24dPNq/
rBfbKqlDefxcCT5cozYrN4Ay6Kf2X0qe5rI6LIr0CfZsh2DqMsLoz/vhevKK+60C
sNMYQ3l2fFt3f211ODqCrPe8gOZ4cNdAndCbRPHE9pxz89G0+8udjfjcrSE7Ez3V
/srjBSrZT4zpdY9dQi+iNg==
`protect END_PROTECTED
