`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oU4i5vBBkariK2j63nwAmkf3btUyNPnLVryRGNrv1RRhfa0VKcsGSHxGDGILI7gJ
IBDO4Owh7O5lrelco1gt6kTAs/7bZ4F4ac278zdb20lcQEGzcnAosLxuXA4fSeNX
ntLIngLuOVt6xGpRqbSz7nMNlJwgIC7A+B0gR3cQNbyYY2tX1/wcj4STBF4J3QG4
OU4/30nXUoWMq1WIFvhqzrwsLbcR0w0bjGSiJey36yqQvaBKw7H/y3LT41rKOVKj
tRMZw1q2Co+NfDWf27CujTL/D+ab6yyws9Ar7SuFOBPWklUV1BHqOx1fzMTZE/0p
palcVBk5cBFzoMieGi5QJFKX2pB3StKdT40NOOW/Y0iSXFErKxomuc+5pYUrefZp
1Ya2eGycHYB3iHionMmIvsVhsL9vSZQmC1G+Q3B6NDYOLlUB3tFMYdxgf18s9ViL
yURsSJolt6otRGaPGn1ntYLrj2OOzQsds1rMseHcfD1KnZRRJUJUYd3AtkXqSkfA
9wQB35cdvT8/hxZeWSau741HRET356lk1ENscEmTUNihM737j4ombdCd2xxMnYj+
YCcU7bMMwNPXKFfCY9yHLnUfwyZIYv92obqyoAC1SH1cuhS5xCyp0P2TzT3sZzeJ
+ym8vr8R9601ekH82HnScHlj3Y2+lrw2ZcEKO086uH2LOhCB+50I7mqtwIRoI1FG
uwis6znaueXqDWsx3jU8A0WQ2VvxNjNeDuQv0O5aEQSuSlcPufzPX4uI4mxlBkjH
+3Gwx0NTRjBdyXlP5mqwFG6HcYvPDGjLMb2CxSR8im9aNA/BAxP8UWIJHeCOFlpc
iWDw85qBkCZyv4UOPlWTCBuYywNqcVaIRjyF4JI/gss=
`protect END_PROTECTED
