`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bTYiYGdL4ETihrIZ4Gbp0b2RXMMQAl54W/genOe92hkM8ZXjH8PDFD7/Ih9SK1jz
Em4LYIKY0OVV+lHAj3CmbUcmw4zkamJIdWJZDBfOoVa6BHdQ4vjcgMm1EEQ242lW
6smpTvfppbO8X3om3VgvzG1JST99RR8+jINo3hjuWq7XZUHsolStqgR6/3+UFWzZ
v9CAgp8nxmHl0izdW2pIpgytxJ668wCpgcbJfIu8xBfcZ7eDcG+mN+f0ff1Qc326
KVqn+bR3wg/3ap1o8FfRZP0oolgI/wzmuwu4iax/bnIwiHszsA7JLGPs3vv2g2Ih
YqIDzxPinlVndcINWnIcMHXCHKisb25N3YGrhItq6O0nmPo25IOixZpkXihY3n0i
Fnk+v5vrP3FQSINoJVzzOIeMWwJUrDsqPE75+UhEEON5Gd+ckoahnb51f54nd24T
qd0Y7gMlm5i+haJYv04WcDVCEVFVyNTZfaMB0TbfTkt96wgmVY2s/3bRMCXibEfc
zS2YPeVn4hPbF734QIHG08wqq042HRLKHuzwygMcsahtBfF5UQYC4m7j/aSW6ijs
RoewTLGh+1p9ISgzeGwJOnfR4GBKSmhCj5VEJaEXufg=
`protect END_PROTECTED
