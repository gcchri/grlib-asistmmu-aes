`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Grel1Fn728RyW/yd3tT/D17rV6n4crwwZ3OQQi795PdN2ww6w8cpDSgeTJhiTlBe
Zj683LEBg/LG2cJ99CvLHnAQxqc2+eK0JY74lpaLy/3Ar5fKbjGi0LWQL+1AdYuF
dzcmXefh2lmPgjMNc2TCtsHt8LpjQBdVaHIvjV4DF014vngogK7bVpfumT2alB48
/C2bn6xU6Ag0WVumIm8MfpTINqXVfmkVP0HTpWDi9TEdMsRJ/QTbgpJyq8fazPEm
GBnSucl3yI6WNHnRWjxtzUIs3si99EyPmDvAmCHY9HGTJQE9T/RPrUWaMddjN/sG
oaaKhOmEFuQGPWafVPgr4Kx+y+IAhM62roJ2Xs+rvyhz+yi6J+G+aA9L/XAxFIxC
gLspsGaH9vLaEaun+2+m1AYYzDB2u2V5UkoHQwiCnKKMj2VSJ/TV/ZO+mNqlW9AX
YmtYOdZPb/r7OxaAk7YueR0PWnkc7D3MNvYMvDxnU47tLz27nZMz7qc6ufHsJR+n
y8P5OE7BIJU1fW7NP3B5dbWb1RQ6dUS42SY6aoa4fqn3M+IxzwdM+zB1ww/2sTdt
`protect END_PROTECTED
