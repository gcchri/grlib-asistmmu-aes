`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V7wBXSeIUSM5uX5osSqBypGZm8Umf9afl4ZhO5ly6p+24X8PHki0J5GpgJT7n1ZA
WC3+PHYB4M6g7o8Cmz4GJ5sPi3vmBBpOuzODuc4COBDpouI0+KCQMJYF5G3380wp
hGFNAQzhaEyORs+3CjtSND9xiqcTeYHCkJk5+7iymcMgZANe1FfLcIw634XELGvO
rULFxoxyGJFy4adAUEXZuwAY+FpJxKcGPCS+X29J1pSKBTLL3LzfD+wc/c3z9kaA
ZxOI+12xD+csMDJ6Zp4gE9Ny1KJpyVG2ygrOTH2rEZAhQmM7vggk32Qn59IB5Cio
ZtzJvC+fr5MdjSKUwEBfUqK7oCJWoz780nSjTXuD2CCjr1jTR7wSaMx2ikCMU/JF
/b/vi87bNlpfj29dtQB2yEqJMRjGytm2j8dEoUncVVa2zzGcIzuGwkLHOVWiAjhz
tMtwFe/lHwb6xakz9HqZxaR4K7RL9Rlny5lL5NmQh7gnLnqLlLNSCGhfSbriTOxs
`protect END_PROTECTED
