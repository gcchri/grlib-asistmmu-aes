`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zv67Dsz5XX6SnKvzMK3jEuby2B2/O2NEng0jo9rOUd5ti+5WoBseuZ74ZY1uPQSn
VQtyuxXlOH2Oyz+0T827MhfKd4yMgx7PREuwqaZr8Wr/pZMMRpNg0NlJB6QFNDua
e5zxASvmikPyUqE89CEdL9jti4C09cfiIxU6iyHbcS33qlJxwZWcYbwEBgpRJCOv
YKn4RB0GWvAr8T0CMa7uo3izwQpJ9tIPyEDI+P1lWPH7T/iNLunfCPQgdCLU41ZO
`protect END_PROTECTED
