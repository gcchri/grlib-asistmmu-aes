`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IVFpw0fseAFBzaLpWUMbq882reY63ox6jsp6U2ylgQXVVLsIUJ1CqHi8dQ5obbDN
WFIUPas82sSyqgKAgJfewIa7EgPTn+2nEJmxTEvNorQZyMA4AeupYhU0JPqViFN6
jpMI2yKNQERtHRbdujCaDRuyV3+3tWsrCpSZWykbiqVnl92a2/+AQCobvEjDOcy+
Mra+M/eW4t8odfajDkFnLA9l/xV/S28VAyoj15mbWtZnUZaaPeIWd/V24YhHCoYA
`protect END_PROTECTED
