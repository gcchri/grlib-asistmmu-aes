`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wf6hAzfjiVVsicOCUvgfgQsCkc+3db8U4o7hmX7aR8zNF58O9y38by3oU2ZokdPl
G6Xlh580PclvQI58ELqwR0VceT/h6LGl5VPOnIa3r6mhYiMZEK/9fJ5gztqhIYZ+
AJ2ukpIdep6xNePHcU2Ft3qBOvAa6WFg85B23oxrPc6tPFAgsvEAWFfQ4zfEh/0N
oyZdjDWmpAHZE47HL8HwjoTj62TDYOWzo+g6Jpz8aiVgSwghDBCyo1h/4AOsnFBS
SWfuBDZe4FWy+QHcBodPh4L2zGXCyAOGhp0uiYQ9CwvbXL/90+Hv5QDt8lqPc6mT
fNOMWME0BgWhnTj8iV2T0NQLGRb2VRmvkmZLF3zriGgzM3w4VjUtYvBcrIJS6vhP
Gb6vkKDNIHWZNmUIsfJCF+gfpn49EJe9YO2hRh3bhx1hFK+BjGRa/5SrxJaSv3Jx
QRoHdPIib12EtPyytJgTfqzDxcUye7pMyvD/mJ0TsYYLd5/X7ArSj6zmmSHoXK6G
`protect END_PROTECTED
