`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yLYlVGNHf8VAtHtpt7onQx5ZyItkDHzU91nmSovJJyz8aRF+pmU/bSrtyIsNGqna
QlwxKN3qEGmEKiDAtRvNqbAo+eMAU7+x7oQgNqPefZxEi3HykruQ1ve5vzm1C7EJ
ydPbwVEhTxXF4YcmxIfrnD8hLQFTTlSNKoEVSl1XOqFTe9CnRufGjQ9aWHcVNTK/
IuSJ6xIHdRPtJ67aGKseL0RLLD2fxyoxzFlrGx0T5lYbK74aASpdw3MgFuumW232
2Y6nC4UQcf5JkTfxIhkUiRvXK7zt//5K5vGTDIh7e+4bjG6Cq++PgyUmmvhE8TaC
mqvi5ui/DdmERLAx2BnpX1L9WdrYLKl8zzPDAOazntxJPjVGbTrw3n+wnuiAcG1u
4x3rNSro2PzMIb+KpqXMKN4NKJi37S4MA1qpo/9YWyGoOgZP8aEZVoovql1lL2vN
Lm85h1PKkLaBMCWYl42SKdMAdCCtW8A39OZStMLo1ycG1/dpWYlAeNaoJmGK6s+b
XnbNjuTY3N9kbL2O73oqvWWg2otuNf/l9qQUCKGucWKe1lKPbe7grPnS2jnRCtVJ
CB/AI00mopXV6fUwwm2kULsMZxQE5Lp/CvVQGCvH/akiqQysirSu4DFZ0Degi3sS
9IgkBWFzH1sz3PaHcKfBl2nJfbb32EQTj6YlSKB2sp2bYPowU7sosIbCMbU4kCCi
cjfDSZNZjs/iTQNAA4MzDEav3F0yeTQCWuWxySKxx5xi2onD6Wug7xmQYhVuNHwz
roPidBu2b9V8wWxEZ3nnrzK81jqDaqevjQej/PyJYgZWIEj7q62YF8x5fFhs6kkX
8eQeo1NALXKRB4fYVnAWiZqprhR7plH3Xexvm9SFuSGWqcqQ02VMKmHBJOm10ibq
kZ6XVgPyhcvjbCTK6wcXLXtRdJFw8C1XPCAoSaDPiRaS+cfduPwbLlQt0+LzXTfs
9IUY4qkdU6ViC2b+rkNKLaXV67PACBfTdd3JXTG67pEAY1gQt52aWI4/FTWX1tO0
ZjF3bUNRwh2QFsDGsD+pkskP4mUgrW0c2GDnBbLZIPAccJoo393JpLt+JFA7yniR
xgL3FnpuNeAOLLjRIjTZm1ltFBA91znHgvVKt3jv01SdYPs15S4mBdPXTSkmcN0G
VLYp7J4SVAqiPKOlXDYthCWPnAzlDwCQy42eKfsBAPlmM76CFUlx1IIdEJ03J2uK
Mln676rb1QLR+gnUQIE/DIcSKS+2NbQDP2ixag+fhfwkc1k7umyGhfHUJt5tdBtr
wb1I7YuqjOqDT0zSIcxbEAMDDX+P1Dyp9UtpvqonQ/5dZb8cHDRGZn5DpLYjy1gJ
jDLaxGSHQ2yHHA+2CRPoDo2RoACBQ7m9dFR/1EC4Th39m2ag6S7sO9mC9NtRIvOB
P/nCya6/iIupaz2ijHoMm5q+mNFuhRBVqVFgT4byTUoeLRxL1nz88DDfZRzg5QSP
33NfavuB8YhTqnS2g9nKaKJbWmGjg50bhlqR7W2KyJZQjtMoxpCCX5xNm1BzKS3S
k+ObIXCz1fQ/yv3wrnmDsyJ6TiUd8F4GTvrZrIDP5shtRBY0S9Qmzef0XXvuiIrq
CHxj5d8nvVnEqju8yVDLHJGnDkuY806BAxn30ClUtMKd8BPahBJrmlVvMkKtrQa5
Wu5oQZaVdJBdH2vJ0liGO6LVqOkkSnnQ643i7cO8xFh/KhSDMYs8Zf0p4lJbFRhs
UN1aJjUJaaXXkGhpUwI3GbhvfqB7Nlj0jLoqAEB8hm2lhRKrJsXPqg5Ll/PWJdvm
gzdA2h3WvGYIvTVHLI2f2txQ6/iewxCuYygaD8m3RZxHljHaosGDvyjTEFgPUkXw
Ix1s3KlZL1o1z9ZfGm5QhjI7nK/inTqA2/xWh2RDHL18R+vycZPz6Csa7k9IDY5d
oe/dGYV7y6H5G12KT++yCDVy/L9fjtdc/h6LDj/mnGf1cAxSxLdtXEPmOKoQtcrf
e/RQs+yoNslVwBkIpcbhiKEWQpYEEhTHcXZl25gp+kBCay/ae68dqMwGEveQb4IL
cfd4bCFTciXcAa/Eo2Jf/A+8/xoo+9gaJPj/FbBiNe89qu3m+jWoL0lKnOn+Qucw
ry7q9Ukuacped2QASygBQIrHKtb07OK50GZ6lxDgQOzhlabc2dfmtjoU2iXrPRmx
`protect END_PROTECTED
