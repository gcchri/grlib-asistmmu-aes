`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HJC53KPKeooqwvYJ41yxKAmtp0QlglB8yCKKLfbB8v2PU/wdDtWLBknnmvjawFC5
lqEWN16dxZPIhP3wkAFbyeoKRZuMbLcsxVGpctrqDAx7I49yhnvKc2RmC02gVqlA
JEZuN67Q2zW9SxwN9SCyb3xZzUIaudPMSSEURxHutj1Vng4JXxGXqD2E7MNvMd94
7CKNzMKO5eBcJLI0iLTrPsSAIDeMoi3kFIKY8i5gsGETx0jM+2bsAuz0x3D8ziYg
SCEsv88h+JJq9n85lJMgs5m7UiuuWZmySFFE9vIHV8urT6cNzOmqtmHCgE+snrRz
bkkICZb77GSP/N1dRrn5Z1uWbkC6paieIcgNQHD5Ag1pPCh5k9VO8nHOSde4WJYX
cAL8e5IILvsNGfIejyq1mroWWbMiu1hJH/Ai46DNMdvOrPihTfldwAQitMUMjaPB
VEgDlCX5nB6PLXFLLLWuV7rCfkXfO5bRCzHBEN0/lvi2pFroZLEBK0MAmC5PDy/t
vnpeNiumWY5PcbxWc3DjPQbxaL+rdJjFoDkP/zYfELv/cRAUmk/hniDp5cvngSde
/QhRoYXI8XH8DMMKGCnsQceKNKd9o+yE58PHxnpdkZtG2pOEqnu3RTm/II6S+0F6
sJuiTr5o36EXoCW7a8mULzUaKog0tB5+VLUXJVKpeQ/u5OO0iYeaKX/ammyqqHLT
i3C3E2LKrmFn3DgIDIlFuTmktgRL4mS8jEl6bIShf+CBMF9vpnWYDK1WjwwjaWRa
EeNZgpdLMiH/yMtSDiza/QgGl3ZQz7rOqgA0+DF+vD2tfYxnQjYORr09FZmV+Dkz
SuiqjnJzUe4CIRIJokYrSTzLsTO2/CQMbpzQjdyI13jJGv/H6+zSf2P6nMXiohX+
crHDrU92tMAJ8uoEVvxxjlQzVU+Cl1bSshL5PZhaTBs=
`protect END_PROTECTED
