`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oNed7AyE+emYfCtOQPri5F01EOFk5fgGEULqSX0e+K8jbi39AXhtFgeuK1d6xu+Z
VV0qaSyUC5enHWzXGsGmay28+xsU1txd/HcsSzHrnOMrCxt6ReXsKgnu0NZ9xKsQ
rGUyOMiYP1QDR/J+nK4xY0Vdk0Kz3M3Ly1stdQzuFSH2P3fx2GE/+xCg6xTulOD7
+mp6PusRnZf/tmKXdkhG8McDRs/Z4uomI1ImrSsbY5kKoMZoot+op1KIB1PSqWeg
mh/OPyarw3SzsIJasrwXtPfUoVMV+W9e9hAPNuqM/7ryjD1Fbd/5OliwI/EREAfS
NmWL/i/vGiaIalc41/6zkw==
`protect END_PROTECTED
