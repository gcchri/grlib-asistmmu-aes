`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bd66CJfkGPVqYf1IDx7/xUeRViqVHipdvn+3h7pOm5pFqU8LL5pvwMLshMKeW/2O
Xmm+zCDmfJpeyZYc7fxtHcdryGahNYseWDnrwr5Nq5We97V0MmZAcF3mBbzr+KF8
wDDeP7ThLnnqNNg+8YzRaZLWPEQQfKhaAE5YRdIRQPOs8JCzUhmrn/5vLTOT7BOj
7MtaUcR/hlLFX7/pXWjadgxxX9ruPIPN1I6eLjb8zQDT9tn6Fw5f5+XWDgUiDfCA
l2H+y+HLCV/ESpK/gXUJvMGpePXd252U2NN3EUyQU/1KDJbLQpG6a0Bex1MCIuUD
Ut66gErE7G66SoPhK4jcmo5rmMgUY9DWJu46tSwA75IMfJYolJGWVF8SWuNhj4yW
NmFpBF+Sq4a89cTJZXQS7OMlf2xQK3CPA0bOlctjW5h1n9UpNhHMGdaTFSfl3h+E
WDESxlN7h6nDPi4V3BidhBFHOI9kwCiBAjDvribrazPJwE0A01ihG5GxzY7Q9gz4
iibB+6MwNcQTk3yshcUJTTEStaMnhMrYKq6amTZTQbiRBRFF9NL3zvS/2naWUEWi
LGUG2bQ4XwjEw5x4+o40v2Oo0/JE9YSrx8PTB36iYx8Uk1qX2xx5nyn9UrdEzAu3
Iaq/85dHHV4wkeDwEBqnrGDCWMB/myGhRy5YU/ihVb8q67zW2pySqAQ2dm40yDBx
NkeY88ul/Af3DEfPvvQQlsOCR2+ubsz36DPDm/IERiAQTXz8vk8XaHJE2ddfuDjZ
BxAUv0k0+eAhTp9FTn9eFA==
`protect END_PROTECTED
