`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DDltP5uqWEF2BfzcVPUzLm9X8YnHxKMMVJlx4EZRAAwg+UqHb4Mm3G+4PtvOgjhr
u18AIm3GTupremBNbPYpL67QKphMBkLFcegl72wD885yhOBPCfQPQTBwJ3OFG5+u
IlPbFDzsGQk8G+oRKEVzlWgaa1oCxvXfNcKwcefOsL5+6ju/ihCaO5+UMsfdm9y0
M+kwpNCfO2bdU6CkzJ1ViTDhM/Z34uAD6hH8Oy4kGOAZ8iQi0zmcevOBPsu1KHXO
/p8hy0UJ2aKlb23EESscZ2/zbB0n4AQ5bPg7n2IdMrkabwvH33Cezw8d9xGaumhv
ohAte69Y1I5lHc49/JGR7+WByREY5PrPM0dZV9vy+rD8jXa2ZCQxj6t2Vhb5yBhQ
RJBWQHJY2hitxoi9IWvlLBo5bnyXR94EFed0GoBlix6tNTIGL/6SePt0NEZHvl+k
46CyDI3AbjJkeTeyQe5Mce/EEXNbgIGrJrtFcV8M6Hw1teOd5kw8D9O1HMFQCGKw
WiJQDWlZ/8asfAbvBHz5fzasLrT5fB9vJFh7wiQTRwSZiZJKRuvH0NQoMx9HWXIi
9WZXGaNgFZON4JpDJHCOIlWsHxGgZG8oBbVkCk7HCQUwE601MeIvzh3tg6FyeyI/
xdcMe2h7xV00tukLwCi2EBQOcZWLHJDqF40wmX92yueepsRhHjPcea2g3C4UzZzt
sEQ3rb//53ZyPhClrKTLFIVi+3P2sEcvhN8htknuMQYiUpvR9SO6l98Ux3cXjLbE
B3SgkKVFDGDtGVroO95q4qNUGUVH1M6bXxABRtwluKGUsgsYUjVbiSdsYYzR00+n
PGukT/CmR1CAtrcMPW3U02eBpxvBGLHOzgu4aRbl3VBtjOJ6xU+44U+DpqwILEbB
RJTK9sH+GW/lJPkKIcjy2yzkmmvYwzFVH7o2cSfWpAnF/y0MnyA9wtcthBQ7bpTS
rFmU4dI+OOGBp2+74bnpohe7SUq1evdwTVQ0FFXuTx/7jOMzPqWR++C7ME6maS5f
ulXaGHHzo1Lyn8wfCOcDIFDoprshfYGu+DkTKce5UE9G9UCZB4ieW4g166UxY5qg
8PwU0wr4FXup39t1mC2J9U1L4UWb4CxQXQkfgdUx4zbczHQzjp2lGybIzy00+QFK
Nt7D8lR077lgvi92Iqrx3phpzcXZPTPy8a6ch6u5Eb92jGWDBEdxZom0orbwBJr1
V7VnRdh6ZSkDC+XkNajjQxKbgSa1TRKQ4G6mLupZo8+koqiof31Z3LuKPKi6VlLo
PT6r4AUcvjZcaSp8IKjHlchWCW/LH5s6flJr0nt7cnnMcmxZgbz7Uv8BIVMxv5Dp
e4wgibGO/J/urR2bs954BSzeUJP0OIuhJJX/6ntkvoPbjgYUiPQOMt4o7VYZTCr3
D8akiJ3qjOVU9Nk/STSCTRjf70egx9WPXZgHVAGWuMJoRQEznEQsiRCzV+KoKIUk
DK5FeCzVKILDPc3Tql02KROBxWt28oHVOcv5f2V+38uVGWAg6TLUaugofBgD+GID
W7dPb5N8D5T1SkyWmmjefLrwS7og8pl39Ujef3KBjjGZcCIe3a6XwHRthgjW8YQg
gD7nWybXkwlKOmRrGvlo6Xs9Kmj0zik9Ok+t5DQkiTO44nXxEpMCiVS8GcGSWeOo
2XZ2HKOTbv7I2pVrjvFYFG7beyQN5WH+L2zVFRmgfKbRYwHfPa7e3vGyyDV9s9Mr
iL0GpNK74xvyJNFaq6NejJVF/RSaMbFVcNI1ejdVD0pncqXuPzkBJptbLTxu7hJr
aIYe5iSnXunJkhBnQhlMPt9a+QZsW0gKjk3bn/iez7807926Gl3cfIEZb1efhzbv
ki1mghVZBcCCJFIkvEJ2X+twukTl6mdntFLo4En+/c8e5fzFheojJIusClAU4q6T
Wzyro7ay0V70ggRMJ3HlRBaWFO1/uCIGKsADj7VOI77j84DJjNnkBoFhsPGkK467
/qj32s14RNMWYq6bwYnuJ6T3UU5Ri69Q4hgUuTILq/sFFatvY8uDhcu9X+oqyFIp
8Jvmn+6lqF8iopN4iDknhzWZR4gQSRzje54c0hSt67TclhDNTUKgTlRvkclQdbvk
DmqCy6wYZnI1HibY9NJaX7xwnGE9op2Y1kIJnkr1gyvsOJQi6/CbPLUU48p78kXf
52ucw7UwK4rYnufyMqwNtajtnTMng93w5EtzPX30jAHODfKmzX6qBBNrCaBDUoci
ZnUnRUmSso4rFOV/WasB5POQqon+mTDLQoPtD5iU/wt22gqETBfDgId8Z5gNYrQh
pikO+sy82zALlgx0n1FLK4IND6DzUajNRrqc8ICORv6eeWEcYYZnrwEq+1KzzyQE
C1w+qiefzyNsSrSlj/RbMyhpZ1+CtfesXJxGfmMfZ2mk+AVIoUlVFMvnC5DAGwxe
SjvQ1WxPQYw3SxpfIALH/wYcRfvdQG/1Xs5x/x4SzriRcVHq7Po2kPybuWksAbHN
O5yOxSXYboTfTyjNEIPfScCaaf+/RIMPTCLPFYH13KM7UsA3qgkmxRGNoF/36AZQ
pIF9VwY4W+urPPhNEB/WdUynqJis3sDRDm4EtId6mD3ZsukyPEJ94oYmdnHa4CHi
pax19vspWG8sjKygdCP7OO/rOnI+JxB93sYxCaCf50bFQaG20iyi6VqeDV6OaPHf
Zrb8MV9etTsvPMYbpGF3OtBgaKNIqsOhSuDCvgkeczu6h4Gk4qYdKYHIvOzZnAH3
jPH7iLJ9KjJW909fAuaKN/uQjEY2iKtDECgUUWxpizeZqr59UmwRNXqna0og/5/e
nb6UfcBU0Dnx+U9QHA83ad0UTU4Pp59vyvxYH2w5vwylQli87tdKNRspJspK/N5t
x7A3gBCHoxHvYrQgUcfgE71MHlxxq5s0X+wvCAYFWMlMxQIQnZwXRRTfQrKj4jKD
WpAYGfaDn4drnJ9zpk2bOurJ7BuD87Gqh2T/00AFJzruiju/vH5tTf57UNODA2dy
rWzpQeig0FRR7YEZJ1Eys7TXqkzBxkScqBfj9rGNvTxuwTDhRvZWpTSgoWQ63d4a
WthSLly6m5JGaTqgUDqvovGKuRSfiFtdVOtCt47yqhcw2d6rzfDzTg5H5+mA/vNn
3gHyR7Mn5gwwhwz2oA3dxEoLZEc1CegBL6AcwJKHCyqusnc1fG1rYDGvSwb7ZOOn
lhEIobeDSG4VtjP5H5bGPRJAo9N33WUmkV2Riz64ywU7nwSyEBdnUSlKF6ZUTDr/
I5++bFCeRMxQC1eeJ/4TOInB4wu7kWE5/kHeicxoIMNWMdIM3F1TBoHd0hG0nfGJ
n+XnTrZ9QraCdjJydlu1THPm/9qaWmlQyBMd7l2RmQI/JQqXa9NtHqIeSq9p8cp+
c0Olf7GVfEuIaTVfhJz02WR2c4oLhZZw/fB5zQCptgJeKaYz1iloFTSltZyV7tlc
WeLbu/BaVjZ42hb5eqnjpt8ME5BQxLVZBa4jXAMM5mA7J1F1azd6MYA18yOZn2GR
4bTq/8Q+mVqLkhbpEoDd15S6+Mg/6kNFzEYYkkxuOCfJXmbJs+P29bevydhS6Dw7
YbDk3cnlXKpMoUBUFMNlcimxRRNfHQdMj7JV02V3Ei+aXUGCuximA/rIJOHFmnbM
gEGffXcz+hGDfxocOzS1dn6/b5M9mAmOH7ms8zF/4e8ty4lyPJlbBB2b/Rl9ROBm
ysjh42FxH5HpwGLGg1bXZ1ySsFexA5ckonIamtz1FW4=
`protect END_PROTECTED
