`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qPdKVY2FTk6uVmeFVV1LWO8hBx4/MEUFIKibFVd2PiavDtxyq4szZ8LaCoumCT3F
yGaybjYGCof01G62qii7hnLq8rzZQgMR6Z6K4AiamrlEzvoTEHmjxk6og5lGVZzD
Gafij0DBhQ7I9gCyo7ZJIJ4PQ9rYSkxDpdrUAPB9uFK08PdsCq8+ce4w/iJ2dPXi
epctoUYTwl/GpBFSwk/81Xi+8wpMNRox98us24/48e8cQYA+UXMS9g0bxEuYhczY
aBsam7NpkilFgLaEU/39VFSh3mUuS/DcLXFivCQNcJQuZZvM/UNOxkSXhziKbDgu
ImmgZT8WPvAUEf/X2UllS6uQQkyCr3Tsin9YNvoYGmr9w96N6/Ik7iifg+e1S6EC
JD3Dn4WclOzxztLNmcrV5F5KwYZfUnaZJSdlDtO2IXc39F0Dl5eOW/0ygf8Fl7Ow
hZrvsvLXJTcf9VI5t5K4oC0aRqeqXjl/utv3sJUN6lSymGBKhi7OLsISc8pQDy+b
MTBYuXDo13hx4AJZxhuFro/hZ6uopMDMFRRsrpTtZOCVEG8eCfr6CH/ELrf6q22z
pSQ9tRp4nleNmVQVAwBnSO/rBazzpY2g/3tDSid4k/jHfdzqS+LyHT38SuaepmW+
O14aeWThNxoEWMUQ1CyK2Myl/4S+C0/zAsbmWhuv5qIkuIL2lbF8f+B5ppUoWn0l
/Tb0olvvqa5vXpC6jIxX37AU02kdw4FKK8CmaBj/zL76m+k3f/QIAg7I3z1HQDjG
6U8nu5Mc1rYx+8HtDA4ruiQNWagKjCCgei6/9SBKBNF9ZCLKgA985O8PZz2HxdC+
3zHMqxnAQ6Wjpd5M7FBPI340wcLGLCBLLh/4/3XhR7WTdC4OdvbLNlJaJeJVv+3v
ZejVwa0Qxwtigti56YaYfEBSS4BvlSCSarll1QnIqjrz9LqMXe1aKzkz0G857HD2
S7lr78z4OjL6rucBfiNoIkD1fJFDRjxodyubddVna6LKmSe0gEBMEgFdt49a4koL
gieL2vP44t+GaD+2JYom3lOe7wrwkUxIaMYAJXNR4ns0qhxmfqmkFSjbLJItQI4d
wAHG/S020jwd1vLhSVJ1Fak71I5O6mB+eRRdHM0HVUUpBO8Mpd8A0SyTWxUMH0LF
wkcw+/ZR1CUW45qIJqOEqNoGf2VyV6zNPsvyJfHX8BcBMT4wJ4F2a3MJk5ql1ZH7
d1WU6GoK613VFEVzIfH5B3ze+YFhMaFSdOVb29DV4qpoxUuXZGtwm3QfiDbE6vLh
3QPW8GDJioUmtnfK4juJJ6v05yQAiCIqPtucVc62Qk//EQNYbcEV5/iekMzY00b5
dy/bpnz2fz6t6Y7OzgGVfcef67WFqOhmOPDR8H9NpP4pnZG05vI56qAVKq5aCTy2
vovLjLk0TjsZ5zwHymAAb9ngiQt+nyfc+0P5eCbFa1ePIScax9QOlkMj2jf+USDK
rSwg5gNdBXU3AAOksj6+Aqhng50e7qP1fK+AQKWn4kZGUUfwR8s4qf4URnhqUc0y
6ktWpyep1v5TsfmCRSrcOYu3eXCXYGDMuZIFtoJB+cR3mgUWxIDi7bFNg/Sg2coT
OqWNKF5a8l558sm1RM1ItXUQhXw/A8owssOOdmgerxlT7hSp7gCQHUIPug4yMVOY
901Oxx6nSHQL23v98en+77UddaIMhMSrgBdgMrzkNEEFBufT1yIRHcXN8Pxprql5
uh/AONhbz3JgIsSCuCjGK401BKvd9pwxIE0pHUiNJLxtJkZebPubbIzoNsEvL0g/
BY02Qu+z+a4O0OkhtlXeDVpPJiv9eMlb4xek2gKYPihd/83D39pfxXXO7sS+Ekqq
sjvDtZzhbSfdyDoGCiHS2sgnNdxIfvVdegvqpRb+rBDmQt4jMUlpUwvhpx+MvIWX
hcudkunGTbOUkV0BBWRqBAeKC4BJFcR8jDKScPkUHJmZIM5+abme+smO1crAwT0i
Dh4zaKE+FrD4yA4csoy79885PYisWqdbBrtdJHmr/zDedDC2vyZFSStUR5UoKGv9
EGahGzCUSkfsppenVDqu9ve8SdbShYUntke1eN2/93HK4CEEXmEk9Qcyd2WNPBL2
e3AXyG7CIMGJlxsY9z4PmSGDooJbATaAOIahfX1DtIre8ua/NNJGFENXQ7vJ62q4
IVTDz8rc1M6bsH7MHGTtM/HhAlJmHr4X6AuWWR+zfaVUUvLNQ1C0ORXLodnnDEJt
TjOv8YL5XM8ZF3GUxsVpuenyFnfnsp04cEsi05xmLvVlde/2ILeZiSVqGfDdQ/d7
B/inSdcLVGVocgrw+K8cLhZFrKXCzW8ujZ+tPgMnbFXzMtmv6ZLRQTTCYF/hPFFw
Xd8MLnRlm2Gb08RkBx5j79n7j8a+UiePZF2LkPuP7avDBkxKkBJaCMBFwBIUcFj5
nMFDsS/rmL+X9YtCjr44/BTMXjvapgy2IwigC2JjEmGdtidl6Jn1ePG+sH8EY8vX
6Pu3S7qL89lKtyHyLNaA/6c332veihbfKtL0iPZgLjWUDAOffmPTs+vcXuxdN7qW
OtTQt6MdVgO/FVLsa2Kmx2DMKA2BG577YbKvEd8EVkKVjyN7CqmBGZL8ualKiJaR
WegDdUFcmPgUdwInR8pKwu/nyjc6D+6KHtSxU5grLvThgHKVYat1SflP8T5clBAC
/7AP+yCTllk8KDOgGWBXoqPoLSdQ7oU2smZEqkkYRcYs8oLVelN51RGLQqUI3qWE
Ry5pYERlRrKxI0ybxA7WXBJbe/liOXtuv8GtfW3fuQxYPn8rlvuFfYpOkzvMwgIP
lpJGppb7/rWyZYRGkxRFkbO6qtGOdWEWcxpsuyJ8+kHX+piV6FQiyA3SyWrcDYaD
Qd3iXnZZAuXkos8KHo4gTMekEAndYVOj+OLh7vPouaRz/QglzLGejhl9Ly22thuG
PrJfPVExklL5/NZ4KYeMWDMTiEscrXeSE8LxS8Ybc6SGV6XS6YTJO8BinjqXTtZP
/yaPHl17s2t5twVlMAGlm5/PYe0Oc/2oxGlwZET0hiE1sp9/BNN8qb1i+NF4qGaj
8nD3HZd0EXYvcbrgAGpUKuc4+gp3S8fxAbVuv9wlo3bQngKexh5vEzehoawYQhcl
i1QG9S1i3QBS8DNtoqeO8oSXZaQsdbyzf2+Wq1HZiIsSTje+i+bIevH5ZMhZL7mm
gJ1njIGFhCm2zNQU5iUSOpLrMo9mBQSN5CGAH1ONZPFqKDaw+GMJo3RW0bSHtJfr
rmDkcFZpoG47Cxfo1fOG/qA14zLcj/SgG65+SsPlVQ0oFjDrCMRvflE3aV60Whzp
vWjE66BSEH9DR9ClxPeolvfasU/+uZxtr9iTFl9RD+He6uutBiqegLEtmgc3QUd8
IZRF4HMvIB20gqEK6jaXaqCpdtM1OtHHS60+0xjSJrao1+ycTjW8TwENgtCsxHPR
VBx/KPlsAqyeDQNEaYRxxHW9kd8p2BZqgNhm2zJLGxlOMqFNuNarxTO08sfGYoMZ
DocXqJB5dNliUN4ZebNo01YpleLoDHnkFk5DCrnGXmI/Jy+RXhs+0molHJdEcOjH
nmyKI0jymUL5b1RGYMlrLKSaOgHxEP6kZL7v8Lv4a5YNxGJDmh15476pYMk5fkt+
V/niDNjrfEl/1M2y7MVfdowyLpN75jBz7WfLIBTyW68tt+natTQgJoqFm7eX9sEH
tQl/vz2bXoCbKgMU+ntedKmILCKGNf5Tv7o0bX2oz7+w3eOdaDZ2meV1uG/pc8qX
K2wc6USggQkG/U79bEeVEeCyOsnDqFAYCTpIS3dG8d8RSddcNcM3EEiEvvQr9uyS
BfbdlOSGnOGTh0FRfhc5jnhT/HkC2G53g+5gosj0qLDM9xDjz5ZrceEOTWe4I1rt
Bg40TdtqnrN6AfK8G8WOJ5Do6oafxUumutZTiCGGrNnvcFPKJnJAMJ71mljz4N21
KHE60iyFqaB7AOeie5HiP0MyRRp0JRVO7ziw1hBH60oJF/KGtHSjPOdp8KFEq3Wh
FFNM6p2DFvMNy4e08zBUmkxsooVvEe3f/iWADhKEQ7N+K9vYo2S1TGZBwOSt7Hs6
/q3rE+A8e5q5HmUx393ehqNgOL2blRXYjfoCxIo68kv/5iqmqAAnifoWnXF53Kos
JxkMHZbMB8i7brNNAS8sKdX1oG3cMmrdHoURbstgZnPAzwW1wWca0uj1Y3AYjOUl
/hdiJ+qz8IaufY1hTptoOiP8jf3YQd9wOXDwGsZN8gS4waPlRbOIcfysJOCmeIzf
2biEf3vyiIIBxuiu7XmWGcDITI+EQVSKA90FEuwtWSShQjLWV8MTj/vYy+Fpb74a
xobV/mvHsYvHOhNT84Fjo0PtMtgtYoSLX7OA/jX5O47d5oFM3umJJwNSFNBS3Ob2
6es9bzu2f/7OfSfLdadTZ5bQdJEyIDzpGv4kn+QROsf24f4ZphHpYt3or0XyQ1PC
HMkkiH7essXgDI2cB//WK7z1FLFO33+11OqxWJwql7d0C886ARpOaX+G3vLmZN4w
No55YncJ/MBt43h5SBtqJ+znOS6IEbxehedXSqVXW/xomc3kg+ES1A1UjcRb5/RQ
P2SaKkziPLix5cg0HbOJiN3sRO1uzrXNfDTtAVEBbek+E0jr8i3iMDmyz9b7NVPT
iLkaOA7jEWDNyw2TRHZAmamU4PmKLKnDz4rQ5gLepQM1opPWBL7hpf5ORKnlDLnr
2t3q4F6KUEDFBVO/YLFw2e3I7/+a3MFLfzcFfU/IKPvGXp3ouX++gSHCEs7qV/hM
DDJnJhZ6gUxw9ogvKtET+Egx4HUK3HuF2x2Gq7GBq7EzHvAiliaB6R2esJOXzHYP
PLdq25tMNWu7y0eiTV90I+Vvou1xYHrrBEvVOb4qK/miciFm34Boryhrh+JDaDOu
0iZKJXT1uc10cttgbqtaNTtEDVeJs8dihbGzQOvfOvP9Zk2yKwvNQEk2pVBCO8hG
aIBXcFQVqsDFlNgj2OBSno0Jd7HyEEli+hXUlBAW12LLRRCXgjXJKQIbqeITKo+Q
H85Y3VBqtbOOlORf4QpW08vjY/ADhuyV5BTPAcvqU4l/kxnCpirkFt8nsVumwX6W
2F+lC1euYkhl/INeAfsD96h1yz0ExBjFkNE0fGFP7qeac2NsPKzzsVFUoNkcI387
O5RZREm3Et6m4UzE1B/gPpQM+8njOLXZhGrw7KvOD6TpI3bc2V97X8eK3BtSZHz0
Q2R0Up+krONLZ4I8jjBhjWceQq/8c4lHtfj2mFT3IDkOCfmMAwOCtwYge/r05Fc3
z8fL5MnYWYkmupWMsr6jrBwyXWdm7k2ITZrB7WukfIIvDBK+mxyGLx0qLApndLYK
pIZ9xC3ivmTjPRpo03QH6Ztwjt4EPqtQcz/uDxmfPwccqgMt8aLdJ6DuHD7pEUft
22M6KTiih2XEhsZMESpZHzJ1oUhHWc11/mwJJc/kpXMC/ClTutH82/Ch8HkHjYuI
jMObsZ45qIo4aBbcupMjDYpYdw+b2E0Y2vo6vamXH5aS/jpynxvU6XONJGiMX1NA
Jvb4/ZBd9E+sLB924lP0o3iLWyJYHmO0MCauwSE0HFg4W9f5m958f5joejgtqJGn
xOYt/4r11/9UnrY2cmB15F0tX62ochMhyaAI4XaN22jCU2eq6ORntj216a9g/E66
wtl29wyuJatBdPj0IPmHmgEiD1ywdLPUsifxy6mHlOCVVt+5EteaKFgQRIp39BEz
uYXPFyIHERN9QwSv+BqpBpR1h6U2Ff9U+0K7Jypd2McqKUvUL5jOMEj0mUqZrEMV
b5V9DxPYbAyk6SPbodyhrbgABFjYnWBGCuFoCZHZSwUGwDEQ97ZqYWaEBjUwOEAX
pIDbJDQ7wqnZPGyN6Qb7uTx6XLtfFrNPrsGo5uSweQCvszcWqn2pzFQ+0+KZoZb1
JTbsm5T3+k/yrZJS20c/Y+G2b4TIaA7GAKbt9EAydBB52j7w8RcnCNJ5AdTESAzQ
LsQmNORl1fY1coTkQzrZ2lzUP6G7JEWOROCbzYeyW3ngDnulTqjtFgoOJA0dFK0G
YJhZwyLeI1pJTp5G5PK2Nuxo7xAdrylt1QUQJDIeujK87bXVMt3MOm0iHObYyvv5
Q4LC0JRjOtOVtXF9KFh/8xgnf2F7voVfNHayzCCsRjgnn9Ec9tgTd4W2M08yo4Ih
`protect END_PROTECTED
