`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1klusn6prB6UagU34lfVguUIEmdbcKJZx+FBEKi3ubwPBfXt7h9yc6tPGrvZPVb6
mqvVcC46NaTHRzbt4/PEX+C0VREKV7lNhxgeJDRAqYlYAj1vNKgRFuKLajcP3MVX
/mhnT4aUspliAiwqsI5VbkYLdPL2A+u703BQK6DfvcTcoEKBCKmtmPRcpZpT+8fT
9cn1EMmoGvDhB2BX4eKmqRNETbRYzqTd0i/ktud/i8/IZZo3lhW+pA1Sq8ZQ5UhP
XyLFNwtNUd9bxnIZvuGcIAZEO51UCDmS7wOR/hhqleNZqWNqGZp7Tp+rre+Uhzsk
D87f/0NfzDADEJ9y3jshRww9s03irK3KrkUx+wUkuZs=
`protect END_PROTECTED
