`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0CwrSgCM8icyoSLbq+m7KcNCDHMZ317jiRrbYcsFSmi6vhYLn2p9Ar+fk3U4hLeO
rBs1hV2DV0aCbcJdwLcc3qsmTYPH1QKIq/xe8hjgq29g4ZcwK4xXUpFWiQ+VRP6t
jiHarBb5Z4ELUVqGJZ4LDnC8rIi6nnhc4iaLvMpDpcSKROsU1rQJ5nQPkiNN3m+e
MbhBfM6KJo89Mk8UwWADN6UDorQY5Rnx+oYfwXrOu15T/budl2PJoaNNwDLVgKVl
kqcJytG3NJHfXLt83lRRPKwa7sRD7I3AGsxQH9Hlq1DTDTTS0iqEqMMMzesMzEC1
wWCxWCCekf3OkgjRKn4ZBEdI9ITbrM32FEybitgFxkbuOCQn0YzhiiaQQQ44XreE
DnnWkuzT6KDwVgvJ0e5f5p9zvtgcSjPd1cdwPJI4M5SF2DZs25RuBMZlm/cGA7Zc
OsgHjL+xBgg04YnnlO2cbnmOGH3tlkF5On8d3PiWr3DKgQ93JUU7sI7tlJFU4pef
nMSYuiZc2/HByxh8MG4j11I0QsbVmpNGU8WfMjzgueu3frzlKkHp/Stjojj4W6BA
w4hYbgH+Nz7h/5nZiHEAUs/L3xwepYPyHHP/DvSBDSs7/IhJ2M7X26BhJ3J0mJAU
pumg7tbjZKDK0COO6I7lZX0LG7hAihfZVXUgpuYMRJ3pV2UClgTcm2Dv9mJa78b1
C7HPrn1qlsmpW2QrDaOqxg==
`protect END_PROTECTED
