`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i9aHNxzrw/j7Nkcean7YdhGlbMLzxHcafb/C3mBBAwcnvAjYPcvWZ3zKQM0Tclsp
DLASPzLpbMt/PWtBn8MZYw/+ki8uWQ3ebplx8rx1P0QoqbMENt5KRtGl9gO46kuF
b+4Rqv8h0ejsSXjfdXawzn3jYpt3IOFpN6SzmfvijGfB1fASAozPDPxL/0RpQ9aJ
eddobaagv7THVkO5Mf2bC0/BSOlrW/Al5SYWB5X97nPJAKmvUKNh/83RpprbVxgQ
YJCym5zwW5dtG69swDueILL1/pw32XWqBvf/o1ZJz6ycH1wEOqGMaRD0yYhq9oag
RftFWYyXbv/YLIq97nkk9LOR4Jw5WA/Q1jwUOdhROSq/+URjlvAk6SkkilZJgwR3
vi5aQvv0LtUVRqRFfl54RMUjShtRtksIQPokYAHeOzsABbc0cW+tZUgq70VUd11k
gBT0x5SJM/EEtTqcCbPz+wl43tqCQ4nZ8hDUqraqIfBCdyPFWBSE/0Ih+XiYGMxL
Q+Qsidix4y/YYvOulsmjMEdPWVJrZpWVB4vFCs1j4+n4xeg+a0AqeJErrci2Ml6c
GPrkLXorZ+sA4Zjyu1DKIIea7/uAZ+YfNDlVEe2VUuBnMIE6PkUjZICbBhp+RljF
GYpGdQpSfrYA2vcjM5V2bbFNY7jhStsQ7GcP+HB38EkDqtMjcOyBKjvY1AxzgbHF
tgxROhegg9AAmfWvKiWH2lEOWPv+LrlV1sdbQKEDP1AbMsDytk/eMN8FeIXtMm5L
hyfcI2Zpi2QQFD7YKkzVKubf7bWromfPf0J492yPU5JeoOMU9npiMof6xQWP+E3r
LsHe2KhZ0kk7UvBuv5/w5S6yft+fwocFs2PlIvCv29/h18zEboGSvNvo09rj+lFT
bn3etejO+8+hxNDLydKo40xg/K968xpulwyv72J5hgPSjSgiuwhjk/eHBbv/SNQa
5fOughZKm2kHF4IA2MOCJkvRgNuXaQnry0MM9GhIvyGAUla60/khTP0Uox2aM7hI
d+0B0JyrCjff4Ww10pOLeyDJvOvXuy1EnYFhecBdzHOiQh8oUpOf3i02yze+F6lQ
zFhaRTfHcT9ujj7cSVZ4nlReK281QrpJCMeEhsZSQh+te26Hk6yD42nliw2f5Z3v
WnWEb8DhB9GK2/uJvr6o7Lk6Co/B6X02rfvXIKUTYG81MPUaje6/C8sA/XEUARJS
RzPJyGuCfEG7bj9PDsn2UH6SMi5sVpupHHUJX2icpQZJYcc63EwjPemKJn6PrTBU
Ik8EMnnm/2eozZ4xWjoHF1Lr7CApaNPrqp+bn0WyAC1MWKRDsv2JloScK8CNqHJG
9hbJoaswAePQkxZIJtpRt0H4GrANHaPG2z90f9g30Un85VNoNraFY1mOIDTV2P2L
mcFSi7KyPkv3SfCXw3+kc7E5FK0W9lsfdElDOpGrTKY=
`protect END_PROTECTED
