`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sFa9p8HiLKO4EdLu7PgxpurMJGmJ1LdATwFnExErfUFvX/UITXc8RjDZlfehgHf1
G4J+YCFxfHvKaEeeAqHCTL7xTk9aYWZj/giNlcP/KoDBvgIDV/f9uuVDiGuSb7iD
pxUoOgrJKtaa+cp5+RDYQNoQPWPN6XCyuRAn8krrz7NhdzHxPy+O+4BcyivhB+Sq
2YEniZpv6MYQRBUXo1rndypEs+7yU+YOT8GDgxNNn1rPHapQJLe1eaHyfY7btuM3
JwPb1tJXuQOWQ6TBOOSjOBtIwq1orqP6mpuPQnbuBfCCwbfT6oQ3OBn7h1mYn+n5
fgwpXUBdLKWOKgRYHMpgCg==
`protect END_PROTECTED
