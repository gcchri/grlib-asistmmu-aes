`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MJi4mpCXsLucXzMcUjouWoFrsNMhfCjHmC08ldHgbivoil027JWHDjMVbm9nnkl6
+cRxpH6LtdeV8lLnfu/y53Ia97wch/GWgSJzwcHmsVHh1t3mpabnatwNQ6MaUbWa
/F+rceXfLD9ZhZRRHQvFUlmHVwvKXVKPpfkdPju7RnvI/9ocSMkS6mNMjpWYm8V2
cmc53ZXc1B/Vr8Ho3jS6ThtwLsKDEwqGPWA7b2VXvH2ZVZr20uEFb5dZilVktu6U
2W7uBEQlc3v7whX7SmHd6pZANk5hAROFRxDXm+FCCk5apWXVNQsAkWhgiwyGxlr9
8DKI89TWW7R9gzefHVUFFMYuTqwe4Db/Mq0zKKvvA8TH5IoejBisxE6C4k2pXI80
RHGAeRSb+5nKnYwfVKGGO9xWdagZhejEpbQNRLfQgz+9N8NUiBZ1BHtL4mHqOF5m
`protect END_PROTECTED
