`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ehJGtrIt3PiA8pqSk9BjuQaTWAQsJrjNObvQe9lMrjz7Qap5kN8G+n2yvvbrN4bJ
+W4Tx2X6zfB6kiGDCFRkQkxDAjQjl1sKaCgbirwUhHFDCNbKIxGKnO0JLyg7F1rk
RhrVMxTvnn0YzaaUtr4jDeNAMiYpfUQyCcK5uUVR4zsLnGtTWNq2BZANyxO7G+2r
FnV1+c8eZ6ZyZoBC3aYOFaldtX88H4E1uSPjm+c6f8PJUNwu9nUv+2+nBxV/nQfR
YGIV6RYyK1JGlOiTfe5CIEWg5LMTBhJRGekh82ZhnFTlILgkwpcUVpT69vHEEbSA
zdXL2lpnZV5TMY/afb9XUwokQOWO6vavT9ShCI3g+f6nvWY0mDXnBHtFCQ51dcAc
`protect END_PROTECTED
