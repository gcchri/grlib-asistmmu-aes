`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e/j5Y3NNuWzz+xeUJMZ8c5N/Chvv//CxLakF4QQkeFkiVMRvLN17zum3wM5NNthw
lc4s33/jt/RN3BAjuohAZjFNo4GBNJOp+al0r9U/O1xAabYdn+KzLV0cdHGV2/f2
pICilfjIo6nRHNMQEyt2BFz2ZsCR6kpmCMA3xMBpk1uUKJHErVx5QSCxfSB6y+Oy
bSqxWvIjxqUu+TKNEzWcEpJ3Q4/ZljJf8+4yWcY+wFkhciP91YR7ls6bxwENLGK5
ucxciP8vlHIWxYKTv85KCOjbnbbSevERvKxqudrfd6A=
`protect END_PROTECTED
