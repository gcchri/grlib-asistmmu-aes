`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TNOi9EzhM0S3wnrtP7+2a0GprFut2GKuoBCLjHDdiJdC6IPe1ca2QK5TmLaOzjdR
4dpZEHjWAyhmYciF+fRMcginyse1dAtbpNlKZjPfDzk75Zpo4ebHqd4jpsXbRPsY
9/nCx2cDIZxfV5egQ62HU05MZiVaBuQAZBrJpT71iDt0hgiIErYEhALY8lFBnXJN
d3C+a/u2VXhdE0rA5C7vBw==
`protect END_PROTECTED
