`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4+bgI6pxwuR5xyB7NP3Yym4Vbngi4EwE13bFowW/G7x8WnHKBKd7RQ/pOa/WOhxQ
/6PKwIT9g/vKEQnd3Ds75YB14bnLe5cjSGWUefsWdwmEyQdBV6FnQQXBaj5EF1Wm
bluWWQ/FNafJduPElCgfqncHME2SmhXwpCBJ09I3ni9ZUZKKooI1eDrJQvbHnyJ3
Hfk4Trrw8TibTZ1XH5LZkv1LriZPjkT5mtbU6M6VbiR1/J20TsmauMtVwUQeOUfd
avlZYUxbQmxplSuyVvr/Dw==
`protect END_PROTECTED
