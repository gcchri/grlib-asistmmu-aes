`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4S8Qm7uD6bzZCHkZJcw0d8WORYRbTaVvN8a7lbvtP8lDTRTEEJPbxnDApHD/z5W+
im/q3wXgnrBsNj3mOf+gkQd4cAt3en6zxblJeQgAgGT8GZBceYrx8ynSretJ3qgt
86obC3kresqJ6ciC8j1yZJ+PgdJbgfkWIgxXy50O1vE/6QU1qFQeHoSSNHk1tNPZ
YOppu3rytqYyt1j7+oJA4QTwf0z2LTzO+irff0j64B8fZUDH5sclIhUuP43pfZWF
g0QxRK/Vrn53JTVWDgfmr3BJFLdlscuJlPzaiz/igi+dfigBogyAK2CG+E7l2Ad/
8JXS8CqDylgbXvJwzyaMc+gxeUkIjXEhThKmFy709kpkUbTmbYIE3Vu3cZ0RKu4a
XcuZLRjIdTuTgVKRSstb+suO6OIrGxCPG0o35SWBvGBWSj+pDs8p4ZY39xj15JEr
gtrmdc/IvWxRlG7FEx590EViD0qF/jKsajAfWVYaFu4tzgUpaQ5VR8FJRN+vvgT5
Evnm2PsJoeEE8twU8pg0xIJXBYykFrPisXrubO+d29umiAcILmykbIqAK9w9Skj3
OgqgJ1ncbL97u8u3jr/MEyVU9OivZDqZt6i/dfJklPeLmVWQTM2sXRX2/NfAC0dE
HYoG9wgv30egs3OnTpsSq7754yvxDFt4KXZVuDTjm2ATes9WyS+jh+2kTmQcExIn
Ch+Ny58lhBWGI2XObFWrI/fHCiOCWDgR9TdewFRPfnWBExgLyYNRu3BtsqSmJO/9
5YDLb97MlQDopwogX49jtjT3dSkv+oiHG9h8cpbF41Si/DDQis3Prwq1USxjlzoL
FjVYso4sl/Lvg1ZztCwd9yUy+7v2/vnM5e2hTFiXAsYOjlR0qyNAn9u1O67Z/QBt
vnZkjl0yF4dJipiU0S1+wZAFj/Z+uTewFduru/hybXTVuUQ2BFtsyGAKehdlCwok
EsAmpv22WPRbLMomHQF+qltuPLQU3+W4cx+VhcBpRURys+/us3x93TjAYJbry5b+
eU5XseL+LcF1rzdCeTAf/brtam+7ikzOrXmMIxwkiFPmnE161sWkTw0Up4JD2OPa
a2wY4dnZMWRx+doTCUsrXplyVXiGX9nNi/vr8u5hHboA2vCZK3mFsMSig6xE41zs
uzdIs/H+yCq4A4H3sm7Ak5CYSSSvsg+yf0VJ9b/GqnRVR5lxFfIQkyD2kqX4Kr/t
Y5qbHf81Ya30maDhUFQezfHF3NAVFcq+kxdfobjQGivsBvWUA7hZE7wd8cuRNDQ0
rFoygFKPR1MRiB/aXxFMySKi58AU+Tmu0bjuPZHWbpp2Zl1S+JvUYz2iNS8B+rmH
IkDC9hDIotf9hKbNnJ/4QcOk653qovsuNDofSwxuZeKmOr2XUZNSsmbetwANuQjw
XJz9d/VhYPN66JVTLKM0LlSyKZkrkkE1vE0iSWOceheVvOfJnZJwqF3QfA32SKP7
LzLhyXxyQqbkluuMXpB/DLZxepBgayCN3uGZEiD9Zlj8M6nV51kb0NM+U9GW104r
qzeCF6ALhm15jIrI2/FfbzLZOec91mMr20DDzhdc6qf4LxtSalTG/bDtJSAEhPI5
Vt2yxMru+FQNY+3bhxCg2jwJThpwgeYdN8K903SbXOH4cCS5Whjv7n0co92SxGjq
3dUWJ4rn8m0Y3vAflFv+A/r8rm43z2bvFd1n/DmfuCUWsW/YtlU+i5VYZi1jW6Gx
LvvNzuhRVQhVQavASf55MDafTqS8haBoHyM1CiJlEu4TBl/nHquleqJN/u6RUwaK
T3O21gblF1ScXRqPHhyfzYQ4zbxx++AcZA4BXOjI0No4Ak3CIRlswXsciS39jXGw
6qzmUbCSWE9N3Wx8E47Cx4XqjSKIlc8w7GW0r5P9yyicyBLZPsAkISZM70nnbbA6
PWE6UIjqT6wlqVsE/js9unakRpJXGPRs8E3u1Rp7G1BJkRa9Z8ENuvtQPEAgU5ge
7npmyrSJSQ/AtvqtyJAbbBmS1qPmqHTOhL3bVni7uaJryaTkuvgTgTA6CwIwajVi
FmQwlpwtYV/NXjYZlccWKHsQubbmcaleZNEwPOslvtk9NVty/Qj/X0WfE5hp3FTu
jAHvvXEPP1SqwMTQUE9LRXN7HYTlQ8BfGIb9UIDUoL7XcV7L2iSgRKKbGIbKB1Qd
VRDvTjAK65oxdjuBTY+LVVG5fYQlQHKyhDmi9nwip3IHLmnuBLmuQ0Q8St5c/X1+
4m7QDy2r3VSUV9+MhrK4CUNI5sXbsnsPNIFp+yoOdDpEM0D32qO9IHzLlnucsUGZ
EB2zlVkopxcMqdX1QHpYSl1o/EAHWeXfg8Kbwbb+LdFpdBy3XbUh7iyYdWktFRiT
03/RTE9+VIiQp+WP34Sh6Ic3Jqv6mbXz4aaNivkVGjrz++RaWoe6oRe7anie2GXt
CfHgS4YlntoQE1OU+9drRcIc6LbQyGyx73vi77DC21QHjmAcmAHZ8pkF5mYEYdO1
NNcarLT/i13pFo3/uAvYjFROxxoVlbHd+gq1qmVrgUkhzdBX8M0NhF2KNXGwsYbi
JnIH1afOK8XlzqDVplWpIsE6rSiP2RidQRgpk/ChB7xRAV76NRyFsWWco5abfhjz
XdWiY67jzfqkJ5BKq4cx8ry2dS7jwZY4NHVIuDPMYwUejw0BqaIr4FHwycCr9kL+
/VR+S8/7uswJzTVB2lsuYyHg60gl88Eu9LxdpW4jeCdpm9Dbxpx/F5j3KIYYhbxW
OXjOaBoES9lOgkgxGD7/Pdd52CIFeKhau4GFuFOxPaSGU87dXES5nJ12/CV3sIYI
9yeOUaMU9OqhtKVE6yo2cuta700Tv/VTS2u00RB/Wghx+fptt6EK5NNiXFW4fGUI
zIzCm+m6RVW/C8ajyoSYHupRbgsXXF3j8aN1/XI9TscfE2ssqmViCGkmGYQ9BHS3
carTF8ND6v2ZrHgm3GAe5HjaUQVWWzVuQp0AQdQaF5rbIpbfLopXV+6Y2A5LjW2h
hqWfeATOMx0FPlesJ0NAyoDp1FhiM7OHFchM3NEt2H7W9iuaeK3fzPv6yHXeRAD3
iSC7PWc3aSR694VJ/79Xv8Hja0DQ8dG9r8hfVuCGnc8gh0eluEsNfRih9TYbniWS
20rjAKJ/VJwYAIxtz36se56AEMeOq04ZQNhVcagsdHSt5I/EL7ICcLUw2tTamr5a
redtJHj4lxDb+Nwjf5zMjN9dK0bkS/2yTQiznS/oULK4z1lPixZJcNZAuVIsn8bg
Cr9tanfi6Yh3EvtXpoNrmISDPL3oLzzhZXWmAMrqaUEksBoEDSWZ+U2D+SDZ1Ifx
x9EucfV9dJOGtRe9yF3Y4TYrmK5QYI1FFaJQ2gNccoc3rYsdACBHYr2eq/h2D/rj
y1Ov+IGmngs/RBhmSlQsY/GxNr1prek0OqgR26ROWK+1uePrEDvVEwIma66L2a7S
v4Wr/4ViKb4UvzKG+bSCWjdcaGNbcWhg326zg8ijOrbYAr3laRywwZJCgu2dAQGc
7uket/nID5q4UhMb1cclTBbTqE9mZulWdehm65C4gbSoB7iFwJ9BcGexdB1KPajQ
DgvWZRlMXrcw0aF3Ig1AcoRfmAK6UPOjxC+meQkAzDXC/d3z4r4fctaoOahJ0H8l
h+q/Qp1c4unF5B7Ix5nY5vO01huOvUB40RoK9h9NXKFFg8vDskNqCfvw40M3aDth
zz6IFhW3V5MN+BIhO9+Q4xY+ROLB7kUDJdf2bUGgwG6fb2ta4ab0tr2pkzmboxJ3
Mge85Wie/zNjj3Qzfn/n5YGbeyxMPCcPUt6ZtjQYKzCRvom1GmSr/4rLaY7tV6cw
/ZadlWxEb1rNxZPNN9KMzduzO5Il4egwIlnWgxPI8iUbgeIp58nR+CAkhWgvVZxp
xIpEgZvKtGghpjIylayLL7kyik8v+mYW+b9eBNwfyVOGm8dDDawJbEGe/qHu5pRL
Aym6rbxESirZrobQfcu2Nuf+3uNxjU6SpNbJWS5etHf9ixVON3Sl6Umqk17rZeKf
NNIy7yDKCuSp4ELOePiWqg797VTxjlvkm1gCWgy2iQKtgdKrRrr/f+BAnDUqMy/A
QnudZEfDsVAMhhrnAwAguoSOOHu60QDtqfdmd29XjR5JCdv7ILkGRWo2E+2EQzQu
URHRxs62l6/7bW3FAgyVxTo3bhZjzxEh8Oe1YU+RyFjefJf66IW68zsDMIa1qARQ
bUNLh0WaqCu/0q8jEzGtNyU0IA+gVluFEugGtj+RDd5PTv6i4k6b2voJV55Aodq4
3oaVCekcMxDP/ki2M+7BCVZzPRqsE1upxgJhE7ocdwMqiOzBNJIlYpwmnilM7V1W
FrvFcwEn+QYZgOYL53In2cYzd4Jhv3acIGo/+MmWwZVfICxU3QjiDJSvRcxfe+kZ
CEI4oqeLuVOpegLcqjQ5gss9dsAuOVcgRdNMMwZpRS6Gj3zPzfDDmsqawmdJZnaT
OCWLNab8CLtChxTIpxd1RZDiC7rH7OCqZd/hw8D4cG0uFlNoDFXBokAwP0a8r9pN
YoRTE7RyGSps9xBRXO7mePupb6m9GdBu/A+4OHaXFPQs2kYxYUGuR6LDGbiKih57
zAG4qtf5eph2p78viKSjq94UVHyh9CDkNL/fUbTL7BBjGcH+DR4GtkDdtdILQFFy
MabNeoDer33ZisYT2jbKocIRLRtXpoI/xHt4vL1GhnCjfSfrwiSmLVWbb5VgtTS/
FQBcLmZ/san2bIG8LV4KVHz+NrzJgqAZ96FnjZoNzimNy+YdIcwQuAZCz7+ol9B4
ErVGY60Fx81l0xLrlOUX0Cm8knXhPimz0e2j2eRKVnMjQ/Wrz86WxyokS1yfDk9u
uWgjU61C9rPbKr4AY3bJvF/cKvOcByRQnWKaIJuIQ74XVCvBjMoHafkselTg+sox
Ly7078luJhpG0GqBceb/0TieCXx99bmDwmqdpXTv0mVRBWC5naR2EEUjgDCGRPfe
UocatwTb/KJt98DmfrHqZBdHYf5JQNABN3Q+CrNuRODWY+zoIshKWj3aV0LleMkg
QSzZVSO9ThkwJPySkM2qpvB91CPknuhMiRqBwOB4SkdXmRjFNKRvchmWbRRazKF8
fG3iQLfSB5IgdYtX52KNlQ3WrK3yU+szV6SQkWFhn+IBNg0ggmagUZMAseoqtZ7I
3GEldKxYCP6Q4Eq2L+4m8LABSxvylaikuX1R7neEM6YL6lpEk7sGJrAf7FkobF2L
SSvHWqalGOCmvIeQkM2hMsqWIJyZPk/PPAZ3CGwN9QesGHHQi5+yd2YH6O1vAnf3
WHaBeSoN59paxb2Tj9L61lSXCXmlBiBXXMinjo0Y6Cimc2EMPDPiCOkA3HI6fdsF
dTph1UYtJttYD9Q6aFGOrtwlKiOatdViNHOQ1ZbjtoucuHiD5yDX5yQglEtm8Vr3
M9eNdc0cDiVPqoC+T7l283e16Pj3rJjivM6Twv36I/OiVZiaTEU7j7pcHyLD5hrf
bplAGASG/fGLK9FcB/50wpKzLGS0pRSiQ3Eoo0Zm73rMQqny2JcMmofK1QHWJKvC
wJ5EfJaqbu2zx4Ew7GKkQQvMCq5pN6dMEC66Z1WLqcm0lYQBdPIpY7O0/b5+63Ho
hphH0sqMvSDT9nnOCqav2uHgA4uQEeu1N3ekWlRBzx9g2grptG3AJ16mf/AbTluo
hazr7hIPR27E2rVkq8F0kVACWY7jD/22hR4w2jkWJDXDyEfIAvrhyQ2vFvYYdLU1
KZ4oWAD2s9pv/6RCxR+xmV7GCBNI8kPq7S7hC47oAHHUE6/31PDiCkGSFtYpINPS
eYpdEgRybmhkC29yfp6l+PcYZUcgU56GVFthb0B9QtCw9AFfef3q9ORPHGLLV7K9
CMrBdR1mifJHvKjmEJdNuQinLfx++8wSknEdXBwqPwF6HoAvHvcycuWat0ZYwX7M
DTmyerkR9kCyKHuCYrYjS+8ZHJbUEboNC0XC+f5bCf5tqeBwZI71dC2TeUmgBhQQ
rLLfLWyTF//FUsJN/wj/PcDU58+iNIwquo1SBCE9v2w032RFJJ5YRKYoNqyg7kve
EJ75S5XxFS8sHJzVAru4aIqVQk61MDp2ZqVrI35mr6n1ZONMcxts4nfUvOx0ySfN
wSCdbAPPP40nQAtrCn6WyJRl+4OhXECuS6kJXRWujTnJxkDz98ejPF7B5xsN1WUg
ZEQTwa8Jrj5kUVdJ9SoOV3qsjhkIyk85h1ARqyOfQUdz4hLgm3NgsA/V/jKiRtDG
hdzokzqOuFB7a9P3lMCVAd0OnHByU+bnGcnzEgNNzfiH2esWsSmzs7YefHEw2MLE
+X9qj/13QIkzNYTnX63XXZBnYmOnFQBhBbDKiNL0DGpIa0KrrB3p6eQ1dCyFruxK
DWE4bhjF/xSGWJ/kAX2OmSuVyKo0tEQD2ndNFKVkXbdHOFTMZWbHvXV6xirfXl1V
BbwQaYYLWTarbPj5FS/rQ6dT37bP7qaFEEmu2zoHjJXVqQ8v07+249pn5WFIkHE6
NJrXbS+bOeaFPnDSmstO5xPHyBVgcw5V1MH8H0Vjn1/+q0+ZhrZ/EgnE0hF9iAvn
u/shZ6SOtYebCjLPK53ydEgJGOxscq3wypCZGWDK6tG5pgxJ2OZuTs4DPQBF/OFy
s8g928jxG4swpQrc0J5Glb+9Y+B5ZfmP44L6tI6bdQkTwRZlgJXm3QcpB8ZmtuwP
27EtNWmoEaxGx4rQHMRbtdeMK0/uo4eTicg8IM8evk8+glit5pfNPaNNinZ52mip
kFR+I75Pwhx9jd379hq0le0SWHYbEo27V/aDm1lDiR6rK9Bwe/BRGEi7R+L+5i05
P5i1zOo+fxEk+QQCg/D5QKoDGC+4A9Ba4M3m0yURXX/E6wihAd+tED2Biz5UwT+z
Fg8re1q2JiZGc5U8hCzZbw==
`protect END_PROTECTED
