`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LTiProTq4ZmO/GsqIJdln/L9rc98d227dcbPlN7dGS3HzqyEHJ9luC3iO7XPD0/E
Xvwh7mudBVp6DnX6qjNwAECTDNWRsVe4bKGk1dIgJ/2DjeUgFjnUmIGSiVmKacyt
7C4Ym15o2gY1xOGF9LBynjVCtV5/h6QX1MJqhbyO1w7zon/sd4A5LZsvmoVFNX9A
0EqDb4Z5yAmG2MEOx48P9Te+sJNqKShdeGjRwOp4gX72EPIIspC9qH9lLc/iKcW6
hPiU4jQ8KD6P0WCnD4KePKuINa0xr5es9hlAIyFHnD856if6fsEHpUCq/Hd9khwR
H/TMO6pZSfXvjzxkeyHek0WI6Jr45rBoCBSuvJc8An2mwoOnCD/B3pAIRhgUAihh
fL0hZ4ExULQ8rjgErPGvJdth60akh+YrFv7+8hi39W8krwR9JQ4/uJFrRKYkdzyj
o+swRklc8HuRU+KWN0fWK1KOfq/pnX7qFypXcyHVDWA=
`protect END_PROTECTED
