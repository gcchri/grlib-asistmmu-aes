`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3qfRaCkKgT1DuYfBFQeumq8K4Eu1SSGv5l1iusNgxVkU7dbFsEprROFYINPquNG5
A7SURJ6EgmdoQo29oi/ciaxXQtorI/6W5yvcbJFXGNbVwU6B1NbDfvinL0zk9ud4
tSGIw1erd6HUT7Mtgih5QpCMyHAYOqUoQer9W2AxpgJx1TLK7Y0zapsQ+WbDbn1v
KXxvF6JZyUEdYg7yM28SoSAms972TRTJ+AA53YQhk4wAmzQ0V+evZQWqo/L2bNsM
Qtyxfr/mJi27LoUkwK1wfPtgVOqPxkkC0N5zxOFZK9xGqORyU47dKHVnUX0XAo9D
s78aX64HlkdbgHMJFXT5iKieYLPup3PBEj6ebybuxxpp33yQItaq6r5GeWCmbXoZ
umbOpD46kbYkth9JsB2EiZA8aFbQOehTKKEUXudSw7rstYTKI2KyOerfoDLBbI60
JnsUjQKMlYnCeLAO6K5SynIw4FJxzlivWUjFK6ooVlQaO8ifZlVKC1MhKhCouHSa
Aa05spQ2hyVPeoFw4M5RnPN7c3IOjhCrdj3DISYEE4FtH0qk0R53osTbs2mozI3+
+zcv8fdyKabc2chMBGKYBwsP0x33askZrhb40zLrEUC/bomwA2jSs9ep9w7VWMtc
LiOv70Vq3MmVv5M3DqWiJvMvcbjGKuy9Ny7cj6lclbHHiIeG0q8+ZkvOEsFa4Ve4
BDhL7TQoTeDtnVmDK3IroOZXyRUDU9GNTDXQP/NmG6eO44TnAg06V/lsbpglANWU
S702yWHhKYb4s1pyZUyH6QSOeal/7LkQTzkZwQ4rlgmtqaNgvVJirtQprgddjrBe
BvGghjlu70gla477v1u0xE7fmsm0+j7n+OSj0559JpjzZZt550sQBcqb/tXKH7Qj
znuhJlQKFEN0T2I9eAUv6MxwD5F1jZYywqaoNTvR9NQEd9qcpuDQmMFblngMwHEX
aFFDQgSo2vIjBtM4Q12kl40823DoGC4Yv5+YKuGlSLZWpND4CjVRUD5A5TMygic/
DbUVxCbc9PXpXdKiWVvN1K1bFnjfDL4DSQ8EEksWiJG+oLGfree6RC0Hk3YkzQaw
iM0GUTWFusEwivY829QfqqCTHWxq3FM8aHrNFJu8pAb1jz37Y7G+GA/Pl51BT1sY
eVujeSnhxRakDskBC/cjaQM8FoomBBey+ujQ+nHfVPjT9BGLfnQHnGWZ66hSEDUu
eJQ/VAnMFbskqxPazIBm6D8wrhnIPiRVMmzximEO2gQQRbY1cu8AZYCYeZ7KDSbc
33JZ1fSvoZe/y++Nu2IYWG+robBdcrgk5mlywDQPesMdQKvc/ZM4emhw5rLMwFmV
ccBkvc8+1B3S6lFwPz2CqKtF/zXpegs5pWRzu7OCW5KCjkQfrEEO/vLTFrUDUyqT
hHM+WqDyMN7YuzDoO0WCQ8LE2inw01LhDPhIIrLYqvSW1yfGmNj/KSwCbTCu6gKe
cpc3U1rzUmqBVZGiSnJVB4fIsODaNSrb4Lgq6faQ3gDt+czeE35fmj4qGSyIY3oE
dz1PS/xePyNd5Gd5UTvzpeb38I8JE3lWFfVgRBQX4zzz7WVjjpoq0sWIrSfAMg3V
KEO7AqCbMzjdYfj6ibxL101PtxvwFlBlzLmfObWEdeajH02w8OFc7a7xYiqAfu6u
GmKYg5xA7hhQahQOyrQDZqVczr5uGcP/SBqQ7+tYbSusKj4W6bT+MZ3idikrlfkH
efIOTrb5BlPlXVjMjWos5auotS2456iH+yPF023C3E44Uackpr9By6S/pyM/H/Hz
WDFY/n167bGso3J+x9CAGSrAQukUiaQM4CmKEMrYprTwOoVnK56qDEdSHzS8xL4y
1WvHsQ/o0EPyI/4fE/Kd2Ug96Sn89xvUFFxdgzSeuUI=
`protect END_PROTECTED
