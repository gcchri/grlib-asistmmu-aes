`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
moQld5HSVxcagsswEaWizQ51Z70iTAFi9EP+lAzJnuTizWq76rLHirq9wNc9Q6uN
taEm7QxOctheUn9OR/gUSXHZpfCuZ1MYaH2SujoXNfHyegM5H+51dDyUn1wc0lAJ
9xXHpZiM1s9l8hyWOMvKR/HTLZYMxY+NhjX6wa9AnRKiSQxtY+3gQx7wOnf4WrDP
z2GtXc0r+lq0Mct4IEaQQErgscn581iqowotVftbcOeU8ckpdkqrAOd5EESdadS1
z/NfW2rZFnuMEfhqUju2/zS+vaaNzVhAczA2yE7lxM4=
`protect END_PROTECTED
