`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3YAPWgFrofHU75UYLJ/c0gPBdGVoxzfUgr+TdMVzwkZkNVp1ylvE3qW6EZGqE+qe
f6LbIOIz8xuWaXVgSWpjRdsn3TYqDWiwgjKtRduvmE8kePSeWk/pqgd/gR88J/d4
3RV3H/CqQeq3eV9mpGU8VIKKQNYiqs1KHOl7En6RSMz8s62ZdF7weVilXtC/UwBU
5RDkquZd1+/n86g3qoXeJyleIh49ykO59Fr74x8pSGH/t430nwHi14kSEytHPYb1
ad0Z7SKiwK+iG25sXnKq0esBqQbz30svmnzMzGJBRMoLaR/Ud/RuPmAWTt8k8VHn
RUuiWmzQzMAUj2RqbRtyXs3EXcPVyljumhwbBVkMP8yAT5JvwtQct67d3rs21efe
Snann5R5XHDqfC+lpPF+OELN7Sv3jq+YqQ4Ne2vq2nhB/tR4PLuaX7bMRHnYIpAB
y2djZ/gU7dKKpJ5mss1Rpw1CVBj+3KQxW36fPHICsMF2Z36aEgUZRWWZBrBypMZ9
s+mRTEvQXXzEhw6sHfPEK9j065ZLMtKaSpJsXL0T1cZcGWHa000Foe+OkNtBKIkZ
+vKwhC4eXMd6GHTepbYeMg==
`protect END_PROTECTED
