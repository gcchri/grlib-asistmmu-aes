`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aYlSVXNfjKGUfFII8is+wHf60mdfch3eba5z+IlaJq5jgkHs9um0x14MUdbb44rz
lS6XYH1PgkCQ1SxH83Bbr8IdGFD99rUTZBsK/QKuIsXACR9ElisUsdUBTte25jaM
Bvt/ZbFSPw+YYY/nQ+HGs36fdsk2jMDKxnQ0b61dzUphwJ6FThqMu5SwVBoorRLz
msaBm8yJrm8ZhW3F0SZdxSk8F2ylLvylcbxnLeRAeDvS2aWUhUU60hoPVkJDG53A
VdkzBzKAeBFx4IoYeGZZMCbNawpeOBCLdKD1pUnmrh9EsgrH3j4Ee3pt2URXyjbn
Rbfmcn7NEIvxmEDZAD4fJzl2wnTtsvuw7Aubn1MKQ+Ewzh0S3PRYAm/O7lMhqF6Z
INWUO3PDtFeCBkykJCp2kRhlzCa82nLNCMS3AVOyuDM3Ken/7S6mHZxiN7o47MKt
ZLBf4DHBCDA6avINLtSYQofioeQTl/fKXfop+G8L+OFqq9eDod3a/nOfBq8OhZ48
pweSRqyVGPJ9yOMWTyGio+YRRoL+FcDEHqbUfyyhLGoQvolw/+edewb2sfeXuxmV
asBeVxOk0x9Yban9E3u4RA==
`protect END_PROTECTED
