`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eyFYwB7ZuHQcx23dT6UgKmz+uA70WYUdU3+wANpdx5VNBp95hRh/gw7vUEljOLE6
aKK0a8HXIXheFD9ScpTCsgUQb/Y8jzRDOfc631LgG1bvSSWNU28af6JwnPv5ZG+G
YACBV8jPONVP9YMCEKjb5VSnGvEp4fth63t/+5EMn3wdlRUJkfrAaup1aV2FPMPI
dPNOYLfCEa8D8Tvl7lehtAWPefDyzQF4ggv/6Hjq2AvGTFRzcs4nDF2uGNkBUjNR
gxbVFx/vJcHQej2FKk6O2ycmJHRZuKn+iOCgkYVBeWmTjkIG07iwcDng8o/bSpTf
9o1cYpf7QMCLvVcX/Dww2lA/Q6wdSIM5Ckk3ZVYkLf+cB8hp5LBd/Mpfmrmf+O9V
`protect END_PROTECTED
