`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zJrzuxXegh0LvoR3vP1+5v3qv4IUta2sliUaU+bx7qJDCnvFFHjJJd+Zzu8sXO8J
+8utd5IJK1HrDgI5at04Ifo9qw+n8yaBQyPPYsqiixrp3pJ+KYcKLT15FcY8/RVC
D1G6/d2bvl8O9u8bJH0fMhmSZ6C/EEjIxMp/GSczOyHQec6oDIfE9bv9fT1+V4LI
nyryGYr5Q87txvUHQpqme2Q/kiSLGajk/hVtJRRYOakqfMg+aaPDtPjFqGcmxNuW
XzDxzAXAZ4X4wL80kiIlK7qid5AYZ6YagBeTh4enE6BsLn7T/k9v0kxMxws+ZYyI
k0TjwX9EVZeqmUQeCfPgF0ohPbq+K9+XSDWOxC+0+n+lFTBFbhoHypwn67puXdw1
6r2+LmQOa6dB+12fTZWsLOWkcCCRT3u80Ju+JSHVB5R582QU2XrpQIS2nKB3zhXO
1/Gr3na7HC5UAmI8+CfJhnsRTpyaGs+TOhfy/vSXcYOBnTMXUgZcflNzvQS4phkL
ecHOBtZUtVGmk+9D/+nPtyGCaaMlxeEgIqmnh9bPY9wkLDG6ocqB25ZiO/JD6qUJ
nU7cjgngJOgP3aGFMuq9Bi6MT2Ntr3Y5lQnqhuL0F9y/gBWjORIid2r+oETgp52L
jkVzqlNVQ8Pj3Vnz9/8uQLVATnEqqrOniuqPqjzbtOq2Wq1Oq8mS+7y1muihAGTY
qpny/hHVRFfBgtJNQu9ynUElfLAfAWKwci6Ohynhvbob6fJ/O8EqcYZmrrNVIb6G
zTMSlvFzaQ2+yqZz5mxV95+lBs6sjgAcKhUoIRuXeKMR0+yNOIJrD13UUjkpuF9m
0wYKfLKwAFPyhqye7TmaprOcmg4l8KeI7A+YpMgv5ocDMPkN3YzeJ0XfanlyjzIa
vWQvNVjGIVGPsj1idAcP2GfJHRY09+TRZ07Vx1uI4zIK9sSayobUmWQ1O0AUXgDR
SwYzL3QQ50XYi/g1mXyIYo0pstEyMVv5OVIy14Q/zcLRyW3QN8ERdcRgrb5zrBnA
muvkqgJOyEsJxg/mvJLHC1eE0lFXh0YSBumYAMbgZJuanHDtYhPP31b7Ro91T49f
OsfdDjEr2MiNl8pcZqO2lG2Om02tW6ewWOI9eL2QjymbIuYtZccX5zbETmWm6PAm
oV/ultnL8I7fUsoL1ZfT7QHHlEnb6DaMsUGS6cqkPbzmO8cPKL2NJP4jO/zIb5ac
Ohr5kNGE0i+0jzymkNnYmLPHfoT9GjRUY/CdGdT5bX2asv3cy0qnKaRuZJZlIaZb
5SITwEi6rmFUj/5oH6AZBpioc3zLBTqal+aR3JtgHkqwy6ydAHmQmojww6KnNWJ6
L1PFrmK3DyWgUb0/XvfNmE/6aWAKqlv6g+w4VABJHlTT6X4e6djjJCyGSaXrB8yB
FnYRozWU1k4Tnzwt5N1tZaxakrMHp0iglVr1vqLwMJnRdkj/2O29XhTp/MeXevaL
R5bzc1Zh6bQvAeNNUrbt2/yxeWtY7XxMrInp77phUTS2ohZjNHjOhnUG5UnXpBG+
uOu8mg6bkSb4ilwE+D/gDSH6+GJMvbLuLfNEWLPZdEjeW1YsFbZtRE6LBZs8QLm6
N1iZICYmuaFLedFZFWSD8e+oEiV9A7SFoQdVv13LjK/gcWOl7Dw0wizy1kmJutdg
A3FnWkh0pOe5N/ykm/LLFEpPTfqlWwuNiw4hDu4mLJZVDv0HguI3XnmhkhEJqZoF
7ca/Q4k1ZGpHQhn9E2W+RojZi/Nk89uPRyilho1ORJ1gEUU2XQYfS7WvDc26F3Qs
en1/b9n0er1vBfxhbsCDZgUSHGKHOXo33y525nrPLomxJHjamjGG01Nb4heroNCg
gTI9fl+8u3zYqNNOHF7nsA==
`protect END_PROTECTED
