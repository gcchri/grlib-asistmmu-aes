`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BZIEJsFlZCfdHjlM7JZdo6v4NYCK3IT4LpIeOnX035WvEQaBaBragwgQ0UZVdLRd
G8eQmcyj6gyRsq9aji//n1eFR4fqt2cHbhcnBBPQkK7EdOrtMrWVZJ1J5S5CEoJY
8XaL9dCfoPgFLfGAEKU3nfSkKxpy+urXxZTPsXaFvi/RvttwozVuBqRtE94RIlOB
cYqI4PBTEkeVvxHCKOLpuw==
`protect END_PROTECTED
