`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qDihPndqnkhv1T3/ljO5W5bxAQTsGRs10YzPDd8XIiKHiFZpICeLWVVYEhvzrlt+
Hr4Tqz5B8UUyYwCVDcALj/nca9G7zOElbuaF5jGQytL4D6EsOLC5HsHjcFS5NvdW
Kj8ojoFPNGv1te7DeSMYJcfa7eex0R92QooqRjGAE5DJxPR/DUF6qnA6RApIFjjE
qryAYCC32xB1o7gCktAbvkG031dG1oNGpKs3cmV4QsWJE4voHHhKQUjRA/aMegOG
hPtOzvrozCzDTTpotW+sWHqRiGCNggrmRrEy1eGewemUvFPM0x3xGmuOOOgGGvKH
npb7io+cKefJfX14aUpMfHZhVzC9OSGC1RIqG2yucaWx5du9kzQJb9hAXJljwY9A
sSAiBRt3xSJeB/8ZuO/LdSZpri/t3q1+Z/nJLYEQTlj/qPGiH5T13OKdfC6OaNy2
`protect END_PROTECTED
